module bar( \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 );
  input \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 ;
  output \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 ;
  wire zero , w136 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w146 , w147 , w148 , w149 , w150 , w151 , w152 , w153 , w154 , w155 , w156 , w157 , w158 , w159 , w160 , w161 , w162 , w163 , w164 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w174 , w175 , w176 , w177 , w178 , w179 , w180 , w181 , w182 , w183 , w184 , w185 , w186 , w187 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w203 , w204 , w205 , w206 , w207 , w208 , w209 , w210 , w211 , w212 , w213 , w214 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w224 , w225 , w226 , w227 , w228 , w229 , w230 , w231 , w232 , w233 , w234 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w250 , w251 , w252 , w253 , w254 , w255 , w256 , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 , w2495 , w2496 , w2497 , w2498 , w2499 , w2500 , w2501 , w2502 , w2503 , w2504 , w2505 , w2506 , w2507 , w2508 , w2509 , w2510 , w2511 , w2512 , w2513 , w2514 , w2515 , w2516 , w2517 , w2518 , w2519 , w2520 , w2521 , w2522 , w2523 , w2524 , w2525 , w2526 , w2527 , w2528 , w2529 , w2530 , w2531 , w2532 , w2533 , w2534 , w2535 , w2536 , w2537 , w2538 , w2539 , w2540 , w2541 , w2542 , w2543 , w2544 , w2545 , w2546 , w2547 , w2548 , w2549 , w2550 , w2551 , w2552 , w2553 , w2554 , w2555 , w2556 , w2557 , w2558 , w2559 , w2560 , w2561 , w2562 , w2563 , w2564 , w2565 , w2566 , w2567 , w2568 , w2569 , w2570 , w2571 , w2572 , w2573 , w2574 , w2575 , w2576 , w2577 , w2578 , w2579 , w2580 , w2581 , w2582 , w2583 , w2584 , w2585 , w2586 , w2587 , w2588 , w2589 , w2590 , w2591 , w2592 , w2593 , w2594 , w2595 , w2596 , w2597 , w2598 , w2599 , w2600 , w2601 , w2602 , w2603 , w2604 , w2605 , w2606 , w2607 , w2608 , w2609 , w2610 , w2611 , w2612 , w2613 , w2614 , w2615 , w2616 , w2617 , w2618 , w2619 , w2620 , w2621 , w2622 , w2623 , w2624 , w2625 , w2626 , w2627 , w2628 , w2629 , w2630 , w2631 , w2632 , w2633 , w2634 , w2635 , w2636 , w2637 , w2638 , w2639 , w2640 , w2641 , w2642 , w2643 , w2644 , w2645 , w2646 , w2647 , w2648 , w2649 , w2650 , w2651 , w2652 , w2653 , w2654 , w2655 , w2656 , w2657 , w2658 , w2659 , w2660 , w2661 , w2662 , w2663 , w2664 , w2665 , w2666 , w2667 , w2668 , w2669 , w2670 , w2671 , w2672 , w2673 , w2674 , w2675 , w2676 , w2677 , w2678 , w2679 , w2680 , w2681 , w2682 , w2683 , w2684 , w2685 , w2686 , w2687 , w2688 , w2689 , w2690 , w2691 , w2692 , w2693 , w2694 , w2695 , w2696 , w2697 , w2698 , w2699 , w2700 , w2701 , w2702 , w2703 , w2704 , w2705 , w2706 , w2707 , w2708 , w2709 , w2710 , w2711 , w2712 , w2713 , w2714 , w2715 , w2716 , w2717 , w2718 , w2719 , w2720 , w2721 , w2722 , w2723 , w2724 , w2725 , w2726 , w2727 , w2728 , w2729 , w2730 , w2731 , w2732 , w2733 , w2734 , w2735 , w2736 , w2737 , w2738 , w2739 , w2740 , w2741 , w2742 , w2743 , w2744 , w2745 , w2746 , w2747 , w2748 , w2749 , w2750 , w2751 , w2752 , w2753 , w2754 , w2755 , w2756 , w2757 , w2758 , w2759 , w2760 , w2761 , w2762 , w2763 , w2764 , w2765 , w2766 , w2767 , w2768 , w2769 , w2770 , w2771 , w2772 , w2773 , w2774 , w2775 , w2776 , w2777 , w2778 , w2779 , w2780 , w2781 , w2782 , w2783 , w2784 , w2785 , w2786 , w2787 , w2788 , w2789 , w2790 , w2791 , w2792 , w2793 , w2794 , w2795 , w2796 , w2797 , w2798 , w2799 , w2800 , w2801 , w2802 , w2803 , w2804 , w2805 , w2806 , w2807 , w2808 , w2809 , w2810 , w2811 , w2812 , w2813 , w2814 , w2815 , w2816 , w2817 , w2818 , w2819 , w2820 , w2821 , w2822 , w2823 , w2824 , w2825 , w2826 , w2827 , w2828 , w2829 , w2830 , w2831 , w2832 , w2833 , w2834 , w2835 , w2836 , w2837 , w2838 , w2839 , w2840 , w2841 , w2842 , w2843 , w2844 , w2845 , w2846 , w2847 , w2848 , w2849 , w2850 , w2851 , w2852 , w2853 , w2854 , w2855 , w2856 , w2857 , w2858 , w2859 , w2860 , w2861 , w2862 , w2863 , w2864 , w2865 , w2866 , w2867 , w2868 , w2869 , w2870 , w2871 , w2872 , w2873 , w2874 , w2875 , w2876 , w2877 , w2878 , w2879 , w2880 , w2881 , w2882 , w2883 , w2884 , w2885 , w2886 , w2887 , w2888 , w2889 , w2890 , w2891 , w2892 , w2893 , w2894 , w2895 , w2896 , w2897 , w2898 , w2899 , w2900 , w2901 , w2902 , w2903 , w2904 , w2905 , w2906 , w2907 , w2908 , w2909 , w2910 , w2911 , w2912 , w2913 , w2914 , w2915 , w2916 , w2917 , w2918 , w2919 , w2920 , w2921 , w2922 , w2923 , w2924 , w2925 , w2926 , w2927 , w2928 , w2929 , w2930 , w2931 , w2932 , w2933 , w2934 , w2935 , w2936 , w2937 , w2938 , w2939 , w2940 , w2941 , w2942 , w2943 , w2944 , w2945 , w2946 , w2947 , w2948 , w2949 , w2950 , w2951 , w2952 , w2953 , w2954 , w2955 , w2956 , w2957 , w2958 , w2959 , w2960 , w2961 , w2962 , w2963 , w2964 , w2965 , w2966 , w2967 , w2968 , w2969 , w2970 , w2971 , w2972 , w2973 , w2974 , w2975 , w2976 , w2977 , w2978 , w2979 , w2980 , w2981 , w2982 , w2983 , w2984 , w2985 , w2986 , w2987 , w2988 , w2989 , w2990 , w2991 , w2992 , w2993 ;
  assign zero = 0;
  assign w136 = \pi077 ^ \pi128 ;
  assign w137 = ( \pi077 & \pi080 ) | ( \pi077 & ~w136 ) | ( \pi080 & ~w136 ) ;
  assign w138 = ( \pi128 & ~\pi129 ) | ( \pi128 & w137 ) | ( ~\pi129 & w137 ) ;
  assign w139 = \pi078 | w138 ;
  assign w140 = \pi079 & w138 ;
  assign w141 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w137 ) | ( \pi129 & w137 ) ;
  assign w142 = ( w139 & w140 ) | ( w139 & w141 ) | ( w140 & w141 ) ;
  assign w143 = \pi073 ^ \pi128 ;
  assign w144 = ( \pi073 & \pi076 ) | ( \pi073 & ~w143 ) | ( \pi076 & ~w143 ) ;
  assign w145 = ( \pi128 & ~\pi129 ) | ( \pi128 & w144 ) | ( ~\pi129 & w144 ) ;
  assign w146 = \pi074 | w145 ;
  assign w147 = \pi075 & w145 ;
  assign w148 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w144 ) | ( \pi129 & w144 ) ;
  assign w149 = ( w146 & w147 ) | ( w146 & w148 ) | ( w147 & w148 ) ;
  assign w150 = \pi065 ^ \pi128 ;
  assign w151 = ( \pi065 & \pi068 ) | ( \pi065 & ~w150 ) | ( \pi068 & ~w150 ) ;
  assign w152 = ( \pi128 & ~\pi129 ) | ( \pi128 & w151 ) | ( ~\pi129 & w151 ) ;
  assign w153 = \pi066 | w152 ;
  assign w154 = \pi067 & w152 ;
  assign w155 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w151 ) | ( \pi129 & w151 ) ;
  assign w156 = ( w153 & w154 ) | ( w153 & w155 ) | ( w154 & w155 ) ;
  assign w157 = \pi069 ^ \pi128 ;
  assign w158 = ( \pi069 & \pi072 ) | ( \pi069 & ~w157 ) | ( \pi072 & ~w157 ) ;
  assign w159 = ( \pi128 & ~\pi129 ) | ( \pi128 & w158 ) | ( ~\pi129 & w158 ) ;
  assign w160 = \pi070 | w159 ;
  assign w161 = \pi071 & w159 ;
  assign w162 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w158 ) | ( \pi129 & w158 ) ;
  assign w163 = ( w160 & w161 ) | ( w160 & w162 ) | ( w161 & w162 ) ;
  assign w164 = \pi130 ^ w142 ;
  assign w165 = ( w142 & w156 ) | ( w142 & w164 ) | ( w156 & w164 ) ;
  assign w166 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w165 ) | ( \pi131 & w165 ) ;
  assign w167 = w149 | w166 ;
  assign w168 = w163 & w166 ;
  assign w169 = ( \pi130 & ~\pi131 ) | ( \pi130 & w165 ) | ( ~\pi131 & w165 ) ;
  assign w170 = ( w167 & w168 ) | ( w167 & w169 ) | ( w168 & w169 ) ;
  assign w171 = \pi093 ^ \pi128 ;
  assign w172 = ( \pi093 & \pi096 ) | ( \pi093 & ~w171 ) | ( \pi096 & ~w171 ) ;
  assign w173 = ( \pi128 & ~\pi129 ) | ( \pi128 & w172 ) | ( ~\pi129 & w172 ) ;
  assign w174 = \pi094 | w173 ;
  assign w175 = \pi095 & w173 ;
  assign w176 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w172 ) | ( \pi129 & w172 ) ;
  assign w177 = ( w174 & w175 ) | ( w174 & w176 ) | ( w175 & w176 ) ;
  assign w178 = \pi089 ^ \pi128 ;
  assign w179 = ( \pi089 & \pi092 ) | ( \pi089 & ~w178 ) | ( \pi092 & ~w178 ) ;
  assign w180 = ( \pi128 & ~\pi129 ) | ( \pi128 & w179 ) | ( ~\pi129 & w179 ) ;
  assign w181 = \pi090 | w180 ;
  assign w182 = \pi091 & w180 ;
  assign w183 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w179 ) | ( \pi129 & w179 ) ;
  assign w184 = ( w181 & w182 ) | ( w181 & w183 ) | ( w182 & w183 ) ;
  assign w185 = \pi081 ^ \pi128 ;
  assign w186 = ( \pi081 & \pi084 ) | ( \pi081 & ~w185 ) | ( \pi084 & ~w185 ) ;
  assign w187 = ( \pi128 & ~\pi129 ) | ( \pi128 & w186 ) | ( ~\pi129 & w186 ) ;
  assign w188 = \pi082 | w187 ;
  assign w189 = \pi083 & w187 ;
  assign w190 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w186 ) | ( \pi129 & w186 ) ;
  assign w191 = ( w188 & w189 ) | ( w188 & w190 ) | ( w189 & w190 ) ;
  assign w192 = \pi085 ^ \pi128 ;
  assign w193 = ( \pi085 & \pi088 ) | ( \pi085 & ~w192 ) | ( \pi088 & ~w192 ) ;
  assign w194 = ( \pi128 & ~\pi129 ) | ( \pi128 & w193 ) | ( ~\pi129 & w193 ) ;
  assign w195 = \pi086 | w194 ;
  assign w196 = \pi087 & w194 ;
  assign w197 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w193 ) | ( \pi129 & w193 ) ;
  assign w198 = ( w195 & w196 ) | ( w195 & w197 ) | ( w196 & w197 ) ;
  assign w199 = \pi130 ^ w177 ;
  assign w200 = ( w177 & w191 ) | ( w177 & w199 ) | ( w191 & w199 ) ;
  assign w201 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w200 ) | ( \pi131 & w200 ) ;
  assign w202 = w184 | w201 ;
  assign w203 = w198 & w201 ;
  assign w204 = ( \pi130 & ~\pi131 ) | ( \pi130 & w200 ) | ( ~\pi131 & w200 ) ;
  assign w205 = ( w202 & w203 ) | ( w202 & w204 ) | ( w203 & w204 ) ;
  assign w206 = \pi000 ^ \pi129 ;
  assign w207 = ( \pi000 & \pi125 ) | ( \pi000 & w206 ) | ( \pi125 & w206 ) ;
  assign w208 = ( \pi128 & ~\pi129 ) | ( \pi128 & w207 ) | ( ~\pi129 & w207 ) ;
  assign w209 = \pi126 | w208 ;
  assign w210 = \pi127 & w208 ;
  assign w211 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w207 ) | ( \pi129 & w207 ) ;
  assign w212 = ( w209 & w210 ) | ( w209 & w211 ) | ( w210 & w211 ) ;
  assign w213 = \pi121 ^ \pi128 ;
  assign w214 = ( \pi121 & \pi124 ) | ( \pi121 & ~w213 ) | ( \pi124 & ~w213 ) ;
  assign w215 = ( \pi128 & ~\pi129 ) | ( \pi128 & w214 ) | ( ~\pi129 & w214 ) ;
  assign w216 = \pi122 | w215 ;
  assign w217 = \pi123 & w215 ;
  assign w218 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w214 ) | ( \pi129 & w214 ) ;
  assign w219 = ( w216 & w217 ) | ( w216 & w218 ) | ( w217 & w218 ) ;
  assign w220 = \pi113 ^ \pi128 ;
  assign w221 = ( \pi113 & \pi116 ) | ( \pi113 & ~w220 ) | ( \pi116 & ~w220 ) ;
  assign w222 = ( \pi128 & ~\pi129 ) | ( \pi128 & w221 ) | ( ~\pi129 & w221 ) ;
  assign w223 = \pi114 | w222 ;
  assign w224 = \pi115 & w222 ;
  assign w225 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w221 ) | ( \pi129 & w221 ) ;
  assign w226 = ( w223 & w224 ) | ( w223 & w225 ) | ( w224 & w225 ) ;
  assign w227 = \pi117 ^ \pi128 ;
  assign w228 = ( \pi117 & \pi120 ) | ( \pi117 & ~w227 ) | ( \pi120 & ~w227 ) ;
  assign w229 = ( \pi128 & ~\pi129 ) | ( \pi128 & w228 ) | ( ~\pi129 & w228 ) ;
  assign w230 = \pi118 | w229 ;
  assign w231 = \pi119 & w229 ;
  assign w232 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w228 ) | ( \pi129 & w228 ) ;
  assign w233 = ( w230 & w231 ) | ( w230 & w232 ) | ( w231 & w232 ) ;
  assign w234 = \pi130 ^ w212 ;
  assign w235 = ( w212 & w226 ) | ( w212 & w234 ) | ( w226 & w234 ) ;
  assign w236 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w235 ) | ( \pi131 & w235 ) ;
  assign w237 = w219 | w236 ;
  assign w238 = w233 & w236 ;
  assign w239 = ( \pi130 & ~\pi131 ) | ( \pi130 & w235 ) | ( ~\pi131 & w235 ) ;
  assign w240 = ( w237 & w238 ) | ( w237 & w239 ) | ( w238 & w239 ) ;
  assign w241 = \pi109 ^ \pi128 ;
  assign w242 = ( \pi109 & \pi112 ) | ( \pi109 & ~w241 ) | ( \pi112 & ~w241 ) ;
  assign w243 = ( \pi128 & ~\pi129 ) | ( \pi128 & w242 ) | ( ~\pi129 & w242 ) ;
  assign w244 = \pi110 | w243 ;
  assign w245 = \pi111 & w243 ;
  assign w246 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w242 ) | ( \pi129 & w242 ) ;
  assign w247 = ( w244 & w245 ) | ( w244 & w246 ) | ( w245 & w246 ) ;
  assign w248 = \pi105 ^ \pi128 ;
  assign w249 = ( \pi105 & \pi108 ) | ( \pi105 & ~w248 ) | ( \pi108 & ~w248 ) ;
  assign w250 = ( \pi128 & ~\pi129 ) | ( \pi128 & w249 ) | ( ~\pi129 & w249 ) ;
  assign w251 = \pi106 | w250 ;
  assign w252 = \pi107 & w250 ;
  assign w253 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w249 ) | ( \pi129 & w249 ) ;
  assign w254 = ( w251 & w252 ) | ( w251 & w253 ) | ( w252 & w253 ) ;
  assign w255 = \pi097 ^ \pi128 ;
  assign w256 = ( \pi097 & \pi100 ) | ( \pi097 & ~w255 ) | ( \pi100 & ~w255 ) ;
  assign w257 = ( \pi128 & ~\pi129 ) | ( \pi128 & w256 ) | ( ~\pi129 & w256 ) ;
  assign w258 = \pi098 | w257 ;
  assign w259 = \pi099 & w257 ;
  assign w260 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w256 ) | ( \pi129 & w256 ) ;
  assign w261 = ( w258 & w259 ) | ( w258 & w260 ) | ( w259 & w260 ) ;
  assign w262 = \pi101 ^ \pi128 ;
  assign w263 = ( \pi101 & \pi104 ) | ( \pi101 & ~w262 ) | ( \pi104 & ~w262 ) ;
  assign w264 = ( \pi128 & ~\pi129 ) | ( \pi128 & w263 ) | ( ~\pi129 & w263 ) ;
  assign w265 = \pi102 | w264 ;
  assign w266 = \pi103 & w264 ;
  assign w267 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w263 ) | ( \pi129 & w263 ) ;
  assign w268 = ( w265 & w266 ) | ( w265 & w267 ) | ( w266 & w267 ) ;
  assign w269 = \pi130 ^ w247 ;
  assign w270 = ( w247 & w261 ) | ( w247 & w269 ) | ( w261 & w269 ) ;
  assign w271 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w270 ) | ( \pi131 & w270 ) ;
  assign w272 = w254 | w271 ;
  assign w273 = w268 & w271 ;
  assign w274 = ( \pi130 & ~\pi131 ) | ( \pi130 & w270 ) | ( ~\pi131 & w270 ) ;
  assign w275 = ( w272 & w273 ) | ( w272 & w274 ) | ( w273 & w274 ) ;
  assign w276 = \pi132 ^ w170 ;
  assign w277 = ( w170 & w240 ) | ( w170 & ~w276 ) | ( w240 & ~w276 ) ;
  assign w278 = ( \pi132 & ~\pi133 ) | ( \pi132 & w277 ) | ( ~\pi133 & w277 ) ;
  assign w279 = w205 | w278 ;
  assign w280 = w275 & w278 ;
  assign w281 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w277 ) | ( \pi133 & w277 ) ;
  assign w282 = ( w279 & w280 ) | ( w279 & w281 ) | ( w280 & w281 ) ;
  assign w283 = \pi013 ^ \pi128 ;
  assign w284 = ( \pi013 & \pi016 ) | ( \pi013 & ~w283 ) | ( \pi016 & ~w283 ) ;
  assign w285 = ( \pi128 & ~\pi129 ) | ( \pi128 & w284 ) | ( ~\pi129 & w284 ) ;
  assign w286 = \pi014 | w285 ;
  assign w287 = \pi015 & w285 ;
  assign w288 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w284 ) | ( \pi129 & w284 ) ;
  assign w289 = ( w286 & w287 ) | ( w286 & w288 ) | ( w287 & w288 ) ;
  assign w290 = \pi009 ^ \pi128 ;
  assign w291 = ( \pi009 & \pi012 ) | ( \pi009 & ~w290 ) | ( \pi012 & ~w290 ) ;
  assign w292 = ( \pi128 & ~\pi129 ) | ( \pi128 & w291 ) | ( ~\pi129 & w291 ) ;
  assign w293 = \pi010 | w292 ;
  assign w294 = \pi011 & w292 ;
  assign w295 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w291 ) | ( \pi129 & w291 ) ;
  assign w296 = ( w293 & w294 ) | ( w293 & w295 ) | ( w294 & w295 ) ;
  assign w297 = \pi001 ^ \pi128 ;
  assign w298 = ( \pi001 & \pi004 ) | ( \pi001 & ~w297 ) | ( \pi004 & ~w297 ) ;
  assign w299 = ( \pi128 & ~\pi129 ) | ( \pi128 & w298 ) | ( ~\pi129 & w298 ) ;
  assign w300 = \pi002 | w299 ;
  assign w301 = \pi003 & w299 ;
  assign w302 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w298 ) | ( \pi129 & w298 ) ;
  assign w303 = ( w300 & w301 ) | ( w300 & w302 ) | ( w301 & w302 ) ;
  assign w304 = \pi005 ^ \pi128 ;
  assign w305 = ( \pi005 & \pi008 ) | ( \pi005 & ~w304 ) | ( \pi008 & ~w304 ) ;
  assign w306 = ( \pi128 & ~\pi129 ) | ( \pi128 & w305 ) | ( ~\pi129 & w305 ) ;
  assign w307 = \pi006 | w306 ;
  assign w308 = \pi007 & w306 ;
  assign w309 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w305 ) | ( \pi129 & w305 ) ;
  assign w310 = ( w307 & w308 ) | ( w307 & w309 ) | ( w308 & w309 ) ;
  assign w311 = \pi130 ^ w289 ;
  assign w312 = ( w289 & w303 ) | ( w289 & w311 ) | ( w303 & w311 ) ;
  assign w313 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w312 ) | ( \pi131 & w312 ) ;
  assign w314 = w296 | w313 ;
  assign w315 = w310 & w313 ;
  assign w316 = ( \pi130 & ~\pi131 ) | ( \pi130 & w312 ) | ( ~\pi131 & w312 ) ;
  assign w317 = ( w314 & w315 ) | ( w314 & w316 ) | ( w315 & w316 ) ;
  assign w318 = \pi029 ^ \pi128 ;
  assign w319 = ( \pi029 & \pi032 ) | ( \pi029 & ~w318 ) | ( \pi032 & ~w318 ) ;
  assign w320 = ( \pi128 & ~\pi129 ) | ( \pi128 & w319 ) | ( ~\pi129 & w319 ) ;
  assign w321 = \pi030 | w320 ;
  assign w322 = \pi031 & w320 ;
  assign w323 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w319 ) | ( \pi129 & w319 ) ;
  assign w324 = ( w321 & w322 ) | ( w321 & w323 ) | ( w322 & w323 ) ;
  assign w325 = \pi025 ^ \pi128 ;
  assign w326 = ( \pi025 & \pi028 ) | ( \pi025 & ~w325 ) | ( \pi028 & ~w325 ) ;
  assign w327 = ( \pi128 & ~\pi129 ) | ( \pi128 & w326 ) | ( ~\pi129 & w326 ) ;
  assign w328 = \pi026 | w327 ;
  assign w329 = \pi027 & w327 ;
  assign w330 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w326 ) | ( \pi129 & w326 ) ;
  assign w331 = ( w328 & w329 ) | ( w328 & w330 ) | ( w329 & w330 ) ;
  assign w332 = \pi017 ^ \pi128 ;
  assign w333 = ( \pi017 & \pi020 ) | ( \pi017 & ~w332 ) | ( \pi020 & ~w332 ) ;
  assign w334 = ( \pi128 & ~\pi129 ) | ( \pi128 & w333 ) | ( ~\pi129 & w333 ) ;
  assign w335 = \pi018 | w334 ;
  assign w336 = \pi019 & w334 ;
  assign w337 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w333 ) | ( \pi129 & w333 ) ;
  assign w338 = ( w335 & w336 ) | ( w335 & w337 ) | ( w336 & w337 ) ;
  assign w339 = \pi021 ^ \pi128 ;
  assign w340 = ( \pi021 & \pi024 ) | ( \pi021 & ~w339 ) | ( \pi024 & ~w339 ) ;
  assign w341 = ( \pi128 & ~\pi129 ) | ( \pi128 & w340 ) | ( ~\pi129 & w340 ) ;
  assign w342 = \pi022 | w341 ;
  assign w343 = \pi023 & w341 ;
  assign w344 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w340 ) | ( \pi129 & w340 ) ;
  assign w345 = ( w342 & w343 ) | ( w342 & w344 ) | ( w343 & w344 ) ;
  assign w346 = \pi130 ^ w324 ;
  assign w347 = ( w324 & w338 ) | ( w324 & w346 ) | ( w338 & w346 ) ;
  assign w348 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w347 ) | ( \pi131 & w347 ) ;
  assign w349 = w331 | w348 ;
  assign w350 = w345 & w348 ;
  assign w351 = ( \pi130 & ~\pi131 ) | ( \pi130 & w347 ) | ( ~\pi131 & w347 ) ;
  assign w352 = ( w349 & w350 ) | ( w349 & w351 ) | ( w350 & w351 ) ;
  assign w353 = \pi061 ^ \pi128 ;
  assign w354 = ( \pi061 & \pi064 ) | ( \pi061 & ~w353 ) | ( \pi064 & ~w353 ) ;
  assign w355 = ( \pi128 & ~\pi129 ) | ( \pi128 & w354 ) | ( ~\pi129 & w354 ) ;
  assign w356 = \pi062 | w355 ;
  assign w357 = \pi063 & w355 ;
  assign w358 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w354 ) | ( \pi129 & w354 ) ;
  assign w359 = ( w356 & w357 ) | ( w356 & w358 ) | ( w357 & w358 ) ;
  assign w360 = \pi057 ^ \pi128 ;
  assign w361 = ( \pi057 & \pi060 ) | ( \pi057 & ~w360 ) | ( \pi060 & ~w360 ) ;
  assign w362 = ( \pi128 & ~\pi129 ) | ( \pi128 & w361 ) | ( ~\pi129 & w361 ) ;
  assign w363 = \pi058 | w362 ;
  assign w364 = \pi059 & w362 ;
  assign w365 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w361 ) | ( \pi129 & w361 ) ;
  assign w366 = ( w363 & w364 ) | ( w363 & w365 ) | ( w364 & w365 ) ;
  assign w367 = \pi049 ^ \pi128 ;
  assign w368 = ( \pi049 & \pi052 ) | ( \pi049 & ~w367 ) | ( \pi052 & ~w367 ) ;
  assign w369 = ( \pi128 & ~\pi129 ) | ( \pi128 & w368 ) | ( ~\pi129 & w368 ) ;
  assign w370 = \pi050 | w369 ;
  assign w371 = \pi051 & w369 ;
  assign w372 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w368 ) | ( \pi129 & w368 ) ;
  assign w373 = ( w370 & w371 ) | ( w370 & w372 ) | ( w371 & w372 ) ;
  assign w374 = \pi053 ^ \pi128 ;
  assign w375 = ( \pi053 & \pi056 ) | ( \pi053 & ~w374 ) | ( \pi056 & ~w374 ) ;
  assign w376 = ( \pi128 & ~\pi129 ) | ( \pi128 & w375 ) | ( ~\pi129 & w375 ) ;
  assign w377 = \pi054 | w376 ;
  assign w378 = \pi055 & w376 ;
  assign w379 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w375 ) | ( \pi129 & w375 ) ;
  assign w380 = ( w377 & w378 ) | ( w377 & w379 ) | ( w378 & w379 ) ;
  assign w381 = \pi130 ^ w359 ;
  assign w382 = ( w359 & w373 ) | ( w359 & w381 ) | ( w373 & w381 ) ;
  assign w383 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w382 ) | ( \pi131 & w382 ) ;
  assign w384 = w366 | w383 ;
  assign w385 = w380 & w383 ;
  assign w386 = ( \pi130 & ~\pi131 ) | ( \pi130 & w382 ) | ( ~\pi131 & w382 ) ;
  assign w387 = ( w384 & w385 ) | ( w384 & w386 ) | ( w385 & w386 ) ;
  assign w388 = \pi045 ^ \pi128 ;
  assign w389 = ( \pi045 & \pi048 ) | ( \pi045 & ~w388 ) | ( \pi048 & ~w388 ) ;
  assign w390 = ( \pi128 & ~\pi129 ) | ( \pi128 & w389 ) | ( ~\pi129 & w389 ) ;
  assign w391 = \pi046 | w390 ;
  assign w392 = \pi047 & w390 ;
  assign w393 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w389 ) | ( \pi129 & w389 ) ;
  assign w394 = ( w391 & w392 ) | ( w391 & w393 ) | ( w392 & w393 ) ;
  assign w395 = \pi041 ^ \pi128 ;
  assign w396 = ( \pi041 & \pi044 ) | ( \pi041 & ~w395 ) | ( \pi044 & ~w395 ) ;
  assign w397 = ( \pi128 & ~\pi129 ) | ( \pi128 & w396 ) | ( ~\pi129 & w396 ) ;
  assign w398 = \pi042 | w397 ;
  assign w399 = \pi043 & w397 ;
  assign w400 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w396 ) | ( \pi129 & w396 ) ;
  assign w401 = ( w398 & w399 ) | ( w398 & w400 ) | ( w399 & w400 ) ;
  assign w402 = \pi033 ^ \pi128 ;
  assign w403 = ( \pi033 & \pi036 ) | ( \pi033 & ~w402 ) | ( \pi036 & ~w402 ) ;
  assign w404 = ( \pi128 & ~\pi129 ) | ( \pi128 & w403 ) | ( ~\pi129 & w403 ) ;
  assign w405 = \pi034 | w404 ;
  assign w406 = \pi035 & w404 ;
  assign w407 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w403 ) | ( \pi129 & w403 ) ;
  assign w408 = ( w405 & w406 ) | ( w405 & w407 ) | ( w406 & w407 ) ;
  assign w409 = \pi037 ^ \pi128 ;
  assign w410 = ( \pi037 & \pi040 ) | ( \pi037 & ~w409 ) | ( \pi040 & ~w409 ) ;
  assign w411 = ( \pi128 & ~\pi129 ) | ( \pi128 & w410 ) | ( ~\pi129 & w410 ) ;
  assign w412 = \pi038 | w411 ;
  assign w413 = \pi039 & w411 ;
  assign w414 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w410 ) | ( \pi129 & w410 ) ;
  assign w415 = ( w412 & w413 ) | ( w412 & w414 ) | ( w413 & w414 ) ;
  assign w416 = \pi130 ^ w394 ;
  assign w417 = ( w394 & w408 ) | ( w394 & w416 ) | ( w408 & w416 ) ;
  assign w418 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w417 ) | ( \pi131 & w417 ) ;
  assign w419 = w401 | w418 ;
  assign w420 = w415 & w418 ;
  assign w421 = ( \pi130 & ~\pi131 ) | ( \pi130 & w417 ) | ( ~\pi131 & w417 ) ;
  assign w422 = ( w419 & w420 ) | ( w419 & w421 ) | ( w420 & w421 ) ;
  assign w423 = \pi132 ^ w317 ;
  assign w424 = ( w317 & w387 ) | ( w317 & ~w423 ) | ( w387 & ~w423 ) ;
  assign w425 = ( \pi132 & ~\pi133 ) | ( \pi132 & w424 ) | ( ~\pi133 & w424 ) ;
  assign w426 = w352 | w425 ;
  assign w427 = w422 & w425 ;
  assign w428 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w424 ) | ( \pi133 & w424 ) ;
  assign w429 = ( w426 & w427 ) | ( w426 & w428 ) | ( w427 & w428 ) ;
  assign w430 = \pi134 ^ w429 ;
  assign w431 = ( w282 & w429 ) | ( w282 & ~w430 ) | ( w429 & ~w430 ) ;
  assign w432 = \pi078 ^ \pi128 ;
  assign w433 = ( \pi078 & \pi081 ) | ( \pi078 & ~w432 ) | ( \pi081 & ~w432 ) ;
  assign w434 = ( \pi128 & ~\pi129 ) | ( \pi128 & w433 ) | ( ~\pi129 & w433 ) ;
  assign w435 = \pi079 | w434 ;
  assign w436 = \pi080 & w434 ;
  assign w437 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w433 ) | ( \pi129 & w433 ) ;
  assign w438 = ( w435 & w436 ) | ( w435 & w437 ) | ( w436 & w437 ) ;
  assign w439 = \pi074 ^ \pi128 ;
  assign w440 = ( \pi074 & \pi077 ) | ( \pi074 & ~w439 ) | ( \pi077 & ~w439 ) ;
  assign w441 = ( \pi128 & ~\pi129 ) | ( \pi128 & w440 ) | ( ~\pi129 & w440 ) ;
  assign w442 = \pi075 | w441 ;
  assign w443 = \pi076 & w441 ;
  assign w444 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w440 ) | ( \pi129 & w440 ) ;
  assign w445 = ( w442 & w443 ) | ( w442 & w444 ) | ( w443 & w444 ) ;
  assign w446 = \pi066 ^ \pi128 ;
  assign w447 = ( \pi066 & \pi069 ) | ( \pi066 & ~w446 ) | ( \pi069 & ~w446 ) ;
  assign w448 = ( \pi128 & ~\pi129 ) | ( \pi128 & w447 ) | ( ~\pi129 & w447 ) ;
  assign w449 = \pi067 | w448 ;
  assign w450 = \pi068 & w448 ;
  assign w451 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w447 ) | ( \pi129 & w447 ) ;
  assign w452 = ( w449 & w450 ) | ( w449 & w451 ) | ( w450 & w451 ) ;
  assign w453 = \pi070 ^ \pi128 ;
  assign w454 = ( \pi070 & \pi073 ) | ( \pi070 & ~w453 ) | ( \pi073 & ~w453 ) ;
  assign w455 = ( \pi128 & ~\pi129 ) | ( \pi128 & w454 ) | ( ~\pi129 & w454 ) ;
  assign w456 = \pi071 | w455 ;
  assign w457 = \pi072 & w455 ;
  assign w458 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w454 ) | ( \pi129 & w454 ) ;
  assign w459 = ( w456 & w457 ) | ( w456 & w458 ) | ( w457 & w458 ) ;
  assign w460 = \pi130 ^ w438 ;
  assign w461 = ( w438 & w452 ) | ( w438 & w460 ) | ( w452 & w460 ) ;
  assign w462 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w461 ) | ( \pi131 & w461 ) ;
  assign w463 = w445 | w462 ;
  assign w464 = w459 & w462 ;
  assign w465 = ( \pi130 & ~\pi131 ) | ( \pi130 & w461 ) | ( ~\pi131 & w461 ) ;
  assign w466 = ( w463 & w464 ) | ( w463 & w465 ) | ( w464 & w465 ) ;
  assign w467 = \pi094 ^ \pi128 ;
  assign w468 = ( \pi094 & \pi097 ) | ( \pi094 & ~w467 ) | ( \pi097 & ~w467 ) ;
  assign w469 = ( \pi128 & ~\pi129 ) | ( \pi128 & w468 ) | ( ~\pi129 & w468 ) ;
  assign w470 = \pi095 | w469 ;
  assign w471 = \pi096 & w469 ;
  assign w472 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w468 ) | ( \pi129 & w468 ) ;
  assign w473 = ( w470 & w471 ) | ( w470 & w472 ) | ( w471 & w472 ) ;
  assign w474 = \pi090 ^ \pi128 ;
  assign w475 = ( \pi090 & \pi093 ) | ( \pi090 & ~w474 ) | ( \pi093 & ~w474 ) ;
  assign w476 = ( \pi128 & ~\pi129 ) | ( \pi128 & w475 ) | ( ~\pi129 & w475 ) ;
  assign w477 = \pi091 | w476 ;
  assign w478 = \pi092 & w476 ;
  assign w479 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w475 ) | ( \pi129 & w475 ) ;
  assign w480 = ( w477 & w478 ) | ( w477 & w479 ) | ( w478 & w479 ) ;
  assign w481 = \pi082 ^ \pi128 ;
  assign w482 = ( \pi082 & \pi085 ) | ( \pi082 & ~w481 ) | ( \pi085 & ~w481 ) ;
  assign w483 = ( \pi128 & ~\pi129 ) | ( \pi128 & w482 ) | ( ~\pi129 & w482 ) ;
  assign w484 = \pi083 | w483 ;
  assign w485 = \pi084 & w483 ;
  assign w486 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w482 ) | ( \pi129 & w482 ) ;
  assign w487 = ( w484 & w485 ) | ( w484 & w486 ) | ( w485 & w486 ) ;
  assign w488 = \pi086 ^ \pi128 ;
  assign w489 = ( \pi086 & \pi089 ) | ( \pi086 & ~w488 ) | ( \pi089 & ~w488 ) ;
  assign w490 = ( \pi128 & ~\pi129 ) | ( \pi128 & w489 ) | ( ~\pi129 & w489 ) ;
  assign w491 = \pi087 | w490 ;
  assign w492 = \pi088 & w490 ;
  assign w493 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w489 ) | ( \pi129 & w489 ) ;
  assign w494 = ( w491 & w492 ) | ( w491 & w493 ) | ( w492 & w493 ) ;
  assign w495 = \pi130 ^ w473 ;
  assign w496 = ( w473 & w487 ) | ( w473 & w495 ) | ( w487 & w495 ) ;
  assign w497 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w496 ) | ( \pi131 & w496 ) ;
  assign w498 = w480 | w497 ;
  assign w499 = w494 & w497 ;
  assign w500 = ( \pi130 & ~\pi131 ) | ( \pi130 & w496 ) | ( ~\pi131 & w496 ) ;
  assign w501 = ( w498 & w499 ) | ( w498 & w500 ) | ( w499 & w500 ) ;
  assign w502 = \pi000 ^ \pi128 ;
  assign w503 = ( \pi000 & \pi127 ) | ( \pi000 & ~w502 ) | ( \pi127 & ~w502 ) ;
  assign w504 = ( \pi128 & \pi129 ) | ( \pi128 & w503 ) | ( \pi129 & w503 ) ;
  assign w505 = \pi001 | w504 ;
  assign w506 = \pi126 & w504 ;
  assign w507 = ( \pi128 & \pi129 ) | ( \pi128 & ~w503 ) | ( \pi129 & ~w503 ) ;
  assign w508 = ( w505 & w506 ) | ( w505 & ~w507 ) | ( w506 & ~w507 ) ;
  assign w509 = \pi122 ^ \pi128 ;
  assign w510 = ( \pi122 & \pi125 ) | ( \pi122 & ~w509 ) | ( \pi125 & ~w509 ) ;
  assign w511 = ( \pi128 & ~\pi129 ) | ( \pi128 & w510 ) | ( ~\pi129 & w510 ) ;
  assign w512 = \pi123 | w511 ;
  assign w513 = \pi124 & w511 ;
  assign w514 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w510 ) | ( \pi129 & w510 ) ;
  assign w515 = ( w512 & w513 ) | ( w512 & w514 ) | ( w513 & w514 ) ;
  assign w516 = \pi114 ^ \pi128 ;
  assign w517 = ( \pi114 & \pi117 ) | ( \pi114 & ~w516 ) | ( \pi117 & ~w516 ) ;
  assign w518 = ( \pi128 & ~\pi129 ) | ( \pi128 & w517 ) | ( ~\pi129 & w517 ) ;
  assign w519 = \pi115 | w518 ;
  assign w520 = \pi116 & w518 ;
  assign w521 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w517 ) | ( \pi129 & w517 ) ;
  assign w522 = ( w519 & w520 ) | ( w519 & w521 ) | ( w520 & w521 ) ;
  assign w523 = \pi118 ^ \pi128 ;
  assign w524 = ( \pi118 & \pi121 ) | ( \pi118 & ~w523 ) | ( \pi121 & ~w523 ) ;
  assign w525 = ( \pi128 & ~\pi129 ) | ( \pi128 & w524 ) | ( ~\pi129 & w524 ) ;
  assign w526 = \pi119 | w525 ;
  assign w527 = \pi120 & w525 ;
  assign w528 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w524 ) | ( \pi129 & w524 ) ;
  assign w529 = ( w526 & w527 ) | ( w526 & w528 ) | ( w527 & w528 ) ;
  assign w530 = \pi130 ^ w508 ;
  assign w531 = ( w508 & w522 ) | ( w508 & w530 ) | ( w522 & w530 ) ;
  assign w532 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w531 ) | ( \pi131 & w531 ) ;
  assign w533 = w515 | w532 ;
  assign w534 = w529 & w532 ;
  assign w535 = ( \pi130 & ~\pi131 ) | ( \pi130 & w531 ) | ( ~\pi131 & w531 ) ;
  assign w536 = ( w533 & w534 ) | ( w533 & w535 ) | ( w534 & w535 ) ;
  assign w537 = \pi110 ^ \pi128 ;
  assign w538 = ( \pi110 & \pi113 ) | ( \pi110 & ~w537 ) | ( \pi113 & ~w537 ) ;
  assign w539 = ( \pi128 & ~\pi129 ) | ( \pi128 & w538 ) | ( ~\pi129 & w538 ) ;
  assign w540 = \pi111 | w539 ;
  assign w541 = \pi112 & w539 ;
  assign w542 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w538 ) | ( \pi129 & w538 ) ;
  assign w543 = ( w540 & w541 ) | ( w540 & w542 ) | ( w541 & w542 ) ;
  assign w544 = \pi106 ^ \pi128 ;
  assign w545 = ( \pi106 & \pi109 ) | ( \pi106 & ~w544 ) | ( \pi109 & ~w544 ) ;
  assign w546 = ( \pi128 & ~\pi129 ) | ( \pi128 & w545 ) | ( ~\pi129 & w545 ) ;
  assign w547 = \pi107 | w546 ;
  assign w548 = \pi108 & w546 ;
  assign w549 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w545 ) | ( \pi129 & w545 ) ;
  assign w550 = ( w547 & w548 ) | ( w547 & w549 ) | ( w548 & w549 ) ;
  assign w551 = \pi098 ^ \pi128 ;
  assign w552 = ( \pi098 & \pi101 ) | ( \pi098 & ~w551 ) | ( \pi101 & ~w551 ) ;
  assign w553 = ( \pi128 & ~\pi129 ) | ( \pi128 & w552 ) | ( ~\pi129 & w552 ) ;
  assign w554 = \pi099 | w553 ;
  assign w555 = \pi100 & w553 ;
  assign w556 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w552 ) | ( \pi129 & w552 ) ;
  assign w557 = ( w554 & w555 ) | ( w554 & w556 ) | ( w555 & w556 ) ;
  assign w558 = \pi102 ^ \pi128 ;
  assign w559 = ( \pi102 & \pi105 ) | ( \pi102 & ~w558 ) | ( \pi105 & ~w558 ) ;
  assign w560 = ( \pi128 & ~\pi129 ) | ( \pi128 & w559 ) | ( ~\pi129 & w559 ) ;
  assign w561 = \pi103 | w560 ;
  assign w562 = \pi104 & w560 ;
  assign w563 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w559 ) | ( \pi129 & w559 ) ;
  assign w564 = ( w561 & w562 ) | ( w561 & w563 ) | ( w562 & w563 ) ;
  assign w565 = \pi130 ^ w543 ;
  assign w566 = ( w543 & w557 ) | ( w543 & w565 ) | ( w557 & w565 ) ;
  assign w567 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w566 ) | ( \pi131 & w566 ) ;
  assign w568 = w550 | w567 ;
  assign w569 = w564 & w567 ;
  assign w570 = ( \pi130 & ~\pi131 ) | ( \pi130 & w566 ) | ( ~\pi131 & w566 ) ;
  assign w571 = ( w568 & w569 ) | ( w568 & w570 ) | ( w569 & w570 ) ;
  assign w572 = \pi132 ^ w466 ;
  assign w573 = ( w466 & w536 ) | ( w466 & ~w572 ) | ( w536 & ~w572 ) ;
  assign w574 = ( \pi132 & ~\pi133 ) | ( \pi132 & w573 ) | ( ~\pi133 & w573 ) ;
  assign w575 = w501 | w574 ;
  assign w576 = w571 & w574 ;
  assign w577 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w573 ) | ( \pi133 & w573 ) ;
  assign w578 = ( w575 & w576 ) | ( w575 & w577 ) | ( w576 & w577 ) ;
  assign w579 = \pi062 ^ \pi128 ;
  assign w580 = ( \pi062 & \pi065 ) | ( \pi062 & ~w579 ) | ( \pi065 & ~w579 ) ;
  assign w581 = ( \pi128 & ~\pi129 ) | ( \pi128 & w580 ) | ( ~\pi129 & w580 ) ;
  assign w582 = \pi063 | w581 ;
  assign w583 = \pi064 & w581 ;
  assign w584 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w580 ) | ( \pi129 & w580 ) ;
  assign w585 = ( w582 & w583 ) | ( w582 & w584 ) | ( w583 & w584 ) ;
  assign w586 = \pi058 ^ \pi128 ;
  assign w587 = ( \pi058 & \pi061 ) | ( \pi058 & ~w586 ) | ( \pi061 & ~w586 ) ;
  assign w588 = ( \pi128 & ~\pi129 ) | ( \pi128 & w587 ) | ( ~\pi129 & w587 ) ;
  assign w589 = \pi059 | w588 ;
  assign w590 = \pi060 & w588 ;
  assign w591 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w587 ) | ( \pi129 & w587 ) ;
  assign w592 = ( w589 & w590 ) | ( w589 & w591 ) | ( w590 & w591 ) ;
  assign w593 = \pi050 ^ \pi128 ;
  assign w594 = ( \pi050 & \pi053 ) | ( \pi050 & ~w593 ) | ( \pi053 & ~w593 ) ;
  assign w595 = ( \pi128 & ~\pi129 ) | ( \pi128 & w594 ) | ( ~\pi129 & w594 ) ;
  assign w596 = \pi051 | w595 ;
  assign w597 = \pi052 & w595 ;
  assign w598 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w594 ) | ( \pi129 & w594 ) ;
  assign w599 = ( w596 & w597 ) | ( w596 & w598 ) | ( w597 & w598 ) ;
  assign w600 = \pi054 ^ \pi128 ;
  assign w601 = ( \pi054 & \pi057 ) | ( \pi054 & ~w600 ) | ( \pi057 & ~w600 ) ;
  assign w602 = ( \pi128 & ~\pi129 ) | ( \pi128 & w601 ) | ( ~\pi129 & w601 ) ;
  assign w603 = \pi055 | w602 ;
  assign w604 = \pi056 & w602 ;
  assign w605 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w601 ) | ( \pi129 & w601 ) ;
  assign w606 = ( w603 & w604 ) | ( w603 & w605 ) | ( w604 & w605 ) ;
  assign w607 = \pi130 ^ w585 ;
  assign w608 = ( w585 & w599 ) | ( w585 & w607 ) | ( w599 & w607 ) ;
  assign w609 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w608 ) | ( \pi131 & w608 ) ;
  assign w610 = w592 | w609 ;
  assign w611 = w606 & w609 ;
  assign w612 = ( \pi130 & ~\pi131 ) | ( \pi130 & w608 ) | ( ~\pi131 & w608 ) ;
  assign w613 = ( w610 & w611 ) | ( w610 & w612 ) | ( w611 & w612 ) ;
  assign w614 = \pi014 ^ \pi128 ;
  assign w615 = ( \pi014 & \pi017 ) | ( \pi014 & ~w614 ) | ( \pi017 & ~w614 ) ;
  assign w616 = ( \pi128 & ~\pi129 ) | ( \pi128 & w615 ) | ( ~\pi129 & w615 ) ;
  assign w617 = \pi015 | w616 ;
  assign w618 = \pi016 & w616 ;
  assign w619 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w615 ) | ( \pi129 & w615 ) ;
  assign w620 = ( w617 & w618 ) | ( w617 & w619 ) | ( w618 & w619 ) ;
  assign w621 = \pi010 ^ \pi128 ;
  assign w622 = ( \pi010 & \pi013 ) | ( \pi010 & ~w621 ) | ( \pi013 & ~w621 ) ;
  assign w623 = ( \pi128 & ~\pi129 ) | ( \pi128 & w622 ) | ( ~\pi129 & w622 ) ;
  assign w624 = \pi011 | w623 ;
  assign w625 = \pi012 & w623 ;
  assign w626 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w622 ) | ( \pi129 & w622 ) ;
  assign w627 = ( w624 & w625 ) | ( w624 & w626 ) | ( w625 & w626 ) ;
  assign w628 = \pi002 ^ \pi128 ;
  assign w629 = ( \pi002 & \pi005 ) | ( \pi002 & ~w628 ) | ( \pi005 & ~w628 ) ;
  assign w630 = ( \pi128 & ~\pi129 ) | ( \pi128 & w629 ) | ( ~\pi129 & w629 ) ;
  assign w631 = \pi003 | w630 ;
  assign w632 = \pi004 & w630 ;
  assign w633 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w629 ) | ( \pi129 & w629 ) ;
  assign w634 = ( w631 & w632 ) | ( w631 & w633 ) | ( w632 & w633 ) ;
  assign w635 = \pi006 ^ \pi128 ;
  assign w636 = ( \pi006 & \pi009 ) | ( \pi006 & ~w635 ) | ( \pi009 & ~w635 ) ;
  assign w637 = ( \pi128 & ~\pi129 ) | ( \pi128 & w636 ) | ( ~\pi129 & w636 ) ;
  assign w638 = \pi007 | w637 ;
  assign w639 = \pi008 & w637 ;
  assign w640 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w636 ) | ( \pi129 & w636 ) ;
  assign w641 = ( w638 & w639 ) | ( w638 & w640 ) | ( w639 & w640 ) ;
  assign w642 = \pi130 ^ w620 ;
  assign w643 = ( w620 & w634 ) | ( w620 & w642 ) | ( w634 & w642 ) ;
  assign w644 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w643 ) | ( \pi131 & w643 ) ;
  assign w645 = w627 | w644 ;
  assign w646 = w641 & w644 ;
  assign w647 = ( \pi130 & ~\pi131 ) | ( \pi130 & w643 ) | ( ~\pi131 & w643 ) ;
  assign w648 = ( w645 & w646 ) | ( w645 & w647 ) | ( w646 & w647 ) ;
  assign w649 = \pi046 ^ \pi128 ;
  assign w650 = ( \pi046 & \pi049 ) | ( \pi046 & ~w649 ) | ( \pi049 & ~w649 ) ;
  assign w651 = ( \pi128 & ~\pi129 ) | ( \pi128 & w650 ) | ( ~\pi129 & w650 ) ;
  assign w652 = \pi047 | w651 ;
  assign w653 = \pi048 & w651 ;
  assign w654 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w650 ) | ( \pi129 & w650 ) ;
  assign w655 = ( w652 & w653 ) | ( w652 & w654 ) | ( w653 & w654 ) ;
  assign w656 = \pi042 ^ \pi128 ;
  assign w657 = ( \pi042 & \pi045 ) | ( \pi042 & ~w656 ) | ( \pi045 & ~w656 ) ;
  assign w658 = ( \pi128 & ~\pi129 ) | ( \pi128 & w657 ) | ( ~\pi129 & w657 ) ;
  assign w659 = \pi043 | w658 ;
  assign w660 = \pi044 & w658 ;
  assign w661 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w657 ) | ( \pi129 & w657 ) ;
  assign w662 = ( w659 & w660 ) | ( w659 & w661 ) | ( w660 & w661 ) ;
  assign w663 = \pi034 ^ \pi128 ;
  assign w664 = ( \pi034 & \pi037 ) | ( \pi034 & ~w663 ) | ( \pi037 & ~w663 ) ;
  assign w665 = ( \pi128 & ~\pi129 ) | ( \pi128 & w664 ) | ( ~\pi129 & w664 ) ;
  assign w666 = \pi035 | w665 ;
  assign w667 = \pi036 & w665 ;
  assign w668 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w664 ) | ( \pi129 & w664 ) ;
  assign w669 = ( w666 & w667 ) | ( w666 & w668 ) | ( w667 & w668 ) ;
  assign w670 = \pi038 ^ \pi128 ;
  assign w671 = ( \pi038 & \pi041 ) | ( \pi038 & ~w670 ) | ( \pi041 & ~w670 ) ;
  assign w672 = ( \pi128 & ~\pi129 ) | ( \pi128 & w671 ) | ( ~\pi129 & w671 ) ;
  assign w673 = \pi039 | w672 ;
  assign w674 = \pi040 & w672 ;
  assign w675 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w671 ) | ( \pi129 & w671 ) ;
  assign w676 = ( w673 & w674 ) | ( w673 & w675 ) | ( w674 & w675 ) ;
  assign w677 = \pi130 ^ w655 ;
  assign w678 = ( w655 & w669 ) | ( w655 & w677 ) | ( w669 & w677 ) ;
  assign w679 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w678 ) | ( \pi131 & w678 ) ;
  assign w680 = w662 | w679 ;
  assign w681 = w676 & w679 ;
  assign w682 = ( \pi130 & ~\pi131 ) | ( \pi130 & w678 ) | ( ~\pi131 & w678 ) ;
  assign w683 = ( w680 & w681 ) | ( w680 & w682 ) | ( w681 & w682 ) ;
  assign w684 = \pi030 ^ \pi128 ;
  assign w685 = ( \pi030 & \pi033 ) | ( \pi030 & ~w684 ) | ( \pi033 & ~w684 ) ;
  assign w686 = ( \pi128 & ~\pi129 ) | ( \pi128 & w685 ) | ( ~\pi129 & w685 ) ;
  assign w687 = \pi031 | w686 ;
  assign w688 = \pi032 & w686 ;
  assign w689 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w685 ) | ( \pi129 & w685 ) ;
  assign w690 = ( w687 & w688 ) | ( w687 & w689 ) | ( w688 & w689 ) ;
  assign w691 = \pi026 ^ \pi128 ;
  assign w692 = ( \pi026 & \pi029 ) | ( \pi026 & ~w691 ) | ( \pi029 & ~w691 ) ;
  assign w693 = ( \pi128 & ~\pi129 ) | ( \pi128 & w692 ) | ( ~\pi129 & w692 ) ;
  assign w694 = \pi027 | w693 ;
  assign w695 = \pi028 & w693 ;
  assign w696 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w692 ) | ( \pi129 & w692 ) ;
  assign w697 = ( w694 & w695 ) | ( w694 & w696 ) | ( w695 & w696 ) ;
  assign w698 = \pi018 ^ \pi128 ;
  assign w699 = ( \pi018 & \pi021 ) | ( \pi018 & ~w698 ) | ( \pi021 & ~w698 ) ;
  assign w700 = ( \pi128 & ~\pi129 ) | ( \pi128 & w699 ) | ( ~\pi129 & w699 ) ;
  assign w701 = \pi019 | w700 ;
  assign w702 = \pi020 & w700 ;
  assign w703 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w699 ) | ( \pi129 & w699 ) ;
  assign w704 = ( w701 & w702 ) | ( w701 & w703 ) | ( w702 & w703 ) ;
  assign w705 = \pi022 ^ \pi128 ;
  assign w706 = ( \pi022 & \pi025 ) | ( \pi022 & ~w705 ) | ( \pi025 & ~w705 ) ;
  assign w707 = ( \pi128 & ~\pi129 ) | ( \pi128 & w706 ) | ( ~\pi129 & w706 ) ;
  assign w708 = \pi023 | w707 ;
  assign w709 = \pi024 & w707 ;
  assign w710 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w706 ) | ( \pi129 & w706 ) ;
  assign w711 = ( w708 & w709 ) | ( w708 & w710 ) | ( w709 & w710 ) ;
  assign w712 = \pi130 ^ w690 ;
  assign w713 = ( w690 & w704 ) | ( w690 & w712 ) | ( w704 & w712 ) ;
  assign w714 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w713 ) | ( \pi131 & w713 ) ;
  assign w715 = w697 | w714 ;
  assign w716 = w711 & w714 ;
  assign w717 = ( \pi130 & ~\pi131 ) | ( \pi130 & w713 ) | ( ~\pi131 & w713 ) ;
  assign w718 = ( w715 & w716 ) | ( w715 & w717 ) | ( w716 & w717 ) ;
  assign w719 = \pi132 ^ w613 ;
  assign w720 = ( w613 & w648 ) | ( w613 & w719 ) | ( w648 & w719 ) ;
  assign w721 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w720 ) | ( \pi133 & w720 ) ;
  assign w722 = w683 | w721 ;
  assign w723 = w718 & w721 ;
  assign w724 = ( \pi132 & ~\pi133 ) | ( \pi132 & w720 ) | ( ~\pi133 & w720 ) ;
  assign w725 = ( w722 & w723 ) | ( w722 & w724 ) | ( w723 & w724 ) ;
  assign w726 = \pi134 ^ w725 ;
  assign w727 = ( w578 & w725 ) | ( w578 & ~w726 ) | ( w725 & ~w726 ) ;
  assign w728 = \pi079 ^ \pi128 ;
  assign w729 = ( \pi079 & \pi082 ) | ( \pi079 & ~w728 ) | ( \pi082 & ~w728 ) ;
  assign w730 = ( \pi128 & ~\pi129 ) | ( \pi128 & w729 ) | ( ~\pi129 & w729 ) ;
  assign w731 = \pi080 | w730 ;
  assign w732 = \pi081 & w730 ;
  assign w733 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w729 ) | ( \pi129 & w729 ) ;
  assign w734 = ( w731 & w732 ) | ( w731 & w733 ) | ( w732 & w733 ) ;
  assign w735 = \pi075 ^ \pi128 ;
  assign w736 = ( \pi075 & \pi078 ) | ( \pi075 & ~w735 ) | ( \pi078 & ~w735 ) ;
  assign w737 = ( \pi128 & ~\pi129 ) | ( \pi128 & w736 ) | ( ~\pi129 & w736 ) ;
  assign w738 = \pi076 | w737 ;
  assign w739 = \pi077 & w737 ;
  assign w740 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w736 ) | ( \pi129 & w736 ) ;
  assign w741 = ( w738 & w739 ) | ( w738 & w740 ) | ( w739 & w740 ) ;
  assign w742 = \pi067 ^ \pi128 ;
  assign w743 = ( \pi067 & \pi070 ) | ( \pi067 & ~w742 ) | ( \pi070 & ~w742 ) ;
  assign w744 = ( \pi128 & ~\pi129 ) | ( \pi128 & w743 ) | ( ~\pi129 & w743 ) ;
  assign w745 = \pi068 | w744 ;
  assign w746 = \pi069 & w744 ;
  assign w747 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w743 ) | ( \pi129 & w743 ) ;
  assign w748 = ( w745 & w746 ) | ( w745 & w747 ) | ( w746 & w747 ) ;
  assign w749 = \pi071 ^ \pi128 ;
  assign w750 = ( \pi071 & \pi074 ) | ( \pi071 & ~w749 ) | ( \pi074 & ~w749 ) ;
  assign w751 = ( \pi128 & ~\pi129 ) | ( \pi128 & w750 ) | ( ~\pi129 & w750 ) ;
  assign w752 = \pi072 | w751 ;
  assign w753 = \pi073 & w751 ;
  assign w754 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w750 ) | ( \pi129 & w750 ) ;
  assign w755 = ( w752 & w753 ) | ( w752 & w754 ) | ( w753 & w754 ) ;
  assign w756 = \pi130 ^ w734 ;
  assign w757 = ( w734 & w748 ) | ( w734 & w756 ) | ( w748 & w756 ) ;
  assign w758 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w757 ) | ( \pi131 & w757 ) ;
  assign w759 = w741 | w758 ;
  assign w760 = w755 & w758 ;
  assign w761 = ( \pi130 & ~\pi131 ) | ( \pi130 & w757 ) | ( ~\pi131 & w757 ) ;
  assign w762 = ( w759 & w760 ) | ( w759 & w761 ) | ( w760 & w761 ) ;
  assign w763 = \pi095 ^ \pi128 ;
  assign w764 = ( \pi095 & \pi098 ) | ( \pi095 & ~w763 ) | ( \pi098 & ~w763 ) ;
  assign w765 = ( \pi128 & ~\pi129 ) | ( \pi128 & w764 ) | ( ~\pi129 & w764 ) ;
  assign w766 = \pi096 | w765 ;
  assign w767 = \pi097 & w765 ;
  assign w768 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w764 ) | ( \pi129 & w764 ) ;
  assign w769 = ( w766 & w767 ) | ( w766 & w768 ) | ( w767 & w768 ) ;
  assign w770 = \pi091 ^ \pi128 ;
  assign w771 = ( \pi091 & \pi094 ) | ( \pi091 & ~w770 ) | ( \pi094 & ~w770 ) ;
  assign w772 = ( \pi128 & ~\pi129 ) | ( \pi128 & w771 ) | ( ~\pi129 & w771 ) ;
  assign w773 = \pi092 | w772 ;
  assign w774 = \pi093 & w772 ;
  assign w775 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w771 ) | ( \pi129 & w771 ) ;
  assign w776 = ( w773 & w774 ) | ( w773 & w775 ) | ( w774 & w775 ) ;
  assign w777 = \pi083 ^ \pi128 ;
  assign w778 = ( \pi083 & \pi086 ) | ( \pi083 & ~w777 ) | ( \pi086 & ~w777 ) ;
  assign w779 = ( \pi128 & ~\pi129 ) | ( \pi128 & w778 ) | ( ~\pi129 & w778 ) ;
  assign w780 = \pi084 | w779 ;
  assign w781 = \pi085 & w779 ;
  assign w782 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w778 ) | ( \pi129 & w778 ) ;
  assign w783 = ( w780 & w781 ) | ( w780 & w782 ) | ( w781 & w782 ) ;
  assign w784 = \pi087 ^ \pi128 ;
  assign w785 = ( \pi087 & \pi090 ) | ( \pi087 & ~w784 ) | ( \pi090 & ~w784 ) ;
  assign w786 = ( \pi128 & ~\pi129 ) | ( \pi128 & w785 ) | ( ~\pi129 & w785 ) ;
  assign w787 = \pi088 | w786 ;
  assign w788 = \pi089 & w786 ;
  assign w789 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w785 ) | ( \pi129 & w785 ) ;
  assign w790 = ( w787 & w788 ) | ( w787 & w789 ) | ( w788 & w789 ) ;
  assign w791 = \pi130 ^ w769 ;
  assign w792 = ( w769 & w783 ) | ( w769 & w791 ) | ( w783 & w791 ) ;
  assign w793 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w792 ) | ( \pi131 & w792 ) ;
  assign w794 = w776 | w793 ;
  assign w795 = w790 & w793 ;
  assign w796 = ( \pi130 & ~\pi131 ) | ( \pi130 & w792 ) | ( ~\pi131 & w792 ) ;
  assign w797 = ( w794 & w795 ) | ( w794 & w796 ) | ( w795 & w796 ) ;
  assign w798 = ( \pi000 & \pi001 ) | ( \pi000 & ~w206 ) | ( \pi001 & ~w206 ) ;
  assign w799 = ( \pi128 & \pi129 ) | ( \pi128 & w798 ) | ( \pi129 & w798 ) ;
  assign w800 = \pi002 | w799 ;
  assign w801 = \pi127 & w799 ;
  assign w802 = ( \pi128 & \pi129 ) | ( \pi128 & ~w798 ) | ( \pi129 & ~w798 ) ;
  assign w803 = ( w800 & w801 ) | ( w800 & ~w802 ) | ( w801 & ~w802 ) ;
  assign w804 = \pi123 ^ \pi128 ;
  assign w805 = ( \pi123 & \pi126 ) | ( \pi123 & ~w804 ) | ( \pi126 & ~w804 ) ;
  assign w806 = ( \pi128 & ~\pi129 ) | ( \pi128 & w805 ) | ( ~\pi129 & w805 ) ;
  assign w807 = \pi124 | w806 ;
  assign w808 = \pi125 & w806 ;
  assign w809 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w805 ) | ( \pi129 & w805 ) ;
  assign w810 = ( w807 & w808 ) | ( w807 & w809 ) | ( w808 & w809 ) ;
  assign w811 = \pi115 ^ \pi128 ;
  assign w812 = ( \pi115 & \pi118 ) | ( \pi115 & ~w811 ) | ( \pi118 & ~w811 ) ;
  assign w813 = ( \pi128 & ~\pi129 ) | ( \pi128 & w812 ) | ( ~\pi129 & w812 ) ;
  assign w814 = \pi116 | w813 ;
  assign w815 = \pi117 & w813 ;
  assign w816 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w812 ) | ( \pi129 & w812 ) ;
  assign w817 = ( w814 & w815 ) | ( w814 & w816 ) | ( w815 & w816 ) ;
  assign w818 = \pi119 ^ \pi128 ;
  assign w819 = ( \pi119 & \pi122 ) | ( \pi119 & ~w818 ) | ( \pi122 & ~w818 ) ;
  assign w820 = ( \pi128 & ~\pi129 ) | ( \pi128 & w819 ) | ( ~\pi129 & w819 ) ;
  assign w821 = \pi120 | w820 ;
  assign w822 = \pi121 & w820 ;
  assign w823 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w819 ) | ( \pi129 & w819 ) ;
  assign w824 = ( w821 & w822 ) | ( w821 & w823 ) | ( w822 & w823 ) ;
  assign w825 = \pi130 ^ w803 ;
  assign w826 = ( w803 & w817 ) | ( w803 & w825 ) | ( w817 & w825 ) ;
  assign w827 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w826 ) | ( \pi131 & w826 ) ;
  assign w828 = w810 | w827 ;
  assign w829 = w824 & w827 ;
  assign w830 = ( \pi130 & ~\pi131 ) | ( \pi130 & w826 ) | ( ~\pi131 & w826 ) ;
  assign w831 = ( w828 & w829 ) | ( w828 & w830 ) | ( w829 & w830 ) ;
  assign w832 = \pi111 ^ \pi128 ;
  assign w833 = ( \pi111 & \pi114 ) | ( \pi111 & ~w832 ) | ( \pi114 & ~w832 ) ;
  assign w834 = ( \pi128 & ~\pi129 ) | ( \pi128 & w833 ) | ( ~\pi129 & w833 ) ;
  assign w835 = \pi112 | w834 ;
  assign w836 = \pi113 & w834 ;
  assign w837 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w833 ) | ( \pi129 & w833 ) ;
  assign w838 = ( w835 & w836 ) | ( w835 & w837 ) | ( w836 & w837 ) ;
  assign w839 = \pi107 ^ \pi128 ;
  assign w840 = ( \pi107 & \pi110 ) | ( \pi107 & ~w839 ) | ( \pi110 & ~w839 ) ;
  assign w841 = ( \pi128 & ~\pi129 ) | ( \pi128 & w840 ) | ( ~\pi129 & w840 ) ;
  assign w842 = \pi108 | w841 ;
  assign w843 = \pi109 & w841 ;
  assign w844 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w840 ) | ( \pi129 & w840 ) ;
  assign w845 = ( w842 & w843 ) | ( w842 & w844 ) | ( w843 & w844 ) ;
  assign w846 = \pi099 ^ \pi128 ;
  assign w847 = ( \pi099 & \pi102 ) | ( \pi099 & ~w846 ) | ( \pi102 & ~w846 ) ;
  assign w848 = ( \pi128 & ~\pi129 ) | ( \pi128 & w847 ) | ( ~\pi129 & w847 ) ;
  assign w849 = \pi100 | w848 ;
  assign w850 = \pi101 & w848 ;
  assign w851 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w847 ) | ( \pi129 & w847 ) ;
  assign w852 = ( w849 & w850 ) | ( w849 & w851 ) | ( w850 & w851 ) ;
  assign w853 = \pi103 ^ \pi128 ;
  assign w854 = ( \pi103 & \pi106 ) | ( \pi103 & ~w853 ) | ( \pi106 & ~w853 ) ;
  assign w855 = ( \pi128 & ~\pi129 ) | ( \pi128 & w854 ) | ( ~\pi129 & w854 ) ;
  assign w856 = \pi104 | w855 ;
  assign w857 = \pi105 & w855 ;
  assign w858 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w854 ) | ( \pi129 & w854 ) ;
  assign w859 = ( w856 & w857 ) | ( w856 & w858 ) | ( w857 & w858 ) ;
  assign w860 = \pi130 ^ w838 ;
  assign w861 = ( w838 & w852 ) | ( w838 & w860 ) | ( w852 & w860 ) ;
  assign w862 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w861 ) | ( \pi131 & w861 ) ;
  assign w863 = w845 | w862 ;
  assign w864 = w859 & w862 ;
  assign w865 = ( \pi130 & ~\pi131 ) | ( \pi130 & w861 ) | ( ~\pi131 & w861 ) ;
  assign w866 = ( w863 & w864 ) | ( w863 & w865 ) | ( w864 & w865 ) ;
  assign w867 = \pi132 ^ w762 ;
  assign w868 = ( w762 & w831 ) | ( w762 & ~w867 ) | ( w831 & ~w867 ) ;
  assign w869 = ( \pi132 & ~\pi133 ) | ( \pi132 & w868 ) | ( ~\pi133 & w868 ) ;
  assign w870 = w797 | w869 ;
  assign w871 = w866 & w869 ;
  assign w872 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w868 ) | ( \pi133 & w868 ) ;
  assign w873 = ( w870 & w871 ) | ( w870 & w872 ) | ( w871 & w872 ) ;
  assign w874 = \pi063 ^ \pi128 ;
  assign w875 = ( \pi063 & \pi066 ) | ( \pi063 & ~w874 ) | ( \pi066 & ~w874 ) ;
  assign w876 = ( \pi128 & ~\pi129 ) | ( \pi128 & w875 ) | ( ~\pi129 & w875 ) ;
  assign w877 = \pi064 | w876 ;
  assign w878 = \pi065 & w876 ;
  assign w879 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w875 ) | ( \pi129 & w875 ) ;
  assign w880 = ( w877 & w878 ) | ( w877 & w879 ) | ( w878 & w879 ) ;
  assign w881 = \pi059 ^ \pi128 ;
  assign w882 = ( \pi059 & \pi062 ) | ( \pi059 & ~w881 ) | ( \pi062 & ~w881 ) ;
  assign w883 = ( \pi128 & ~\pi129 ) | ( \pi128 & w882 ) | ( ~\pi129 & w882 ) ;
  assign w884 = \pi060 | w883 ;
  assign w885 = \pi061 & w883 ;
  assign w886 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w882 ) | ( \pi129 & w882 ) ;
  assign w887 = ( w884 & w885 ) | ( w884 & w886 ) | ( w885 & w886 ) ;
  assign w888 = \pi051 ^ \pi128 ;
  assign w889 = ( \pi051 & \pi054 ) | ( \pi051 & ~w888 ) | ( \pi054 & ~w888 ) ;
  assign w890 = ( \pi128 & ~\pi129 ) | ( \pi128 & w889 ) | ( ~\pi129 & w889 ) ;
  assign w891 = \pi052 | w890 ;
  assign w892 = \pi053 & w890 ;
  assign w893 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w889 ) | ( \pi129 & w889 ) ;
  assign w894 = ( w891 & w892 ) | ( w891 & w893 ) | ( w892 & w893 ) ;
  assign w895 = \pi055 ^ \pi128 ;
  assign w896 = ( \pi055 & \pi058 ) | ( \pi055 & ~w895 ) | ( \pi058 & ~w895 ) ;
  assign w897 = ( \pi128 & ~\pi129 ) | ( \pi128 & w896 ) | ( ~\pi129 & w896 ) ;
  assign w898 = \pi056 | w897 ;
  assign w899 = \pi057 & w897 ;
  assign w900 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w896 ) | ( \pi129 & w896 ) ;
  assign w901 = ( w898 & w899 ) | ( w898 & w900 ) | ( w899 & w900 ) ;
  assign w902 = \pi130 ^ w880 ;
  assign w903 = ( w880 & w894 ) | ( w880 & w902 ) | ( w894 & w902 ) ;
  assign w904 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w903 ) | ( \pi131 & w903 ) ;
  assign w905 = w887 | w904 ;
  assign w906 = w901 & w904 ;
  assign w907 = ( \pi130 & ~\pi131 ) | ( \pi130 & w903 ) | ( ~\pi131 & w903 ) ;
  assign w908 = ( w905 & w906 ) | ( w905 & w907 ) | ( w906 & w907 ) ;
  assign w909 = \pi015 ^ \pi128 ;
  assign w910 = ( \pi015 & \pi018 ) | ( \pi015 & ~w909 ) | ( \pi018 & ~w909 ) ;
  assign w911 = ( \pi128 & ~\pi129 ) | ( \pi128 & w910 ) | ( ~\pi129 & w910 ) ;
  assign w912 = \pi016 | w911 ;
  assign w913 = \pi017 & w911 ;
  assign w914 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w910 ) | ( \pi129 & w910 ) ;
  assign w915 = ( w912 & w913 ) | ( w912 & w914 ) | ( w913 & w914 ) ;
  assign w916 = \pi011 ^ \pi128 ;
  assign w917 = ( \pi011 & \pi014 ) | ( \pi011 & ~w916 ) | ( \pi014 & ~w916 ) ;
  assign w918 = ( \pi128 & ~\pi129 ) | ( \pi128 & w917 ) | ( ~\pi129 & w917 ) ;
  assign w919 = \pi012 | w918 ;
  assign w920 = \pi013 & w918 ;
  assign w921 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w917 ) | ( \pi129 & w917 ) ;
  assign w922 = ( w919 & w920 ) | ( w919 & w921 ) | ( w920 & w921 ) ;
  assign w923 = \pi003 ^ \pi128 ;
  assign w924 = ( \pi003 & \pi006 ) | ( \pi003 & ~w923 ) | ( \pi006 & ~w923 ) ;
  assign w925 = ( \pi128 & ~\pi129 ) | ( \pi128 & w924 ) | ( ~\pi129 & w924 ) ;
  assign w926 = \pi004 | w925 ;
  assign w927 = \pi005 & w925 ;
  assign w928 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w924 ) | ( \pi129 & w924 ) ;
  assign w929 = ( w926 & w927 ) | ( w926 & w928 ) | ( w927 & w928 ) ;
  assign w930 = \pi007 ^ \pi128 ;
  assign w931 = ( \pi007 & \pi010 ) | ( \pi007 & ~w930 ) | ( \pi010 & ~w930 ) ;
  assign w932 = ( \pi128 & ~\pi129 ) | ( \pi128 & w931 ) | ( ~\pi129 & w931 ) ;
  assign w933 = \pi008 | w932 ;
  assign w934 = \pi009 & w932 ;
  assign w935 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w931 ) | ( \pi129 & w931 ) ;
  assign w936 = ( w933 & w934 ) | ( w933 & w935 ) | ( w934 & w935 ) ;
  assign w937 = \pi130 ^ w915 ;
  assign w938 = ( w915 & w929 ) | ( w915 & w937 ) | ( w929 & w937 ) ;
  assign w939 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w938 ) | ( \pi131 & w938 ) ;
  assign w940 = w922 | w939 ;
  assign w941 = w936 & w939 ;
  assign w942 = ( \pi130 & ~\pi131 ) | ( \pi130 & w938 ) | ( ~\pi131 & w938 ) ;
  assign w943 = ( w940 & w941 ) | ( w940 & w942 ) | ( w941 & w942 ) ;
  assign w944 = \pi047 ^ \pi128 ;
  assign w945 = ( \pi047 & \pi050 ) | ( \pi047 & ~w944 ) | ( \pi050 & ~w944 ) ;
  assign w946 = ( \pi128 & ~\pi129 ) | ( \pi128 & w945 ) | ( ~\pi129 & w945 ) ;
  assign w947 = \pi048 | w946 ;
  assign w948 = \pi049 & w946 ;
  assign w949 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w945 ) | ( \pi129 & w945 ) ;
  assign w950 = ( w947 & w948 ) | ( w947 & w949 ) | ( w948 & w949 ) ;
  assign w951 = \pi043 ^ \pi128 ;
  assign w952 = ( \pi043 & \pi046 ) | ( \pi043 & ~w951 ) | ( \pi046 & ~w951 ) ;
  assign w953 = ( \pi128 & ~\pi129 ) | ( \pi128 & w952 ) | ( ~\pi129 & w952 ) ;
  assign w954 = \pi044 | w953 ;
  assign w955 = \pi045 & w953 ;
  assign w956 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w952 ) | ( \pi129 & w952 ) ;
  assign w957 = ( w954 & w955 ) | ( w954 & w956 ) | ( w955 & w956 ) ;
  assign w958 = \pi035 ^ \pi128 ;
  assign w959 = ( \pi035 & \pi038 ) | ( \pi035 & ~w958 ) | ( \pi038 & ~w958 ) ;
  assign w960 = ( \pi128 & ~\pi129 ) | ( \pi128 & w959 ) | ( ~\pi129 & w959 ) ;
  assign w961 = \pi036 | w960 ;
  assign w962 = \pi037 & w960 ;
  assign w963 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w959 ) | ( \pi129 & w959 ) ;
  assign w964 = ( w961 & w962 ) | ( w961 & w963 ) | ( w962 & w963 ) ;
  assign w965 = \pi039 ^ \pi128 ;
  assign w966 = ( \pi039 & \pi042 ) | ( \pi039 & ~w965 ) | ( \pi042 & ~w965 ) ;
  assign w967 = ( \pi128 & ~\pi129 ) | ( \pi128 & w966 ) | ( ~\pi129 & w966 ) ;
  assign w968 = \pi040 | w967 ;
  assign w969 = \pi041 & w967 ;
  assign w970 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w966 ) | ( \pi129 & w966 ) ;
  assign w971 = ( w968 & w969 ) | ( w968 & w970 ) | ( w969 & w970 ) ;
  assign w972 = \pi130 ^ w950 ;
  assign w973 = ( w950 & w964 ) | ( w950 & w972 ) | ( w964 & w972 ) ;
  assign w974 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w973 ) | ( \pi131 & w973 ) ;
  assign w975 = w957 | w974 ;
  assign w976 = w971 & w974 ;
  assign w977 = ( \pi130 & ~\pi131 ) | ( \pi130 & w973 ) | ( ~\pi131 & w973 ) ;
  assign w978 = ( w975 & w976 ) | ( w975 & w977 ) | ( w976 & w977 ) ;
  assign w979 = \pi031 ^ \pi128 ;
  assign w980 = ( \pi031 & \pi034 ) | ( \pi031 & ~w979 ) | ( \pi034 & ~w979 ) ;
  assign w981 = ( \pi128 & ~\pi129 ) | ( \pi128 & w980 ) | ( ~\pi129 & w980 ) ;
  assign w982 = \pi032 | w981 ;
  assign w983 = \pi033 & w981 ;
  assign w984 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w980 ) | ( \pi129 & w980 ) ;
  assign w985 = ( w982 & w983 ) | ( w982 & w984 ) | ( w983 & w984 ) ;
  assign w986 = \pi027 ^ \pi128 ;
  assign w987 = ( \pi027 & \pi030 ) | ( \pi027 & ~w986 ) | ( \pi030 & ~w986 ) ;
  assign w988 = ( \pi128 & ~\pi129 ) | ( \pi128 & w987 ) | ( ~\pi129 & w987 ) ;
  assign w989 = \pi028 | w988 ;
  assign w990 = \pi029 & w988 ;
  assign w991 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w987 ) | ( \pi129 & w987 ) ;
  assign w992 = ( w989 & w990 ) | ( w989 & w991 ) | ( w990 & w991 ) ;
  assign w993 = \pi019 ^ \pi128 ;
  assign w994 = ( \pi019 & \pi022 ) | ( \pi019 & ~w993 ) | ( \pi022 & ~w993 ) ;
  assign w995 = ( \pi128 & ~\pi129 ) | ( \pi128 & w994 ) | ( ~\pi129 & w994 ) ;
  assign w996 = \pi020 | w995 ;
  assign w997 = \pi021 & w995 ;
  assign w998 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w994 ) | ( \pi129 & w994 ) ;
  assign w999 = ( w996 & w997 ) | ( w996 & w998 ) | ( w997 & w998 ) ;
  assign w1000 = \pi023 ^ \pi128 ;
  assign w1001 = ( \pi023 & \pi026 ) | ( \pi023 & ~w1000 ) | ( \pi026 & ~w1000 ) ;
  assign w1002 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1001 ) | ( ~\pi129 & w1001 ) ;
  assign w1003 = \pi024 | w1002 ;
  assign w1004 = \pi025 & w1002 ;
  assign w1005 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1001 ) | ( \pi129 & w1001 ) ;
  assign w1006 = ( w1003 & w1004 ) | ( w1003 & w1005 ) | ( w1004 & w1005 ) ;
  assign w1007 = \pi130 ^ w985 ;
  assign w1008 = ( w985 & w999 ) | ( w985 & w1007 ) | ( w999 & w1007 ) ;
  assign w1009 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1008 ) | ( \pi131 & w1008 ) ;
  assign w1010 = w992 | w1009 ;
  assign w1011 = w1006 & w1009 ;
  assign w1012 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1008 ) | ( ~\pi131 & w1008 ) ;
  assign w1013 = ( w1010 & w1011 ) | ( w1010 & w1012 ) | ( w1011 & w1012 ) ;
  assign w1014 = \pi132 ^ w908 ;
  assign w1015 = ( w908 & w943 ) | ( w908 & w1014 ) | ( w943 & w1014 ) ;
  assign w1016 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1015 ) | ( \pi133 & w1015 ) ;
  assign w1017 = w978 | w1016 ;
  assign w1018 = w1013 & w1016 ;
  assign w1019 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1015 ) | ( ~\pi133 & w1015 ) ;
  assign w1020 = ( w1017 & w1018 ) | ( w1017 & w1019 ) | ( w1018 & w1019 ) ;
  assign w1021 = \pi134 ^ w1020 ;
  assign w1022 = ( w873 & w1020 ) | ( w873 & ~w1021 ) | ( w1020 & ~w1021 ) ;
  assign w1023 = \pi112 ^ \pi128 ;
  assign w1024 = ( \pi112 & \pi115 ) | ( \pi112 & ~w1023 ) | ( \pi115 & ~w1023 ) ;
  assign w1025 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1024 ) | ( ~\pi129 & w1024 ) ;
  assign w1026 = \pi113 | w1025 ;
  assign w1027 = \pi114 & w1025 ;
  assign w1028 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1024 ) | ( \pi129 & w1024 ) ;
  assign w1029 = ( w1026 & w1027 ) | ( w1026 & w1028 ) | ( w1027 & w1028 ) ;
  assign w1030 = \pi108 ^ \pi128 ;
  assign w1031 = ( \pi108 & \pi111 ) | ( \pi108 & ~w1030 ) | ( \pi111 & ~w1030 ) ;
  assign w1032 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1031 ) | ( ~\pi129 & w1031 ) ;
  assign w1033 = \pi109 | w1032 ;
  assign w1034 = \pi110 & w1032 ;
  assign w1035 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1031 ) | ( \pi129 & w1031 ) ;
  assign w1036 = ( w1033 & w1034 ) | ( w1033 & w1035 ) | ( w1034 & w1035 ) ;
  assign w1037 = \pi100 ^ \pi128 ;
  assign w1038 = ( \pi100 & \pi103 ) | ( \pi100 & ~w1037 ) | ( \pi103 & ~w1037 ) ;
  assign w1039 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1038 ) | ( ~\pi129 & w1038 ) ;
  assign w1040 = \pi101 | w1039 ;
  assign w1041 = \pi102 & w1039 ;
  assign w1042 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1038 ) | ( \pi129 & w1038 ) ;
  assign w1043 = ( w1040 & w1041 ) | ( w1040 & w1042 ) | ( w1041 & w1042 ) ;
  assign w1044 = \pi104 ^ \pi128 ;
  assign w1045 = ( \pi104 & \pi107 ) | ( \pi104 & ~w1044 ) | ( \pi107 & ~w1044 ) ;
  assign w1046 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1045 ) | ( ~\pi129 & w1045 ) ;
  assign w1047 = \pi105 | w1046 ;
  assign w1048 = \pi106 & w1046 ;
  assign w1049 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1045 ) | ( \pi129 & w1045 ) ;
  assign w1050 = ( w1047 & w1048 ) | ( w1047 & w1049 ) | ( w1048 & w1049 ) ;
  assign w1051 = \pi130 ^ w1029 ;
  assign w1052 = ( w1029 & w1043 ) | ( w1029 & w1051 ) | ( w1043 & w1051 ) ;
  assign w1053 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1052 ) | ( \pi131 & w1052 ) ;
  assign w1054 = w1036 | w1053 ;
  assign w1055 = w1050 & w1053 ;
  assign w1056 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1052 ) | ( ~\pi131 & w1052 ) ;
  assign w1057 = ( w1054 & w1055 ) | ( w1054 & w1056 ) | ( w1055 & w1056 ) ;
  assign w1058 = \pi096 ^ \pi128 ;
  assign w1059 = ( \pi096 & \pi099 ) | ( \pi096 & ~w1058 ) | ( \pi099 & ~w1058 ) ;
  assign w1060 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1059 ) | ( ~\pi129 & w1059 ) ;
  assign w1061 = \pi097 | w1060 ;
  assign w1062 = \pi098 & w1060 ;
  assign w1063 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1059 ) | ( \pi129 & w1059 ) ;
  assign w1064 = ( w1061 & w1062 ) | ( w1061 & w1063 ) | ( w1062 & w1063 ) ;
  assign w1065 = \pi092 ^ \pi128 ;
  assign w1066 = ( \pi092 & \pi095 ) | ( \pi092 & ~w1065 ) | ( \pi095 & ~w1065 ) ;
  assign w1067 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1066 ) | ( ~\pi129 & w1066 ) ;
  assign w1068 = \pi093 | w1067 ;
  assign w1069 = \pi094 & w1067 ;
  assign w1070 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1066 ) | ( \pi129 & w1066 ) ;
  assign w1071 = ( w1068 & w1069 ) | ( w1068 & w1070 ) | ( w1069 & w1070 ) ;
  assign w1072 = \pi084 ^ \pi128 ;
  assign w1073 = ( \pi084 & \pi087 ) | ( \pi084 & ~w1072 ) | ( \pi087 & ~w1072 ) ;
  assign w1074 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1073 ) | ( ~\pi129 & w1073 ) ;
  assign w1075 = \pi085 | w1074 ;
  assign w1076 = \pi086 & w1074 ;
  assign w1077 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1073 ) | ( \pi129 & w1073 ) ;
  assign w1078 = ( w1075 & w1076 ) | ( w1075 & w1077 ) | ( w1076 & w1077 ) ;
  assign w1079 = \pi088 ^ \pi128 ;
  assign w1080 = ( \pi088 & \pi091 ) | ( \pi088 & ~w1079 ) | ( \pi091 & ~w1079 ) ;
  assign w1081 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1080 ) | ( ~\pi129 & w1080 ) ;
  assign w1082 = \pi089 | w1081 ;
  assign w1083 = \pi090 & w1081 ;
  assign w1084 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1080 ) | ( \pi129 & w1080 ) ;
  assign w1085 = ( w1082 & w1083 ) | ( w1082 & w1084 ) | ( w1083 & w1084 ) ;
  assign w1086 = \pi130 ^ w1064 ;
  assign w1087 = ( w1064 & w1078 ) | ( w1064 & w1086 ) | ( w1078 & w1086 ) ;
  assign w1088 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1087 ) | ( \pi131 & w1087 ) ;
  assign w1089 = w1071 | w1088 ;
  assign w1090 = w1085 & w1088 ;
  assign w1091 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1087 ) | ( ~\pi131 & w1087 ) ;
  assign w1092 = ( w1089 & w1090 ) | ( w1089 & w1091 ) | ( w1090 & w1091 ) ;
  assign w1093 = ( \pi000 & \pi003 ) | ( \pi000 & ~w502 ) | ( \pi003 & ~w502 ) ;
  assign w1094 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1093 ) | ( ~\pi129 & w1093 ) ;
  assign w1095 = \pi001 | w1094 ;
  assign w1096 = \pi002 & w1094 ;
  assign w1097 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1093 ) | ( \pi129 & w1093 ) ;
  assign w1098 = ( w1095 & w1096 ) | ( w1095 & w1097 ) | ( w1096 & w1097 ) ;
  assign w1099 = \pi124 ^ \pi128 ;
  assign w1100 = ( \pi124 & \pi127 ) | ( \pi124 & ~w1099 ) | ( \pi127 & ~w1099 ) ;
  assign w1101 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1100 ) | ( ~\pi129 & w1100 ) ;
  assign w1102 = \pi125 | w1101 ;
  assign w1103 = \pi126 & w1101 ;
  assign w1104 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1100 ) | ( \pi129 & w1100 ) ;
  assign w1105 = ( w1102 & w1103 ) | ( w1102 & w1104 ) | ( w1103 & w1104 ) ;
  assign w1106 = \pi116 ^ \pi128 ;
  assign w1107 = ( \pi116 & \pi119 ) | ( \pi116 & ~w1106 ) | ( \pi119 & ~w1106 ) ;
  assign w1108 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1107 ) | ( ~\pi129 & w1107 ) ;
  assign w1109 = \pi117 | w1108 ;
  assign w1110 = \pi118 & w1108 ;
  assign w1111 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1107 ) | ( \pi129 & w1107 ) ;
  assign w1112 = ( w1109 & w1110 ) | ( w1109 & w1111 ) | ( w1110 & w1111 ) ;
  assign w1113 = \pi120 ^ \pi128 ;
  assign w1114 = ( \pi120 & \pi123 ) | ( \pi120 & ~w1113 ) | ( \pi123 & ~w1113 ) ;
  assign w1115 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1114 ) | ( ~\pi129 & w1114 ) ;
  assign w1116 = \pi121 | w1115 ;
  assign w1117 = \pi122 & w1115 ;
  assign w1118 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1114 ) | ( \pi129 & w1114 ) ;
  assign w1119 = ( w1116 & w1117 ) | ( w1116 & w1118 ) | ( w1117 & w1118 ) ;
  assign w1120 = \pi130 ^ w1098 ;
  assign w1121 = ( w1098 & w1112 ) | ( w1098 & w1120 ) | ( w1112 & w1120 ) ;
  assign w1122 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1121 ) | ( \pi131 & w1121 ) ;
  assign w1123 = w1105 | w1122 ;
  assign w1124 = w1119 & w1122 ;
  assign w1125 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1121 ) | ( ~\pi131 & w1121 ) ;
  assign w1126 = ( w1123 & w1124 ) | ( w1123 & w1125 ) | ( w1124 & w1125 ) ;
  assign w1127 = \pi080 ^ \pi128 ;
  assign w1128 = ( \pi080 & \pi083 ) | ( \pi080 & ~w1127 ) | ( \pi083 & ~w1127 ) ;
  assign w1129 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1128 ) | ( ~\pi129 & w1128 ) ;
  assign w1130 = \pi081 | w1129 ;
  assign w1131 = \pi082 & w1129 ;
  assign w1132 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1128 ) | ( \pi129 & w1128 ) ;
  assign w1133 = ( w1130 & w1131 ) | ( w1130 & w1132 ) | ( w1131 & w1132 ) ;
  assign w1134 = \pi076 ^ \pi128 ;
  assign w1135 = ( \pi076 & \pi079 ) | ( \pi076 & ~w1134 ) | ( \pi079 & ~w1134 ) ;
  assign w1136 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1135 ) | ( ~\pi129 & w1135 ) ;
  assign w1137 = \pi077 | w1136 ;
  assign w1138 = \pi078 & w1136 ;
  assign w1139 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1135 ) | ( \pi129 & w1135 ) ;
  assign w1140 = ( w1137 & w1138 ) | ( w1137 & w1139 ) | ( w1138 & w1139 ) ;
  assign w1141 = \pi068 ^ \pi128 ;
  assign w1142 = ( \pi068 & \pi071 ) | ( \pi068 & ~w1141 ) | ( \pi071 & ~w1141 ) ;
  assign w1143 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1142 ) | ( ~\pi129 & w1142 ) ;
  assign w1144 = \pi069 | w1143 ;
  assign w1145 = \pi070 & w1143 ;
  assign w1146 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1142 ) | ( \pi129 & w1142 ) ;
  assign w1147 = ( w1144 & w1145 ) | ( w1144 & w1146 ) | ( w1145 & w1146 ) ;
  assign w1148 = \pi072 ^ \pi128 ;
  assign w1149 = ( \pi072 & \pi075 ) | ( \pi072 & ~w1148 ) | ( \pi075 & ~w1148 ) ;
  assign w1150 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1149 ) | ( ~\pi129 & w1149 ) ;
  assign w1151 = \pi073 | w1150 ;
  assign w1152 = \pi074 & w1150 ;
  assign w1153 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1149 ) | ( \pi129 & w1149 ) ;
  assign w1154 = ( w1151 & w1152 ) | ( w1151 & w1153 ) | ( w1152 & w1153 ) ;
  assign w1155 = \pi130 ^ w1133 ;
  assign w1156 = ( w1133 & w1147 ) | ( w1133 & w1155 ) | ( w1147 & w1155 ) ;
  assign w1157 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1156 ) | ( \pi131 & w1156 ) ;
  assign w1158 = w1140 | w1157 ;
  assign w1159 = w1154 & w1157 ;
  assign w1160 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1156 ) | ( ~\pi131 & w1156 ) ;
  assign w1161 = ( w1158 & w1159 ) | ( w1158 & w1160 ) | ( w1159 & w1160 ) ;
  assign w1162 = \pi132 ^ w1057 ;
  assign w1163 = ( w1057 & w1092 ) | ( w1057 & ~w1162 ) | ( w1092 & ~w1162 ) ;
  assign w1164 = ( \pi132 & \pi133 ) | ( \pi132 & w1163 ) | ( \pi133 & w1163 ) ;
  assign w1165 = w1126 | w1164 ;
  assign w1166 = w1161 & w1164 ;
  assign w1167 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1163 ) | ( \pi133 & ~w1163 ) ;
  assign w1168 = ( w1165 & w1166 ) | ( w1165 & ~w1167 ) | ( w1166 & ~w1167 ) ;
  assign w1169 = \pi064 ^ \pi128 ;
  assign w1170 = ( \pi064 & \pi067 ) | ( \pi064 & ~w1169 ) | ( \pi067 & ~w1169 ) ;
  assign w1171 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1170 ) | ( ~\pi129 & w1170 ) ;
  assign w1172 = \pi065 | w1171 ;
  assign w1173 = \pi066 & w1171 ;
  assign w1174 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1170 ) | ( \pi129 & w1170 ) ;
  assign w1175 = ( w1172 & w1173 ) | ( w1172 & w1174 ) | ( w1173 & w1174 ) ;
  assign w1176 = \pi060 ^ \pi128 ;
  assign w1177 = ( \pi060 & \pi063 ) | ( \pi060 & ~w1176 ) | ( \pi063 & ~w1176 ) ;
  assign w1178 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1177 ) | ( ~\pi129 & w1177 ) ;
  assign w1179 = \pi061 | w1178 ;
  assign w1180 = \pi062 & w1178 ;
  assign w1181 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1177 ) | ( \pi129 & w1177 ) ;
  assign w1182 = ( w1179 & w1180 ) | ( w1179 & w1181 ) | ( w1180 & w1181 ) ;
  assign w1183 = \pi052 ^ \pi128 ;
  assign w1184 = ( \pi052 & \pi055 ) | ( \pi052 & ~w1183 ) | ( \pi055 & ~w1183 ) ;
  assign w1185 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1184 ) | ( ~\pi129 & w1184 ) ;
  assign w1186 = \pi053 | w1185 ;
  assign w1187 = \pi054 & w1185 ;
  assign w1188 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1184 ) | ( \pi129 & w1184 ) ;
  assign w1189 = ( w1186 & w1187 ) | ( w1186 & w1188 ) | ( w1187 & w1188 ) ;
  assign w1190 = \pi056 ^ \pi128 ;
  assign w1191 = ( \pi056 & \pi059 ) | ( \pi056 & ~w1190 ) | ( \pi059 & ~w1190 ) ;
  assign w1192 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1191 ) | ( ~\pi129 & w1191 ) ;
  assign w1193 = \pi057 | w1192 ;
  assign w1194 = \pi058 & w1192 ;
  assign w1195 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1191 ) | ( \pi129 & w1191 ) ;
  assign w1196 = ( w1193 & w1194 ) | ( w1193 & w1195 ) | ( w1194 & w1195 ) ;
  assign w1197 = \pi130 ^ w1175 ;
  assign w1198 = ( w1175 & w1189 ) | ( w1175 & w1197 ) | ( w1189 & w1197 ) ;
  assign w1199 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1198 ) | ( \pi131 & w1198 ) ;
  assign w1200 = w1182 | w1199 ;
  assign w1201 = w1196 & w1199 ;
  assign w1202 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1198 ) | ( ~\pi131 & w1198 ) ;
  assign w1203 = ( w1200 & w1201 ) | ( w1200 & w1202 ) | ( w1201 & w1202 ) ;
  assign w1204 = \pi048 ^ \pi128 ;
  assign w1205 = ( \pi048 & \pi051 ) | ( \pi048 & ~w1204 ) | ( \pi051 & ~w1204 ) ;
  assign w1206 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1205 ) | ( ~\pi129 & w1205 ) ;
  assign w1207 = \pi049 | w1206 ;
  assign w1208 = \pi050 & w1206 ;
  assign w1209 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1205 ) | ( \pi129 & w1205 ) ;
  assign w1210 = ( w1207 & w1208 ) | ( w1207 & w1209 ) | ( w1208 & w1209 ) ;
  assign w1211 = \pi044 ^ \pi128 ;
  assign w1212 = ( \pi044 & \pi047 ) | ( \pi044 & ~w1211 ) | ( \pi047 & ~w1211 ) ;
  assign w1213 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1212 ) | ( ~\pi129 & w1212 ) ;
  assign w1214 = \pi045 | w1213 ;
  assign w1215 = \pi046 & w1213 ;
  assign w1216 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1212 ) | ( \pi129 & w1212 ) ;
  assign w1217 = ( w1214 & w1215 ) | ( w1214 & w1216 ) | ( w1215 & w1216 ) ;
  assign w1218 = \pi036 ^ \pi128 ;
  assign w1219 = ( \pi036 & \pi039 ) | ( \pi036 & ~w1218 ) | ( \pi039 & ~w1218 ) ;
  assign w1220 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1219 ) | ( ~\pi129 & w1219 ) ;
  assign w1221 = \pi037 | w1220 ;
  assign w1222 = \pi038 & w1220 ;
  assign w1223 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1219 ) | ( \pi129 & w1219 ) ;
  assign w1224 = ( w1221 & w1222 ) | ( w1221 & w1223 ) | ( w1222 & w1223 ) ;
  assign w1225 = \pi040 ^ \pi128 ;
  assign w1226 = ( \pi040 & \pi043 ) | ( \pi040 & ~w1225 ) | ( \pi043 & ~w1225 ) ;
  assign w1227 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1226 ) | ( ~\pi129 & w1226 ) ;
  assign w1228 = \pi041 | w1227 ;
  assign w1229 = \pi042 & w1227 ;
  assign w1230 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1226 ) | ( \pi129 & w1226 ) ;
  assign w1231 = ( w1228 & w1229 ) | ( w1228 & w1230 ) | ( w1229 & w1230 ) ;
  assign w1232 = \pi130 ^ w1210 ;
  assign w1233 = ( w1210 & w1224 ) | ( w1210 & w1232 ) | ( w1224 & w1232 ) ;
  assign w1234 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1233 ) | ( \pi131 & w1233 ) ;
  assign w1235 = w1217 | w1234 ;
  assign w1236 = w1231 & w1234 ;
  assign w1237 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1233 ) | ( ~\pi131 & w1233 ) ;
  assign w1238 = ( w1235 & w1236 ) | ( w1235 & w1237 ) | ( w1236 & w1237 ) ;
  assign w1239 = \pi016 ^ \pi128 ;
  assign w1240 = ( \pi016 & \pi019 ) | ( \pi016 & ~w1239 ) | ( \pi019 & ~w1239 ) ;
  assign w1241 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1240 ) | ( ~\pi129 & w1240 ) ;
  assign w1242 = \pi017 | w1241 ;
  assign w1243 = \pi018 & w1241 ;
  assign w1244 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1240 ) | ( \pi129 & w1240 ) ;
  assign w1245 = ( w1242 & w1243 ) | ( w1242 & w1244 ) | ( w1243 & w1244 ) ;
  assign w1246 = \pi012 ^ \pi128 ;
  assign w1247 = ( \pi012 & \pi015 ) | ( \pi012 & ~w1246 ) | ( \pi015 & ~w1246 ) ;
  assign w1248 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1247 ) | ( ~\pi129 & w1247 ) ;
  assign w1249 = \pi013 | w1248 ;
  assign w1250 = \pi014 & w1248 ;
  assign w1251 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1247 ) | ( \pi129 & w1247 ) ;
  assign w1252 = ( w1249 & w1250 ) | ( w1249 & w1251 ) | ( w1250 & w1251 ) ;
  assign w1253 = \pi004 ^ \pi128 ;
  assign w1254 = ( \pi004 & \pi007 ) | ( \pi004 & ~w1253 ) | ( \pi007 & ~w1253 ) ;
  assign w1255 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1254 ) | ( ~\pi129 & w1254 ) ;
  assign w1256 = \pi005 | w1255 ;
  assign w1257 = \pi006 & w1255 ;
  assign w1258 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1254 ) | ( \pi129 & w1254 ) ;
  assign w1259 = ( w1256 & w1257 ) | ( w1256 & w1258 ) | ( w1257 & w1258 ) ;
  assign w1260 = \pi008 ^ \pi128 ;
  assign w1261 = ( \pi008 & \pi011 ) | ( \pi008 & ~w1260 ) | ( \pi011 & ~w1260 ) ;
  assign w1262 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1261 ) | ( ~\pi129 & w1261 ) ;
  assign w1263 = \pi009 | w1262 ;
  assign w1264 = \pi010 & w1262 ;
  assign w1265 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1261 ) | ( \pi129 & w1261 ) ;
  assign w1266 = ( w1263 & w1264 ) | ( w1263 & w1265 ) | ( w1264 & w1265 ) ;
  assign w1267 = \pi130 ^ w1245 ;
  assign w1268 = ( w1245 & w1259 ) | ( w1245 & w1267 ) | ( w1259 & w1267 ) ;
  assign w1269 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1268 ) | ( \pi131 & w1268 ) ;
  assign w1270 = w1252 | w1269 ;
  assign w1271 = w1266 & w1269 ;
  assign w1272 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1268 ) | ( ~\pi131 & w1268 ) ;
  assign w1273 = ( w1270 & w1271 ) | ( w1270 & w1272 ) | ( w1271 & w1272 ) ;
  assign w1274 = \pi032 ^ \pi128 ;
  assign w1275 = ( \pi032 & \pi035 ) | ( \pi032 & ~w1274 ) | ( \pi035 & ~w1274 ) ;
  assign w1276 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1275 ) | ( ~\pi129 & w1275 ) ;
  assign w1277 = \pi033 | w1276 ;
  assign w1278 = \pi034 & w1276 ;
  assign w1279 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1275 ) | ( \pi129 & w1275 ) ;
  assign w1280 = ( w1277 & w1278 ) | ( w1277 & w1279 ) | ( w1278 & w1279 ) ;
  assign w1281 = \pi028 ^ \pi128 ;
  assign w1282 = ( \pi028 & \pi031 ) | ( \pi028 & ~w1281 ) | ( \pi031 & ~w1281 ) ;
  assign w1283 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1282 ) | ( ~\pi129 & w1282 ) ;
  assign w1284 = \pi029 | w1283 ;
  assign w1285 = \pi030 & w1283 ;
  assign w1286 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1282 ) | ( \pi129 & w1282 ) ;
  assign w1287 = ( w1284 & w1285 ) | ( w1284 & w1286 ) | ( w1285 & w1286 ) ;
  assign w1288 = \pi020 ^ \pi128 ;
  assign w1289 = ( \pi020 & \pi023 ) | ( \pi020 & ~w1288 ) | ( \pi023 & ~w1288 ) ;
  assign w1290 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1289 ) | ( ~\pi129 & w1289 ) ;
  assign w1291 = \pi021 | w1290 ;
  assign w1292 = \pi022 & w1290 ;
  assign w1293 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1289 ) | ( \pi129 & w1289 ) ;
  assign w1294 = ( w1291 & w1292 ) | ( w1291 & w1293 ) | ( w1292 & w1293 ) ;
  assign w1295 = \pi024 ^ \pi128 ;
  assign w1296 = ( \pi024 & \pi027 ) | ( \pi024 & ~w1295 ) | ( \pi027 & ~w1295 ) ;
  assign w1297 = ( \pi128 & ~\pi129 ) | ( \pi128 & w1296 ) | ( ~\pi129 & w1296 ) ;
  assign w1298 = \pi025 | w1297 ;
  assign w1299 = \pi026 & w1297 ;
  assign w1300 = ( ~\pi128 & \pi129 ) | ( ~\pi128 & w1296 ) | ( \pi129 & w1296 ) ;
  assign w1301 = ( w1298 & w1299 ) | ( w1298 & w1300 ) | ( w1299 & w1300 ) ;
  assign w1302 = \pi130 ^ w1280 ;
  assign w1303 = ( w1280 & w1294 ) | ( w1280 & w1302 ) | ( w1294 & w1302 ) ;
  assign w1304 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1303 ) | ( \pi131 & w1303 ) ;
  assign w1305 = w1287 | w1304 ;
  assign w1306 = w1301 & w1304 ;
  assign w1307 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1303 ) | ( ~\pi131 & w1303 ) ;
  assign w1308 = ( w1305 & w1306 ) | ( w1305 & w1307 ) | ( w1306 & w1307 ) ;
  assign w1309 = \pi132 ^ w1203 ;
  assign w1310 = ( w1203 & w1273 ) | ( w1203 & w1309 ) | ( w1273 & w1309 ) ;
  assign w1311 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1310 ) | ( \pi133 & w1310 ) ;
  assign w1312 = w1238 | w1311 ;
  assign w1313 = w1308 & w1311 ;
  assign w1314 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1310 ) | ( ~\pi133 & w1310 ) ;
  assign w1315 = ( w1312 & w1313 ) | ( w1312 & w1314 ) | ( w1313 & w1314 ) ;
  assign w1316 = \pi134 ^ w1315 ;
  assign w1317 = ( w1168 & w1315 ) | ( w1168 & ~w1316 ) | ( w1315 & ~w1316 ) ;
  assign w1318 = \pi131 ^ w142 ;
  assign w1319 = ( w142 & w149 ) | ( w142 & w1318 ) | ( w149 & w1318 ) ;
  assign w1320 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1319 ) | ( \pi131 & ~w1319 ) ;
  assign w1321 = ~w163 & w1320 ;
  assign w1322 = w191 & ~w1320 ;
  assign w1323 = ( \pi130 & \pi131 ) | ( \pi130 & w1319 ) | ( \pi131 & w1319 ) ;
  assign w1324 = ( ~w1321 & w1322 ) | ( ~w1321 & w1323 ) | ( w1322 & w1323 ) ;
  assign w1325 = \pi131 ^ w177 ;
  assign w1326 = ( w177 & w184 ) | ( w177 & w1325 ) | ( w184 & w1325 ) ;
  assign w1327 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1326 ) | ( \pi131 & ~w1326 ) ;
  assign w1328 = ~w198 & w1327 ;
  assign w1329 = w261 & ~w1327 ;
  assign w1330 = ( \pi130 & \pi131 ) | ( \pi130 & w1326 ) | ( \pi131 & w1326 ) ;
  assign w1331 = ( ~w1328 & w1329 ) | ( ~w1328 & w1330 ) | ( w1329 & w1330 ) ;
  assign w1332 = \pi131 ^ w212 ;
  assign w1333 = ( w212 & w219 ) | ( w212 & w1332 ) | ( w219 & w1332 ) ;
  assign w1334 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1333 ) | ( \pi131 & ~w1333 ) ;
  assign w1335 = ~w233 & w1334 ;
  assign w1336 = w303 & ~w1334 ;
  assign w1337 = ( \pi130 & \pi131 ) | ( \pi130 & w1333 ) | ( \pi131 & w1333 ) ;
  assign w1338 = ( ~w1335 & w1336 ) | ( ~w1335 & w1337 ) | ( w1336 & w1337 ) ;
  assign w1339 = \pi130 ^ w226 ;
  assign w1340 = ( w226 & w268 ) | ( w226 & w1339 ) | ( w268 & w1339 ) ;
  assign w1341 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1340 ) | ( \pi131 & w1340 ) ;
  assign w1342 = w247 | w1341 ;
  assign w1343 = w254 & w1341 ;
  assign w1344 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1340 ) | ( ~\pi131 & w1340 ) ;
  assign w1345 = ( w1342 & w1343 ) | ( w1342 & w1344 ) | ( w1343 & w1344 ) ;
  assign w1346 = \pi132 ^ w1324 ;
  assign w1347 = ( w1324 & w1338 ) | ( w1324 & ~w1346 ) | ( w1338 & ~w1346 ) ;
  assign w1348 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1347 ) | ( ~\pi133 & w1347 ) ;
  assign w1349 = w1331 | w1348 ;
  assign w1350 = w1345 & w1348 ;
  assign w1351 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1347 ) | ( \pi133 & w1347 ) ;
  assign w1352 = ( w1349 & w1350 ) | ( w1349 & w1351 ) | ( w1350 & w1351 ) ;
  assign w1353 = \pi130 ^ w373 ;
  assign w1354 = ( w373 & w415 ) | ( w373 & w1353 ) | ( w415 & w1353 ) ;
  assign w1355 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1354 ) | ( \pi131 & w1354 ) ;
  assign w1356 = w394 | w1355 ;
  assign w1357 = w401 & w1355 ;
  assign w1358 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1354 ) | ( ~\pi131 & w1354 ) ;
  assign w1359 = ( w1356 & w1357 ) | ( w1356 & w1358 ) | ( w1357 & w1358 ) ;
  assign w1360 = \pi130 ^ w156 ;
  assign w1361 = ( w156 & w380 ) | ( w156 & w1360 ) | ( w380 & w1360 ) ;
  assign w1362 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1361 ) | ( \pi131 & w1361 ) ;
  assign w1363 = w359 | w1362 ;
  assign w1364 = w366 & w1362 ;
  assign w1365 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1361 ) | ( ~\pi131 & w1361 ) ;
  assign w1366 = ( w1363 & w1364 ) | ( w1363 & w1365 ) | ( w1364 & w1365 ) ;
  assign w1367 = \pi131 ^ w324 ;
  assign w1368 = ( w324 & w331 ) | ( w324 & w1367 ) | ( w331 & w1367 ) ;
  assign w1369 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1368 ) | ( \pi131 & ~w1368 ) ;
  assign w1370 = ~w345 & w1369 ;
  assign w1371 = w408 & ~w1369 ;
  assign w1372 = ( \pi130 & \pi131 ) | ( \pi130 & w1368 ) | ( \pi131 & w1368 ) ;
  assign w1373 = ( ~w1370 & w1371 ) | ( ~w1370 & w1372 ) | ( w1371 & w1372 ) ;
  assign w1374 = \pi131 ^ w289 ;
  assign w1375 = ( w289 & w296 ) | ( w289 & w1374 ) | ( w296 & w1374 ) ;
  assign w1376 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1375 ) | ( \pi131 & ~w1375 ) ;
  assign w1377 = ~w310 & w1376 ;
  assign w1378 = w338 & ~w1376 ;
  assign w1379 = ( \pi130 & \pi131 ) | ( \pi130 & w1375 ) | ( \pi131 & w1375 ) ;
  assign w1380 = ( ~w1377 & w1378 ) | ( ~w1377 & w1379 ) | ( w1378 & w1379 ) ;
  assign w1381 = \pi132 ^ w1359 ;
  assign w1382 = ( w1359 & w1373 ) | ( w1359 & ~w1381 ) | ( w1373 & ~w1381 ) ;
  assign w1383 = ( \pi132 & \pi133 ) | ( \pi132 & w1382 ) | ( \pi133 & w1382 ) ;
  assign w1384 = w1366 | w1383 ;
  assign w1385 = w1380 & w1383 ;
  assign w1386 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1382 ) | ( \pi133 & ~w1382 ) ;
  assign w1387 = ( w1384 & w1385 ) | ( w1384 & ~w1386 ) | ( w1385 & ~w1386 ) ;
  assign w1388 = \pi134 ^ w1387 ;
  assign w1389 = ( w1352 & w1387 ) | ( w1352 & ~w1388 ) | ( w1387 & ~w1388 ) ;
  assign w1390 = \pi131 ^ w438 ;
  assign w1391 = ( w438 & w445 ) | ( w438 & w1390 ) | ( w445 & w1390 ) ;
  assign w1392 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1391 ) | ( \pi131 & ~w1391 ) ;
  assign w1393 = ~w459 & w1392 ;
  assign w1394 = w487 & ~w1392 ;
  assign w1395 = ( \pi130 & \pi131 ) | ( \pi130 & w1391 ) | ( \pi131 & w1391 ) ;
  assign w1396 = ( ~w1393 & w1394 ) | ( ~w1393 & w1395 ) | ( w1394 & w1395 ) ;
  assign w1397 = \pi131 ^ w473 ;
  assign w1398 = ( w473 & w480 ) | ( w473 & w1397 ) | ( w480 & w1397 ) ;
  assign w1399 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1398 ) | ( \pi131 & ~w1398 ) ;
  assign w1400 = ~w494 & w1399 ;
  assign w1401 = w557 & ~w1399 ;
  assign w1402 = ( \pi130 & \pi131 ) | ( \pi130 & w1398 ) | ( \pi131 & w1398 ) ;
  assign w1403 = ( ~w1400 & w1401 ) | ( ~w1400 & w1402 ) | ( w1401 & w1402 ) ;
  assign w1404 = \pi131 ^ w508 ;
  assign w1405 = ( w508 & w515 ) | ( w508 & w1404 ) | ( w515 & w1404 ) ;
  assign w1406 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1405 ) | ( \pi131 & ~w1405 ) ;
  assign w1407 = ~w529 & w1406 ;
  assign w1408 = w634 & ~w1406 ;
  assign w1409 = ( \pi130 & \pi131 ) | ( \pi130 & w1405 ) | ( \pi131 & w1405 ) ;
  assign w1410 = ( ~w1407 & w1408 ) | ( ~w1407 & w1409 ) | ( w1408 & w1409 ) ;
  assign w1411 = \pi130 ^ w522 ;
  assign w1412 = ( w522 & w564 ) | ( w522 & w1411 ) | ( w564 & w1411 ) ;
  assign w1413 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1412 ) | ( \pi131 & w1412 ) ;
  assign w1414 = w543 | w1413 ;
  assign w1415 = w550 & w1413 ;
  assign w1416 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1412 ) | ( ~\pi131 & w1412 ) ;
  assign w1417 = ( w1414 & w1415 ) | ( w1414 & w1416 ) | ( w1415 & w1416 ) ;
  assign w1418 = \pi132 ^ w1396 ;
  assign w1419 = ( w1396 & w1410 ) | ( w1396 & ~w1418 ) | ( w1410 & ~w1418 ) ;
  assign w1420 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1419 ) | ( ~\pi133 & w1419 ) ;
  assign w1421 = w1403 | w1420 ;
  assign w1422 = w1417 & w1420 ;
  assign w1423 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1419 ) | ( \pi133 & w1419 ) ;
  assign w1424 = ( w1421 & w1422 ) | ( w1421 & w1423 ) | ( w1422 & w1423 ) ;
  assign w1425 = \pi130 ^ w599 ;
  assign w1426 = ( w599 & w676 ) | ( w599 & w1425 ) | ( w676 & w1425 ) ;
  assign w1427 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1426 ) | ( \pi131 & w1426 ) ;
  assign w1428 = w655 | w1427 ;
  assign w1429 = w662 & w1427 ;
  assign w1430 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1426 ) | ( ~\pi131 & w1426 ) ;
  assign w1431 = ( w1428 & w1429 ) | ( w1428 & w1430 ) | ( w1429 & w1430 ) ;
  assign w1432 = \pi130 ^ w452 ;
  assign w1433 = ( w452 & w606 ) | ( w452 & w1432 ) | ( w606 & w1432 ) ;
  assign w1434 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1433 ) | ( \pi131 & w1433 ) ;
  assign w1435 = w585 | w1434 ;
  assign w1436 = w592 & w1434 ;
  assign w1437 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1433 ) | ( ~\pi131 & w1433 ) ;
  assign w1438 = ( w1435 & w1436 ) | ( w1435 & w1437 ) | ( w1436 & w1437 ) ;
  assign w1439 = \pi130 ^ w669 ;
  assign w1440 = ( w669 & w711 ) | ( w669 & w1439 ) | ( w711 & w1439 ) ;
  assign w1441 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1440 ) | ( \pi131 & w1440 ) ;
  assign w1442 = w690 | w1441 ;
  assign w1443 = w697 & w1441 ;
  assign w1444 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1440 ) | ( ~\pi131 & w1440 ) ;
  assign w1445 = ( w1442 & w1443 ) | ( w1442 & w1444 ) | ( w1443 & w1444 ) ;
  assign w1446 = \pi131 ^ w620 ;
  assign w1447 = ( w620 & w627 ) | ( w620 & w1446 ) | ( w627 & w1446 ) ;
  assign w1448 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1447 ) | ( \pi131 & ~w1447 ) ;
  assign w1449 = ~w641 & w1448 ;
  assign w1450 = w704 & ~w1448 ;
  assign w1451 = ( \pi130 & \pi131 ) | ( \pi130 & w1447 ) | ( \pi131 & w1447 ) ;
  assign w1452 = ( ~w1449 & w1450 ) | ( ~w1449 & w1451 ) | ( w1450 & w1451 ) ;
  assign w1453 = \pi132 ^ w1431 ;
  assign w1454 = ( w1431 & w1445 ) | ( w1431 & ~w1453 ) | ( w1445 & ~w1453 ) ;
  assign w1455 = ( \pi132 & \pi133 ) | ( \pi132 & w1454 ) | ( \pi133 & w1454 ) ;
  assign w1456 = w1438 | w1455 ;
  assign w1457 = w1452 & w1455 ;
  assign w1458 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1454 ) | ( \pi133 & ~w1454 ) ;
  assign w1459 = ( w1456 & w1457 ) | ( w1456 & ~w1458 ) | ( w1457 & ~w1458 ) ;
  assign w1460 = \pi134 ^ w1459 ;
  assign w1461 = ( w1424 & w1459 ) | ( w1424 & ~w1460 ) | ( w1459 & ~w1460 ) ;
  assign w1462 = \pi131 ^ w734 ;
  assign w1463 = ( w734 & w741 ) | ( w734 & w1462 ) | ( w741 & w1462 ) ;
  assign w1464 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1463 ) | ( \pi131 & ~w1463 ) ;
  assign w1465 = ~w755 & w1464 ;
  assign w1466 = w783 & ~w1464 ;
  assign w1467 = ( \pi130 & \pi131 ) | ( \pi130 & w1463 ) | ( \pi131 & w1463 ) ;
  assign w1468 = ( ~w1465 & w1466 ) | ( ~w1465 & w1467 ) | ( w1466 & w1467 ) ;
  assign w1469 = \pi131 ^ w769 ;
  assign w1470 = ( w769 & w776 ) | ( w769 & w1469 ) | ( w776 & w1469 ) ;
  assign w1471 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1470 ) | ( \pi131 & ~w1470 ) ;
  assign w1472 = ~w790 & w1471 ;
  assign w1473 = w852 & ~w1471 ;
  assign w1474 = ( \pi130 & \pi131 ) | ( \pi130 & w1470 ) | ( \pi131 & w1470 ) ;
  assign w1475 = ( ~w1472 & w1473 ) | ( ~w1472 & w1474 ) | ( w1473 & w1474 ) ;
  assign w1476 = \pi131 ^ w803 ;
  assign w1477 = ( w803 & w810 ) | ( w803 & w1476 ) | ( w810 & w1476 ) ;
  assign w1478 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1477 ) | ( \pi131 & ~w1477 ) ;
  assign w1479 = ~w824 & w1478 ;
  assign w1480 = w929 & ~w1478 ;
  assign w1481 = ( \pi130 & \pi131 ) | ( \pi130 & w1477 ) | ( \pi131 & w1477 ) ;
  assign w1482 = ( ~w1479 & w1480 ) | ( ~w1479 & w1481 ) | ( w1480 & w1481 ) ;
  assign w1483 = \pi130 ^ w817 ;
  assign w1484 = ( w817 & w859 ) | ( w817 & w1483 ) | ( w859 & w1483 ) ;
  assign w1485 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1484 ) | ( \pi131 & w1484 ) ;
  assign w1486 = w838 | w1485 ;
  assign w1487 = w845 & w1485 ;
  assign w1488 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1484 ) | ( ~\pi131 & w1484 ) ;
  assign w1489 = ( w1486 & w1487 ) | ( w1486 & w1488 ) | ( w1487 & w1488 ) ;
  assign w1490 = \pi132 ^ w1468 ;
  assign w1491 = ( w1468 & w1482 ) | ( w1468 & ~w1490 ) | ( w1482 & ~w1490 ) ;
  assign w1492 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1491 ) | ( ~\pi133 & w1491 ) ;
  assign w1493 = w1475 | w1492 ;
  assign w1494 = w1489 & w1492 ;
  assign w1495 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1491 ) | ( \pi133 & w1491 ) ;
  assign w1496 = ( w1493 & w1494 ) | ( w1493 & w1495 ) | ( w1494 & w1495 ) ;
  assign w1497 = \pi130 ^ w894 ;
  assign w1498 = ( w894 & w971 ) | ( w894 & w1497 ) | ( w971 & w1497 ) ;
  assign w1499 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1498 ) | ( \pi131 & w1498 ) ;
  assign w1500 = w950 | w1499 ;
  assign w1501 = w957 & w1499 ;
  assign w1502 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1498 ) | ( ~\pi131 & w1498 ) ;
  assign w1503 = ( w1500 & w1501 ) | ( w1500 & w1502 ) | ( w1501 & w1502 ) ;
  assign w1504 = \pi130 ^ w748 ;
  assign w1505 = ( w748 & w901 ) | ( w748 & w1504 ) | ( w901 & w1504 ) ;
  assign w1506 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1505 ) | ( \pi131 & w1505 ) ;
  assign w1507 = w880 | w1506 ;
  assign w1508 = w887 & w1506 ;
  assign w1509 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1505 ) | ( ~\pi131 & w1505 ) ;
  assign w1510 = ( w1507 & w1508 ) | ( w1507 & w1509 ) | ( w1508 & w1509 ) ;
  assign w1511 = \pi130 ^ w964 ;
  assign w1512 = ( w964 & w1006 ) | ( w964 & w1511 ) | ( w1006 & w1511 ) ;
  assign w1513 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1512 ) | ( \pi131 & w1512 ) ;
  assign w1514 = w985 | w1513 ;
  assign w1515 = w992 & w1513 ;
  assign w1516 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1512 ) | ( ~\pi131 & w1512 ) ;
  assign w1517 = ( w1514 & w1515 ) | ( w1514 & w1516 ) | ( w1515 & w1516 ) ;
  assign w1518 = \pi131 ^ w915 ;
  assign w1519 = ( w915 & w922 ) | ( w915 & w1518 ) | ( w922 & w1518 ) ;
  assign w1520 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1519 ) | ( \pi131 & ~w1519 ) ;
  assign w1521 = ~w936 & w1520 ;
  assign w1522 = w999 & ~w1520 ;
  assign w1523 = ( \pi130 & \pi131 ) | ( \pi130 & w1519 ) | ( \pi131 & w1519 ) ;
  assign w1524 = ( ~w1521 & w1522 ) | ( ~w1521 & w1523 ) | ( w1522 & w1523 ) ;
  assign w1525 = \pi132 ^ w1503 ;
  assign w1526 = ( w1503 & w1517 ) | ( w1503 & ~w1525 ) | ( w1517 & ~w1525 ) ;
  assign w1527 = ( \pi132 & \pi133 ) | ( \pi132 & w1526 ) | ( \pi133 & w1526 ) ;
  assign w1528 = w1510 | w1527 ;
  assign w1529 = w1524 & w1527 ;
  assign w1530 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1526 ) | ( \pi133 & ~w1526 ) ;
  assign w1531 = ( w1528 & w1529 ) | ( w1528 & ~w1530 ) | ( w1529 & ~w1530 ) ;
  assign w1532 = \pi134 ^ w1531 ;
  assign w1533 = ( w1496 & w1531 ) | ( w1496 & ~w1532 ) | ( w1531 & ~w1532 ) ;
  assign w1534 = \pi130 ^ w1078 ;
  assign w1535 = ( w1078 & w1154 ) | ( w1078 & w1534 ) | ( w1154 & w1534 ) ;
  assign w1536 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1535 ) | ( \pi131 & w1535 ) ;
  assign w1537 = w1133 | w1536 ;
  assign w1538 = w1140 & w1536 ;
  assign w1539 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1535 ) | ( ~\pi131 & w1535 ) ;
  assign w1540 = ( w1537 & w1538 ) | ( w1537 & w1539 ) | ( w1538 & w1539 ) ;
  assign w1541 = \pi130 ^ w1043 ;
  assign w1542 = ( w1043 & w1085 ) | ( w1043 & w1541 ) | ( w1085 & w1541 ) ;
  assign w1543 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1542 ) | ( \pi131 & w1542 ) ;
  assign w1544 = w1064 | w1543 ;
  assign w1545 = w1071 & w1543 ;
  assign w1546 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1542 ) | ( ~\pi131 & w1542 ) ;
  assign w1547 = ( w1544 & w1545 ) | ( w1544 & w1546 ) | ( w1545 & w1546 ) ;
  assign w1548 = \pi131 ^ w1098 ;
  assign w1549 = ( w1098 & w1105 ) | ( w1098 & w1548 ) | ( w1105 & w1548 ) ;
  assign w1550 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1549 ) | ( \pi131 & ~w1549 ) ;
  assign w1551 = ~w1119 & w1550 ;
  assign w1552 = w1259 & ~w1550 ;
  assign w1553 = ( \pi130 & \pi131 ) | ( \pi130 & w1549 ) | ( \pi131 & w1549 ) ;
  assign w1554 = ( ~w1551 & w1552 ) | ( ~w1551 & w1553 ) | ( w1552 & w1553 ) ;
  assign w1555 = \pi131 ^ w1029 ;
  assign w1556 = ( w1029 & w1036 ) | ( w1029 & w1555 ) | ( w1036 & w1555 ) ;
  assign w1557 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1556 ) | ( \pi131 & ~w1556 ) ;
  assign w1558 = ~w1050 & w1557 ;
  assign w1559 = w1112 & ~w1557 ;
  assign w1560 = ( \pi130 & \pi131 ) | ( \pi130 & w1556 ) | ( \pi131 & w1556 ) ;
  assign w1561 = ( ~w1558 & w1559 ) | ( ~w1558 & w1560 ) | ( w1559 & w1560 ) ;
  assign w1562 = \pi132 ^ w1540 ;
  assign w1563 = ( w1540 & w1554 ) | ( w1540 & ~w1562 ) | ( w1554 & ~w1562 ) ;
  assign w1564 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1563 ) | ( ~\pi133 & w1563 ) ;
  assign w1565 = w1547 | w1564 ;
  assign w1566 = w1561 & w1564 ;
  assign w1567 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1563 ) | ( \pi133 & w1563 ) ;
  assign w1568 = ( w1565 & w1566 ) | ( w1565 & w1567 ) | ( w1566 & w1567 ) ;
  assign w1569 = \pi130 ^ w1189 ;
  assign w1570 = ( w1189 & w1231 ) | ( w1189 & w1569 ) | ( w1231 & w1569 ) ;
  assign w1571 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1570 ) | ( \pi131 & w1570 ) ;
  assign w1572 = w1210 | w1571 ;
  assign w1573 = w1217 & w1571 ;
  assign w1574 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1570 ) | ( ~\pi131 & w1570 ) ;
  assign w1575 = ( w1572 & w1573 ) | ( w1572 & w1574 ) | ( w1573 & w1574 ) ;
  assign w1576 = \pi130 ^ w1147 ;
  assign w1577 = ( w1147 & w1196 ) | ( w1147 & w1576 ) | ( w1196 & w1576 ) ;
  assign w1578 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1577 ) | ( \pi131 & w1577 ) ;
  assign w1579 = w1175 | w1578 ;
  assign w1580 = w1182 & w1578 ;
  assign w1581 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1577 ) | ( ~\pi131 & w1577 ) ;
  assign w1582 = ( w1579 & w1580 ) | ( w1579 & w1581 ) | ( w1580 & w1581 ) ;
  assign w1583 = \pi130 ^ w1224 ;
  assign w1584 = ( w1224 & w1301 ) | ( w1224 & w1583 ) | ( w1301 & w1583 ) ;
  assign w1585 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1584 ) | ( \pi131 & w1584 ) ;
  assign w1586 = w1280 | w1585 ;
  assign w1587 = w1287 & w1585 ;
  assign w1588 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1584 ) | ( ~\pi131 & w1584 ) ;
  assign w1589 = ( w1586 & w1587 ) | ( w1586 & w1588 ) | ( w1587 & w1588 ) ;
  assign w1590 = \pi131 ^ w1245 ;
  assign w1591 = ( w1245 & w1252 ) | ( w1245 & w1590 ) | ( w1252 & w1590 ) ;
  assign w1592 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1591 ) | ( \pi131 & ~w1591 ) ;
  assign w1593 = ~w1266 & w1592 ;
  assign w1594 = w1294 & ~w1592 ;
  assign w1595 = ( \pi130 & \pi131 ) | ( \pi130 & w1591 ) | ( \pi131 & w1591 ) ;
  assign w1596 = ( ~w1593 & w1594 ) | ( ~w1593 & w1595 ) | ( w1594 & w1595 ) ;
  assign w1597 = \pi132 ^ w1575 ;
  assign w1598 = ( w1575 & w1589 ) | ( w1575 & ~w1597 ) | ( w1589 & ~w1597 ) ;
  assign w1599 = ( \pi132 & \pi133 ) | ( \pi132 & w1598 ) | ( \pi133 & w1598 ) ;
  assign w1600 = w1582 | w1599 ;
  assign w1601 = w1596 & w1599 ;
  assign w1602 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1598 ) | ( \pi133 & ~w1598 ) ;
  assign w1603 = ( w1600 & w1601 ) | ( w1600 & ~w1602 ) | ( w1601 & ~w1602 ) ;
  assign w1604 = \pi134 ^ w1603 ;
  assign w1605 = ( w1568 & w1603 ) | ( w1568 & ~w1604 ) | ( w1603 & ~w1604 ) ;
  assign w1606 = ( w142 & w164 ) | ( w142 & w191 ) | ( w164 & w191 ) ;
  assign w1607 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1606 ) | ( \pi131 & ~w1606 ) ;
  assign w1608 = ~w149 & w1607 ;
  assign w1609 = w198 & ~w1607 ;
  assign w1610 = ( \pi130 & \pi131 ) | ( \pi130 & w1606 ) | ( \pi131 & w1606 ) ;
  assign w1611 = ( ~w1608 & w1609 ) | ( ~w1608 & w1610 ) | ( w1609 & w1610 ) ;
  assign w1612 = ( w177 & w199 ) | ( w177 & w261 ) | ( w199 & w261 ) ;
  assign w1613 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1612 ) | ( \pi131 & ~w1612 ) ;
  assign w1614 = ~w184 & w1613 ;
  assign w1615 = w268 & ~w1613 ;
  assign w1616 = ( \pi130 & \pi131 ) | ( \pi130 & w1612 ) | ( \pi131 & w1612 ) ;
  assign w1617 = ( ~w1614 & w1615 ) | ( ~w1614 & w1616 ) | ( w1615 & w1616 ) ;
  assign w1618 = ( w212 & w234 ) | ( w212 & w303 ) | ( w234 & w303 ) ;
  assign w1619 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1618 ) | ( \pi131 & ~w1618 ) ;
  assign w1620 = ~w219 & w1619 ;
  assign w1621 = w310 & ~w1619 ;
  assign w1622 = ( \pi130 & \pi131 ) | ( \pi130 & w1618 ) | ( \pi131 & w1618 ) ;
  assign w1623 = ( ~w1620 & w1621 ) | ( ~w1620 & w1622 ) | ( w1621 & w1622 ) ;
  assign w1624 = ( w226 & w247 ) | ( w226 & ~w1339 ) | ( w247 & ~w1339 ) ;
  assign w1625 = ( \pi130 & \pi131 ) | ( \pi130 & w1624 ) | ( \pi131 & w1624 ) ;
  assign w1626 = w233 | w1625 ;
  assign w1627 = w254 & w1625 ;
  assign w1628 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1624 ) | ( \pi131 & ~w1624 ) ;
  assign w1629 = ( w1626 & w1627 ) | ( w1626 & ~w1628 ) | ( w1627 & ~w1628 ) ;
  assign w1630 = \pi132 ^ w1611 ;
  assign w1631 = ( w1611 & w1623 ) | ( w1611 & ~w1630 ) | ( w1623 & ~w1630 ) ;
  assign w1632 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1631 ) | ( ~\pi133 & w1631 ) ;
  assign w1633 = w1617 | w1632 ;
  assign w1634 = w1629 & w1632 ;
  assign w1635 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1631 ) | ( \pi133 & w1631 ) ;
  assign w1636 = ( w1633 & w1634 ) | ( w1633 & w1635 ) | ( w1634 & w1635 ) ;
  assign w1637 = ( w373 & w394 ) | ( w373 & ~w1353 ) | ( w394 & ~w1353 ) ;
  assign w1638 = ( \pi130 & \pi131 ) | ( \pi130 & w1637 ) | ( \pi131 & w1637 ) ;
  assign w1639 = w380 | w1638 ;
  assign w1640 = w401 & w1638 ;
  assign w1641 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1637 ) | ( \pi131 & ~w1637 ) ;
  assign w1642 = ( w1639 & w1640 ) | ( w1639 & ~w1641 ) | ( w1640 & ~w1641 ) ;
  assign w1643 = ( w156 & w359 ) | ( w156 & ~w1360 ) | ( w359 & ~w1360 ) ;
  assign w1644 = ( \pi130 & \pi131 ) | ( \pi130 & w1643 ) | ( \pi131 & w1643 ) ;
  assign w1645 = w163 | w1644 ;
  assign w1646 = w366 & w1644 ;
  assign w1647 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1643 ) | ( \pi131 & ~w1643 ) ;
  assign w1648 = ( w1645 & w1646 ) | ( w1645 & ~w1647 ) | ( w1646 & ~w1647 ) ;
  assign w1649 = ( w324 & w346 ) | ( w324 & w408 ) | ( w346 & w408 ) ;
  assign w1650 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1649 ) | ( \pi131 & ~w1649 ) ;
  assign w1651 = ~w331 & w1650 ;
  assign w1652 = w415 & ~w1650 ;
  assign w1653 = ( \pi130 & \pi131 ) | ( \pi130 & w1649 ) | ( \pi131 & w1649 ) ;
  assign w1654 = ( ~w1651 & w1652 ) | ( ~w1651 & w1653 ) | ( w1652 & w1653 ) ;
  assign w1655 = ( w289 & w311 ) | ( w289 & w338 ) | ( w311 & w338 ) ;
  assign w1656 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1655 ) | ( \pi131 & ~w1655 ) ;
  assign w1657 = ~w296 & w1656 ;
  assign w1658 = w345 & ~w1656 ;
  assign w1659 = ( \pi130 & \pi131 ) | ( \pi130 & w1655 ) | ( \pi131 & w1655 ) ;
  assign w1660 = ( ~w1657 & w1658 ) | ( ~w1657 & w1659 ) | ( w1658 & w1659 ) ;
  assign w1661 = \pi132 ^ w1642 ;
  assign w1662 = ( w1642 & w1654 ) | ( w1642 & ~w1661 ) | ( w1654 & ~w1661 ) ;
  assign w1663 = ( \pi132 & \pi133 ) | ( \pi132 & w1662 ) | ( \pi133 & w1662 ) ;
  assign w1664 = w1648 | w1663 ;
  assign w1665 = w1660 & w1663 ;
  assign w1666 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1662 ) | ( \pi133 & ~w1662 ) ;
  assign w1667 = ( w1664 & w1665 ) | ( w1664 & ~w1666 ) | ( w1665 & ~w1666 ) ;
  assign w1668 = \pi134 ^ w1667 ;
  assign w1669 = ( w1636 & w1667 ) | ( w1636 & ~w1668 ) | ( w1667 & ~w1668 ) ;
  assign w1670 = ( w438 & w460 ) | ( w438 & w487 ) | ( w460 & w487 ) ;
  assign w1671 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1670 ) | ( \pi131 & ~w1670 ) ;
  assign w1672 = ~w445 & w1671 ;
  assign w1673 = w494 & ~w1671 ;
  assign w1674 = ( \pi130 & \pi131 ) | ( \pi130 & w1670 ) | ( \pi131 & w1670 ) ;
  assign w1675 = ( ~w1672 & w1673 ) | ( ~w1672 & w1674 ) | ( w1673 & w1674 ) ;
  assign w1676 = ( w473 & w495 ) | ( w473 & w557 ) | ( w495 & w557 ) ;
  assign w1677 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1676 ) | ( \pi131 & ~w1676 ) ;
  assign w1678 = ~w480 & w1677 ;
  assign w1679 = w564 & ~w1677 ;
  assign w1680 = ( \pi130 & \pi131 ) | ( \pi130 & w1676 ) | ( \pi131 & w1676 ) ;
  assign w1681 = ( ~w1678 & w1679 ) | ( ~w1678 & w1680 ) | ( w1679 & w1680 ) ;
  assign w1682 = ( w508 & w530 ) | ( w508 & w634 ) | ( w530 & w634 ) ;
  assign w1683 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1682 ) | ( \pi131 & ~w1682 ) ;
  assign w1684 = ~w515 & w1683 ;
  assign w1685 = w641 & ~w1683 ;
  assign w1686 = ( \pi130 & \pi131 ) | ( \pi130 & w1682 ) | ( \pi131 & w1682 ) ;
  assign w1687 = ( ~w1684 & w1685 ) | ( ~w1684 & w1686 ) | ( w1685 & w1686 ) ;
  assign w1688 = ( w522 & w543 ) | ( w522 & ~w1411 ) | ( w543 & ~w1411 ) ;
  assign w1689 = ( \pi130 & \pi131 ) | ( \pi130 & w1688 ) | ( \pi131 & w1688 ) ;
  assign w1690 = w529 | w1689 ;
  assign w1691 = w550 & w1689 ;
  assign w1692 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1688 ) | ( \pi131 & ~w1688 ) ;
  assign w1693 = ( w1690 & w1691 ) | ( w1690 & ~w1692 ) | ( w1691 & ~w1692 ) ;
  assign w1694 = \pi132 ^ w1675 ;
  assign w1695 = ( w1675 & w1687 ) | ( w1675 & ~w1694 ) | ( w1687 & ~w1694 ) ;
  assign w1696 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1695 ) | ( ~\pi133 & w1695 ) ;
  assign w1697 = w1681 | w1696 ;
  assign w1698 = w1693 & w1696 ;
  assign w1699 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1695 ) | ( \pi133 & w1695 ) ;
  assign w1700 = ( w1697 & w1698 ) | ( w1697 & w1699 ) | ( w1698 & w1699 ) ;
  assign w1701 = ( w599 & w655 ) | ( w599 & ~w1425 ) | ( w655 & ~w1425 ) ;
  assign w1702 = ( \pi130 & \pi131 ) | ( \pi130 & w1701 ) | ( \pi131 & w1701 ) ;
  assign w1703 = w606 | w1702 ;
  assign w1704 = w662 & w1702 ;
  assign w1705 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1701 ) | ( \pi131 & ~w1701 ) ;
  assign w1706 = ( w1703 & w1704 ) | ( w1703 & ~w1705 ) | ( w1704 & ~w1705 ) ;
  assign w1707 = ( w452 & w585 ) | ( w452 & ~w1432 ) | ( w585 & ~w1432 ) ;
  assign w1708 = ( \pi130 & \pi131 ) | ( \pi130 & w1707 ) | ( \pi131 & w1707 ) ;
  assign w1709 = w459 | w1708 ;
  assign w1710 = w592 & w1708 ;
  assign w1711 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1707 ) | ( \pi131 & ~w1707 ) ;
  assign w1712 = ( w1709 & w1710 ) | ( w1709 & ~w1711 ) | ( w1710 & ~w1711 ) ;
  assign w1713 = ( w669 & w690 ) | ( w669 & ~w1439 ) | ( w690 & ~w1439 ) ;
  assign w1714 = ( \pi130 & \pi131 ) | ( \pi130 & w1713 ) | ( \pi131 & w1713 ) ;
  assign w1715 = w676 | w1714 ;
  assign w1716 = w697 & w1714 ;
  assign w1717 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1713 ) | ( \pi131 & ~w1713 ) ;
  assign w1718 = ( w1715 & w1716 ) | ( w1715 & ~w1717 ) | ( w1716 & ~w1717 ) ;
  assign w1719 = ( w620 & w642 ) | ( w620 & w704 ) | ( w642 & w704 ) ;
  assign w1720 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1719 ) | ( \pi131 & ~w1719 ) ;
  assign w1721 = ~w627 & w1720 ;
  assign w1722 = w711 & ~w1720 ;
  assign w1723 = ( \pi130 & \pi131 ) | ( \pi130 & w1719 ) | ( \pi131 & w1719 ) ;
  assign w1724 = ( ~w1721 & w1722 ) | ( ~w1721 & w1723 ) | ( w1722 & w1723 ) ;
  assign w1725 = \pi132 ^ w1706 ;
  assign w1726 = ( w1706 & w1718 ) | ( w1706 & ~w1725 ) | ( w1718 & ~w1725 ) ;
  assign w1727 = ( \pi132 & \pi133 ) | ( \pi132 & w1726 ) | ( \pi133 & w1726 ) ;
  assign w1728 = w1712 | w1727 ;
  assign w1729 = w1724 & w1727 ;
  assign w1730 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1726 ) | ( \pi133 & ~w1726 ) ;
  assign w1731 = ( w1728 & w1729 ) | ( w1728 & ~w1730 ) | ( w1729 & ~w1730 ) ;
  assign w1732 = \pi134 ^ w1731 ;
  assign w1733 = ( w1700 & w1731 ) | ( w1700 & ~w1732 ) | ( w1731 & ~w1732 ) ;
  assign w1734 = ( w734 & w756 ) | ( w734 & w783 ) | ( w756 & w783 ) ;
  assign w1735 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1734 ) | ( \pi131 & ~w1734 ) ;
  assign w1736 = ~w741 & w1735 ;
  assign w1737 = w790 & ~w1735 ;
  assign w1738 = ( \pi130 & \pi131 ) | ( \pi130 & w1734 ) | ( \pi131 & w1734 ) ;
  assign w1739 = ( ~w1736 & w1737 ) | ( ~w1736 & w1738 ) | ( w1737 & w1738 ) ;
  assign w1740 = ( w769 & w791 ) | ( w769 & w852 ) | ( w791 & w852 ) ;
  assign w1741 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1740 ) | ( \pi131 & ~w1740 ) ;
  assign w1742 = ~w776 & w1741 ;
  assign w1743 = w859 & ~w1741 ;
  assign w1744 = ( \pi130 & \pi131 ) | ( \pi130 & w1740 ) | ( \pi131 & w1740 ) ;
  assign w1745 = ( ~w1742 & w1743 ) | ( ~w1742 & w1744 ) | ( w1743 & w1744 ) ;
  assign w1746 = ( w803 & w825 ) | ( w803 & w929 ) | ( w825 & w929 ) ;
  assign w1747 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1746 ) | ( \pi131 & ~w1746 ) ;
  assign w1748 = ~w810 & w1747 ;
  assign w1749 = w936 & ~w1747 ;
  assign w1750 = ( \pi130 & \pi131 ) | ( \pi130 & w1746 ) | ( \pi131 & w1746 ) ;
  assign w1751 = ( ~w1748 & w1749 ) | ( ~w1748 & w1750 ) | ( w1749 & w1750 ) ;
  assign w1752 = ( w817 & w838 ) | ( w817 & ~w1483 ) | ( w838 & ~w1483 ) ;
  assign w1753 = ( \pi130 & \pi131 ) | ( \pi130 & w1752 ) | ( \pi131 & w1752 ) ;
  assign w1754 = w824 | w1753 ;
  assign w1755 = w845 & w1753 ;
  assign w1756 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1752 ) | ( \pi131 & ~w1752 ) ;
  assign w1757 = ( w1754 & w1755 ) | ( w1754 & ~w1756 ) | ( w1755 & ~w1756 ) ;
  assign w1758 = \pi132 ^ w1739 ;
  assign w1759 = ( w1739 & w1751 ) | ( w1739 & ~w1758 ) | ( w1751 & ~w1758 ) ;
  assign w1760 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1759 ) | ( ~\pi133 & w1759 ) ;
  assign w1761 = w1745 | w1760 ;
  assign w1762 = w1757 & w1760 ;
  assign w1763 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1759 ) | ( \pi133 & w1759 ) ;
  assign w1764 = ( w1761 & w1762 ) | ( w1761 & w1763 ) | ( w1762 & w1763 ) ;
  assign w1765 = ( w894 & w950 ) | ( w894 & ~w1497 ) | ( w950 & ~w1497 ) ;
  assign w1766 = ( \pi130 & \pi131 ) | ( \pi130 & w1765 ) | ( \pi131 & w1765 ) ;
  assign w1767 = w901 | w1766 ;
  assign w1768 = w957 & w1766 ;
  assign w1769 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1765 ) | ( \pi131 & ~w1765 ) ;
  assign w1770 = ( w1767 & w1768 ) | ( w1767 & ~w1769 ) | ( w1768 & ~w1769 ) ;
  assign w1771 = ( w748 & w880 ) | ( w748 & ~w1504 ) | ( w880 & ~w1504 ) ;
  assign w1772 = ( \pi130 & \pi131 ) | ( \pi130 & w1771 ) | ( \pi131 & w1771 ) ;
  assign w1773 = w755 | w1772 ;
  assign w1774 = w887 & w1772 ;
  assign w1775 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1771 ) | ( \pi131 & ~w1771 ) ;
  assign w1776 = ( w1773 & w1774 ) | ( w1773 & ~w1775 ) | ( w1774 & ~w1775 ) ;
  assign w1777 = ( w964 & w985 ) | ( w964 & ~w1511 ) | ( w985 & ~w1511 ) ;
  assign w1778 = ( \pi130 & \pi131 ) | ( \pi130 & w1777 ) | ( \pi131 & w1777 ) ;
  assign w1779 = w971 | w1778 ;
  assign w1780 = w992 & w1778 ;
  assign w1781 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1777 ) | ( \pi131 & ~w1777 ) ;
  assign w1782 = ( w1779 & w1780 ) | ( w1779 & ~w1781 ) | ( w1780 & ~w1781 ) ;
  assign w1783 = ( w915 & w937 ) | ( w915 & w999 ) | ( w937 & w999 ) ;
  assign w1784 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1783 ) | ( \pi131 & ~w1783 ) ;
  assign w1785 = ~w922 & w1784 ;
  assign w1786 = w1006 & ~w1784 ;
  assign w1787 = ( \pi130 & \pi131 ) | ( \pi130 & w1783 ) | ( \pi131 & w1783 ) ;
  assign w1788 = ( ~w1785 & w1786 ) | ( ~w1785 & w1787 ) | ( w1786 & w1787 ) ;
  assign w1789 = \pi132 ^ w1770 ;
  assign w1790 = ( w1770 & w1782 ) | ( w1770 & ~w1789 ) | ( w1782 & ~w1789 ) ;
  assign w1791 = ( \pi132 & \pi133 ) | ( \pi132 & w1790 ) | ( \pi133 & w1790 ) ;
  assign w1792 = w1776 | w1791 ;
  assign w1793 = w1788 & w1791 ;
  assign w1794 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1790 ) | ( \pi133 & ~w1790 ) ;
  assign w1795 = ( w1792 & w1793 ) | ( w1792 & ~w1794 ) | ( w1793 & ~w1794 ) ;
  assign w1796 = \pi134 ^ w1795 ;
  assign w1797 = ( w1764 & w1795 ) | ( w1764 & ~w1796 ) | ( w1795 & ~w1796 ) ;
  assign w1798 = ( w1078 & w1133 ) | ( w1078 & ~w1534 ) | ( w1133 & ~w1534 ) ;
  assign w1799 = ( \pi130 & \pi131 ) | ( \pi130 & w1798 ) | ( \pi131 & w1798 ) ;
  assign w1800 = w1085 | w1799 ;
  assign w1801 = w1140 & w1799 ;
  assign w1802 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1798 ) | ( \pi131 & ~w1798 ) ;
  assign w1803 = ( w1800 & w1801 ) | ( w1800 & ~w1802 ) | ( w1801 & ~w1802 ) ;
  assign w1804 = ( w1043 & w1064 ) | ( w1043 & ~w1541 ) | ( w1064 & ~w1541 ) ;
  assign w1805 = ( \pi130 & \pi131 ) | ( \pi130 & w1804 ) | ( \pi131 & w1804 ) ;
  assign w1806 = w1050 | w1805 ;
  assign w1807 = w1071 & w1805 ;
  assign w1808 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1804 ) | ( \pi131 & ~w1804 ) ;
  assign w1809 = ( w1806 & w1807 ) | ( w1806 & ~w1808 ) | ( w1807 & ~w1808 ) ;
  assign w1810 = ( w1098 & w1120 ) | ( w1098 & w1259 ) | ( w1120 & w1259 ) ;
  assign w1811 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1810 ) | ( \pi131 & ~w1810 ) ;
  assign w1812 = ~w1105 & w1811 ;
  assign w1813 = w1266 & ~w1811 ;
  assign w1814 = ( \pi130 & \pi131 ) | ( \pi130 & w1810 ) | ( \pi131 & w1810 ) ;
  assign w1815 = ( ~w1812 & w1813 ) | ( ~w1812 & w1814 ) | ( w1813 & w1814 ) ;
  assign w1816 = ( w1029 & w1051 ) | ( w1029 & w1112 ) | ( w1051 & w1112 ) ;
  assign w1817 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1816 ) | ( \pi131 & ~w1816 ) ;
  assign w1818 = ~w1036 & w1817 ;
  assign w1819 = w1119 & ~w1817 ;
  assign w1820 = ( \pi130 & \pi131 ) | ( \pi130 & w1816 ) | ( \pi131 & w1816 ) ;
  assign w1821 = ( ~w1818 & w1819 ) | ( ~w1818 & w1820 ) | ( w1819 & w1820 ) ;
  assign w1822 = \pi132 ^ w1803 ;
  assign w1823 = ( w1803 & w1815 ) | ( w1803 & ~w1822 ) | ( w1815 & ~w1822 ) ;
  assign w1824 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1823 ) | ( ~\pi133 & w1823 ) ;
  assign w1825 = w1809 | w1824 ;
  assign w1826 = w1821 & w1824 ;
  assign w1827 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1823 ) | ( \pi133 & w1823 ) ;
  assign w1828 = ( w1825 & w1826 ) | ( w1825 & w1827 ) | ( w1826 & w1827 ) ;
  assign w1829 = ( w1189 & w1210 ) | ( w1189 & ~w1569 ) | ( w1210 & ~w1569 ) ;
  assign w1830 = ( \pi130 & \pi131 ) | ( \pi130 & w1829 ) | ( \pi131 & w1829 ) ;
  assign w1831 = w1196 | w1830 ;
  assign w1832 = w1217 & w1830 ;
  assign w1833 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1829 ) | ( \pi131 & ~w1829 ) ;
  assign w1834 = ( w1831 & w1832 ) | ( w1831 & ~w1833 ) | ( w1832 & ~w1833 ) ;
  assign w1835 = ( w1147 & w1175 ) | ( w1147 & ~w1576 ) | ( w1175 & ~w1576 ) ;
  assign w1836 = ( \pi130 & \pi131 ) | ( \pi130 & w1835 ) | ( \pi131 & w1835 ) ;
  assign w1837 = w1154 | w1836 ;
  assign w1838 = w1182 & w1836 ;
  assign w1839 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1835 ) | ( \pi131 & ~w1835 ) ;
  assign w1840 = ( w1837 & w1838 ) | ( w1837 & ~w1839 ) | ( w1838 & ~w1839 ) ;
  assign w1841 = ( w1224 & w1280 ) | ( w1224 & ~w1583 ) | ( w1280 & ~w1583 ) ;
  assign w1842 = ( \pi130 & \pi131 ) | ( \pi130 & w1841 ) | ( \pi131 & w1841 ) ;
  assign w1843 = w1231 | w1842 ;
  assign w1844 = w1287 & w1842 ;
  assign w1845 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1841 ) | ( \pi131 & ~w1841 ) ;
  assign w1846 = ( w1843 & w1844 ) | ( w1843 & ~w1845 ) | ( w1844 & ~w1845 ) ;
  assign w1847 = ( w1245 & w1267 ) | ( w1245 & w1294 ) | ( w1267 & w1294 ) ;
  assign w1848 = ( \pi130 & \pi131 ) | ( \pi130 & ~w1847 ) | ( \pi131 & ~w1847 ) ;
  assign w1849 = ~w1252 & w1848 ;
  assign w1850 = w1301 & ~w1848 ;
  assign w1851 = ( \pi130 & \pi131 ) | ( \pi130 & w1847 ) | ( \pi131 & w1847 ) ;
  assign w1852 = ( ~w1849 & w1850 ) | ( ~w1849 & w1851 ) | ( w1850 & w1851 ) ;
  assign w1853 = \pi132 ^ w1834 ;
  assign w1854 = ( w1834 & w1846 ) | ( w1834 & ~w1853 ) | ( w1846 & ~w1853 ) ;
  assign w1855 = ( \pi132 & \pi133 ) | ( \pi132 & w1854 ) | ( \pi133 & w1854 ) ;
  assign w1856 = w1840 | w1855 ;
  assign w1857 = w1852 & w1855 ;
  assign w1858 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1854 ) | ( \pi133 & ~w1854 ) ;
  assign w1859 = ( w1856 & w1857 ) | ( w1856 & ~w1858 ) | ( w1857 & ~w1858 ) ;
  assign w1860 = \pi134 ^ w1859 ;
  assign w1861 = ( w1828 & w1859 ) | ( w1828 & ~w1860 ) | ( w1859 & ~w1860 ) ;
  assign w1862 = ( w142 & ~w164 ) | ( w142 & w184 ) | ( ~w164 & w184 ) ;
  assign w1863 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1862 ) | ( ~\pi131 & w1862 ) ;
  assign w1864 = w191 | w1863 ;
  assign w1865 = w198 & w1863 ;
  assign w1866 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1862 ) | ( \pi131 & w1862 ) ;
  assign w1867 = ( w1864 & w1865 ) | ( w1864 & w1866 ) | ( w1865 & w1866 ) ;
  assign w1868 = ( w177 & ~w199 ) | ( w177 & w254 ) | ( ~w199 & w254 ) ;
  assign w1869 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1868 ) | ( ~\pi131 & w1868 ) ;
  assign w1870 = w261 | w1869 ;
  assign w1871 = w268 & w1869 ;
  assign w1872 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1868 ) | ( \pi131 & w1868 ) ;
  assign w1873 = ( w1870 & w1871 ) | ( w1870 & w1872 ) | ( w1871 & w1872 ) ;
  assign w1874 = ( w212 & ~w234 ) | ( w212 & w296 ) | ( ~w234 & w296 ) ;
  assign w1875 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1874 ) | ( ~\pi131 & w1874 ) ;
  assign w1876 = w303 | w1875 ;
  assign w1877 = w310 & w1875 ;
  assign w1878 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1874 ) | ( \pi131 & w1874 ) ;
  assign w1879 = ( w1876 & w1877 ) | ( w1876 & w1878 ) | ( w1877 & w1878 ) ;
  assign w1880 = \pi131 ^ w219 ;
  assign w1881 = ( w219 & w247 ) | ( w219 & w1880 ) | ( w247 & w1880 ) ;
  assign w1882 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1881 ) | ( ~\pi131 & w1881 ) ;
  assign w1883 = w226 | w1882 ;
  assign w1884 = w233 & w1882 ;
  assign w1885 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1881 ) | ( \pi131 & w1881 ) ;
  assign w1886 = ( w1883 & w1884 ) | ( w1883 & w1885 ) | ( w1884 & w1885 ) ;
  assign w1887 = \pi132 ^ w1867 ;
  assign w1888 = ( w1867 & w1879 ) | ( w1867 & ~w1887 ) | ( w1879 & ~w1887 ) ;
  assign w1889 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1888 ) | ( ~\pi133 & w1888 ) ;
  assign w1890 = w1873 | w1889 ;
  assign w1891 = w1886 & w1889 ;
  assign w1892 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1888 ) | ( \pi133 & w1888 ) ;
  assign w1893 = ( w1890 & w1891 ) | ( w1890 & w1892 ) | ( w1891 & w1892 ) ;
  assign w1894 = \pi131 ^ w366 ;
  assign w1895 = ( w366 & w394 ) | ( w366 & w1894 ) | ( w394 & w1894 ) ;
  assign w1896 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1895 ) | ( ~\pi131 & w1895 ) ;
  assign w1897 = w373 | w1896 ;
  assign w1898 = w380 & w1896 ;
  assign w1899 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1895 ) | ( \pi131 & w1895 ) ;
  assign w1900 = ( w1897 & w1898 ) | ( w1897 & w1899 ) | ( w1898 & w1899 ) ;
  assign w1901 = \pi131 ^ w149 ;
  assign w1902 = ( w149 & w359 ) | ( w149 & w1901 ) | ( w359 & w1901 ) ;
  assign w1903 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1902 ) | ( ~\pi131 & w1902 ) ;
  assign w1904 = w156 | w1903 ;
  assign w1905 = w163 & w1903 ;
  assign w1906 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1902 ) | ( \pi131 & w1902 ) ;
  assign w1907 = ( w1904 & w1905 ) | ( w1904 & w1906 ) | ( w1905 & w1906 ) ;
  assign w1908 = ( w324 & ~w346 ) | ( w324 & w401 ) | ( ~w346 & w401 ) ;
  assign w1909 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1908 ) | ( ~\pi131 & w1908 ) ;
  assign w1910 = w408 | w1909 ;
  assign w1911 = w415 & w1909 ;
  assign w1912 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1908 ) | ( \pi131 & w1908 ) ;
  assign w1913 = ( w1910 & w1911 ) | ( w1910 & w1912 ) | ( w1911 & w1912 ) ;
  assign w1914 = ( w289 & ~w311 ) | ( w289 & w331 ) | ( ~w311 & w331 ) ;
  assign w1915 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1914 ) | ( ~\pi131 & w1914 ) ;
  assign w1916 = w338 | w1915 ;
  assign w1917 = w345 & w1915 ;
  assign w1918 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1914 ) | ( \pi131 & w1914 ) ;
  assign w1919 = ( w1916 & w1917 ) | ( w1916 & w1918 ) | ( w1917 & w1918 ) ;
  assign w1920 = \pi132 ^ w1900 ;
  assign w1921 = ( w1900 & w1913 ) | ( w1900 & ~w1920 ) | ( w1913 & ~w1920 ) ;
  assign w1922 = ( \pi132 & \pi133 ) | ( \pi132 & w1921 ) | ( \pi133 & w1921 ) ;
  assign w1923 = w1907 | w1922 ;
  assign w1924 = w1919 & w1922 ;
  assign w1925 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1921 ) | ( \pi133 & ~w1921 ) ;
  assign w1926 = ( w1923 & w1924 ) | ( w1923 & ~w1925 ) | ( w1924 & ~w1925 ) ;
  assign w1927 = \pi134 ^ w1926 ;
  assign w1928 = ( w1893 & w1926 ) | ( w1893 & ~w1927 ) | ( w1926 & ~w1927 ) ;
  assign w1929 = ( w438 & ~w460 ) | ( w438 & w480 ) | ( ~w460 & w480 ) ;
  assign w1930 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1929 ) | ( ~\pi131 & w1929 ) ;
  assign w1931 = w487 | w1930 ;
  assign w1932 = w494 & w1930 ;
  assign w1933 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1929 ) | ( \pi131 & w1929 ) ;
  assign w1934 = ( w1931 & w1932 ) | ( w1931 & w1933 ) | ( w1932 & w1933 ) ;
  assign w1935 = ( w473 & ~w495 ) | ( w473 & w550 ) | ( ~w495 & w550 ) ;
  assign w1936 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1935 ) | ( ~\pi131 & w1935 ) ;
  assign w1937 = w557 | w1936 ;
  assign w1938 = w564 & w1936 ;
  assign w1939 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1935 ) | ( \pi131 & w1935 ) ;
  assign w1940 = ( w1937 & w1938 ) | ( w1937 & w1939 ) | ( w1938 & w1939 ) ;
  assign w1941 = ( w508 & ~w530 ) | ( w508 & w627 ) | ( ~w530 & w627 ) ;
  assign w1942 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1941 ) | ( ~\pi131 & w1941 ) ;
  assign w1943 = w634 | w1942 ;
  assign w1944 = w641 & w1942 ;
  assign w1945 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1941 ) | ( \pi131 & w1941 ) ;
  assign w1946 = ( w1943 & w1944 ) | ( w1943 & w1945 ) | ( w1944 & w1945 ) ;
  assign w1947 = \pi131 ^ w515 ;
  assign w1948 = ( w515 & w543 ) | ( w515 & w1947 ) | ( w543 & w1947 ) ;
  assign w1949 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1948 ) | ( ~\pi131 & w1948 ) ;
  assign w1950 = w522 | w1949 ;
  assign w1951 = w529 & w1949 ;
  assign w1952 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1948 ) | ( \pi131 & w1948 ) ;
  assign w1953 = ( w1950 & w1951 ) | ( w1950 & w1952 ) | ( w1951 & w1952 ) ;
  assign w1954 = \pi132 ^ w1934 ;
  assign w1955 = ( w1934 & w1946 ) | ( w1934 & ~w1954 ) | ( w1946 & ~w1954 ) ;
  assign w1956 = ( \pi132 & ~\pi133 ) | ( \pi132 & w1955 ) | ( ~\pi133 & w1955 ) ;
  assign w1957 = w1940 | w1956 ;
  assign w1958 = w1953 & w1956 ;
  assign w1959 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w1955 ) | ( \pi133 & w1955 ) ;
  assign w1960 = ( w1957 & w1958 ) | ( w1957 & w1959 ) | ( w1958 & w1959 ) ;
  assign w1961 = \pi131 ^ w592 ;
  assign w1962 = ( w592 & w655 ) | ( w592 & w1961 ) | ( w655 & w1961 ) ;
  assign w1963 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1962 ) | ( ~\pi131 & w1962 ) ;
  assign w1964 = w599 | w1963 ;
  assign w1965 = w606 & w1963 ;
  assign w1966 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1962 ) | ( \pi131 & w1962 ) ;
  assign w1967 = ( w1964 & w1965 ) | ( w1964 & w1966 ) | ( w1965 & w1966 ) ;
  assign w1968 = \pi131 ^ w445 ;
  assign w1969 = ( w445 & w585 ) | ( w445 & w1968 ) | ( w585 & w1968 ) ;
  assign w1970 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1969 ) | ( ~\pi131 & w1969 ) ;
  assign w1971 = w452 | w1970 ;
  assign w1972 = w459 & w1970 ;
  assign w1973 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1969 ) | ( \pi131 & w1969 ) ;
  assign w1974 = ( w1971 & w1972 ) | ( w1971 & w1973 ) | ( w1972 & w1973 ) ;
  assign w1975 = \pi131 ^ w662 ;
  assign w1976 = ( w662 & w690 ) | ( w662 & w1975 ) | ( w690 & w1975 ) ;
  assign w1977 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1976 ) | ( ~\pi131 & w1976 ) ;
  assign w1978 = w669 | w1977 ;
  assign w1979 = w676 & w1977 ;
  assign w1980 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1976 ) | ( \pi131 & w1976 ) ;
  assign w1981 = ( w1978 & w1979 ) | ( w1978 & w1980 ) | ( w1979 & w1980 ) ;
  assign w1982 = ( w620 & ~w642 ) | ( w620 & w697 ) | ( ~w642 & w697 ) ;
  assign w1983 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1982 ) | ( ~\pi131 & w1982 ) ;
  assign w1984 = w704 | w1983 ;
  assign w1985 = w711 & w1983 ;
  assign w1986 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1982 ) | ( \pi131 & w1982 ) ;
  assign w1987 = ( w1984 & w1985 ) | ( w1984 & w1986 ) | ( w1985 & w1986 ) ;
  assign w1988 = \pi132 ^ w1967 ;
  assign w1989 = ( w1967 & w1981 ) | ( w1967 & ~w1988 ) | ( w1981 & ~w1988 ) ;
  assign w1990 = ( \pi132 & \pi133 ) | ( \pi132 & w1989 ) | ( \pi133 & w1989 ) ;
  assign w1991 = w1974 | w1990 ;
  assign w1992 = w1987 & w1990 ;
  assign w1993 = ( \pi132 & \pi133 ) | ( \pi132 & ~w1989 ) | ( \pi133 & ~w1989 ) ;
  assign w1994 = ( w1991 & w1992 ) | ( w1991 & ~w1993 ) | ( w1992 & ~w1993 ) ;
  assign w1995 = \pi134 ^ w1994 ;
  assign w1996 = ( w1960 & w1994 ) | ( w1960 & ~w1995 ) | ( w1994 & ~w1995 ) ;
  assign w1997 = ( w734 & ~w756 ) | ( w734 & w776 ) | ( ~w756 & w776 ) ;
  assign w1998 = ( \pi130 & ~\pi131 ) | ( \pi130 & w1997 ) | ( ~\pi131 & w1997 ) ;
  assign w1999 = w783 | w1998 ;
  assign w2000 = w790 & w1998 ;
  assign w2001 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w1997 ) | ( \pi131 & w1997 ) ;
  assign w2002 = ( w1999 & w2000 ) | ( w1999 & w2001 ) | ( w2000 & w2001 ) ;
  assign w2003 = ( w769 & ~w791 ) | ( w769 & w845 ) | ( ~w791 & w845 ) ;
  assign w2004 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2003 ) | ( ~\pi131 & w2003 ) ;
  assign w2005 = w852 | w2004 ;
  assign w2006 = w859 & w2004 ;
  assign w2007 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2003 ) | ( \pi131 & w2003 ) ;
  assign w2008 = ( w2005 & w2006 ) | ( w2005 & w2007 ) | ( w2006 & w2007 ) ;
  assign w2009 = ( w803 & ~w825 ) | ( w803 & w922 ) | ( ~w825 & w922 ) ;
  assign w2010 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2009 ) | ( ~\pi131 & w2009 ) ;
  assign w2011 = w929 | w2010 ;
  assign w2012 = w936 & w2010 ;
  assign w2013 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2009 ) | ( \pi131 & w2009 ) ;
  assign w2014 = ( w2011 & w2012 ) | ( w2011 & w2013 ) | ( w2012 & w2013 ) ;
  assign w2015 = \pi131 ^ w810 ;
  assign w2016 = ( w810 & w838 ) | ( w810 & w2015 ) | ( w838 & w2015 ) ;
  assign w2017 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2016 ) | ( ~\pi131 & w2016 ) ;
  assign w2018 = w817 | w2017 ;
  assign w2019 = w824 & w2017 ;
  assign w2020 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2016 ) | ( \pi131 & w2016 ) ;
  assign w2021 = ( w2018 & w2019 ) | ( w2018 & w2020 ) | ( w2019 & w2020 ) ;
  assign w2022 = \pi132 ^ w2002 ;
  assign w2023 = ( w2002 & w2014 ) | ( w2002 & ~w2022 ) | ( w2014 & ~w2022 ) ;
  assign w2024 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2023 ) | ( ~\pi133 & w2023 ) ;
  assign w2025 = w2008 | w2024 ;
  assign w2026 = w2021 & w2024 ;
  assign w2027 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2023 ) | ( \pi133 & w2023 ) ;
  assign w2028 = ( w2025 & w2026 ) | ( w2025 & w2027 ) | ( w2026 & w2027 ) ;
  assign w2029 = \pi131 ^ w887 ;
  assign w2030 = ( w887 & w950 ) | ( w887 & w2029 ) | ( w950 & w2029 ) ;
  assign w2031 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2030 ) | ( ~\pi131 & w2030 ) ;
  assign w2032 = w894 | w2031 ;
  assign w2033 = w901 & w2031 ;
  assign w2034 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2030 ) | ( \pi131 & w2030 ) ;
  assign w2035 = ( w2032 & w2033 ) | ( w2032 & w2034 ) | ( w2033 & w2034 ) ;
  assign w2036 = \pi131 ^ w741 ;
  assign w2037 = ( w741 & w880 ) | ( w741 & w2036 ) | ( w880 & w2036 ) ;
  assign w2038 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2037 ) | ( ~\pi131 & w2037 ) ;
  assign w2039 = w748 | w2038 ;
  assign w2040 = w755 & w2038 ;
  assign w2041 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2037 ) | ( \pi131 & w2037 ) ;
  assign w2042 = ( w2039 & w2040 ) | ( w2039 & w2041 ) | ( w2040 & w2041 ) ;
  assign w2043 = \pi131 ^ w957 ;
  assign w2044 = ( w957 & w985 ) | ( w957 & w2043 ) | ( w985 & w2043 ) ;
  assign w2045 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2044 ) | ( ~\pi131 & w2044 ) ;
  assign w2046 = w964 | w2045 ;
  assign w2047 = w971 & w2045 ;
  assign w2048 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2044 ) | ( \pi131 & w2044 ) ;
  assign w2049 = ( w2046 & w2047 ) | ( w2046 & w2048 ) | ( w2047 & w2048 ) ;
  assign w2050 = ( w915 & ~w937 ) | ( w915 & w992 ) | ( ~w937 & w992 ) ;
  assign w2051 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2050 ) | ( ~\pi131 & w2050 ) ;
  assign w2052 = w999 | w2051 ;
  assign w2053 = w1006 & w2051 ;
  assign w2054 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2050 ) | ( \pi131 & w2050 ) ;
  assign w2055 = ( w2052 & w2053 ) | ( w2052 & w2054 ) | ( w2053 & w2054 ) ;
  assign w2056 = \pi132 ^ w2035 ;
  assign w2057 = ( w2035 & w2049 ) | ( w2035 & ~w2056 ) | ( w2049 & ~w2056 ) ;
  assign w2058 = ( \pi132 & \pi133 ) | ( \pi132 & w2057 ) | ( \pi133 & w2057 ) ;
  assign w2059 = w2042 | w2058 ;
  assign w2060 = w2055 & w2058 ;
  assign w2061 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2057 ) | ( \pi133 & ~w2057 ) ;
  assign w2062 = ( w2059 & w2060 ) | ( w2059 & ~w2061 ) | ( w2060 & ~w2061 ) ;
  assign w2063 = \pi134 ^ w2062 ;
  assign w2064 = ( w2028 & w2062 ) | ( w2028 & ~w2063 ) | ( w2062 & ~w2063 ) ;
  assign w2065 = \pi131 ^ w1071 ;
  assign w2066 = ( w1071 & w1133 ) | ( w1071 & w2065 ) | ( w1133 & w2065 ) ;
  assign w2067 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2066 ) | ( ~\pi131 & w2066 ) ;
  assign w2068 = w1078 | w2067 ;
  assign w2069 = w1085 & w2067 ;
  assign w2070 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2066 ) | ( \pi131 & w2066 ) ;
  assign w2071 = ( w2068 & w2069 ) | ( w2068 & w2070 ) | ( w2069 & w2070 ) ;
  assign w2072 = \pi131 ^ w1036 ;
  assign w2073 = ( w1036 & w1064 ) | ( w1036 & w2072 ) | ( w1064 & w2072 ) ;
  assign w2074 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2073 ) | ( ~\pi131 & w2073 ) ;
  assign w2075 = w1043 | w2074 ;
  assign w2076 = w1050 & w2074 ;
  assign w2077 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2073 ) | ( \pi131 & w2073 ) ;
  assign w2078 = ( w2075 & w2076 ) | ( w2075 & w2077 ) | ( w2076 & w2077 ) ;
  assign w2079 = ( w1098 & ~w1120 ) | ( w1098 & w1252 ) | ( ~w1120 & w1252 ) ;
  assign w2080 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2079 ) | ( ~\pi131 & w2079 ) ;
  assign w2081 = w1259 | w2080 ;
  assign w2082 = w1266 & w2080 ;
  assign w2083 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2079 ) | ( \pi131 & w2079 ) ;
  assign w2084 = ( w2081 & w2082 ) | ( w2081 & w2083 ) | ( w2082 & w2083 ) ;
  assign w2085 = ( w1029 & ~w1051 ) | ( w1029 & w1105 ) | ( ~w1051 & w1105 ) ;
  assign w2086 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2085 ) | ( ~\pi131 & w2085 ) ;
  assign w2087 = w1112 | w2086 ;
  assign w2088 = w1119 & w2086 ;
  assign w2089 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2085 ) | ( \pi131 & w2085 ) ;
  assign w2090 = ( w2087 & w2088 ) | ( w2087 & w2089 ) | ( w2088 & w2089 ) ;
  assign w2091 = \pi132 ^ w2071 ;
  assign w2092 = ( w2071 & w2084 ) | ( w2071 & ~w2091 ) | ( w2084 & ~w2091 ) ;
  assign w2093 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2092 ) | ( ~\pi133 & w2092 ) ;
  assign w2094 = w2078 | w2093 ;
  assign w2095 = w2090 & w2093 ;
  assign w2096 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2092 ) | ( \pi133 & w2092 ) ;
  assign w2097 = ( w2094 & w2095 ) | ( w2094 & w2096 ) | ( w2095 & w2096 ) ;
  assign w2098 = \pi131 ^ w1182 ;
  assign w2099 = ( w1182 & w1210 ) | ( w1182 & w2098 ) | ( w1210 & w2098 ) ;
  assign w2100 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2099 ) | ( ~\pi131 & w2099 ) ;
  assign w2101 = w1189 | w2100 ;
  assign w2102 = w1196 & w2100 ;
  assign w2103 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2099 ) | ( \pi131 & w2099 ) ;
  assign w2104 = ( w2101 & w2102 ) | ( w2101 & w2103 ) | ( w2102 & w2103 ) ;
  assign w2105 = \pi131 ^ w1140 ;
  assign w2106 = ( w1140 & w1175 ) | ( w1140 & w2105 ) | ( w1175 & w2105 ) ;
  assign w2107 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2106 ) | ( ~\pi131 & w2106 ) ;
  assign w2108 = w1147 | w2107 ;
  assign w2109 = w1154 & w2107 ;
  assign w2110 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2106 ) | ( \pi131 & w2106 ) ;
  assign w2111 = ( w2108 & w2109 ) | ( w2108 & w2110 ) | ( w2109 & w2110 ) ;
  assign w2112 = \pi131 ^ w1217 ;
  assign w2113 = ( w1217 & w1280 ) | ( w1217 & w2112 ) | ( w1280 & w2112 ) ;
  assign w2114 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2113 ) | ( ~\pi131 & w2113 ) ;
  assign w2115 = w1224 | w2114 ;
  assign w2116 = w1231 & w2114 ;
  assign w2117 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2113 ) | ( \pi131 & w2113 ) ;
  assign w2118 = ( w2115 & w2116 ) | ( w2115 & w2117 ) | ( w2116 & w2117 ) ;
  assign w2119 = ( w1245 & ~w1267 ) | ( w1245 & w1287 ) | ( ~w1267 & w1287 ) ;
  assign w2120 = ( \pi130 & ~\pi131 ) | ( \pi130 & w2119 ) | ( ~\pi131 & w2119 ) ;
  assign w2121 = w1294 | w2120 ;
  assign w2122 = w1301 & w2120 ;
  assign w2123 = ( ~\pi130 & \pi131 ) | ( ~\pi130 & w2119 ) | ( \pi131 & w2119 ) ;
  assign w2124 = ( w2121 & w2122 ) | ( w2121 & w2123 ) | ( w2122 & w2123 ) ;
  assign w2125 = \pi132 ^ w2104 ;
  assign w2126 = ( w2104 & w2118 ) | ( w2104 & ~w2125 ) | ( w2118 & ~w2125 ) ;
  assign w2127 = ( \pi132 & \pi133 ) | ( \pi132 & w2126 ) | ( \pi133 & w2126 ) ;
  assign w2128 = w2111 | w2127 ;
  assign w2129 = w2124 & w2127 ;
  assign w2130 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2126 ) | ( \pi133 & ~w2126 ) ;
  assign w2131 = ( w2128 & w2129 ) | ( w2128 & ~w2130 ) | ( w2129 & ~w2130 ) ;
  assign w2132 = \pi134 ^ w2131 ;
  assign w2133 = ( w2097 & w2131 ) | ( w2097 & ~w2132 ) | ( w2131 & ~w2132 ) ;
  assign w2134 = \pi133 ^ w205 ;
  assign w2135 = ( w205 & w317 ) | ( w205 & ~w2134 ) | ( w317 & ~w2134 ) ;
  assign w2136 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2135 ) | ( \pi133 & w2135 ) ;
  assign w2137 = w240 | w2136 ;
  assign w2138 = w275 & w2136 ;
  assign w2139 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2135 ) | ( ~\pi133 & w2135 ) ;
  assign w2140 = ( w2137 & w2138 ) | ( w2137 & w2139 ) | ( w2138 & w2139 ) ;
  assign w2141 = ( w170 & w276 ) | ( w170 & w352 ) | ( w276 & w352 ) ;
  assign w2142 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2141 ) | ( \pi133 & w2141 ) ;
  assign w2143 = w387 | w2142 ;
  assign w2144 = w422 & w2142 ;
  assign w2145 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2141 ) | ( ~\pi133 & w2141 ) ;
  assign w2146 = ( w2143 & w2144 ) | ( w2143 & w2145 ) | ( w2144 & w2145 ) ;
  assign w2147 = \pi134 ^ w2146 ;
  assign w2148 = ( w2140 & w2146 ) | ( w2140 & ~w2147 ) | ( w2146 & ~w2147 ) ;
  assign w2149 = \pi133 ^ w501 ;
  assign w2150 = ( w501 & w648 ) | ( w501 & ~w2149 ) | ( w648 & ~w2149 ) ;
  assign w2151 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2150 ) | ( \pi133 & w2150 ) ;
  assign w2152 = w536 | w2151 ;
  assign w2153 = w571 & w2151 ;
  assign w2154 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2150 ) | ( ~\pi133 & w2150 ) ;
  assign w2155 = ( w2152 & w2153 ) | ( w2152 & w2154 ) | ( w2153 & w2154 ) ;
  assign w2156 = ( w466 & w572 ) | ( w466 & w718 ) | ( w572 & w718 ) ;
  assign w2157 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2156 ) | ( \pi133 & w2156 ) ;
  assign w2158 = w613 | w2157 ;
  assign w2159 = w683 & w2157 ;
  assign w2160 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2156 ) | ( ~\pi133 & w2156 ) ;
  assign w2161 = ( w2158 & w2159 ) | ( w2158 & w2160 ) | ( w2159 & w2160 ) ;
  assign w2162 = \pi134 ^ w2161 ;
  assign w2163 = ( w2155 & w2161 ) | ( w2155 & ~w2162 ) | ( w2161 & ~w2162 ) ;
  assign w2164 = \pi133 ^ w797 ;
  assign w2165 = ( w797 & w943 ) | ( w797 & ~w2164 ) | ( w943 & ~w2164 ) ;
  assign w2166 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2165 ) | ( \pi133 & w2165 ) ;
  assign w2167 = w831 | w2166 ;
  assign w2168 = w866 & w2166 ;
  assign w2169 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2165 ) | ( ~\pi133 & w2165 ) ;
  assign w2170 = ( w2167 & w2168 ) | ( w2167 & w2169 ) | ( w2168 & w2169 ) ;
  assign w2171 = ( w762 & w867 ) | ( w762 & w1013 ) | ( w867 & w1013 ) ;
  assign w2172 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2171 ) | ( \pi133 & w2171 ) ;
  assign w2173 = w908 | w2172 ;
  assign w2174 = w978 & w2172 ;
  assign w2175 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2171 ) | ( ~\pi133 & w2171 ) ;
  assign w2176 = ( w2173 & w2174 ) | ( w2173 & w2175 ) | ( w2174 & w2175 ) ;
  assign w2177 = \pi134 ^ w2176 ;
  assign w2178 = ( w2170 & w2176 ) | ( w2170 & ~w2177 ) | ( w2176 & ~w2177 ) ;
  assign w2179 = ( w1057 & w1126 ) | ( w1057 & w1162 ) | ( w1126 & w1162 ) ;
  assign w2180 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2179 ) | ( \pi133 & ~w2179 ) ;
  assign w2181 = ~w1092 & w2180 ;
  assign w2182 = w1273 & ~w2180 ;
  assign w2183 = ( \pi132 & \pi133 ) | ( \pi132 & w2179 ) | ( \pi133 & w2179 ) ;
  assign w2184 = ( ~w2181 & w2182 ) | ( ~w2181 & w2183 ) | ( w2182 & w2183 ) ;
  assign w2185 = \pi132 ^ w1161 ;
  assign w2186 = ( w1161 & w1308 ) | ( w1161 & w2185 ) | ( w1308 & w2185 ) ;
  assign w2187 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2186 ) | ( \pi133 & w2186 ) ;
  assign w2188 = w1203 | w2187 ;
  assign w2189 = w1238 & w2187 ;
  assign w2190 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2186 ) | ( ~\pi133 & w2186 ) ;
  assign w2191 = ( w2188 & w2189 ) | ( w2188 & w2190 ) | ( w2189 & w2190 ) ;
  assign w2192 = \pi134 ^ w2191 ;
  assign w2193 = ( w2184 & w2191 ) | ( w2184 & ~w2192 ) | ( w2191 & ~w2192 ) ;
  assign w2194 = \pi133 ^ w1331 ;
  assign w2195 = ( w1331 & w1380 ) | ( w1331 & ~w2194 ) | ( w1380 & ~w2194 ) ;
  assign w2196 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2195 ) | ( \pi133 & w2195 ) ;
  assign w2197 = w1338 | w2196 ;
  assign w2198 = w1345 & w2196 ;
  assign w2199 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2195 ) | ( ~\pi133 & w2195 ) ;
  assign w2200 = ( w2197 & w2198 ) | ( w2197 & w2199 ) | ( w2198 & w2199 ) ;
  assign w2201 = \pi133 ^ w1324 ;
  assign w2202 = ( w1324 & w1373 ) | ( w1324 & w2201 ) | ( w1373 & w2201 ) ;
  assign w2203 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2202 ) | ( ~\pi133 & w2202 ) ;
  assign w2204 = w1359 | w2203 ;
  assign w2205 = w1366 & w2203 ;
  assign w2206 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2202 ) | ( \pi133 & w2202 ) ;
  assign w2207 = ( w2204 & w2205 ) | ( w2204 & w2206 ) | ( w2205 & w2206 ) ;
  assign w2208 = \pi134 ^ w2207 ;
  assign w2209 = ( w2200 & w2207 ) | ( w2200 & ~w2208 ) | ( w2207 & ~w2208 ) ;
  assign w2210 = \pi133 ^ w1403 ;
  assign w2211 = ( w1403 & w1452 ) | ( w1403 & ~w2210 ) | ( w1452 & ~w2210 ) ;
  assign w2212 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2211 ) | ( \pi133 & w2211 ) ;
  assign w2213 = w1410 | w2212 ;
  assign w2214 = w1417 & w2212 ;
  assign w2215 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2211 ) | ( ~\pi133 & w2211 ) ;
  assign w2216 = ( w2213 & w2214 ) | ( w2213 & w2215 ) | ( w2214 & w2215 ) ;
  assign w2217 = \pi133 ^ w1396 ;
  assign w2218 = ( w1396 & w1445 ) | ( w1396 & w2217 ) | ( w1445 & w2217 ) ;
  assign w2219 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2218 ) | ( ~\pi133 & w2218 ) ;
  assign w2220 = w1431 | w2219 ;
  assign w2221 = w1438 & w2219 ;
  assign w2222 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2218 ) | ( \pi133 & w2218 ) ;
  assign w2223 = ( w2220 & w2221 ) | ( w2220 & w2222 ) | ( w2221 & w2222 ) ;
  assign w2224 = \pi134 ^ w2223 ;
  assign w2225 = ( w2216 & w2223 ) | ( w2216 & ~w2224 ) | ( w2223 & ~w2224 ) ;
  assign w2226 = \pi133 ^ w1475 ;
  assign w2227 = ( w1475 & w1524 ) | ( w1475 & ~w2226 ) | ( w1524 & ~w2226 ) ;
  assign w2228 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2227 ) | ( \pi133 & w2227 ) ;
  assign w2229 = w1482 | w2228 ;
  assign w2230 = w1489 & w2228 ;
  assign w2231 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2227 ) | ( ~\pi133 & w2227 ) ;
  assign w2232 = ( w2229 & w2230 ) | ( w2229 & w2231 ) | ( w2230 & w2231 ) ;
  assign w2233 = \pi133 ^ w1468 ;
  assign w2234 = ( w1468 & w1517 ) | ( w1468 & w2233 ) | ( w1517 & w2233 ) ;
  assign w2235 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2234 ) | ( ~\pi133 & w2234 ) ;
  assign w2236 = w1503 | w2235 ;
  assign w2237 = w1510 & w2235 ;
  assign w2238 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2234 ) | ( \pi133 & w2234 ) ;
  assign w2239 = ( w2236 & w2237 ) | ( w2236 & w2238 ) | ( w2237 & w2238 ) ;
  assign w2240 = \pi134 ^ w2239 ;
  assign w2241 = ( w2232 & w2239 ) | ( w2232 & ~w2240 ) | ( w2239 & ~w2240 ) ;
  assign w2242 = \pi133 ^ w1547 ;
  assign w2243 = ( w1547 & w1596 ) | ( w1547 & ~w2242 ) | ( w1596 & ~w2242 ) ;
  assign w2244 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2243 ) | ( \pi133 & w2243 ) ;
  assign w2245 = w1554 | w2244 ;
  assign w2246 = w1561 & w2244 ;
  assign w2247 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2243 ) | ( ~\pi133 & w2243 ) ;
  assign w2248 = ( w2245 & w2246 ) | ( w2245 & w2247 ) | ( w2246 & w2247 ) ;
  assign w2249 = \pi133 ^ w1540 ;
  assign w2250 = ( w1540 & w1589 ) | ( w1540 & w2249 ) | ( w1589 & w2249 ) ;
  assign w2251 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2250 ) | ( ~\pi133 & w2250 ) ;
  assign w2252 = w1575 | w2251 ;
  assign w2253 = w1582 & w2251 ;
  assign w2254 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2250 ) | ( \pi133 & w2250 ) ;
  assign w2255 = ( w2252 & w2253 ) | ( w2252 & w2254 ) | ( w2253 & w2254 ) ;
  assign w2256 = \pi134 ^ w2255 ;
  assign w2257 = ( w2248 & w2255 ) | ( w2248 & ~w2256 ) | ( w2255 & ~w2256 ) ;
  assign w2258 = \pi133 ^ w1617 ;
  assign w2259 = ( w1617 & w1660 ) | ( w1617 & ~w2258 ) | ( w1660 & ~w2258 ) ;
  assign w2260 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2259 ) | ( \pi133 & w2259 ) ;
  assign w2261 = w1623 | w2260 ;
  assign w2262 = w1629 & w2260 ;
  assign w2263 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2259 ) | ( ~\pi133 & w2259 ) ;
  assign w2264 = ( w2261 & w2262 ) | ( w2261 & w2263 ) | ( w2262 & w2263 ) ;
  assign w2265 = \pi133 ^ w1611 ;
  assign w2266 = ( w1611 & w1654 ) | ( w1611 & w2265 ) | ( w1654 & w2265 ) ;
  assign w2267 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2266 ) | ( ~\pi133 & w2266 ) ;
  assign w2268 = w1642 | w2267 ;
  assign w2269 = w1648 & w2267 ;
  assign w2270 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2266 ) | ( \pi133 & w2266 ) ;
  assign w2271 = ( w2268 & w2269 ) | ( w2268 & w2270 ) | ( w2269 & w2270 ) ;
  assign w2272 = \pi134 ^ w2271 ;
  assign w2273 = ( w2264 & w2271 ) | ( w2264 & ~w2272 ) | ( w2271 & ~w2272 ) ;
  assign w2274 = \pi133 ^ w1681 ;
  assign w2275 = ( w1681 & w1724 ) | ( w1681 & ~w2274 ) | ( w1724 & ~w2274 ) ;
  assign w2276 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2275 ) | ( \pi133 & w2275 ) ;
  assign w2277 = w1687 | w2276 ;
  assign w2278 = w1693 & w2276 ;
  assign w2279 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2275 ) | ( ~\pi133 & w2275 ) ;
  assign w2280 = ( w2277 & w2278 ) | ( w2277 & w2279 ) | ( w2278 & w2279 ) ;
  assign w2281 = \pi133 ^ w1675 ;
  assign w2282 = ( w1675 & w1718 ) | ( w1675 & w2281 ) | ( w1718 & w2281 ) ;
  assign w2283 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2282 ) | ( ~\pi133 & w2282 ) ;
  assign w2284 = w1706 | w2283 ;
  assign w2285 = w1712 & w2283 ;
  assign w2286 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2282 ) | ( \pi133 & w2282 ) ;
  assign w2287 = ( w2284 & w2285 ) | ( w2284 & w2286 ) | ( w2285 & w2286 ) ;
  assign w2288 = \pi134 ^ w2287 ;
  assign w2289 = ( w2280 & w2287 ) | ( w2280 & ~w2288 ) | ( w2287 & ~w2288 ) ;
  assign w2290 = \pi133 ^ w1745 ;
  assign w2291 = ( w1745 & w1788 ) | ( w1745 & ~w2290 ) | ( w1788 & ~w2290 ) ;
  assign w2292 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2291 ) | ( \pi133 & w2291 ) ;
  assign w2293 = w1751 | w2292 ;
  assign w2294 = w1757 & w2292 ;
  assign w2295 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2291 ) | ( ~\pi133 & w2291 ) ;
  assign w2296 = ( w2293 & w2294 ) | ( w2293 & w2295 ) | ( w2294 & w2295 ) ;
  assign w2297 = \pi133 ^ w1739 ;
  assign w2298 = ( w1739 & w1782 ) | ( w1739 & w2297 ) | ( w1782 & w2297 ) ;
  assign w2299 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2298 ) | ( ~\pi133 & w2298 ) ;
  assign w2300 = w1770 | w2299 ;
  assign w2301 = w1776 & w2299 ;
  assign w2302 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2298 ) | ( \pi133 & w2298 ) ;
  assign w2303 = ( w2300 & w2301 ) | ( w2300 & w2302 ) | ( w2301 & w2302 ) ;
  assign w2304 = \pi134 ^ w2303 ;
  assign w2305 = ( w2296 & w2303 ) | ( w2296 & ~w2304 ) | ( w2303 & ~w2304 ) ;
  assign w2306 = \pi133 ^ w1809 ;
  assign w2307 = ( w1809 & w1852 ) | ( w1809 & ~w2306 ) | ( w1852 & ~w2306 ) ;
  assign w2308 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2307 ) | ( \pi133 & w2307 ) ;
  assign w2309 = w1815 | w2308 ;
  assign w2310 = w1821 & w2308 ;
  assign w2311 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2307 ) | ( ~\pi133 & w2307 ) ;
  assign w2312 = ( w2309 & w2310 ) | ( w2309 & w2311 ) | ( w2310 & w2311 ) ;
  assign w2313 = \pi133 ^ w1803 ;
  assign w2314 = ( w1803 & w1846 ) | ( w1803 & w2313 ) | ( w1846 & w2313 ) ;
  assign w2315 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2314 ) | ( ~\pi133 & w2314 ) ;
  assign w2316 = w1834 | w2315 ;
  assign w2317 = w1840 & w2315 ;
  assign w2318 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2314 ) | ( \pi133 & w2314 ) ;
  assign w2319 = ( w2316 & w2317 ) | ( w2316 & w2318 ) | ( w2317 & w2318 ) ;
  assign w2320 = \pi134 ^ w2319 ;
  assign w2321 = ( w2312 & w2319 ) | ( w2312 & ~w2320 ) | ( w2319 & ~w2320 ) ;
  assign w2322 = \pi133 ^ w1873 ;
  assign w2323 = ( w1873 & w1919 ) | ( w1873 & ~w2322 ) | ( w1919 & ~w2322 ) ;
  assign w2324 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2323 ) | ( \pi133 & w2323 ) ;
  assign w2325 = w1879 | w2324 ;
  assign w2326 = w1886 & w2324 ;
  assign w2327 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2323 ) | ( ~\pi133 & w2323 ) ;
  assign w2328 = ( w2325 & w2326 ) | ( w2325 & w2327 ) | ( w2326 & w2327 ) ;
  assign w2329 = \pi133 ^ w1867 ;
  assign w2330 = ( w1867 & w1913 ) | ( w1867 & w2329 ) | ( w1913 & w2329 ) ;
  assign w2331 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2330 ) | ( ~\pi133 & w2330 ) ;
  assign w2332 = w1900 | w2331 ;
  assign w2333 = w1907 & w2331 ;
  assign w2334 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2330 ) | ( \pi133 & w2330 ) ;
  assign w2335 = ( w2332 & w2333 ) | ( w2332 & w2334 ) | ( w2333 & w2334 ) ;
  assign w2336 = \pi134 ^ w2335 ;
  assign w2337 = ( w2328 & w2335 ) | ( w2328 & ~w2336 ) | ( w2335 & ~w2336 ) ;
  assign w2338 = \pi133 ^ w1940 ;
  assign w2339 = ( w1940 & w1987 ) | ( w1940 & ~w2338 ) | ( w1987 & ~w2338 ) ;
  assign w2340 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2339 ) | ( \pi133 & w2339 ) ;
  assign w2341 = w1946 | w2340 ;
  assign w2342 = w1953 & w2340 ;
  assign w2343 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2339 ) | ( ~\pi133 & w2339 ) ;
  assign w2344 = ( w2341 & w2342 ) | ( w2341 & w2343 ) | ( w2342 & w2343 ) ;
  assign w2345 = \pi133 ^ w1934 ;
  assign w2346 = ( w1934 & w1981 ) | ( w1934 & w2345 ) | ( w1981 & w2345 ) ;
  assign w2347 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2346 ) | ( ~\pi133 & w2346 ) ;
  assign w2348 = w1967 | w2347 ;
  assign w2349 = w1974 & w2347 ;
  assign w2350 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2346 ) | ( \pi133 & w2346 ) ;
  assign w2351 = ( w2348 & w2349 ) | ( w2348 & w2350 ) | ( w2349 & w2350 ) ;
  assign w2352 = \pi134 ^ w2351 ;
  assign w2353 = ( w2344 & w2351 ) | ( w2344 & ~w2352 ) | ( w2351 & ~w2352 ) ;
  assign w2354 = \pi133 ^ w2008 ;
  assign w2355 = ( w2008 & w2055 ) | ( w2008 & ~w2354 ) | ( w2055 & ~w2354 ) ;
  assign w2356 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2355 ) | ( \pi133 & w2355 ) ;
  assign w2357 = w2014 | w2356 ;
  assign w2358 = w2021 & w2356 ;
  assign w2359 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2355 ) | ( ~\pi133 & w2355 ) ;
  assign w2360 = ( w2357 & w2358 ) | ( w2357 & w2359 ) | ( w2358 & w2359 ) ;
  assign w2361 = \pi133 ^ w2002 ;
  assign w2362 = ( w2002 & w2049 ) | ( w2002 & w2361 ) | ( w2049 & w2361 ) ;
  assign w2363 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2362 ) | ( ~\pi133 & w2362 ) ;
  assign w2364 = w2035 | w2363 ;
  assign w2365 = w2042 & w2363 ;
  assign w2366 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2362 ) | ( \pi133 & w2362 ) ;
  assign w2367 = ( w2364 & w2365 ) | ( w2364 & w2366 ) | ( w2365 & w2366 ) ;
  assign w2368 = \pi134 ^ w2367 ;
  assign w2369 = ( w2360 & w2367 ) | ( w2360 & ~w2368 ) | ( w2367 & ~w2368 ) ;
  assign w2370 = \pi133 ^ w2078 ;
  assign w2371 = ( w2078 & w2124 ) | ( w2078 & ~w2370 ) | ( w2124 & ~w2370 ) ;
  assign w2372 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2371 ) | ( \pi133 & w2371 ) ;
  assign w2373 = w2084 | w2372 ;
  assign w2374 = w2090 & w2372 ;
  assign w2375 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2371 ) | ( ~\pi133 & w2371 ) ;
  assign w2376 = ( w2373 & w2374 ) | ( w2373 & w2375 ) | ( w2374 & w2375 ) ;
  assign w2377 = \pi133 ^ w2071 ;
  assign w2378 = ( w2071 & w2118 ) | ( w2071 & w2377 ) | ( w2118 & w2377 ) ;
  assign w2379 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2378 ) | ( ~\pi133 & w2378 ) ;
  assign w2380 = w2104 | w2379 ;
  assign w2381 = w2111 & w2379 ;
  assign w2382 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2378 ) | ( \pi133 & w2378 ) ;
  assign w2383 = ( w2380 & w2381 ) | ( w2380 & w2382 ) | ( w2381 & w2382 ) ;
  assign w2384 = \pi134 ^ w2383 ;
  assign w2385 = ( w2376 & w2383 ) | ( w2376 & ~w2384 ) | ( w2383 & ~w2384 ) ;
  assign w2386 = \pi132 ^ w240 ;
  assign w2387 = ( w240 & w317 ) | ( w240 & w2386 ) | ( w317 & w2386 ) ;
  assign w2388 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2387 ) | ( \pi133 & ~w2387 ) ;
  assign w2389 = ~w275 & w2388 ;
  assign w2390 = w352 & ~w2388 ;
  assign w2391 = ( \pi132 & \pi133 ) | ( \pi132 & w2387 ) | ( \pi133 & w2387 ) ;
  assign w2392 = ( ~w2389 & w2390 ) | ( ~w2389 & w2391 ) | ( w2390 & w2391 ) ;
  assign w2393 = ( w170 & ~w276 ) | ( w170 & w387 ) | ( ~w276 & w387 ) ;
  assign w2394 = ( \pi132 & \pi133 ) | ( \pi132 & w2393 ) | ( \pi133 & w2393 ) ;
  assign w2395 = w205 | w2394 ;
  assign w2396 = w422 & w2394 ;
  assign w2397 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2393 ) | ( \pi133 & ~w2393 ) ;
  assign w2398 = ( w2395 & w2396 ) | ( w2395 & ~w2397 ) | ( w2396 & ~w2397 ) ;
  assign w2399 = \pi134 ^ w2398 ;
  assign w2400 = ( w2392 & w2398 ) | ( w2392 & ~w2399 ) | ( w2398 & ~w2399 ) ;
  assign w2401 = \pi132 ^ w536 ;
  assign w2402 = ( w536 & w648 ) | ( w536 & w2401 ) | ( w648 & w2401 ) ;
  assign w2403 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2402 ) | ( \pi133 & ~w2402 ) ;
  assign w2404 = ~w571 & w2403 ;
  assign w2405 = w718 & ~w2403 ;
  assign w2406 = ( \pi132 & \pi133 ) | ( \pi132 & w2402 ) | ( \pi133 & w2402 ) ;
  assign w2407 = ( ~w2404 & w2405 ) | ( ~w2404 & w2406 ) | ( w2405 & w2406 ) ;
  assign w2408 = ( w466 & ~w572 ) | ( w466 & w613 ) | ( ~w572 & w613 ) ;
  assign w2409 = ( \pi132 & \pi133 ) | ( \pi132 & w2408 ) | ( \pi133 & w2408 ) ;
  assign w2410 = w501 | w2409 ;
  assign w2411 = w683 & w2409 ;
  assign w2412 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2408 ) | ( \pi133 & ~w2408 ) ;
  assign w2413 = ( w2410 & w2411 ) | ( w2410 & ~w2412 ) | ( w2411 & ~w2412 ) ;
  assign w2414 = \pi134 ^ w2413 ;
  assign w2415 = ( w2407 & w2413 ) | ( w2407 & ~w2414 ) | ( w2413 & ~w2414 ) ;
  assign w2416 = \pi132 ^ w831 ;
  assign w2417 = ( w831 & w943 ) | ( w831 & w2416 ) | ( w943 & w2416 ) ;
  assign w2418 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2417 ) | ( \pi133 & ~w2417 ) ;
  assign w2419 = ~w866 & w2418 ;
  assign w2420 = w1013 & ~w2418 ;
  assign w2421 = ( \pi132 & \pi133 ) | ( \pi132 & w2417 ) | ( \pi133 & w2417 ) ;
  assign w2422 = ( ~w2419 & w2420 ) | ( ~w2419 & w2421 ) | ( w2420 & w2421 ) ;
  assign w2423 = ( w762 & ~w867 ) | ( w762 & w908 ) | ( ~w867 & w908 ) ;
  assign w2424 = ( \pi132 & \pi133 ) | ( \pi132 & w2423 ) | ( \pi133 & w2423 ) ;
  assign w2425 = w797 | w2424 ;
  assign w2426 = w978 & w2424 ;
  assign w2427 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2423 ) | ( \pi133 & ~w2423 ) ;
  assign w2428 = ( w2425 & w2426 ) | ( w2425 & ~w2427 ) | ( w2426 & ~w2427 ) ;
  assign w2429 = \pi134 ^ w2428 ;
  assign w2430 = ( w2422 & w2428 ) | ( w2422 & ~w2429 ) | ( w2428 & ~w2429 ) ;
  assign w2431 = ( w1057 & ~w1162 ) | ( w1057 & w1308 ) | ( ~w1162 & w1308 ) ;
  assign w2432 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2431 ) | ( ~\pi133 & w2431 ) ;
  assign w2433 = w1126 | w2432 ;
  assign w2434 = w1273 & w2432 ;
  assign w2435 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2431 ) | ( \pi133 & w2431 ) ;
  assign w2436 = ( w2433 & w2434 ) | ( w2433 & w2435 ) | ( w2434 & w2435 ) ;
  assign w2437 = \pi132 ^ w1092 ;
  assign w2438 = ( w1092 & w1238 ) | ( w1092 & w2437 ) | ( w1238 & w2437 ) ;
  assign w2439 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2438 ) | ( \pi133 & w2438 ) ;
  assign w2440 = w1161 | w2439 ;
  assign w2441 = w1203 & w2439 ;
  assign w2442 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2438 ) | ( ~\pi133 & w2438 ) ;
  assign w2443 = ( w2440 & w2441 ) | ( w2440 & w2442 ) | ( w2441 & w2442 ) ;
  assign w2444 = \pi134 ^ w2443 ;
  assign w2445 = ( w2436 & w2443 ) | ( w2436 & ~w2444 ) | ( w2443 & ~w2444 ) ;
  assign w2446 = \pi132 ^ w1338 ;
  assign w2447 = ( w1338 & w1380 ) | ( w1338 & w2446 ) | ( w1380 & w2446 ) ;
  assign w2448 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2447 ) | ( \pi133 & ~w2447 ) ;
  assign w2449 = ~w1345 & w2448 ;
  assign w2450 = w1373 & ~w2448 ;
  assign w2451 = ( \pi132 & \pi133 ) | ( \pi132 & w2447 ) | ( \pi133 & w2447 ) ;
  assign w2452 = ( ~w2449 & w2450 ) | ( ~w2449 & w2451 ) | ( w2450 & w2451 ) ;
  assign w2453 = ( w1324 & ~w1346 ) | ( w1324 & w1366 ) | ( ~w1346 & w1366 ) ;
  assign w2454 = ( \pi132 & \pi133 ) | ( \pi132 & w2453 ) | ( \pi133 & w2453 ) ;
  assign w2455 = w1331 | w2454 ;
  assign w2456 = w1359 & w2454 ;
  assign w2457 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2453 ) | ( \pi133 & ~w2453 ) ;
  assign w2458 = ( w2455 & w2456 ) | ( w2455 & ~w2457 ) | ( w2456 & ~w2457 ) ;
  assign w2459 = \pi134 ^ w2458 ;
  assign w2460 = ( w2452 & w2458 ) | ( w2452 & ~w2459 ) | ( w2458 & ~w2459 ) ;
  assign w2461 = \pi132 ^ w1410 ;
  assign w2462 = ( w1410 & w1452 ) | ( w1410 & w2461 ) | ( w1452 & w2461 ) ;
  assign w2463 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2462 ) | ( \pi133 & ~w2462 ) ;
  assign w2464 = ~w1417 & w2463 ;
  assign w2465 = w1445 & ~w2463 ;
  assign w2466 = ( \pi132 & \pi133 ) | ( \pi132 & w2462 ) | ( \pi133 & w2462 ) ;
  assign w2467 = ( ~w2464 & w2465 ) | ( ~w2464 & w2466 ) | ( w2465 & w2466 ) ;
  assign w2468 = ( w1396 & ~w1418 ) | ( w1396 & w1438 ) | ( ~w1418 & w1438 ) ;
  assign w2469 = ( \pi132 & \pi133 ) | ( \pi132 & w2468 ) | ( \pi133 & w2468 ) ;
  assign w2470 = w1403 | w2469 ;
  assign w2471 = w1431 & w2469 ;
  assign w2472 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2468 ) | ( \pi133 & ~w2468 ) ;
  assign w2473 = ( w2470 & w2471 ) | ( w2470 & ~w2472 ) | ( w2471 & ~w2472 ) ;
  assign w2474 = \pi134 ^ w2473 ;
  assign w2475 = ( w2467 & w2473 ) | ( w2467 & ~w2474 ) | ( w2473 & ~w2474 ) ;
  assign w2476 = \pi132 ^ w1482 ;
  assign w2477 = ( w1482 & w1524 ) | ( w1482 & w2476 ) | ( w1524 & w2476 ) ;
  assign w2478 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2477 ) | ( \pi133 & ~w2477 ) ;
  assign w2479 = ~w1489 & w2478 ;
  assign w2480 = w1517 & ~w2478 ;
  assign w2481 = ( \pi132 & \pi133 ) | ( \pi132 & w2477 ) | ( \pi133 & w2477 ) ;
  assign w2482 = ( ~w2479 & w2480 ) | ( ~w2479 & w2481 ) | ( w2480 & w2481 ) ;
  assign w2483 = ( w1468 & ~w1490 ) | ( w1468 & w1510 ) | ( ~w1490 & w1510 ) ;
  assign w2484 = ( \pi132 & \pi133 ) | ( \pi132 & w2483 ) | ( \pi133 & w2483 ) ;
  assign w2485 = w1475 | w2484 ;
  assign w2486 = w1503 & w2484 ;
  assign w2487 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2483 ) | ( \pi133 & ~w2483 ) ;
  assign w2488 = ( w2485 & w2486 ) | ( w2485 & ~w2487 ) | ( w2486 & ~w2487 ) ;
  assign w2489 = \pi134 ^ w2488 ;
  assign w2490 = ( w2482 & w2488 ) | ( w2482 & ~w2489 ) | ( w2488 & ~w2489 ) ;
  assign w2491 = \pi132 ^ w1554 ;
  assign w2492 = ( w1554 & w1596 ) | ( w1554 & w2491 ) | ( w1596 & w2491 ) ;
  assign w2493 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2492 ) | ( \pi133 & ~w2492 ) ;
  assign w2494 = ~w1561 & w2493 ;
  assign w2495 = w1589 & ~w2493 ;
  assign w2496 = ( \pi132 & \pi133 ) | ( \pi132 & w2492 ) | ( \pi133 & w2492 ) ;
  assign w2497 = ( ~w2494 & w2495 ) | ( ~w2494 & w2496 ) | ( w2495 & w2496 ) ;
  assign w2498 = ( w1540 & ~w1562 ) | ( w1540 & w1582 ) | ( ~w1562 & w1582 ) ;
  assign w2499 = ( \pi132 & \pi133 ) | ( \pi132 & w2498 ) | ( \pi133 & w2498 ) ;
  assign w2500 = w1547 | w2499 ;
  assign w2501 = w1575 & w2499 ;
  assign w2502 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2498 ) | ( \pi133 & ~w2498 ) ;
  assign w2503 = ( w2500 & w2501 ) | ( w2500 & ~w2502 ) | ( w2501 & ~w2502 ) ;
  assign w2504 = \pi134 ^ w2503 ;
  assign w2505 = ( w2497 & w2503 ) | ( w2497 & ~w2504 ) | ( w2503 & ~w2504 ) ;
  assign w2506 = \pi132 ^ w1623 ;
  assign w2507 = ( w1623 & w1660 ) | ( w1623 & w2506 ) | ( w1660 & w2506 ) ;
  assign w2508 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2507 ) | ( \pi133 & ~w2507 ) ;
  assign w2509 = ~w1629 & w2508 ;
  assign w2510 = w1654 & ~w2508 ;
  assign w2511 = ( \pi132 & \pi133 ) | ( \pi132 & w2507 ) | ( \pi133 & w2507 ) ;
  assign w2512 = ( ~w2509 & w2510 ) | ( ~w2509 & w2511 ) | ( w2510 & w2511 ) ;
  assign w2513 = ( w1611 & ~w1630 ) | ( w1611 & w1648 ) | ( ~w1630 & w1648 ) ;
  assign w2514 = ( \pi132 & \pi133 ) | ( \pi132 & w2513 ) | ( \pi133 & w2513 ) ;
  assign w2515 = w1617 | w2514 ;
  assign w2516 = w1642 & w2514 ;
  assign w2517 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2513 ) | ( \pi133 & ~w2513 ) ;
  assign w2518 = ( w2515 & w2516 ) | ( w2515 & ~w2517 ) | ( w2516 & ~w2517 ) ;
  assign w2519 = \pi134 ^ w2518 ;
  assign w2520 = ( w2512 & w2518 ) | ( w2512 & ~w2519 ) | ( w2518 & ~w2519 ) ;
  assign w2521 = \pi132 ^ w1687 ;
  assign w2522 = ( w1687 & w1724 ) | ( w1687 & w2521 ) | ( w1724 & w2521 ) ;
  assign w2523 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2522 ) | ( \pi133 & ~w2522 ) ;
  assign w2524 = ~w1693 & w2523 ;
  assign w2525 = w1718 & ~w2523 ;
  assign w2526 = ( \pi132 & \pi133 ) | ( \pi132 & w2522 ) | ( \pi133 & w2522 ) ;
  assign w2527 = ( ~w2524 & w2525 ) | ( ~w2524 & w2526 ) | ( w2525 & w2526 ) ;
  assign w2528 = ( w1675 & ~w1694 ) | ( w1675 & w1712 ) | ( ~w1694 & w1712 ) ;
  assign w2529 = ( \pi132 & \pi133 ) | ( \pi132 & w2528 ) | ( \pi133 & w2528 ) ;
  assign w2530 = w1681 | w2529 ;
  assign w2531 = w1706 & w2529 ;
  assign w2532 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2528 ) | ( \pi133 & ~w2528 ) ;
  assign w2533 = ( w2530 & w2531 ) | ( w2530 & ~w2532 ) | ( w2531 & ~w2532 ) ;
  assign w2534 = \pi134 ^ w2533 ;
  assign w2535 = ( w2527 & w2533 ) | ( w2527 & ~w2534 ) | ( w2533 & ~w2534 ) ;
  assign w2536 = \pi132 ^ w1751 ;
  assign w2537 = ( w1751 & w1788 ) | ( w1751 & w2536 ) | ( w1788 & w2536 ) ;
  assign w2538 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2537 ) | ( \pi133 & ~w2537 ) ;
  assign w2539 = ~w1757 & w2538 ;
  assign w2540 = w1782 & ~w2538 ;
  assign w2541 = ( \pi132 & \pi133 ) | ( \pi132 & w2537 ) | ( \pi133 & w2537 ) ;
  assign w2542 = ( ~w2539 & w2540 ) | ( ~w2539 & w2541 ) | ( w2540 & w2541 ) ;
  assign w2543 = ( w1739 & ~w1758 ) | ( w1739 & w1776 ) | ( ~w1758 & w1776 ) ;
  assign w2544 = ( \pi132 & \pi133 ) | ( \pi132 & w2543 ) | ( \pi133 & w2543 ) ;
  assign w2545 = w1745 | w2544 ;
  assign w2546 = w1770 & w2544 ;
  assign w2547 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2543 ) | ( \pi133 & ~w2543 ) ;
  assign w2548 = ( w2545 & w2546 ) | ( w2545 & ~w2547 ) | ( w2546 & ~w2547 ) ;
  assign w2549 = \pi134 ^ w2548 ;
  assign w2550 = ( w2542 & w2548 ) | ( w2542 & ~w2549 ) | ( w2548 & ~w2549 ) ;
  assign w2551 = \pi132 ^ w1815 ;
  assign w2552 = ( w1815 & w1852 ) | ( w1815 & w2551 ) | ( w1852 & w2551 ) ;
  assign w2553 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2552 ) | ( \pi133 & ~w2552 ) ;
  assign w2554 = ~w1821 & w2553 ;
  assign w2555 = w1846 & ~w2553 ;
  assign w2556 = ( \pi132 & \pi133 ) | ( \pi132 & w2552 ) | ( \pi133 & w2552 ) ;
  assign w2557 = ( ~w2554 & w2555 ) | ( ~w2554 & w2556 ) | ( w2555 & w2556 ) ;
  assign w2558 = ( w1803 & ~w1822 ) | ( w1803 & w1840 ) | ( ~w1822 & w1840 ) ;
  assign w2559 = ( \pi132 & \pi133 ) | ( \pi132 & w2558 ) | ( \pi133 & w2558 ) ;
  assign w2560 = w1809 | w2559 ;
  assign w2561 = w1834 & w2559 ;
  assign w2562 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2558 ) | ( \pi133 & ~w2558 ) ;
  assign w2563 = ( w2560 & w2561 ) | ( w2560 & ~w2562 ) | ( w2561 & ~w2562 ) ;
  assign w2564 = \pi134 ^ w2563 ;
  assign w2565 = ( w2557 & w2563 ) | ( w2557 & ~w2564 ) | ( w2563 & ~w2564 ) ;
  assign w2566 = \pi132 ^ w1879 ;
  assign w2567 = ( w1879 & w1919 ) | ( w1879 & w2566 ) | ( w1919 & w2566 ) ;
  assign w2568 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2567 ) | ( \pi133 & ~w2567 ) ;
  assign w2569 = ~w1886 & w2568 ;
  assign w2570 = w1913 & ~w2568 ;
  assign w2571 = ( \pi132 & \pi133 ) | ( \pi132 & w2567 ) | ( \pi133 & w2567 ) ;
  assign w2572 = ( ~w2569 & w2570 ) | ( ~w2569 & w2571 ) | ( w2570 & w2571 ) ;
  assign w2573 = ( w1867 & ~w1887 ) | ( w1867 & w1907 ) | ( ~w1887 & w1907 ) ;
  assign w2574 = ( \pi132 & \pi133 ) | ( \pi132 & w2573 ) | ( \pi133 & w2573 ) ;
  assign w2575 = w1873 | w2574 ;
  assign w2576 = w1900 & w2574 ;
  assign w2577 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2573 ) | ( \pi133 & ~w2573 ) ;
  assign w2578 = ( w2575 & w2576 ) | ( w2575 & ~w2577 ) | ( w2576 & ~w2577 ) ;
  assign w2579 = \pi134 ^ w2578 ;
  assign w2580 = ( w2572 & w2578 ) | ( w2572 & ~w2579 ) | ( w2578 & ~w2579 ) ;
  assign w2581 = \pi132 ^ w1946 ;
  assign w2582 = ( w1946 & w1987 ) | ( w1946 & w2581 ) | ( w1987 & w2581 ) ;
  assign w2583 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2582 ) | ( \pi133 & ~w2582 ) ;
  assign w2584 = ~w1953 & w2583 ;
  assign w2585 = w1981 & ~w2583 ;
  assign w2586 = ( \pi132 & \pi133 ) | ( \pi132 & w2582 ) | ( \pi133 & w2582 ) ;
  assign w2587 = ( ~w2584 & w2585 ) | ( ~w2584 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2588 = ( w1934 & ~w1954 ) | ( w1934 & w1974 ) | ( ~w1954 & w1974 ) ;
  assign w2589 = ( \pi132 & \pi133 ) | ( \pi132 & w2588 ) | ( \pi133 & w2588 ) ;
  assign w2590 = w1940 | w2589 ;
  assign w2591 = w1967 & w2589 ;
  assign w2592 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2588 ) | ( \pi133 & ~w2588 ) ;
  assign w2593 = ( w2590 & w2591 ) | ( w2590 & ~w2592 ) | ( w2591 & ~w2592 ) ;
  assign w2594 = \pi134 ^ w2593 ;
  assign w2595 = ( w2587 & w2593 ) | ( w2587 & ~w2594 ) | ( w2593 & ~w2594 ) ;
  assign w2596 = \pi132 ^ w2014 ;
  assign w2597 = ( w2014 & w2055 ) | ( w2014 & w2596 ) | ( w2055 & w2596 ) ;
  assign w2598 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2597 ) | ( \pi133 & ~w2597 ) ;
  assign w2599 = ~w2021 & w2598 ;
  assign w2600 = w2049 & ~w2598 ;
  assign w2601 = ( \pi132 & \pi133 ) | ( \pi132 & w2597 ) | ( \pi133 & w2597 ) ;
  assign w2602 = ( ~w2599 & w2600 ) | ( ~w2599 & w2601 ) | ( w2600 & w2601 ) ;
  assign w2603 = ( w2002 & ~w2022 ) | ( w2002 & w2042 ) | ( ~w2022 & w2042 ) ;
  assign w2604 = ( \pi132 & \pi133 ) | ( \pi132 & w2603 ) | ( \pi133 & w2603 ) ;
  assign w2605 = w2008 | w2604 ;
  assign w2606 = w2035 & w2604 ;
  assign w2607 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2603 ) | ( \pi133 & ~w2603 ) ;
  assign w2608 = ( w2605 & w2606 ) | ( w2605 & ~w2607 ) | ( w2606 & ~w2607 ) ;
  assign w2609 = \pi134 ^ w2608 ;
  assign w2610 = ( w2602 & w2608 ) | ( w2602 & ~w2609 ) | ( w2608 & ~w2609 ) ;
  assign w2611 = \pi132 ^ w2084 ;
  assign w2612 = ( w2084 & w2124 ) | ( w2084 & w2611 ) | ( w2124 & w2611 ) ;
  assign w2613 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2612 ) | ( \pi133 & ~w2612 ) ;
  assign w2614 = ~w2090 & w2613 ;
  assign w2615 = w2118 & ~w2613 ;
  assign w2616 = ( \pi132 & \pi133 ) | ( \pi132 & w2612 ) | ( \pi133 & w2612 ) ;
  assign w2617 = ( ~w2614 & w2615 ) | ( ~w2614 & w2616 ) | ( w2615 & w2616 ) ;
  assign w2618 = ( w2071 & ~w2091 ) | ( w2071 & w2111 ) | ( ~w2091 & w2111 ) ;
  assign w2619 = ( \pi132 & \pi133 ) | ( \pi132 & w2618 ) | ( \pi133 & w2618 ) ;
  assign w2620 = w2078 | w2619 ;
  assign w2621 = w2104 & w2619 ;
  assign w2622 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2618 ) | ( \pi133 & ~w2618 ) ;
  assign w2623 = ( w2620 & w2621 ) | ( w2620 & ~w2622 ) | ( w2621 & ~w2622 ) ;
  assign w2624 = \pi134 ^ w2623 ;
  assign w2625 = ( w2617 & w2623 ) | ( w2617 & ~w2624 ) | ( w2623 & ~w2624 ) ;
  assign w2626 = ( w240 & w422 ) | ( w240 & ~w2386 ) | ( w422 & ~w2386 ) ;
  assign w2627 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2626 ) | ( ~\pi133 & w2626 ) ;
  assign w2628 = w317 | w2627 ;
  assign w2629 = w352 & w2627 ;
  assign w2630 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2626 ) | ( \pi133 & w2626 ) ;
  assign w2631 = ( w2628 & w2629 ) | ( w2628 & w2630 ) | ( w2629 & w2630 ) ;
  assign w2632 = \pi133 ^ w170 ;
  assign w2633 = ( w170 & w205 ) | ( w170 & ~w2632 ) | ( w205 & ~w2632 ) ;
  assign w2634 = ( \pi132 & \pi133 ) | ( \pi132 & w2633 ) | ( \pi133 & w2633 ) ;
  assign w2635 = w275 | w2634 ;
  assign w2636 = w387 & w2634 ;
  assign w2637 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2633 ) | ( \pi133 & ~w2633 ) ;
  assign w2638 = ( w2635 & w2636 ) | ( w2635 & ~w2637 ) | ( w2636 & ~w2637 ) ;
  assign w2639 = \pi134 ^ w2638 ;
  assign w2640 = ( w2631 & w2638 ) | ( w2631 & ~w2639 ) | ( w2638 & ~w2639 ) ;
  assign w2641 = ( w536 & w683 ) | ( w536 & ~w2401 ) | ( w683 & ~w2401 ) ;
  assign w2642 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2641 ) | ( ~\pi133 & w2641 ) ;
  assign w2643 = w648 | w2642 ;
  assign w2644 = w718 & w2642 ;
  assign w2645 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2641 ) | ( \pi133 & w2641 ) ;
  assign w2646 = ( w2643 & w2644 ) | ( w2643 & w2645 ) | ( w2644 & w2645 ) ;
  assign w2647 = \pi133 ^ w466 ;
  assign w2648 = ( w466 & w501 ) | ( w466 & ~w2647 ) | ( w501 & ~w2647 ) ;
  assign w2649 = ( \pi132 & \pi133 ) | ( \pi132 & w2648 ) | ( \pi133 & w2648 ) ;
  assign w2650 = w571 | w2649 ;
  assign w2651 = w613 & w2649 ;
  assign w2652 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2648 ) | ( \pi133 & ~w2648 ) ;
  assign w2653 = ( w2650 & w2651 ) | ( w2650 & ~w2652 ) | ( w2651 & ~w2652 ) ;
  assign w2654 = \pi134 ^ w2653 ;
  assign w2655 = ( w2646 & w2653 ) | ( w2646 & ~w2654 ) | ( w2653 & ~w2654 ) ;
  assign w2656 = ( w831 & w978 ) | ( w831 & ~w2416 ) | ( w978 & ~w2416 ) ;
  assign w2657 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2656 ) | ( ~\pi133 & w2656 ) ;
  assign w2658 = w943 | w2657 ;
  assign w2659 = w1013 & w2657 ;
  assign w2660 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2656 ) | ( \pi133 & w2656 ) ;
  assign w2661 = ( w2658 & w2659 ) | ( w2658 & w2660 ) | ( w2659 & w2660 ) ;
  assign w2662 = \pi133 ^ w762 ;
  assign w2663 = ( w762 & w797 ) | ( w762 & ~w2662 ) | ( w797 & ~w2662 ) ;
  assign w2664 = ( \pi132 & \pi133 ) | ( \pi132 & w2663 ) | ( \pi133 & w2663 ) ;
  assign w2665 = w866 | w2664 ;
  assign w2666 = w908 & w2664 ;
  assign w2667 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2663 ) | ( \pi133 & ~w2663 ) ;
  assign w2668 = ( w2665 & w2666 ) | ( w2665 & ~w2667 ) | ( w2666 & ~w2667 ) ;
  assign w2669 = \pi134 ^ w2668 ;
  assign w2670 = ( w2661 & w2668 ) | ( w2661 & ~w2669 ) | ( w2668 & ~w2669 ) ;
  assign w2671 = \pi132 ^ w1126 ;
  assign w2672 = ( w1126 & w1238 ) | ( w1126 & ~w2671 ) | ( w1238 & ~w2671 ) ;
  assign w2673 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2672 ) | ( ~\pi133 & w2672 ) ;
  assign w2674 = w1273 | w2673 ;
  assign w2675 = w1308 & w2673 ;
  assign w2676 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2672 ) | ( \pi133 & w2672 ) ;
  assign w2677 = ( w2674 & w2675 ) | ( w2674 & w2676 ) | ( w2675 & w2676 ) ;
  assign w2678 = ( w1057 & w1162 ) | ( w1057 & w1203 ) | ( w1162 & w1203 ) ;
  assign w2679 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2678 ) | ( \pi133 & w2678 ) ;
  assign w2680 = w1092 | w2679 ;
  assign w2681 = w1161 & w2679 ;
  assign w2682 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2678 ) | ( ~\pi133 & w2678 ) ;
  assign w2683 = ( w2680 & w2681 ) | ( w2680 & w2682 ) | ( w2681 & w2682 ) ;
  assign w2684 = \pi134 ^ w2683 ;
  assign w2685 = ( w2677 & w2683 ) | ( w2677 & ~w2684 ) | ( w2683 & ~w2684 ) ;
  assign w2686 = \pi133 ^ w1338 ;
  assign w2687 = ( w1338 & w1359 ) | ( w1338 & ~w2686 ) | ( w1359 & ~w2686 ) ;
  assign w2688 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2687 ) | ( \pi133 & w2687 ) ;
  assign w2689 = w1373 | w2688 ;
  assign w2690 = w1380 & w2688 ;
  assign w2691 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2687 ) | ( ~\pi133 & w2687 ) ;
  assign w2692 = ( w2689 & w2690 ) | ( w2689 & w2691 ) | ( w2690 & w2691 ) ;
  assign w2693 = ( w1324 & w1331 ) | ( w1324 & ~w2201 ) | ( w1331 & ~w2201 ) ;
  assign w2694 = ( \pi132 & \pi133 ) | ( \pi132 & w2693 ) | ( \pi133 & w2693 ) ;
  assign w2695 = w1345 | w2694 ;
  assign w2696 = w1366 & w2694 ;
  assign w2697 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2693 ) | ( \pi133 & ~w2693 ) ;
  assign w2698 = ( w2695 & w2696 ) | ( w2695 & ~w2697 ) | ( w2696 & ~w2697 ) ;
  assign w2699 = \pi134 ^ w2698 ;
  assign w2700 = ( w2692 & w2698 ) | ( w2692 & ~w2699 ) | ( w2698 & ~w2699 ) ;
  assign w2701 = \pi133 ^ w1410 ;
  assign w2702 = ( w1410 & w1431 ) | ( w1410 & ~w2701 ) | ( w1431 & ~w2701 ) ;
  assign w2703 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2702 ) | ( \pi133 & w2702 ) ;
  assign w2704 = w1445 | w2703 ;
  assign w2705 = w1452 & w2703 ;
  assign w2706 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2702 ) | ( ~\pi133 & w2702 ) ;
  assign w2707 = ( w2704 & w2705 ) | ( w2704 & w2706 ) | ( w2705 & w2706 ) ;
  assign w2708 = ( w1396 & w1403 ) | ( w1396 & ~w2217 ) | ( w1403 & ~w2217 ) ;
  assign w2709 = ( \pi132 & \pi133 ) | ( \pi132 & w2708 ) | ( \pi133 & w2708 ) ;
  assign w2710 = w1417 | w2709 ;
  assign w2711 = w1438 & w2709 ;
  assign w2712 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2708 ) | ( \pi133 & ~w2708 ) ;
  assign w2713 = ( w2710 & w2711 ) | ( w2710 & ~w2712 ) | ( w2711 & ~w2712 ) ;
  assign w2714 = \pi134 ^ w2713 ;
  assign w2715 = ( w2707 & w2713 ) | ( w2707 & ~w2714 ) | ( w2713 & ~w2714 ) ;
  assign w2716 = \pi133 ^ w1482 ;
  assign w2717 = ( w1482 & w1503 ) | ( w1482 & ~w2716 ) | ( w1503 & ~w2716 ) ;
  assign w2718 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2717 ) | ( \pi133 & w2717 ) ;
  assign w2719 = w1517 | w2718 ;
  assign w2720 = w1524 & w2718 ;
  assign w2721 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2717 ) | ( ~\pi133 & w2717 ) ;
  assign w2722 = ( w2719 & w2720 ) | ( w2719 & w2721 ) | ( w2720 & w2721 ) ;
  assign w2723 = ( w1468 & w1475 ) | ( w1468 & ~w2233 ) | ( w1475 & ~w2233 ) ;
  assign w2724 = ( \pi132 & \pi133 ) | ( \pi132 & w2723 ) | ( \pi133 & w2723 ) ;
  assign w2725 = w1489 | w2724 ;
  assign w2726 = w1510 & w2724 ;
  assign w2727 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2723 ) | ( \pi133 & ~w2723 ) ;
  assign w2728 = ( w2725 & w2726 ) | ( w2725 & ~w2727 ) | ( w2726 & ~w2727 ) ;
  assign w2729 = \pi134 ^ w2728 ;
  assign w2730 = ( w2722 & w2728 ) | ( w2722 & ~w2729 ) | ( w2728 & ~w2729 ) ;
  assign w2731 = \pi133 ^ w1554 ;
  assign w2732 = ( w1554 & w1575 ) | ( w1554 & ~w2731 ) | ( w1575 & ~w2731 ) ;
  assign w2733 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2732 ) | ( \pi133 & w2732 ) ;
  assign w2734 = w1589 | w2733 ;
  assign w2735 = w1596 & w2733 ;
  assign w2736 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2732 ) | ( ~\pi133 & w2732 ) ;
  assign w2737 = ( w2734 & w2735 ) | ( w2734 & w2736 ) | ( w2735 & w2736 ) ;
  assign w2738 = ( w1540 & w1547 ) | ( w1540 & ~w2249 ) | ( w1547 & ~w2249 ) ;
  assign w2739 = ( \pi132 & \pi133 ) | ( \pi132 & w2738 ) | ( \pi133 & w2738 ) ;
  assign w2740 = w1561 | w2739 ;
  assign w2741 = w1582 & w2739 ;
  assign w2742 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2738 ) | ( \pi133 & ~w2738 ) ;
  assign w2743 = ( w2740 & w2741 ) | ( w2740 & ~w2742 ) | ( w2741 & ~w2742 ) ;
  assign w2744 = \pi134 ^ w2743 ;
  assign w2745 = ( w2737 & w2743 ) | ( w2737 & ~w2744 ) | ( w2743 & ~w2744 ) ;
  assign w2746 = \pi133 ^ w1623 ;
  assign w2747 = ( w1623 & w1642 ) | ( w1623 & ~w2746 ) | ( w1642 & ~w2746 ) ;
  assign w2748 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2747 ) | ( \pi133 & w2747 ) ;
  assign w2749 = w1654 | w2748 ;
  assign w2750 = w1660 & w2748 ;
  assign w2751 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2747 ) | ( ~\pi133 & w2747 ) ;
  assign w2752 = ( w2749 & w2750 ) | ( w2749 & w2751 ) | ( w2750 & w2751 ) ;
  assign w2753 = ( w1611 & w1617 ) | ( w1611 & ~w2265 ) | ( w1617 & ~w2265 ) ;
  assign w2754 = ( \pi132 & \pi133 ) | ( \pi132 & w2753 ) | ( \pi133 & w2753 ) ;
  assign w2755 = w1629 | w2754 ;
  assign w2756 = w1648 & w2754 ;
  assign w2757 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2753 ) | ( \pi133 & ~w2753 ) ;
  assign w2758 = ( w2755 & w2756 ) | ( w2755 & ~w2757 ) | ( w2756 & ~w2757 ) ;
  assign w2759 = \pi134 ^ w2758 ;
  assign w2760 = ( w2752 & w2758 ) | ( w2752 & ~w2759 ) | ( w2758 & ~w2759 ) ;
  assign w2761 = \pi133 ^ w1687 ;
  assign w2762 = ( w1687 & w1706 ) | ( w1687 & ~w2761 ) | ( w1706 & ~w2761 ) ;
  assign w2763 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2762 ) | ( \pi133 & w2762 ) ;
  assign w2764 = w1718 | w2763 ;
  assign w2765 = w1724 & w2763 ;
  assign w2766 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2762 ) | ( ~\pi133 & w2762 ) ;
  assign w2767 = ( w2764 & w2765 ) | ( w2764 & w2766 ) | ( w2765 & w2766 ) ;
  assign w2768 = ( w1675 & w1681 ) | ( w1675 & ~w2281 ) | ( w1681 & ~w2281 ) ;
  assign w2769 = ( \pi132 & \pi133 ) | ( \pi132 & w2768 ) | ( \pi133 & w2768 ) ;
  assign w2770 = w1693 | w2769 ;
  assign w2771 = w1712 & w2769 ;
  assign w2772 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2768 ) | ( \pi133 & ~w2768 ) ;
  assign w2773 = ( w2770 & w2771 ) | ( w2770 & ~w2772 ) | ( w2771 & ~w2772 ) ;
  assign w2774 = \pi134 ^ w2773 ;
  assign w2775 = ( w2767 & w2773 ) | ( w2767 & ~w2774 ) | ( w2773 & ~w2774 ) ;
  assign w2776 = \pi133 ^ w1751 ;
  assign w2777 = ( w1751 & w1770 ) | ( w1751 & ~w2776 ) | ( w1770 & ~w2776 ) ;
  assign w2778 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2777 ) | ( \pi133 & w2777 ) ;
  assign w2779 = w1782 | w2778 ;
  assign w2780 = w1788 & w2778 ;
  assign w2781 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2777 ) | ( ~\pi133 & w2777 ) ;
  assign w2782 = ( w2779 & w2780 ) | ( w2779 & w2781 ) | ( w2780 & w2781 ) ;
  assign w2783 = ( w1739 & w1745 ) | ( w1739 & ~w2297 ) | ( w1745 & ~w2297 ) ;
  assign w2784 = ( \pi132 & \pi133 ) | ( \pi132 & w2783 ) | ( \pi133 & w2783 ) ;
  assign w2785 = w1757 | w2784 ;
  assign w2786 = w1776 & w2784 ;
  assign w2787 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2783 ) | ( \pi133 & ~w2783 ) ;
  assign w2788 = ( w2785 & w2786 ) | ( w2785 & ~w2787 ) | ( w2786 & ~w2787 ) ;
  assign w2789 = \pi134 ^ w2788 ;
  assign w2790 = ( w2782 & w2788 ) | ( w2782 & ~w2789 ) | ( w2788 & ~w2789 ) ;
  assign w2791 = \pi133 ^ w1815 ;
  assign w2792 = ( w1815 & w1834 ) | ( w1815 & ~w2791 ) | ( w1834 & ~w2791 ) ;
  assign w2793 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2792 ) | ( \pi133 & w2792 ) ;
  assign w2794 = w1846 | w2793 ;
  assign w2795 = w1852 & w2793 ;
  assign w2796 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2792 ) | ( ~\pi133 & w2792 ) ;
  assign w2797 = ( w2794 & w2795 ) | ( w2794 & w2796 ) | ( w2795 & w2796 ) ;
  assign w2798 = ( w1803 & w1809 ) | ( w1803 & ~w2313 ) | ( w1809 & ~w2313 ) ;
  assign w2799 = ( \pi132 & \pi133 ) | ( \pi132 & w2798 ) | ( \pi133 & w2798 ) ;
  assign w2800 = w1821 | w2799 ;
  assign w2801 = w1840 & w2799 ;
  assign w2802 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2798 ) | ( \pi133 & ~w2798 ) ;
  assign w2803 = ( w2800 & w2801 ) | ( w2800 & ~w2802 ) | ( w2801 & ~w2802 ) ;
  assign w2804 = \pi134 ^ w2803 ;
  assign w2805 = ( w2797 & w2803 ) | ( w2797 & ~w2804 ) | ( w2803 & ~w2804 ) ;
  assign w2806 = \pi133 ^ w1879 ;
  assign w2807 = ( w1879 & w1900 ) | ( w1879 & ~w2806 ) | ( w1900 & ~w2806 ) ;
  assign w2808 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2807 ) | ( \pi133 & w2807 ) ;
  assign w2809 = w1913 | w2808 ;
  assign w2810 = w1919 & w2808 ;
  assign w2811 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2807 ) | ( ~\pi133 & w2807 ) ;
  assign w2812 = ( w2809 & w2810 ) | ( w2809 & w2811 ) | ( w2810 & w2811 ) ;
  assign w2813 = ( w1867 & w1873 ) | ( w1867 & ~w2329 ) | ( w1873 & ~w2329 ) ;
  assign w2814 = ( \pi132 & \pi133 ) | ( \pi132 & w2813 ) | ( \pi133 & w2813 ) ;
  assign w2815 = w1886 | w2814 ;
  assign w2816 = w1907 & w2814 ;
  assign w2817 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2813 ) | ( \pi133 & ~w2813 ) ;
  assign w2818 = ( w2815 & w2816 ) | ( w2815 & ~w2817 ) | ( w2816 & ~w2817 ) ;
  assign w2819 = \pi134 ^ w2818 ;
  assign w2820 = ( w2812 & w2818 ) | ( w2812 & ~w2819 ) | ( w2818 & ~w2819 ) ;
  assign w2821 = \pi133 ^ w1946 ;
  assign w2822 = ( w1946 & w1967 ) | ( w1946 & ~w2821 ) | ( w1967 & ~w2821 ) ;
  assign w2823 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2822 ) | ( \pi133 & w2822 ) ;
  assign w2824 = w1981 | w2823 ;
  assign w2825 = w1987 & w2823 ;
  assign w2826 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2822 ) | ( ~\pi133 & w2822 ) ;
  assign w2827 = ( w2824 & w2825 ) | ( w2824 & w2826 ) | ( w2825 & w2826 ) ;
  assign w2828 = ( w1934 & w1940 ) | ( w1934 & ~w2345 ) | ( w1940 & ~w2345 ) ;
  assign w2829 = ( \pi132 & \pi133 ) | ( \pi132 & w2828 ) | ( \pi133 & w2828 ) ;
  assign w2830 = w1953 | w2829 ;
  assign w2831 = w1974 & w2829 ;
  assign w2832 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2828 ) | ( \pi133 & ~w2828 ) ;
  assign w2833 = ( w2830 & w2831 ) | ( w2830 & ~w2832 ) | ( w2831 & ~w2832 ) ;
  assign w2834 = \pi134 ^ w2833 ;
  assign w2835 = ( w2827 & w2833 ) | ( w2827 & ~w2834 ) | ( w2833 & ~w2834 ) ;
  assign w2836 = \pi133 ^ w2014 ;
  assign w2837 = ( w2014 & w2035 ) | ( w2014 & ~w2836 ) | ( w2035 & ~w2836 ) ;
  assign w2838 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2837 ) | ( \pi133 & w2837 ) ;
  assign w2839 = w2049 | w2838 ;
  assign w2840 = w2055 & w2838 ;
  assign w2841 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2837 ) | ( ~\pi133 & w2837 ) ;
  assign w2842 = ( w2839 & w2840 ) | ( w2839 & w2841 ) | ( w2840 & w2841 ) ;
  assign w2843 = ( w2002 & w2008 ) | ( w2002 & ~w2361 ) | ( w2008 & ~w2361 ) ;
  assign w2844 = ( \pi132 & \pi133 ) | ( \pi132 & w2843 ) | ( \pi133 & w2843 ) ;
  assign w2845 = w2021 | w2844 ;
  assign w2846 = w2042 & w2844 ;
  assign w2847 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2843 ) | ( \pi133 & ~w2843 ) ;
  assign w2848 = ( w2845 & w2846 ) | ( w2845 & ~w2847 ) | ( w2846 & ~w2847 ) ;
  assign w2849 = \pi134 ^ w2848 ;
  assign w2850 = ( w2842 & w2848 ) | ( w2842 & ~w2849 ) | ( w2848 & ~w2849 ) ;
  assign w2851 = \pi133 ^ w2084 ;
  assign w2852 = ( w2084 & w2104 ) | ( w2084 & ~w2851 ) | ( w2104 & ~w2851 ) ;
  assign w2853 = ( ~\pi132 & \pi133 ) | ( ~\pi132 & w2852 ) | ( \pi133 & w2852 ) ;
  assign w2854 = w2118 | w2853 ;
  assign w2855 = w2124 & w2853 ;
  assign w2856 = ( \pi132 & ~\pi133 ) | ( \pi132 & w2852 ) | ( ~\pi133 & w2852 ) ;
  assign w2857 = ( w2854 & w2855 ) | ( w2854 & w2856 ) | ( w2855 & w2856 ) ;
  assign w2858 = ( w2071 & w2078 ) | ( w2071 & ~w2377 ) | ( w2078 & ~w2377 ) ;
  assign w2859 = ( \pi132 & \pi133 ) | ( \pi132 & w2858 ) | ( \pi133 & w2858 ) ;
  assign w2860 = w2090 | w2859 ;
  assign w2861 = w2111 & w2859 ;
  assign w2862 = ( \pi132 & \pi133 ) | ( \pi132 & ~w2858 ) | ( \pi133 & ~w2858 ) ;
  assign w2863 = ( w2860 & w2861 ) | ( w2860 & ~w2862 ) | ( w2861 & ~w2862 ) ;
  assign w2864 = \pi134 ^ w2863 ;
  assign w2865 = ( w2857 & w2863 ) | ( w2857 & ~w2864 ) | ( w2863 & ~w2864 ) ;
  assign w2866 = \pi134 ^ w282 ;
  assign w2867 = ( w282 & w429 ) | ( w282 & ~w2866 ) | ( w429 & ~w2866 ) ;
  assign w2868 = \pi134 ^ w578 ;
  assign w2869 = ( w578 & w725 ) | ( w578 & ~w2868 ) | ( w725 & ~w2868 ) ;
  assign w2870 = \pi134 ^ w873 ;
  assign w2871 = ( w873 & w1020 ) | ( w873 & ~w2870 ) | ( w1020 & ~w2870 ) ;
  assign w2872 = \pi134 ^ w1168 ;
  assign w2873 = ( w1168 & w1315 ) | ( w1168 & ~w2872 ) | ( w1315 & ~w2872 ) ;
  assign w2874 = \pi134 ^ w1352 ;
  assign w2875 = ( w1352 & w1387 ) | ( w1352 & ~w2874 ) | ( w1387 & ~w2874 ) ;
  assign w2876 = \pi134 ^ w1424 ;
  assign w2877 = ( w1424 & w1459 ) | ( w1424 & ~w2876 ) | ( w1459 & ~w2876 ) ;
  assign w2878 = \pi134 ^ w1496 ;
  assign w2879 = ( w1496 & w1531 ) | ( w1496 & ~w2878 ) | ( w1531 & ~w2878 ) ;
  assign w2880 = \pi134 ^ w1568 ;
  assign w2881 = ( w1568 & w1603 ) | ( w1568 & ~w2880 ) | ( w1603 & ~w2880 ) ;
  assign w2882 = \pi134 ^ w1636 ;
  assign w2883 = ( w1636 & w1667 ) | ( w1636 & ~w2882 ) | ( w1667 & ~w2882 ) ;
  assign w2884 = \pi134 ^ w1700 ;
  assign w2885 = ( w1700 & w1731 ) | ( w1700 & ~w2884 ) | ( w1731 & ~w2884 ) ;
  assign w2886 = \pi134 ^ w1764 ;
  assign w2887 = ( w1764 & w1795 ) | ( w1764 & ~w2886 ) | ( w1795 & ~w2886 ) ;
  assign w2888 = \pi134 ^ w1828 ;
  assign w2889 = ( w1828 & w1859 ) | ( w1828 & ~w2888 ) | ( w1859 & ~w2888 ) ;
  assign w2890 = \pi134 ^ w1893 ;
  assign w2891 = ( w1893 & w1926 ) | ( w1893 & ~w2890 ) | ( w1926 & ~w2890 ) ;
  assign w2892 = \pi134 ^ w1960 ;
  assign w2893 = ( w1960 & w1994 ) | ( w1960 & ~w2892 ) | ( w1994 & ~w2892 ) ;
  assign w2894 = \pi134 ^ w2028 ;
  assign w2895 = ( w2028 & w2062 ) | ( w2028 & ~w2894 ) | ( w2062 & ~w2894 ) ;
  assign w2896 = \pi134 ^ w2097 ;
  assign w2897 = ( w2097 & w2131 ) | ( w2097 & ~w2896 ) | ( w2131 & ~w2896 ) ;
  assign w2898 = \pi134 ^ w2140 ;
  assign w2899 = ( w2140 & w2146 ) | ( w2140 & ~w2898 ) | ( w2146 & ~w2898 ) ;
  assign w2900 = \pi134 ^ w2155 ;
  assign w2901 = ( w2155 & w2161 ) | ( w2155 & ~w2900 ) | ( w2161 & ~w2900 ) ;
  assign w2902 = \pi134 ^ w2170 ;
  assign w2903 = ( w2170 & w2176 ) | ( w2170 & ~w2902 ) | ( w2176 & ~w2902 ) ;
  assign w2904 = \pi134 ^ w2184 ;
  assign w2905 = ( w2184 & w2191 ) | ( w2184 & ~w2904 ) | ( w2191 & ~w2904 ) ;
  assign w2906 = \pi134 ^ w2200 ;
  assign w2907 = ( w2200 & w2207 ) | ( w2200 & ~w2906 ) | ( w2207 & ~w2906 ) ;
  assign w2908 = \pi134 ^ w2216 ;
  assign w2909 = ( w2216 & w2223 ) | ( w2216 & ~w2908 ) | ( w2223 & ~w2908 ) ;
  assign w2910 = \pi134 ^ w2232 ;
  assign w2911 = ( w2232 & w2239 ) | ( w2232 & ~w2910 ) | ( w2239 & ~w2910 ) ;
  assign w2912 = \pi134 ^ w2248 ;
  assign w2913 = ( w2248 & w2255 ) | ( w2248 & ~w2912 ) | ( w2255 & ~w2912 ) ;
  assign w2914 = \pi134 ^ w2264 ;
  assign w2915 = ( w2264 & w2271 ) | ( w2264 & ~w2914 ) | ( w2271 & ~w2914 ) ;
  assign w2916 = \pi134 ^ w2280 ;
  assign w2917 = ( w2280 & w2287 ) | ( w2280 & ~w2916 ) | ( w2287 & ~w2916 ) ;
  assign w2918 = \pi134 ^ w2296 ;
  assign w2919 = ( w2296 & w2303 ) | ( w2296 & ~w2918 ) | ( w2303 & ~w2918 ) ;
  assign w2920 = \pi134 ^ w2312 ;
  assign w2921 = ( w2312 & w2319 ) | ( w2312 & ~w2920 ) | ( w2319 & ~w2920 ) ;
  assign w2922 = \pi134 ^ w2328 ;
  assign w2923 = ( w2328 & w2335 ) | ( w2328 & ~w2922 ) | ( w2335 & ~w2922 ) ;
  assign w2924 = \pi134 ^ w2344 ;
  assign w2925 = ( w2344 & w2351 ) | ( w2344 & ~w2924 ) | ( w2351 & ~w2924 ) ;
  assign w2926 = \pi134 ^ w2360 ;
  assign w2927 = ( w2360 & w2367 ) | ( w2360 & ~w2926 ) | ( w2367 & ~w2926 ) ;
  assign w2928 = \pi134 ^ w2376 ;
  assign w2929 = ( w2376 & w2383 ) | ( w2376 & ~w2928 ) | ( w2383 & ~w2928 ) ;
  assign w2930 = \pi134 ^ w2392 ;
  assign w2931 = ( w2392 & w2398 ) | ( w2392 & ~w2930 ) | ( w2398 & ~w2930 ) ;
  assign w2932 = \pi134 ^ w2407 ;
  assign w2933 = ( w2407 & w2413 ) | ( w2407 & ~w2932 ) | ( w2413 & ~w2932 ) ;
  assign w2934 = \pi134 ^ w2422 ;
  assign w2935 = ( w2422 & w2428 ) | ( w2422 & ~w2934 ) | ( w2428 & ~w2934 ) ;
  assign w2936 = \pi134 ^ w2436 ;
  assign w2937 = ( w2436 & w2443 ) | ( w2436 & ~w2936 ) | ( w2443 & ~w2936 ) ;
  assign w2938 = \pi134 ^ w2452 ;
  assign w2939 = ( w2452 & w2458 ) | ( w2452 & ~w2938 ) | ( w2458 & ~w2938 ) ;
  assign w2940 = \pi134 ^ w2467 ;
  assign w2941 = ( w2467 & w2473 ) | ( w2467 & ~w2940 ) | ( w2473 & ~w2940 ) ;
  assign w2942 = \pi134 ^ w2482 ;
  assign w2943 = ( w2482 & w2488 ) | ( w2482 & ~w2942 ) | ( w2488 & ~w2942 ) ;
  assign w2944 = \pi134 ^ w2497 ;
  assign w2945 = ( w2497 & w2503 ) | ( w2497 & ~w2944 ) | ( w2503 & ~w2944 ) ;
  assign w2946 = \pi134 ^ w2512 ;
  assign w2947 = ( w2512 & w2518 ) | ( w2512 & ~w2946 ) | ( w2518 & ~w2946 ) ;
  assign w2948 = \pi134 ^ w2527 ;
  assign w2949 = ( w2527 & w2533 ) | ( w2527 & ~w2948 ) | ( w2533 & ~w2948 ) ;
  assign w2950 = \pi134 ^ w2542 ;
  assign w2951 = ( w2542 & w2548 ) | ( w2542 & ~w2950 ) | ( w2548 & ~w2950 ) ;
  assign w2952 = \pi134 ^ w2557 ;
  assign w2953 = ( w2557 & w2563 ) | ( w2557 & ~w2952 ) | ( w2563 & ~w2952 ) ;
  assign w2954 = \pi134 ^ w2572 ;
  assign w2955 = ( w2572 & w2578 ) | ( w2572 & ~w2954 ) | ( w2578 & ~w2954 ) ;
  assign w2956 = \pi134 ^ w2587 ;
  assign w2957 = ( w2587 & w2593 ) | ( w2587 & ~w2956 ) | ( w2593 & ~w2956 ) ;
  assign w2958 = \pi134 ^ w2602 ;
  assign w2959 = ( w2602 & w2608 ) | ( w2602 & ~w2958 ) | ( w2608 & ~w2958 ) ;
  assign w2960 = \pi134 ^ w2617 ;
  assign w2961 = ( w2617 & w2623 ) | ( w2617 & ~w2960 ) | ( w2623 & ~w2960 ) ;
  assign w2962 = \pi134 ^ w2631 ;
  assign w2963 = ( w2631 & w2638 ) | ( w2631 & ~w2962 ) | ( w2638 & ~w2962 ) ;
  assign w2964 = \pi134 ^ w2646 ;
  assign w2965 = ( w2646 & w2653 ) | ( w2646 & ~w2964 ) | ( w2653 & ~w2964 ) ;
  assign w2966 = \pi134 ^ w2661 ;
  assign w2967 = ( w2661 & w2668 ) | ( w2661 & ~w2966 ) | ( w2668 & ~w2966 ) ;
  assign w2968 = \pi134 ^ w2677 ;
  assign w2969 = ( w2677 & w2683 ) | ( w2677 & ~w2968 ) | ( w2683 & ~w2968 ) ;
  assign w2970 = \pi134 ^ w2692 ;
  assign w2971 = ( w2692 & w2698 ) | ( w2692 & ~w2970 ) | ( w2698 & ~w2970 ) ;
  assign w2972 = \pi134 ^ w2707 ;
  assign w2973 = ( w2707 & w2713 ) | ( w2707 & ~w2972 ) | ( w2713 & ~w2972 ) ;
  assign w2974 = \pi134 ^ w2722 ;
  assign w2975 = ( w2722 & w2728 ) | ( w2722 & ~w2974 ) | ( w2728 & ~w2974 ) ;
  assign w2976 = \pi134 ^ w2737 ;
  assign w2977 = ( w2737 & w2743 ) | ( w2737 & ~w2976 ) | ( w2743 & ~w2976 ) ;
  assign w2978 = \pi134 ^ w2752 ;
  assign w2979 = ( w2752 & w2758 ) | ( w2752 & ~w2978 ) | ( w2758 & ~w2978 ) ;
  assign w2980 = \pi134 ^ w2767 ;
  assign w2981 = ( w2767 & w2773 ) | ( w2767 & ~w2980 ) | ( w2773 & ~w2980 ) ;
  assign w2982 = \pi134 ^ w2782 ;
  assign w2983 = ( w2782 & w2788 ) | ( w2782 & ~w2982 ) | ( w2788 & ~w2982 ) ;
  assign w2984 = \pi134 ^ w2797 ;
  assign w2985 = ( w2797 & w2803 ) | ( w2797 & ~w2984 ) | ( w2803 & ~w2984 ) ;
  assign w2986 = \pi134 ^ w2812 ;
  assign w2987 = ( w2812 & w2818 ) | ( w2812 & ~w2986 ) | ( w2818 & ~w2986 ) ;
  assign w2988 = \pi134 ^ w2827 ;
  assign w2989 = ( w2827 & w2833 ) | ( w2827 & ~w2988 ) | ( w2833 & ~w2988 ) ;
  assign w2990 = \pi134 ^ w2842 ;
  assign w2991 = ( w2842 & w2848 ) | ( w2842 & ~w2990 ) | ( w2848 & ~w2990 ) ;
  assign w2992 = \pi134 ^ w2857 ;
  assign w2993 = ( w2857 & w2863 ) | ( w2857 & ~w2992 ) | ( w2863 & ~w2992 ) ;
  assign \po000 = w431 ;
  assign \po001 = w727 ;
  assign \po002 = w1022 ;
  assign \po003 = w1317 ;
  assign \po004 = w1389 ;
  assign \po005 = w1461 ;
  assign \po006 = w1533 ;
  assign \po007 = w1605 ;
  assign \po008 = w1669 ;
  assign \po009 = w1733 ;
  assign \po010 = w1797 ;
  assign \po011 = w1861 ;
  assign \po012 = w1928 ;
  assign \po013 = w1996 ;
  assign \po014 = w2064 ;
  assign \po015 = w2133 ;
  assign \po016 = w2148 ;
  assign \po017 = w2163 ;
  assign \po018 = w2178 ;
  assign \po019 = w2193 ;
  assign \po020 = w2209 ;
  assign \po021 = w2225 ;
  assign \po022 = w2241 ;
  assign \po023 = w2257 ;
  assign \po024 = w2273 ;
  assign \po025 = w2289 ;
  assign \po026 = w2305 ;
  assign \po027 = w2321 ;
  assign \po028 = w2337 ;
  assign \po029 = w2353 ;
  assign \po030 = w2369 ;
  assign \po031 = w2385 ;
  assign \po032 = w2400 ;
  assign \po033 = w2415 ;
  assign \po034 = w2430 ;
  assign \po035 = w2445 ;
  assign \po036 = w2460 ;
  assign \po037 = w2475 ;
  assign \po038 = w2490 ;
  assign \po039 = w2505 ;
  assign \po040 = w2520 ;
  assign \po041 = w2535 ;
  assign \po042 = w2550 ;
  assign \po043 = w2565 ;
  assign \po044 = w2580 ;
  assign \po045 = w2595 ;
  assign \po046 = w2610 ;
  assign \po047 = w2625 ;
  assign \po048 = w2640 ;
  assign \po049 = w2655 ;
  assign \po050 = w2670 ;
  assign \po051 = w2685 ;
  assign \po052 = w2700 ;
  assign \po053 = w2715 ;
  assign \po054 = w2730 ;
  assign \po055 = w2745 ;
  assign \po056 = w2760 ;
  assign \po057 = w2775 ;
  assign \po058 = w2790 ;
  assign \po059 = w2805 ;
  assign \po060 = w2820 ;
  assign \po061 = w2835 ;
  assign \po062 = w2850 ;
  assign \po063 = w2865 ;
  assign \po064 = w2867 ;
  assign \po065 = w2869 ;
  assign \po066 = w2871 ;
  assign \po067 = w2873 ;
  assign \po068 = w2875 ;
  assign \po069 = w2877 ;
  assign \po070 = w2879 ;
  assign \po071 = w2881 ;
  assign \po072 = w2883 ;
  assign \po073 = w2885 ;
  assign \po074 = w2887 ;
  assign \po075 = w2889 ;
  assign \po076 = w2891 ;
  assign \po077 = w2893 ;
  assign \po078 = w2895 ;
  assign \po079 = w2897 ;
  assign \po080 = w2899 ;
  assign \po081 = w2901 ;
  assign \po082 = w2903 ;
  assign \po083 = w2905 ;
  assign \po084 = w2907 ;
  assign \po085 = w2909 ;
  assign \po086 = w2911 ;
  assign \po087 = w2913 ;
  assign \po088 = w2915 ;
  assign \po089 = w2917 ;
  assign \po090 = w2919 ;
  assign \po091 = w2921 ;
  assign \po092 = w2923 ;
  assign \po093 = w2925 ;
  assign \po094 = w2927 ;
  assign \po095 = w2929 ;
  assign \po096 = w2931 ;
  assign \po097 = w2933 ;
  assign \po098 = w2935 ;
  assign \po099 = w2937 ;
  assign \po100 = w2939 ;
  assign \po101 = w2941 ;
  assign \po102 = w2943 ;
  assign \po103 = w2945 ;
  assign \po104 = w2947 ;
  assign \po105 = w2949 ;
  assign \po106 = w2951 ;
  assign \po107 = w2953 ;
  assign \po108 = w2955 ;
  assign \po109 = w2957 ;
  assign \po110 = w2959 ;
  assign \po111 = w2961 ;
  assign \po112 = w2963 ;
  assign \po113 = w2965 ;
  assign \po114 = w2967 ;
  assign \po115 = w2969 ;
  assign \po116 = w2971 ;
  assign \po117 = w2973 ;
  assign \po118 = w2975 ;
  assign \po119 = w2977 ;
  assign \po120 = w2979 ;
  assign \po121 = w2981 ;
  assign \po122 = w2983 ;
  assign \po123 = w2985 ;
  assign \po124 = w2987 ;
  assign \po125 = w2989 ;
  assign \po126 = w2991 ;
  assign \po127 = w2993 ;
endmodule
