module max( \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 , \pi135 , \pi136 , \pi137 , \pi138 , \pi139 , \pi140 , \pi141 , \pi142 , \pi143 , \pi144 , \pi145 , \pi146 , \pi147 , \pi148 , \pi149 , \pi150 , \pi151 , \pi152 , \pi153 , \pi154 , \pi155 , \pi156 , \pi157 , \pi158 , \pi159 , \pi160 , \pi161 , \pi162 , \pi163 , \pi164 , \pi165 , \pi166 , \pi167 , \pi168 , \pi169 , \pi170 , \pi171 , \pi172 , \pi173 , \pi174 , \pi175 , \pi176 , \pi177 , \pi178 , \pi179 , \pi180 , \pi181 , \pi182 , \pi183 , \pi184 , \pi185 , \pi186 , \pi187 , \pi188 , \pi189 , \pi190 , \pi191 , \pi192 , \pi193 , \pi194 , \pi195 , \pi196 , \pi197 , \pi198 , \pi199 , \pi200 , \pi201 , \pi202 , \pi203 , \pi204 , \pi205 , \pi206 , \pi207 , \pi208 , \pi209 , \pi210 , \pi211 , \pi212 , \pi213 , \pi214 , \pi215 , \pi216 , \pi217 , \pi218 , \pi219 , \pi220 , \pi221 , \pi222 , \pi223 , \pi224 , \pi225 , \pi226 , \pi227 , \pi228 , \pi229 , \pi230 , \pi231 , \pi232 , \pi233 , \pi234 , \pi235 , \pi236 , \pi237 , \pi238 , \pi239 , \pi240 , \pi241 , \pi242 , \pi243 , \pi244 , \pi245 , \pi246 , \pi247 , \pi248 , \pi249 , \pi250 , \pi251 , \pi252 , \pi253 , \pi254 , \pi255 , \pi256 , \pi257 , \pi258 , \pi259 , \pi260 , \pi261 , \pi262 , \pi263 , \pi264 , \pi265 , \pi266 , \pi267 , \pi268 , \pi269 , \pi270 , \pi271 , \pi272 , \pi273 , \pi274 , \pi275 , \pi276 , \pi277 , \pi278 , \pi279 , \pi280 , \pi281 , \pi282 , \pi283 , \pi284 , \pi285 , \pi286 , \pi287 , \pi288 , \pi289 , \pi290 , \pi291 , \pi292 , \pi293 , \pi294 , \pi295 , \pi296 , \pi297 , \pi298 , \pi299 , \pi300 , \pi301 , \pi302 , \pi303 , \pi304 , \pi305 , \pi306 , \pi307 , \pi308 , \pi309 , \pi310 , \pi311 , \pi312 , \pi313 , \pi314 , \pi315 , \pi316 , \pi317 , \pi318 , \pi319 , \pi320 , \pi321 , \pi322 , \pi323 , \pi324 , \pi325 , \pi326 , \pi327 , \pi328 , \pi329 , \pi330 , \pi331 , \pi332 , \pi333 , \pi334 , \pi335 , \pi336 , \pi337 , \pi338 , \pi339 , \pi340 , \pi341 , \pi342 , \pi343 , \pi344 , \pi345 , \pi346 , \pi347 , \pi348 , \pi349 , \pi350 , \pi351 , \pi352 , \pi353 , \pi354 , \pi355 , \pi356 , \pi357 , \pi358 , \pi359 , \pi360 , \pi361 , \pi362 , \pi363 , \pi364 , \pi365 , \pi366 , \pi367 , \pi368 , \pi369 , \pi370 , \pi371 , \pi372 , \pi373 , \pi374 , \pi375 , \pi376 , \pi377 , \pi378 , \pi379 , \pi380 , \pi381 , \pi382 , \pi383 , \pi384 , \pi385 , \pi386 , \pi387 , \pi388 , \pi389 , \pi390 , \pi391 , \pi392 , \pi393 , \pi394 , \pi395 , \pi396 , \pi397 , \pi398 , \pi399 , \pi400 , \pi401 , \pi402 , \pi403 , \pi404 , \pi405 , \pi406 , \pi407 , \pi408 , \pi409 , \pi410 , \pi411 , \pi412 , \pi413 , \pi414 , \pi415 , \pi416 , \pi417 , \pi418 , \pi419 , \pi420 , \pi421 , \pi422 , \pi423 , \pi424 , \pi425 , \pi426 , \pi427 , \pi428 , \pi429 , \pi430 , \pi431 , \pi432 , \pi433 , \pi434 , \pi435 , \pi436 , \pi437 , \pi438 , \pi439 , \pi440 , \pi441 , \pi442 , \pi443 , \pi444 , \pi445 , \pi446 , \pi447 , \pi448 , \pi449 , \pi450 , \pi451 , \pi452 , \pi453 , \pi454 , \pi455 , \pi456 , \pi457 , \pi458 , \pi459 , \pi460 , \pi461 , \pi462 , \pi463 , \pi464 , \pi465 , \pi466 , \pi467 , \pi468 , \pi469 , \pi470 , \pi471 , \pi472 , \pi473 , \pi474 , \pi475 , \pi476 , \pi477 , \pi478 , \pi479 , \pi480 , \pi481 , \pi482 , \pi483 , \pi484 , \pi485 , \pi486 , \pi487 , \pi488 , \pi489 , \pi490 , \pi491 , \pi492 , \pi493 , \pi494 , \pi495 , \pi496 , \pi497 , \pi498 , \pi499 , \pi500 , \pi501 , \pi502 , \pi503 , \pi504 , \pi505 , \pi506 , \pi507 , \pi508 , \pi509 , \pi510 , \pi511 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 , \po128 , \po129 );
  input \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 , \pi135 , \pi136 , \pi137 , \pi138 , \pi139 , \pi140 , \pi141 , \pi142 , \pi143 , \pi144 , \pi145 , \pi146 , \pi147 , \pi148 , \pi149 , \pi150 , \pi151 , \pi152 , \pi153 , \pi154 , \pi155 , \pi156 , \pi157 , \pi158 , \pi159 , \pi160 , \pi161 , \pi162 , \pi163 , \pi164 , \pi165 , \pi166 , \pi167 , \pi168 , \pi169 , \pi170 , \pi171 , \pi172 , \pi173 , \pi174 , \pi175 , \pi176 , \pi177 , \pi178 , \pi179 , \pi180 , \pi181 , \pi182 , \pi183 , \pi184 , \pi185 , \pi186 , \pi187 , \pi188 , \pi189 , \pi190 , \pi191 , \pi192 , \pi193 , \pi194 , \pi195 , \pi196 , \pi197 , \pi198 , \pi199 , \pi200 , \pi201 , \pi202 , \pi203 , \pi204 , \pi205 , \pi206 , \pi207 , \pi208 , \pi209 , \pi210 , \pi211 , \pi212 , \pi213 , \pi214 , \pi215 , \pi216 , \pi217 , \pi218 , \pi219 , \pi220 , \pi221 , \pi222 , \pi223 , \pi224 , \pi225 , \pi226 , \pi227 , \pi228 , \pi229 , \pi230 , \pi231 , \pi232 , \pi233 , \pi234 , \pi235 , \pi236 , \pi237 , \pi238 , \pi239 , \pi240 , \pi241 , \pi242 , \pi243 , \pi244 , \pi245 , \pi246 , \pi247 , \pi248 , \pi249 , \pi250 , \pi251 , \pi252 , \pi253 , \pi254 , \pi255 , \pi256 , \pi257 , \pi258 , \pi259 , \pi260 , \pi261 , \pi262 , \pi263 , \pi264 , \pi265 , \pi266 , \pi267 , \pi268 , \pi269 , \pi270 , \pi271 , \pi272 , \pi273 , \pi274 , \pi275 , \pi276 , \pi277 , \pi278 , \pi279 , \pi280 , \pi281 , \pi282 , \pi283 , \pi284 , \pi285 , \pi286 , \pi287 , \pi288 , \pi289 , \pi290 , \pi291 , \pi292 , \pi293 , \pi294 , \pi295 , \pi296 , \pi297 , \pi298 , \pi299 , \pi300 , \pi301 , \pi302 , \pi303 , \pi304 , \pi305 , \pi306 , \pi307 , \pi308 , \pi309 , \pi310 , \pi311 , \pi312 , \pi313 , \pi314 , \pi315 , \pi316 , \pi317 , \pi318 , \pi319 , \pi320 , \pi321 , \pi322 , \pi323 , \pi324 , \pi325 , \pi326 , \pi327 , \pi328 , \pi329 , \pi330 , \pi331 , \pi332 , \pi333 , \pi334 , \pi335 , \pi336 , \pi337 , \pi338 , \pi339 , \pi340 , \pi341 , \pi342 , \pi343 , \pi344 , \pi345 , \pi346 , \pi347 , \pi348 , \pi349 , \pi350 , \pi351 , \pi352 , \pi353 , \pi354 , \pi355 , \pi356 , \pi357 , \pi358 , \pi359 , \pi360 , \pi361 , \pi362 , \pi363 , \pi364 , \pi365 , \pi366 , \pi367 , \pi368 , \pi369 , \pi370 , \pi371 , \pi372 , \pi373 , \pi374 , \pi375 , \pi376 , \pi377 , \pi378 , \pi379 , \pi380 , \pi381 , \pi382 , \pi383 , \pi384 , \pi385 , \pi386 , \pi387 , \pi388 , \pi389 , \pi390 , \pi391 , \pi392 , \pi393 , \pi394 , \pi395 , \pi396 , \pi397 , \pi398 , \pi399 , \pi400 , \pi401 , \pi402 , \pi403 , \pi404 , \pi405 , \pi406 , \pi407 , \pi408 , \pi409 , \pi410 , \pi411 , \pi412 , \pi413 , \pi414 , \pi415 , \pi416 , \pi417 , \pi418 , \pi419 , \pi420 , \pi421 , \pi422 , \pi423 , \pi424 , \pi425 , \pi426 , \pi427 , \pi428 , \pi429 , \pi430 , \pi431 , \pi432 , \pi433 , \pi434 , \pi435 , \pi436 , \pi437 , \pi438 , \pi439 , \pi440 , \pi441 , \pi442 , \pi443 , \pi444 , \pi445 , \pi446 , \pi447 , \pi448 , \pi449 , \pi450 , \pi451 , \pi452 , \pi453 , \pi454 , \pi455 , \pi456 , \pi457 , \pi458 , \pi459 , \pi460 , \pi461 , \pi462 , \pi463 , \pi464 , \pi465 , \pi466 , \pi467 , \pi468 , \pi469 , \pi470 , \pi471 , \pi472 , \pi473 , \pi474 , \pi475 , \pi476 , \pi477 , \pi478 , \pi479 , \pi480 , \pi481 , \pi482 , \pi483 , \pi484 , \pi485 , \pi486 , \pi487 , \pi488 , \pi489 , \pi490 , \pi491 , \pi492 , \pi493 , \pi494 , \pi495 , \pi496 , \pi497 , \pi498 , \pi499 , \pi500 , \pi501 , \pi502 , \pi503 , \pi504 , \pi505 , \pi506 , \pi507 , \pi508 , \pi509 , \pi510 , \pi511 ;
  output \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 , \po128 , \po129 ;
  wire zero , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 ;
  assign zero = 0;
  assign w513 = \pi374 | \pi502 ;
  assign w514 = ~\pi375 & \pi503 ;
  assign w515 = ( ~\pi374 & w513 ) | ( ~\pi374 & w514 ) | ( w513 & w514 ) ;
  assign w516 = \pi372 & ~\pi500 ;
  assign w517 = ( \pi373 & ~\pi501 ) | ( \pi373 & w516 ) | ( ~\pi501 & w516 ) ;
  assign w518 = \pi366 | \pi494 ;
  assign w519 = ~\pi367 & \pi495 ;
  assign w520 = ( ~\pi366 & w518 ) | ( ~\pi366 & w519 ) | ( w518 & w519 ) ;
  assign w521 = \pi358 | \pi486 ;
  assign w522 = ~\pi359 & \pi487 ;
  assign w523 = ( ~\pi358 & w521 ) | ( ~\pi358 & w522 ) | ( w521 & w522 ) ;
  assign w524 = \pi356 & ~\pi484 ;
  assign w525 = ( \pi357 & ~\pi485 ) | ( \pi357 & w524 ) | ( ~\pi485 & w524 ) ;
  assign w526 = \pi350 | \pi478 ;
  assign w527 = ~\pi351 & \pi479 ;
  assign w528 = ( ~\pi350 & w526 ) | ( ~\pi350 & w527 ) | ( w526 & w527 ) ;
  assign w529 = \pi342 | \pi470 ;
  assign w530 = ~\pi343 & \pi471 ;
  assign w531 = ( ~\pi342 & w529 ) | ( ~\pi342 & w530 ) | ( w529 & w530 ) ;
  assign w532 = \pi340 & ~\pi468 ;
  assign w533 = ( \pi341 & ~\pi469 ) | ( \pi341 & w532 ) | ( ~\pi469 & w532 ) ;
  assign w534 = \pi334 | \pi462 ;
  assign w535 = ~\pi335 & \pi463 ;
  assign w536 = ( ~\pi334 & w534 ) | ( ~\pi334 & w535 ) | ( w534 & w535 ) ;
  assign w537 = \pi326 | \pi454 ;
  assign w538 = ~\pi327 & \pi455 ;
  assign w539 = ( ~\pi326 & w537 ) | ( ~\pi326 & w538 ) | ( w537 & w538 ) ;
  assign w540 = \pi324 & ~\pi452 ;
  assign w541 = ( \pi325 & ~\pi453 ) | ( \pi325 & w540 ) | ( ~\pi453 & w540 ) ;
  assign w542 = \pi318 | \pi446 ;
  assign w543 = ~\pi319 & \pi447 ;
  assign w544 = ( ~\pi318 & w542 ) | ( ~\pi318 & w543 ) | ( w542 & w543 ) ;
  assign w545 = \pi316 & \pi444 ;
  assign w546 = \pi317 & \pi445 ;
  assign w547 = ( \pi445 & w544 ) | ( \pi445 & ~w546 ) | ( w544 & ~w546 ) ;
  assign w548 = ( \pi444 & ~w545 ) | ( \pi444 & w547 ) | ( ~w545 & w547 ) ;
  assign w549 = \pi312 & ~\pi440 ;
  assign w550 = ( \pi313 & ~\pi441 ) | ( \pi313 & w549 ) | ( ~\pi441 & w549 ) ;
  assign w551 = \pi315 & ~w548 ;
  assign w552 = ( \pi314 & ~\pi442 ) | ( \pi314 & w550 ) | ( ~\pi442 & w550 ) ;
  assign w553 = \pi443 | w548 ;
  assign w554 = ( w551 & w552 ) | ( w551 & ~w553 ) | ( w552 & ~w553 ) ;
  assign w555 = \pi316 & ~\pi444 ;
  assign w556 = ( \pi317 & ~\pi445 ) | ( \pi317 & w555 ) | ( ~\pi445 & w555 ) ;
  assign w557 = \pi303 & ~\pi431 ;
  assign w558 = \pi302 | \pi430 ;
  assign w559 = ~\pi303 & \pi431 ;
  assign w560 = ( ~\pi302 & w558 ) | ( ~\pi302 & w559 ) | ( w558 & w559 ) ;
  assign w561 = \pi300 & \pi428 ;
  assign w562 = \pi301 & \pi429 ;
  assign w563 = ( \pi429 & w560 ) | ( \pi429 & ~w562 ) | ( w560 & ~w562 ) ;
  assign w564 = ( \pi428 & ~w561 ) | ( \pi428 & w563 ) | ( ~w561 & w563 ) ;
  assign w565 = \pi298 | \pi426 ;
  assign w566 = ~\pi299 & \pi427 ;
  assign w567 = ( ~\pi298 & w565 ) | ( ~\pi298 & w566 ) | ( w565 & w566 ) ;
  assign w568 = \pi296 & ~\pi424 ;
  assign w569 = ( \pi297 & ~\pi425 ) | ( \pi297 & w568 ) | ( ~\pi425 & w568 ) ;
  assign w570 = \pi299 & ~w564 ;
  assign w571 = ( \pi298 & ~\pi426 ) | ( \pi298 & w569 ) | ( ~\pi426 & w569 ) ;
  assign w572 = \pi427 | w564 ;
  assign w573 = ( w570 & w571 ) | ( w570 & ~w572 ) | ( w571 & ~w572 ) ;
  assign w574 = \pi300 & ~\pi428 ;
  assign w575 = ( \pi301 & ~\pi429 ) | ( \pi301 & w574 ) | ( ~\pi429 & w574 ) ;
  assign w576 = \pi256 & ~\pi384 ;
  assign w577 = ( \pi257 & ~\pi385 ) | ( \pi257 & w576 ) | ( ~\pi385 & w576 ) ;
  assign w578 = ( \pi258 & ~\pi386 ) | ( \pi258 & w577 ) | ( ~\pi386 & w577 ) ;
  assign w579 = ( \pi259 & ~\pi387 ) | ( \pi259 & w578 ) | ( ~\pi387 & w578 ) ;
  assign w580 = ( \pi260 & ~\pi388 ) | ( \pi260 & w579 ) | ( ~\pi388 & w579 ) ;
  assign w581 = ( \pi261 & ~\pi389 ) | ( \pi261 & w580 ) | ( ~\pi389 & w580 ) ;
  assign w582 = ( \pi262 & ~\pi390 ) | ( \pi262 & w581 ) | ( ~\pi390 & w581 ) ;
  assign w583 = ( \pi263 & ~\pi391 ) | ( \pi263 & w582 ) | ( ~\pi391 & w582 ) ;
  assign w584 = ( \pi264 & ~\pi392 ) | ( \pi264 & w583 ) | ( ~\pi392 & w583 ) ;
  assign w585 = ( \pi265 & ~\pi393 ) | ( \pi265 & w584 ) | ( ~\pi393 & w584 ) ;
  assign w586 = ( \pi266 & ~\pi394 ) | ( \pi266 & w585 ) | ( ~\pi394 & w585 ) ;
  assign w587 = ( \pi267 & ~\pi395 ) | ( \pi267 & w586 ) | ( ~\pi395 & w586 ) ;
  assign w588 = ( \pi268 & ~\pi396 ) | ( \pi268 & w587 ) | ( ~\pi396 & w587 ) ;
  assign w589 = ( \pi269 & ~\pi397 ) | ( \pi269 & w588 ) | ( ~\pi397 & w588 ) ;
  assign w590 = ( \pi270 & ~\pi398 ) | ( \pi270 & w589 ) | ( ~\pi398 & w589 ) ;
  assign w591 = ( \pi271 & ~\pi399 ) | ( \pi271 & w590 ) | ( ~\pi399 & w590 ) ;
  assign w592 = ( \pi272 & ~\pi400 ) | ( \pi272 & w591 ) | ( ~\pi400 & w591 ) ;
  assign w593 = ( \pi273 & ~\pi401 ) | ( \pi273 & w592 ) | ( ~\pi401 & w592 ) ;
  assign w594 = ( \pi274 & ~\pi402 ) | ( \pi274 & w593 ) | ( ~\pi402 & w593 ) ;
  assign w595 = ( \pi275 & ~\pi403 ) | ( \pi275 & w594 ) | ( ~\pi403 & w594 ) ;
  assign w596 = ( \pi276 & ~\pi404 ) | ( \pi276 & w595 ) | ( ~\pi404 & w595 ) ;
  assign w597 = ( \pi277 & ~\pi405 ) | ( \pi277 & w596 ) | ( ~\pi405 & w596 ) ;
  assign w598 = ( \pi278 & ~\pi406 ) | ( \pi278 & w597 ) | ( ~\pi406 & w597 ) ;
  assign w599 = ( \pi279 & ~\pi407 ) | ( \pi279 & w598 ) | ( ~\pi407 & w598 ) ;
  assign w600 = ( \pi280 & ~\pi408 ) | ( \pi280 & w599 ) | ( ~\pi408 & w599 ) ;
  assign w601 = ( \pi281 & ~\pi409 ) | ( \pi281 & w600 ) | ( ~\pi409 & w600 ) ;
  assign w602 = ( \pi282 & ~\pi410 ) | ( \pi282 & w601 ) | ( ~\pi410 & w601 ) ;
  assign w603 = ( \pi283 & ~\pi411 ) | ( \pi283 & w602 ) | ( ~\pi411 & w602 ) ;
  assign w604 = ( \pi284 & ~\pi412 ) | ( \pi284 & w603 ) | ( ~\pi412 & w603 ) ;
  assign w605 = ( \pi285 & ~\pi413 ) | ( \pi285 & w604 ) | ( ~\pi413 & w604 ) ;
  assign w606 = ( \pi286 & ~\pi414 ) | ( \pi286 & w605 ) | ( ~\pi414 & w605 ) ;
  assign w607 = ( \pi287 & ~\pi415 ) | ( \pi287 & w606 ) | ( ~\pi415 & w606 ) ;
  assign w608 = \pi294 | \pi422 ;
  assign w609 = ~\pi295 & \pi423 ;
  assign w610 = ( ~\pi294 & w608 ) | ( ~\pi294 & w609 ) | ( w608 & w609 ) ;
  assign w611 = \pi292 & \pi420 ;
  assign w612 = \pi293 & \pi421 ;
  assign w613 = ( \pi421 & w610 ) | ( \pi421 & ~w612 ) | ( w610 & ~w612 ) ;
  assign w614 = ( \pi420 & ~w611 ) | ( \pi420 & w613 ) | ( ~w611 & w613 ) ;
  assign w615 = \pi290 | \pi418 ;
  assign w616 = ~\pi291 & \pi419 ;
  assign w617 = ( ~\pi290 & w615 ) | ( ~\pi290 & w616 ) | ( w615 & w616 ) ;
  assign w618 = w607 & ~w614 ;
  assign w619 = ( \pi289 & ~\pi417 ) | ( \pi289 & w618 ) | ( ~\pi417 & w618 ) ;
  assign w620 = ( w617 & w618 ) | ( w617 & ~w619 ) | ( w618 & ~w619 ) ;
  assign w621 = w618 & ~w620 ;
  assign w622 = \pi292 & ~\pi420 ;
  assign w623 = ( \pi293 & ~\pi421 ) | ( \pi293 & w622 ) | ( ~\pi421 & w622 ) ;
  assign w624 = \pi288 & ~\pi416 ;
  assign w625 = ( \pi289 & ~\pi417 ) | ( \pi289 & w624 ) | ( ~\pi417 & w624 ) ;
  assign w626 = \pi291 & ~w614 ;
  assign w627 = ( \pi290 & ~\pi418 ) | ( \pi290 & w625 ) | ( ~\pi418 & w625 ) ;
  assign w628 = \pi419 | w614 ;
  assign w629 = ( w626 & w627 ) | ( w626 & ~w628 ) | ( w627 & ~w628 ) ;
  assign w630 = \pi295 | w629 ;
  assign w631 = ( \pi294 & ~\pi422 ) | ( \pi294 & w623 ) | ( ~\pi422 & w623 ) ;
  assign w632 = \pi423 & ~w629 ;
  assign w633 = ( w630 & w631 ) | ( w630 & ~w632 ) | ( w631 & ~w632 ) ;
  assign w634 = \pi296 & \pi424 ;
  assign w635 = \pi297 & \pi425 ;
  assign w636 = ( \pi425 & w567 ) | ( \pi425 & ~w635 ) | ( w567 & ~w635 ) ;
  assign w637 = ( \pi424 & ~w634 ) | ( \pi424 & w636 ) | ( ~w634 & w636 ) ;
  assign w638 = ( ~w564 & w633 ) | ( ~w564 & w637 ) | ( w633 & w637 ) ;
  assign w639 = ( \pi288 & \pi416 ) | ( \pi288 & w638 ) | ( \pi416 & w638 ) ;
  assign w640 = ( ~w564 & w621 ) | ( ~w564 & w638 ) | ( w621 & w638 ) ;
  assign w641 = ( ~\pi416 & w639 ) | ( ~\pi416 & w640 ) | ( w639 & w640 ) ;
  assign w642 = ~w637 & w641 ;
  assign w643 = ( ~\pi303 & \pi431 ) | ( ~\pi303 & w642 ) | ( \pi431 & w642 ) ;
  assign w644 = ~w642 & w643 ;
  assign w645 = ( \pi302 & ~\pi430 ) | ( \pi302 & w575 ) | ( ~\pi430 & w575 ) ;
  assign w646 = ( w642 & ~w644 ) | ( w642 & w645 ) | ( ~w644 & w645 ) ;
  assign w647 = \pi310 | \pi438 ;
  assign w648 = ~\pi311 & \pi439 ;
  assign w649 = ( ~\pi310 & w647 ) | ( ~\pi310 & w648 ) | ( w647 & w648 ) ;
  assign w650 = \pi308 & \pi436 ;
  assign w651 = \pi309 & \pi437 ;
  assign w652 = ( \pi437 & w649 ) | ( \pi437 & ~w651 ) | ( w649 & ~w651 ) ;
  assign w653 = ( \pi436 & ~w650 ) | ( \pi436 & w652 ) | ( ~w650 & w652 ) ;
  assign w654 = ~\pi305 & \pi433 ;
  assign w655 = ( ~\pi307 & \pi435 ) | ( ~\pi307 & w654 ) | ( \pi435 & w654 ) ;
  assign w656 = \pi434 | w655 ;
  assign w657 = ( ~\pi306 & w655 ) | ( ~\pi306 & w656 ) | ( w655 & w656 ) ;
  assign w658 = w654 | w657 ;
  assign w659 = w653 | w658 ;
  assign w660 = ( ~\pi304 & \pi432 ) | ( ~\pi304 & w658 ) | ( \pi432 & w658 ) ;
  assign w661 = w659 | w660 ;
  assign w662 = \pi304 & ~\pi432 ;
  assign w663 = ( \pi305 & ~\pi433 ) | ( \pi305 & w662 ) | ( ~\pi433 & w662 ) ;
  assign w664 = \pi307 & ~w653 ;
  assign w665 = ( \pi306 & ~\pi434 ) | ( \pi306 & w663 ) | ( ~\pi434 & w663 ) ;
  assign w666 = \pi435 | w653 ;
  assign w667 = ( w664 & w665 ) | ( w664 & ~w666 ) | ( w665 & ~w666 ) ;
  assign w668 = \pi308 & ~\pi436 ;
  assign w669 = ( \pi309 & ~\pi437 ) | ( \pi309 & w668 ) | ( ~\pi437 & w668 ) ;
  assign w670 = \pi311 | w667 ;
  assign w671 = ( \pi310 & ~\pi438 ) | ( \pi310 & w669 ) | ( ~\pi438 & w669 ) ;
  assign w672 = \pi439 & ~w667 ;
  assign w673 = ( w670 & w671 ) | ( w670 & ~w672 ) | ( w671 & ~w672 ) ;
  assign w674 = \pi312 & \pi440 ;
  assign w675 = \pi313 & \pi441 ;
  assign w676 = ( \pi441 & w548 ) | ( \pi441 & ~w675 ) | ( w548 & ~w675 ) ;
  assign w677 = ( \pi440 & ~w674 ) | ( \pi440 & w676 ) | ( ~w674 & w676 ) ;
  assign w678 = \pi314 & \pi442 ;
  assign w679 = \pi315 & \pi443 ;
  assign w680 = ( \pi443 & w677 ) | ( \pi443 & ~w679 ) | ( w677 & ~w679 ) ;
  assign w681 = ( \pi442 & ~w678 ) | ( \pi442 & w680 ) | ( ~w678 & w680 ) ;
  assign w682 = w673 & ~w681 ;
  assign w683 = ( w661 & w681 ) | ( w661 & ~w682 ) | ( w681 & ~w682 ) ;
  assign w684 = ( ~w557 & w646 ) | ( ~w557 & w682 ) | ( w646 & w682 ) ;
  assign w685 = ( w573 & ~w683 ) | ( w573 & w684 ) | ( ~w683 & w684 ) ;
  assign w686 = ( w557 & ~w683 ) | ( w557 & w685 ) | ( ~w683 & w685 ) ;
  assign w687 = ( ~\pi319 & \pi447 ) | ( ~\pi319 & w686 ) | ( \pi447 & w686 ) ;
  assign w688 = ~w686 & w687 ;
  assign w689 = ( \pi318 & ~\pi446 ) | ( \pi318 & w556 ) | ( ~\pi446 & w556 ) ;
  assign w690 = ( w686 & ~w688 ) | ( w686 & w689 ) | ( ~w688 & w689 ) ;
  assign w691 = ~\pi320 & \pi448 ;
  assign w692 = ( \pi319 & ~\pi447 ) | ( \pi319 & w690 ) | ( ~\pi447 & w690 ) ;
  assign w693 = ~w691 & w692 ;
  assign w694 = ( w690 & ~w691 ) | ( w690 & w693 ) | ( ~w691 & w693 ) ;
  assign w695 = ( w554 & ~w691 ) | ( w554 & w694 ) | ( ~w691 & w694 ) ;
  assign w696 = ( \pi321 & ~\pi449 ) | ( \pi321 & w695 ) | ( ~\pi449 & w695 ) ;
  assign w697 = w695 & w696 ;
  assign w698 = \pi320 & ~\pi448 ;
  assign w699 = ( \pi321 & ~\pi449 ) | ( \pi321 & w698 ) | ( ~\pi449 & w698 ) ;
  assign w700 = w697 | w699 ;
  assign w701 = ( \pi322 & ~\pi450 ) | ( \pi322 & w700 ) | ( ~\pi450 & w700 ) ;
  assign w702 = ( \pi323 & ~\pi451 ) | ( \pi323 & w701 ) | ( ~\pi451 & w701 ) ;
  assign w703 = \pi324 | \pi452 ;
  assign w704 = ( \pi325 & \pi453 ) | ( \pi325 & ~w539 ) | ( \pi453 & ~w539 ) ;
  assign w705 = ( \pi325 & w702 ) | ( \pi325 & ~w704 ) | ( w702 & ~w704 ) ;
  assign w706 = ~w539 & w705 ;
  assign w707 = ( \pi324 & ~w703 ) | ( \pi324 & w706 ) | ( ~w703 & w706 ) ;
  assign w708 = \pi327 | w707 ;
  assign w709 = ( \pi326 & ~\pi454 ) | ( \pi326 & w541 ) | ( ~\pi454 & w541 ) ;
  assign w710 = \pi455 & ~w707 ;
  assign w711 = ( w708 & w709 ) | ( w708 & ~w710 ) | ( w709 & ~w710 ) ;
  assign w712 = \pi330 | \pi458 ;
  assign w713 = ~\pi331 & \pi459 ;
  assign w714 = ( ~\pi330 & w712 ) | ( ~\pi330 & w713 ) | ( w712 & w713 ) ;
  assign w715 = \pi328 | \pi456 ;
  assign w716 = ( \pi329 & \pi457 ) | ( \pi329 & ~w714 ) | ( \pi457 & ~w714 ) ;
  assign w717 = ( \pi329 & w711 ) | ( \pi329 & ~w716 ) | ( w711 & ~w716 ) ;
  assign w718 = ~w714 & w717 ;
  assign w719 = ( \pi328 & ~w715 ) | ( \pi328 & w718 ) | ( ~w715 & w718 ) ;
  assign w720 = \pi328 & ~\pi456 ;
  assign w721 = ( \pi329 & ~\pi457 ) | ( \pi329 & w720 ) | ( ~\pi457 & w720 ) ;
  assign w722 = \pi331 | w719 ;
  assign w723 = ( \pi330 & ~\pi458 ) | ( \pi330 & w721 ) | ( ~\pi458 & w721 ) ;
  assign w724 = \pi459 & ~w719 ;
  assign w725 = ( w722 & w723 ) | ( w722 & ~w724 ) | ( w723 & ~w724 ) ;
  assign w726 = \pi332 | \pi460 ;
  assign w727 = ~\pi333 & \pi461 ;
  assign w728 = ( ~\pi332 & w726 ) | ( ~\pi332 & w727 ) | ( w726 & w727 ) ;
  assign w729 = ( w535 & w725 ) | ( w535 & ~w728 ) | ( w725 & ~w728 ) ;
  assign w730 = ( \pi334 & ~\pi462 ) | ( \pi334 & w729 ) | ( ~\pi462 & w729 ) ;
  assign w731 = ~w535 & w730 ;
  assign w732 = w536 & ~w731 ;
  assign w733 = ( \pi332 & ~\pi460 ) | ( \pi332 & w732 ) | ( ~\pi460 & w732 ) ;
  assign w734 = ( \pi333 & ~\pi461 ) | ( \pi333 & w733 ) | ( ~\pi461 & w733 ) ;
  assign w735 = ( w731 & ~w732 ) | ( w731 & w734 ) | ( ~w732 & w734 ) ;
  assign w736 = \pi335 | w735 ;
  assign w737 = ( ~\pi463 & w735 ) | ( ~\pi463 & w736 ) | ( w735 & w736 ) ;
  assign w738 = ~\pi337 & \pi465 ;
  assign w739 = w737 & ~w738 ;
  assign w740 = \pi338 & \pi466 ;
  assign w741 = \pi339 & \pi467 ;
  assign w742 = ( ~\pi467 & w739 ) | ( ~\pi467 & w741 ) | ( w739 & w741 ) ;
  assign w743 = ( ~\pi466 & w740 ) | ( ~\pi466 & w742 ) | ( w740 & w742 ) ;
  assign w744 = \pi336 & ~\pi464 ;
  assign w745 = ( \pi337 & ~\pi465 ) | ( \pi337 & w744 ) | ( ~\pi465 & w744 ) ;
  assign w746 = ( \pi338 & ~\pi466 ) | ( \pi338 & w745 ) | ( ~\pi466 & w745 ) ;
  assign w747 = ( \pi339 & ~\pi467 ) | ( \pi339 & w746 ) | ( ~\pi467 & w746 ) ;
  assign w748 = \pi340 & \pi468 ;
  assign w749 = \pi341 & \pi469 ;
  assign w750 = ( \pi469 & w531 ) | ( \pi469 & ~w749 ) | ( w531 & ~w749 ) ;
  assign w751 = ( \pi468 & ~w748 ) | ( \pi468 & w750 ) | ( ~w748 & w750 ) ;
  assign w752 = w747 & ~w751 ;
  assign w753 = ( w743 & ~w751 ) | ( w743 & w752 ) | ( ~w751 & w752 ) ;
  assign w754 = ~\pi336 & \pi464 ;
  assign w755 = ( w752 & w753 ) | ( w752 & ~w754 ) | ( w753 & ~w754 ) ;
  assign w756 = \pi343 | w755 ;
  assign w757 = ( \pi342 & ~\pi470 ) | ( \pi342 & w533 ) | ( ~\pi470 & w533 ) ;
  assign w758 = \pi471 & ~w755 ;
  assign w759 = ( w756 & w757 ) | ( w756 & ~w758 ) | ( w757 & ~w758 ) ;
  assign w760 = \pi346 | \pi474 ;
  assign w761 = ~\pi347 & \pi475 ;
  assign w762 = ( ~\pi346 & w760 ) | ( ~\pi346 & w761 ) | ( w760 & w761 ) ;
  assign w763 = \pi344 | \pi472 ;
  assign w764 = ( \pi345 & \pi473 ) | ( \pi345 & ~w762 ) | ( \pi473 & ~w762 ) ;
  assign w765 = ( \pi345 & w759 ) | ( \pi345 & ~w764 ) | ( w759 & ~w764 ) ;
  assign w766 = ~w762 & w765 ;
  assign w767 = ( \pi344 & ~w763 ) | ( \pi344 & w766 ) | ( ~w763 & w766 ) ;
  assign w768 = \pi344 & ~\pi472 ;
  assign w769 = ( \pi345 & ~\pi473 ) | ( \pi345 & w768 ) | ( ~\pi473 & w768 ) ;
  assign w770 = \pi347 | w767 ;
  assign w771 = ( \pi346 & ~\pi474 ) | ( \pi346 & w769 ) | ( ~\pi474 & w769 ) ;
  assign w772 = \pi475 & ~w767 ;
  assign w773 = ( w770 & w771 ) | ( w770 & ~w772 ) | ( w771 & ~w772 ) ;
  assign w774 = \pi348 | \pi476 ;
  assign w775 = ~\pi349 & \pi477 ;
  assign w776 = ( ~\pi348 & w774 ) | ( ~\pi348 & w775 ) | ( w774 & w775 ) ;
  assign w777 = ( w527 & w773 ) | ( w527 & ~w776 ) | ( w773 & ~w776 ) ;
  assign w778 = ( \pi350 & ~\pi478 ) | ( \pi350 & w777 ) | ( ~\pi478 & w777 ) ;
  assign w779 = ~w527 & w778 ;
  assign w780 = w528 & ~w779 ;
  assign w781 = ( \pi348 & ~\pi476 ) | ( \pi348 & w780 ) | ( ~\pi476 & w780 ) ;
  assign w782 = ( \pi349 & ~\pi477 ) | ( \pi349 & w781 ) | ( ~\pi477 & w781 ) ;
  assign w783 = ( w779 & ~w780 ) | ( w779 & w782 ) | ( ~w780 & w782 ) ;
  assign w784 = \pi351 | w783 ;
  assign w785 = ( ~\pi479 & w783 ) | ( ~\pi479 & w784 ) | ( w783 & w784 ) ;
  assign w786 = ~\pi353 & \pi481 ;
  assign w787 = w785 & ~w786 ;
  assign w788 = \pi354 & \pi482 ;
  assign w789 = \pi355 & \pi483 ;
  assign w790 = ( ~\pi483 & w787 ) | ( ~\pi483 & w789 ) | ( w787 & w789 ) ;
  assign w791 = ( ~\pi482 & w788 ) | ( ~\pi482 & w790 ) | ( w788 & w790 ) ;
  assign w792 = \pi352 & ~\pi480 ;
  assign w793 = ( \pi353 & ~\pi481 ) | ( \pi353 & w792 ) | ( ~\pi481 & w792 ) ;
  assign w794 = ( \pi354 & ~\pi482 ) | ( \pi354 & w793 ) | ( ~\pi482 & w793 ) ;
  assign w795 = ( \pi355 & ~\pi483 ) | ( \pi355 & w794 ) | ( ~\pi483 & w794 ) ;
  assign w796 = \pi356 & \pi484 ;
  assign w797 = \pi357 & \pi485 ;
  assign w798 = ( \pi485 & w523 ) | ( \pi485 & ~w797 ) | ( w523 & ~w797 ) ;
  assign w799 = ( \pi484 & ~w796 ) | ( \pi484 & w798 ) | ( ~w796 & w798 ) ;
  assign w800 = w795 & ~w799 ;
  assign w801 = ( w791 & ~w799 ) | ( w791 & w800 ) | ( ~w799 & w800 ) ;
  assign w802 = ~\pi352 & \pi480 ;
  assign w803 = ( w800 & w801 ) | ( w800 & ~w802 ) | ( w801 & ~w802 ) ;
  assign w804 = \pi359 | w803 ;
  assign w805 = ( \pi358 & ~\pi486 ) | ( \pi358 & w525 ) | ( ~\pi486 & w525 ) ;
  assign w806 = \pi487 & ~w803 ;
  assign w807 = ( w804 & w805 ) | ( w804 & ~w806 ) | ( w805 & ~w806 ) ;
  assign w808 = \pi362 | \pi490 ;
  assign w809 = ~\pi363 & \pi491 ;
  assign w810 = ( ~\pi362 & w808 ) | ( ~\pi362 & w809 ) | ( w808 & w809 ) ;
  assign w811 = \pi360 | \pi488 ;
  assign w812 = ( \pi361 & \pi489 ) | ( \pi361 & ~w810 ) | ( \pi489 & ~w810 ) ;
  assign w813 = ( \pi361 & w807 ) | ( \pi361 & ~w812 ) | ( w807 & ~w812 ) ;
  assign w814 = ~w810 & w813 ;
  assign w815 = ( \pi360 & ~w811 ) | ( \pi360 & w814 ) | ( ~w811 & w814 ) ;
  assign w816 = \pi360 & ~\pi488 ;
  assign w817 = ( \pi361 & ~\pi489 ) | ( \pi361 & w816 ) | ( ~\pi489 & w816 ) ;
  assign w818 = \pi363 | w815 ;
  assign w819 = ( \pi362 & ~\pi490 ) | ( \pi362 & w817 ) | ( ~\pi490 & w817 ) ;
  assign w820 = \pi491 & ~w815 ;
  assign w821 = ( w818 & w819 ) | ( w818 & ~w820 ) | ( w819 & ~w820 ) ;
  assign w822 = \pi364 | \pi492 ;
  assign w823 = ~\pi365 & \pi493 ;
  assign w824 = ( ~\pi364 & w822 ) | ( ~\pi364 & w823 ) | ( w822 & w823 ) ;
  assign w825 = ( w519 & w821 ) | ( w519 & ~w824 ) | ( w821 & ~w824 ) ;
  assign w826 = ( \pi366 & ~\pi494 ) | ( \pi366 & w825 ) | ( ~\pi494 & w825 ) ;
  assign w827 = ~w519 & w826 ;
  assign w828 = w520 & ~w827 ;
  assign w829 = ( \pi364 & ~\pi492 ) | ( \pi364 & w828 ) | ( ~\pi492 & w828 ) ;
  assign w830 = ( \pi365 & ~\pi493 ) | ( \pi365 & w829 ) | ( ~\pi493 & w829 ) ;
  assign w831 = ( w827 & ~w828 ) | ( w827 & w830 ) | ( ~w828 & w830 ) ;
  assign w832 = \pi367 | w831 ;
  assign w833 = ( ~\pi495 & w831 ) | ( ~\pi495 & w832 ) | ( w831 & w832 ) ;
  assign w834 = ~\pi369 & \pi497 ;
  assign w835 = w833 & ~w834 ;
  assign w836 = \pi370 & \pi498 ;
  assign w837 = \pi371 & \pi499 ;
  assign w838 = ( ~\pi499 & w835 ) | ( ~\pi499 & w837 ) | ( w835 & w837 ) ;
  assign w839 = ( ~\pi498 & w836 ) | ( ~\pi498 & w838 ) | ( w836 & w838 ) ;
  assign w840 = \pi368 & ~\pi496 ;
  assign w841 = ( \pi369 & ~\pi497 ) | ( \pi369 & w840 ) | ( ~\pi497 & w840 ) ;
  assign w842 = ( \pi370 & ~\pi498 ) | ( \pi370 & w841 ) | ( ~\pi498 & w841 ) ;
  assign w843 = ( \pi371 & ~\pi499 ) | ( \pi371 & w842 ) | ( ~\pi499 & w842 ) ;
  assign w844 = \pi372 & \pi500 ;
  assign w845 = \pi373 & \pi501 ;
  assign w846 = ( \pi501 & w515 ) | ( \pi501 & ~w845 ) | ( w515 & ~w845 ) ;
  assign w847 = ( \pi500 & ~w844 ) | ( \pi500 & w846 ) | ( ~w844 & w846 ) ;
  assign w848 = w843 & ~w847 ;
  assign w849 = ( w839 & ~w847 ) | ( w839 & w848 ) | ( ~w847 & w848 ) ;
  assign w850 = ~\pi368 & \pi496 ;
  assign w851 = ( w848 & w849 ) | ( w848 & ~w850 ) | ( w849 & ~w850 ) ;
  assign w852 = \pi375 | w851 ;
  assign w853 = ( \pi374 & ~\pi502 ) | ( \pi374 & w517 ) | ( ~\pi502 & w517 ) ;
  assign w854 = \pi503 & ~w851 ;
  assign w855 = ( w852 & w853 ) | ( w852 & ~w854 ) | ( w853 & ~w854 ) ;
  assign w856 = \pi378 | \pi506 ;
  assign w857 = ~\pi379 & \pi507 ;
  assign w858 = ( ~\pi378 & w856 ) | ( ~\pi378 & w857 ) | ( w856 & w857 ) ;
  assign w859 = \pi376 | \pi504 ;
  assign w860 = ( \pi377 & \pi505 ) | ( \pi377 & ~w858 ) | ( \pi505 & ~w858 ) ;
  assign w861 = ( \pi377 & w855 ) | ( \pi377 & ~w860 ) | ( w855 & ~w860 ) ;
  assign w862 = ~w858 & w861 ;
  assign w863 = ( \pi376 & ~w859 ) | ( \pi376 & w862 ) | ( ~w859 & w862 ) ;
  assign w864 = \pi376 & ~\pi504 ;
  assign w865 = ( \pi377 & ~\pi505 ) | ( \pi377 & w864 ) | ( ~\pi505 & w864 ) ;
  assign w866 = \pi379 | w863 ;
  assign w867 = ( \pi378 & ~\pi506 ) | ( \pi378 & w865 ) | ( ~\pi506 & w865 ) ;
  assign w868 = \pi507 & ~w863 ;
  assign w869 = ( w866 & w867 ) | ( w866 & ~w868 ) | ( w867 & ~w868 ) ;
  assign w870 = \pi383 & ~\pi511 ;
  assign w871 = \pi381 | \pi509 ;
  assign w872 = ~\pi382 & \pi510 ;
  assign w873 = ( ~\pi381 & w871 ) | ( ~\pi381 & w872 ) | ( w871 & w872 ) ;
  assign w874 = \pi380 & ~\pi508 ;
  assign w875 = ( \pi381 & ~\pi509 ) | ( \pi381 & w874 ) | ( ~\pi509 & w874 ) ;
  assign w876 = ( \pi382 & ~\pi510 ) | ( \pi382 & w875 ) | ( ~\pi510 & w875 ) ;
  assign w877 = ~w870 & w876 ;
  assign w878 = ( \pi380 & \pi508 ) | ( \pi380 & w877 ) | ( \pi508 & w877 ) ;
  assign w879 = ( ~\pi508 & w869 ) | ( ~\pi508 & w878 ) | ( w869 & w878 ) ;
  assign w880 = ( w870 & w873 ) | ( w870 & ~w877 ) | ( w873 & ~w877 ) ;
  assign w881 = ( w877 & w879 ) | ( w877 & ~w880 ) | ( w879 & ~w880 ) ;
  assign w882 = ( \pi383 & \pi511 ) | ( \pi383 & w881 ) | ( \pi511 & w881 ) ;
  assign w883 = \pi383 & w882 ;
  assign w884 = \pi118 | \pi246 ;
  assign w885 = ~\pi119 & \pi247 ;
  assign w886 = ( ~\pi118 & w884 ) | ( ~\pi118 & w885 ) | ( w884 & w885 ) ;
  assign w887 = \pi116 & ~\pi244 ;
  assign w888 = ( \pi117 & ~\pi245 ) | ( \pi117 & w887 ) | ( ~\pi245 & w887 ) ;
  assign w889 = \pi110 | \pi238 ;
  assign w890 = ~\pi111 & \pi239 ;
  assign w891 = ( ~\pi110 & w889 ) | ( ~\pi110 & w890 ) | ( w889 & w890 ) ;
  assign w892 = \pi102 | \pi230 ;
  assign w893 = ~\pi103 & \pi231 ;
  assign w894 = ( ~\pi102 & w892 ) | ( ~\pi102 & w893 ) | ( w892 & w893 ) ;
  assign w895 = \pi100 & ~\pi228 ;
  assign w896 = ( \pi101 & ~\pi229 ) | ( \pi101 & w895 ) | ( ~\pi229 & w895 ) ;
  assign w897 = \pi094 | \pi222 ;
  assign w898 = ~\pi095 & \pi223 ;
  assign w899 = ( ~\pi094 & w897 ) | ( ~\pi094 & w898 ) | ( w897 & w898 ) ;
  assign w900 = \pi086 | \pi214 ;
  assign w901 = ~\pi087 & \pi215 ;
  assign w902 = ( ~\pi086 & w900 ) | ( ~\pi086 & w901 ) | ( w900 & w901 ) ;
  assign w903 = \pi084 & ~\pi212 ;
  assign w904 = ( \pi085 & ~\pi213 ) | ( \pi085 & w903 ) | ( ~\pi213 & w903 ) ;
  assign w905 = \pi078 | \pi206 ;
  assign w906 = ~\pi079 & \pi207 ;
  assign w907 = ( ~\pi078 & w905 ) | ( ~\pi078 & w906 ) | ( w905 & w906 ) ;
  assign w908 = \pi070 | \pi198 ;
  assign w909 = ~\pi071 & \pi199 ;
  assign w910 = ( ~\pi070 & w908 ) | ( ~\pi070 & w909 ) | ( w908 & w909 ) ;
  assign w911 = \pi068 & ~\pi196 ;
  assign w912 = ( \pi069 & ~\pi197 ) | ( \pi069 & w911 ) | ( ~\pi197 & w911 ) ;
  assign w913 = \pi062 | \pi190 ;
  assign w914 = ~\pi063 & \pi191 ;
  assign w915 = ( ~\pi062 & w913 ) | ( ~\pi062 & w914 ) | ( w913 & w914 ) ;
  assign w916 = \pi060 & \pi188 ;
  assign w917 = \pi061 & \pi189 ;
  assign w918 = ( \pi189 & w915 ) | ( \pi189 & ~w917 ) | ( w915 & ~w917 ) ;
  assign w919 = ( \pi188 & ~w916 ) | ( \pi188 & w918 ) | ( ~w916 & w918 ) ;
  assign w920 = \pi056 & ~\pi184 ;
  assign w921 = ( \pi057 & ~\pi185 ) | ( \pi057 & w920 ) | ( ~\pi185 & w920 ) ;
  assign w922 = \pi059 & ~w919 ;
  assign w923 = ( \pi058 & ~\pi186 ) | ( \pi058 & w921 ) | ( ~\pi186 & w921 ) ;
  assign w924 = \pi187 | w919 ;
  assign w925 = ( w922 & w923 ) | ( w922 & ~w924 ) | ( w923 & ~w924 ) ;
  assign w926 = \pi060 & ~\pi188 ;
  assign w927 = ( \pi061 & ~\pi189 ) | ( \pi061 & w926 ) | ( ~\pi189 & w926 ) ;
  assign w928 = \pi047 & ~\pi175 ;
  assign w929 = \pi046 | \pi174 ;
  assign w930 = ~\pi047 & \pi175 ;
  assign w931 = ( ~\pi046 & w929 ) | ( ~\pi046 & w930 ) | ( w929 & w930 ) ;
  assign w932 = \pi044 & \pi172 ;
  assign w933 = \pi045 & \pi173 ;
  assign w934 = ( \pi173 & w931 ) | ( \pi173 & ~w933 ) | ( w931 & ~w933 ) ;
  assign w935 = ( \pi172 & ~w932 ) | ( \pi172 & w934 ) | ( ~w932 & w934 ) ;
  assign w936 = \pi042 | \pi170 ;
  assign w937 = ~\pi043 & \pi171 ;
  assign w938 = ( ~\pi042 & w936 ) | ( ~\pi042 & w937 ) | ( w936 & w937 ) ;
  assign w939 = \pi040 & ~\pi168 ;
  assign w940 = ( \pi041 & ~\pi169 ) | ( \pi041 & w939 ) | ( ~\pi169 & w939 ) ;
  assign w941 = \pi043 & ~w935 ;
  assign w942 = ( \pi042 & ~\pi170 ) | ( \pi042 & w940 ) | ( ~\pi170 & w940 ) ;
  assign w943 = \pi171 | w935 ;
  assign w944 = ( w941 & w942 ) | ( w941 & ~w943 ) | ( w942 & ~w943 ) ;
  assign w945 = \pi044 & ~\pi172 ;
  assign w946 = ( \pi045 & ~\pi173 ) | ( \pi045 & w945 ) | ( ~\pi173 & w945 ) ;
  assign w947 = \pi000 & ~\pi128 ;
  assign w948 = ( \pi001 & ~\pi129 ) | ( \pi001 & w947 ) | ( ~\pi129 & w947 ) ;
  assign w949 = ( \pi002 & ~\pi130 ) | ( \pi002 & w948 ) | ( ~\pi130 & w948 ) ;
  assign w950 = ( \pi003 & ~\pi131 ) | ( \pi003 & w949 ) | ( ~\pi131 & w949 ) ;
  assign w951 = ( \pi004 & ~\pi132 ) | ( \pi004 & w950 ) | ( ~\pi132 & w950 ) ;
  assign w952 = ( \pi005 & ~\pi133 ) | ( \pi005 & w951 ) | ( ~\pi133 & w951 ) ;
  assign w953 = ( \pi006 & ~\pi134 ) | ( \pi006 & w952 ) | ( ~\pi134 & w952 ) ;
  assign w954 = ( \pi007 & ~\pi135 ) | ( \pi007 & w953 ) | ( ~\pi135 & w953 ) ;
  assign w955 = ( \pi008 & ~\pi136 ) | ( \pi008 & w954 ) | ( ~\pi136 & w954 ) ;
  assign w956 = ( \pi009 & ~\pi137 ) | ( \pi009 & w955 ) | ( ~\pi137 & w955 ) ;
  assign w957 = ( \pi010 & ~\pi138 ) | ( \pi010 & w956 ) | ( ~\pi138 & w956 ) ;
  assign w958 = ( \pi011 & ~\pi139 ) | ( \pi011 & w957 ) | ( ~\pi139 & w957 ) ;
  assign w959 = ( \pi012 & ~\pi140 ) | ( \pi012 & w958 ) | ( ~\pi140 & w958 ) ;
  assign w960 = ( \pi013 & ~\pi141 ) | ( \pi013 & w959 ) | ( ~\pi141 & w959 ) ;
  assign w961 = ( \pi014 & ~\pi142 ) | ( \pi014 & w960 ) | ( ~\pi142 & w960 ) ;
  assign w962 = ( \pi015 & ~\pi143 ) | ( \pi015 & w961 ) | ( ~\pi143 & w961 ) ;
  assign w963 = ( \pi016 & ~\pi144 ) | ( \pi016 & w962 ) | ( ~\pi144 & w962 ) ;
  assign w964 = ( \pi017 & ~\pi145 ) | ( \pi017 & w963 ) | ( ~\pi145 & w963 ) ;
  assign w965 = ( \pi018 & ~\pi146 ) | ( \pi018 & w964 ) | ( ~\pi146 & w964 ) ;
  assign w966 = ( \pi019 & ~\pi147 ) | ( \pi019 & w965 ) | ( ~\pi147 & w965 ) ;
  assign w967 = ( \pi020 & ~\pi148 ) | ( \pi020 & w966 ) | ( ~\pi148 & w966 ) ;
  assign w968 = ( \pi021 & ~\pi149 ) | ( \pi021 & w967 ) | ( ~\pi149 & w967 ) ;
  assign w969 = ( \pi022 & ~\pi150 ) | ( \pi022 & w968 ) | ( ~\pi150 & w968 ) ;
  assign w970 = ( \pi023 & ~\pi151 ) | ( \pi023 & w969 ) | ( ~\pi151 & w969 ) ;
  assign w971 = ( \pi024 & ~\pi152 ) | ( \pi024 & w970 ) | ( ~\pi152 & w970 ) ;
  assign w972 = ( \pi025 & ~\pi153 ) | ( \pi025 & w971 ) | ( ~\pi153 & w971 ) ;
  assign w973 = ( \pi026 & ~\pi154 ) | ( \pi026 & w972 ) | ( ~\pi154 & w972 ) ;
  assign w974 = ( \pi027 & ~\pi155 ) | ( \pi027 & w973 ) | ( ~\pi155 & w973 ) ;
  assign w975 = ( \pi028 & ~\pi156 ) | ( \pi028 & w974 ) | ( ~\pi156 & w974 ) ;
  assign w976 = ( \pi029 & ~\pi157 ) | ( \pi029 & w975 ) | ( ~\pi157 & w975 ) ;
  assign w977 = ( \pi030 & ~\pi158 ) | ( \pi030 & w976 ) | ( ~\pi158 & w976 ) ;
  assign w978 = ( \pi031 & ~\pi159 ) | ( \pi031 & w977 ) | ( ~\pi159 & w977 ) ;
  assign w979 = \pi038 | \pi166 ;
  assign w980 = ~\pi039 & \pi167 ;
  assign w981 = ( ~\pi038 & w979 ) | ( ~\pi038 & w980 ) | ( w979 & w980 ) ;
  assign w982 = \pi036 & \pi164 ;
  assign w983 = \pi037 & \pi165 ;
  assign w984 = ( \pi165 & w981 ) | ( \pi165 & ~w983 ) | ( w981 & ~w983 ) ;
  assign w985 = ( \pi164 & ~w982 ) | ( \pi164 & w984 ) | ( ~w982 & w984 ) ;
  assign w986 = \pi034 | \pi162 ;
  assign w987 = ~\pi035 & \pi163 ;
  assign w988 = ( ~\pi034 & w986 ) | ( ~\pi034 & w987 ) | ( w986 & w987 ) ;
  assign w989 = w978 & ~w985 ;
  assign w990 = ( \pi033 & ~\pi161 ) | ( \pi033 & w989 ) | ( ~\pi161 & w989 ) ;
  assign w991 = ( w988 & w989 ) | ( w988 & ~w990 ) | ( w989 & ~w990 ) ;
  assign w992 = w989 & ~w991 ;
  assign w993 = \pi036 & ~\pi164 ;
  assign w994 = ( \pi037 & ~\pi165 ) | ( \pi037 & w993 ) | ( ~\pi165 & w993 ) ;
  assign w995 = \pi032 & ~\pi160 ;
  assign w996 = ( \pi033 & ~\pi161 ) | ( \pi033 & w995 ) | ( ~\pi161 & w995 ) ;
  assign w997 = \pi035 & ~w985 ;
  assign w998 = ( \pi034 & ~\pi162 ) | ( \pi034 & w996 ) | ( ~\pi162 & w996 ) ;
  assign w999 = \pi163 | w985 ;
  assign w1000 = ( w997 & w998 ) | ( w997 & ~w999 ) | ( w998 & ~w999 ) ;
  assign w1001 = \pi039 | w1000 ;
  assign w1002 = ( \pi038 & ~\pi166 ) | ( \pi038 & w994 ) | ( ~\pi166 & w994 ) ;
  assign w1003 = \pi167 & ~w1000 ;
  assign w1004 = ( w1001 & w1002 ) | ( w1001 & ~w1003 ) | ( w1002 & ~w1003 ) ;
  assign w1005 = \pi040 & \pi168 ;
  assign w1006 = \pi041 & \pi169 ;
  assign w1007 = ( \pi169 & w938 ) | ( \pi169 & ~w1006 ) | ( w938 & ~w1006 ) ;
  assign w1008 = ( \pi168 & ~w1005 ) | ( \pi168 & w1007 ) | ( ~w1005 & w1007 ) ;
  assign w1009 = ( ~w935 & w1004 ) | ( ~w935 & w1008 ) | ( w1004 & w1008 ) ;
  assign w1010 = ( \pi032 & \pi160 ) | ( \pi032 & w1009 ) | ( \pi160 & w1009 ) ;
  assign w1011 = ( ~w935 & w992 ) | ( ~w935 & w1009 ) | ( w992 & w1009 ) ;
  assign w1012 = ( ~\pi160 & w1010 ) | ( ~\pi160 & w1011 ) | ( w1010 & w1011 ) ;
  assign w1013 = ~w1008 & w1012 ;
  assign w1014 = ( ~\pi047 & \pi175 ) | ( ~\pi047 & w1013 ) | ( \pi175 & w1013 ) ;
  assign w1015 = ~w1013 & w1014 ;
  assign w1016 = ( \pi046 & ~\pi174 ) | ( \pi046 & w946 ) | ( ~\pi174 & w946 ) ;
  assign w1017 = ( w1013 & ~w1015 ) | ( w1013 & w1016 ) | ( ~w1015 & w1016 ) ;
  assign w1018 = \pi054 | \pi182 ;
  assign w1019 = ~\pi055 & \pi183 ;
  assign w1020 = ( ~\pi054 & w1018 ) | ( ~\pi054 & w1019 ) | ( w1018 & w1019 ) ;
  assign w1021 = \pi052 & \pi180 ;
  assign w1022 = \pi053 & \pi181 ;
  assign w1023 = ( \pi181 & w1020 ) | ( \pi181 & ~w1022 ) | ( w1020 & ~w1022 ) ;
  assign w1024 = ( \pi180 & ~w1021 ) | ( \pi180 & w1023 ) | ( ~w1021 & w1023 ) ;
  assign w1025 = ~\pi049 & \pi177 ;
  assign w1026 = ( ~\pi051 & \pi179 ) | ( ~\pi051 & w1025 ) | ( \pi179 & w1025 ) ;
  assign w1027 = \pi178 | w1026 ;
  assign w1028 = ( ~\pi050 & w1026 ) | ( ~\pi050 & w1027 ) | ( w1026 & w1027 ) ;
  assign w1029 = w1025 | w1028 ;
  assign w1030 = w1024 | w1029 ;
  assign w1031 = ( ~\pi048 & \pi176 ) | ( ~\pi048 & w1029 ) | ( \pi176 & w1029 ) ;
  assign w1032 = w1030 | w1031 ;
  assign w1033 = \pi048 & ~\pi176 ;
  assign w1034 = ( \pi049 & ~\pi177 ) | ( \pi049 & w1033 ) | ( ~\pi177 & w1033 ) ;
  assign w1035 = \pi051 & ~w1024 ;
  assign w1036 = ( \pi050 & ~\pi178 ) | ( \pi050 & w1034 ) | ( ~\pi178 & w1034 ) ;
  assign w1037 = \pi179 | w1024 ;
  assign w1038 = ( w1035 & w1036 ) | ( w1035 & ~w1037 ) | ( w1036 & ~w1037 ) ;
  assign w1039 = \pi052 & ~\pi180 ;
  assign w1040 = ( \pi053 & ~\pi181 ) | ( \pi053 & w1039 ) | ( ~\pi181 & w1039 ) ;
  assign w1041 = \pi055 | w1038 ;
  assign w1042 = ( \pi054 & ~\pi182 ) | ( \pi054 & w1040 ) | ( ~\pi182 & w1040 ) ;
  assign w1043 = \pi183 & ~w1038 ;
  assign w1044 = ( w1041 & w1042 ) | ( w1041 & ~w1043 ) | ( w1042 & ~w1043 ) ;
  assign w1045 = \pi056 & \pi184 ;
  assign w1046 = \pi057 & \pi185 ;
  assign w1047 = ( \pi185 & w919 ) | ( \pi185 & ~w1046 ) | ( w919 & ~w1046 ) ;
  assign w1048 = ( \pi184 & ~w1045 ) | ( \pi184 & w1047 ) | ( ~w1045 & w1047 ) ;
  assign w1049 = \pi058 & \pi186 ;
  assign w1050 = \pi059 & \pi187 ;
  assign w1051 = ( \pi187 & w1048 ) | ( \pi187 & ~w1050 ) | ( w1048 & ~w1050 ) ;
  assign w1052 = ( \pi186 & ~w1049 ) | ( \pi186 & w1051 ) | ( ~w1049 & w1051 ) ;
  assign w1053 = w1044 & ~w1052 ;
  assign w1054 = ( w1032 & w1052 ) | ( w1032 & ~w1053 ) | ( w1052 & ~w1053 ) ;
  assign w1055 = ( ~w928 & w1017 ) | ( ~w928 & w1053 ) | ( w1017 & w1053 ) ;
  assign w1056 = ( w944 & ~w1054 ) | ( w944 & w1055 ) | ( ~w1054 & w1055 ) ;
  assign w1057 = ( w928 & ~w1054 ) | ( w928 & w1056 ) | ( ~w1054 & w1056 ) ;
  assign w1058 = ( ~\pi063 & \pi191 ) | ( ~\pi063 & w1057 ) | ( \pi191 & w1057 ) ;
  assign w1059 = ~w1057 & w1058 ;
  assign w1060 = ( \pi062 & ~\pi190 ) | ( \pi062 & w927 ) | ( ~\pi190 & w927 ) ;
  assign w1061 = ( w1057 & ~w1059 ) | ( w1057 & w1060 ) | ( ~w1059 & w1060 ) ;
  assign w1062 = ~\pi064 & \pi192 ;
  assign w1063 = ( \pi063 & ~\pi191 ) | ( \pi063 & w1061 ) | ( ~\pi191 & w1061 ) ;
  assign w1064 = ~w1062 & w1063 ;
  assign w1065 = ( w1061 & ~w1062 ) | ( w1061 & w1064 ) | ( ~w1062 & w1064 ) ;
  assign w1066 = ( w925 & ~w1062 ) | ( w925 & w1065 ) | ( ~w1062 & w1065 ) ;
  assign w1067 = ( \pi065 & ~\pi193 ) | ( \pi065 & w1066 ) | ( ~\pi193 & w1066 ) ;
  assign w1068 = w1066 & w1067 ;
  assign w1069 = \pi064 & ~\pi192 ;
  assign w1070 = ( \pi065 & ~\pi193 ) | ( \pi065 & w1069 ) | ( ~\pi193 & w1069 ) ;
  assign w1071 = w1068 | w1070 ;
  assign w1072 = ( \pi066 & ~\pi194 ) | ( \pi066 & w1071 ) | ( ~\pi194 & w1071 ) ;
  assign w1073 = ( \pi067 & ~\pi195 ) | ( \pi067 & w1072 ) | ( ~\pi195 & w1072 ) ;
  assign w1074 = \pi068 | \pi196 ;
  assign w1075 = ( \pi069 & \pi197 ) | ( \pi069 & ~w910 ) | ( \pi197 & ~w910 ) ;
  assign w1076 = ( \pi069 & w1073 ) | ( \pi069 & ~w1075 ) | ( w1073 & ~w1075 ) ;
  assign w1077 = ~w910 & w1076 ;
  assign w1078 = ( \pi068 & ~w1074 ) | ( \pi068 & w1077 ) | ( ~w1074 & w1077 ) ;
  assign w1079 = \pi071 | w1078 ;
  assign w1080 = ( \pi070 & ~\pi198 ) | ( \pi070 & w912 ) | ( ~\pi198 & w912 ) ;
  assign w1081 = \pi199 & ~w1078 ;
  assign w1082 = ( w1079 & w1080 ) | ( w1079 & ~w1081 ) | ( w1080 & ~w1081 ) ;
  assign w1083 = \pi074 | \pi202 ;
  assign w1084 = ~\pi075 & \pi203 ;
  assign w1085 = ( ~\pi074 & w1083 ) | ( ~\pi074 & w1084 ) | ( w1083 & w1084 ) ;
  assign w1086 = \pi072 | \pi200 ;
  assign w1087 = ( \pi073 & \pi201 ) | ( \pi073 & ~w1085 ) | ( \pi201 & ~w1085 ) ;
  assign w1088 = ( \pi073 & w1082 ) | ( \pi073 & ~w1087 ) | ( w1082 & ~w1087 ) ;
  assign w1089 = ~w1085 & w1088 ;
  assign w1090 = ( \pi072 & ~w1086 ) | ( \pi072 & w1089 ) | ( ~w1086 & w1089 ) ;
  assign w1091 = \pi072 & ~\pi200 ;
  assign w1092 = ( \pi073 & ~\pi201 ) | ( \pi073 & w1091 ) | ( ~\pi201 & w1091 ) ;
  assign w1093 = \pi075 | w1090 ;
  assign w1094 = ( \pi074 & ~\pi202 ) | ( \pi074 & w1092 ) | ( ~\pi202 & w1092 ) ;
  assign w1095 = \pi203 & ~w1090 ;
  assign w1096 = ( w1093 & w1094 ) | ( w1093 & ~w1095 ) | ( w1094 & ~w1095 ) ;
  assign w1097 = \pi076 | \pi204 ;
  assign w1098 = ~\pi077 & \pi205 ;
  assign w1099 = ( ~\pi076 & w1097 ) | ( ~\pi076 & w1098 ) | ( w1097 & w1098 ) ;
  assign w1100 = ( w906 & w1096 ) | ( w906 & ~w1099 ) | ( w1096 & ~w1099 ) ;
  assign w1101 = ( \pi078 & ~\pi206 ) | ( \pi078 & w1100 ) | ( ~\pi206 & w1100 ) ;
  assign w1102 = ~w906 & w1101 ;
  assign w1103 = w907 & ~w1102 ;
  assign w1104 = ( \pi076 & ~\pi204 ) | ( \pi076 & w1103 ) | ( ~\pi204 & w1103 ) ;
  assign w1105 = ( \pi077 & ~\pi205 ) | ( \pi077 & w1104 ) | ( ~\pi205 & w1104 ) ;
  assign w1106 = ( w1102 & ~w1103 ) | ( w1102 & w1105 ) | ( ~w1103 & w1105 ) ;
  assign w1107 = \pi079 | w1106 ;
  assign w1108 = ( ~\pi207 & w1106 ) | ( ~\pi207 & w1107 ) | ( w1106 & w1107 ) ;
  assign w1109 = ~\pi081 & \pi209 ;
  assign w1110 = w1108 & ~w1109 ;
  assign w1111 = \pi082 & \pi210 ;
  assign w1112 = \pi083 & \pi211 ;
  assign w1113 = ( ~\pi211 & w1110 ) | ( ~\pi211 & w1112 ) | ( w1110 & w1112 ) ;
  assign w1114 = ( ~\pi210 & w1111 ) | ( ~\pi210 & w1113 ) | ( w1111 & w1113 ) ;
  assign w1115 = \pi080 & ~\pi208 ;
  assign w1116 = ( \pi081 & ~\pi209 ) | ( \pi081 & w1115 ) | ( ~\pi209 & w1115 ) ;
  assign w1117 = ( \pi082 & ~\pi210 ) | ( \pi082 & w1116 ) | ( ~\pi210 & w1116 ) ;
  assign w1118 = ( \pi083 & ~\pi211 ) | ( \pi083 & w1117 ) | ( ~\pi211 & w1117 ) ;
  assign w1119 = \pi084 & \pi212 ;
  assign w1120 = \pi085 & \pi213 ;
  assign w1121 = ( \pi213 & w902 ) | ( \pi213 & ~w1120 ) | ( w902 & ~w1120 ) ;
  assign w1122 = ( \pi212 & ~w1119 ) | ( \pi212 & w1121 ) | ( ~w1119 & w1121 ) ;
  assign w1123 = w1118 & ~w1122 ;
  assign w1124 = ( w1114 & ~w1122 ) | ( w1114 & w1123 ) | ( ~w1122 & w1123 ) ;
  assign w1125 = ~\pi080 & \pi208 ;
  assign w1126 = ( w1123 & w1124 ) | ( w1123 & ~w1125 ) | ( w1124 & ~w1125 ) ;
  assign w1127 = \pi087 | w1126 ;
  assign w1128 = ( \pi086 & ~\pi214 ) | ( \pi086 & w904 ) | ( ~\pi214 & w904 ) ;
  assign w1129 = \pi215 & ~w1126 ;
  assign w1130 = ( w1127 & w1128 ) | ( w1127 & ~w1129 ) | ( w1128 & ~w1129 ) ;
  assign w1131 = \pi090 | \pi218 ;
  assign w1132 = ~\pi091 & \pi219 ;
  assign w1133 = ( ~\pi090 & w1131 ) | ( ~\pi090 & w1132 ) | ( w1131 & w1132 ) ;
  assign w1134 = \pi088 | \pi216 ;
  assign w1135 = ( \pi089 & \pi217 ) | ( \pi089 & ~w1133 ) | ( \pi217 & ~w1133 ) ;
  assign w1136 = ( \pi089 & w1130 ) | ( \pi089 & ~w1135 ) | ( w1130 & ~w1135 ) ;
  assign w1137 = ~w1133 & w1136 ;
  assign w1138 = ( \pi088 & ~w1134 ) | ( \pi088 & w1137 ) | ( ~w1134 & w1137 ) ;
  assign w1139 = \pi088 & ~\pi216 ;
  assign w1140 = ( \pi089 & ~\pi217 ) | ( \pi089 & w1139 ) | ( ~\pi217 & w1139 ) ;
  assign w1141 = \pi091 | w1138 ;
  assign w1142 = ( \pi090 & ~\pi218 ) | ( \pi090 & w1140 ) | ( ~\pi218 & w1140 ) ;
  assign w1143 = \pi219 & ~w1138 ;
  assign w1144 = ( w1141 & w1142 ) | ( w1141 & ~w1143 ) | ( w1142 & ~w1143 ) ;
  assign w1145 = \pi092 | \pi220 ;
  assign w1146 = ~\pi093 & \pi221 ;
  assign w1147 = ( ~\pi092 & w1145 ) | ( ~\pi092 & w1146 ) | ( w1145 & w1146 ) ;
  assign w1148 = ( w898 & w1144 ) | ( w898 & ~w1147 ) | ( w1144 & ~w1147 ) ;
  assign w1149 = ( \pi094 & ~\pi222 ) | ( \pi094 & w1148 ) | ( ~\pi222 & w1148 ) ;
  assign w1150 = ~w898 & w1149 ;
  assign w1151 = w899 & ~w1150 ;
  assign w1152 = ( \pi092 & ~\pi220 ) | ( \pi092 & w1151 ) | ( ~\pi220 & w1151 ) ;
  assign w1153 = ( \pi093 & ~\pi221 ) | ( \pi093 & w1152 ) | ( ~\pi221 & w1152 ) ;
  assign w1154 = ( w1150 & ~w1151 ) | ( w1150 & w1153 ) | ( ~w1151 & w1153 ) ;
  assign w1155 = \pi095 | w1154 ;
  assign w1156 = ( ~\pi223 & w1154 ) | ( ~\pi223 & w1155 ) | ( w1154 & w1155 ) ;
  assign w1157 = ~\pi097 & \pi225 ;
  assign w1158 = w1156 & ~w1157 ;
  assign w1159 = \pi098 & \pi226 ;
  assign w1160 = \pi099 & \pi227 ;
  assign w1161 = ( ~\pi227 & w1158 ) | ( ~\pi227 & w1160 ) | ( w1158 & w1160 ) ;
  assign w1162 = ( ~\pi226 & w1159 ) | ( ~\pi226 & w1161 ) | ( w1159 & w1161 ) ;
  assign w1163 = \pi096 & ~\pi224 ;
  assign w1164 = ( \pi097 & ~\pi225 ) | ( \pi097 & w1163 ) | ( ~\pi225 & w1163 ) ;
  assign w1165 = ( \pi098 & ~\pi226 ) | ( \pi098 & w1164 ) | ( ~\pi226 & w1164 ) ;
  assign w1166 = ( \pi099 & ~\pi227 ) | ( \pi099 & w1165 ) | ( ~\pi227 & w1165 ) ;
  assign w1167 = \pi100 & \pi228 ;
  assign w1168 = \pi101 & \pi229 ;
  assign w1169 = ( \pi229 & w894 ) | ( \pi229 & ~w1168 ) | ( w894 & ~w1168 ) ;
  assign w1170 = ( \pi228 & ~w1167 ) | ( \pi228 & w1169 ) | ( ~w1167 & w1169 ) ;
  assign w1171 = w1166 & ~w1170 ;
  assign w1172 = ( w1162 & ~w1170 ) | ( w1162 & w1171 ) | ( ~w1170 & w1171 ) ;
  assign w1173 = ~\pi096 & \pi224 ;
  assign w1174 = ( w1171 & w1172 ) | ( w1171 & ~w1173 ) | ( w1172 & ~w1173 ) ;
  assign w1175 = \pi103 | w1174 ;
  assign w1176 = ( \pi102 & ~\pi230 ) | ( \pi102 & w896 ) | ( ~\pi230 & w896 ) ;
  assign w1177 = \pi231 & ~w1174 ;
  assign w1178 = ( w1175 & w1176 ) | ( w1175 & ~w1177 ) | ( w1176 & ~w1177 ) ;
  assign w1179 = \pi106 | \pi234 ;
  assign w1180 = ~\pi107 & \pi235 ;
  assign w1181 = ( ~\pi106 & w1179 ) | ( ~\pi106 & w1180 ) | ( w1179 & w1180 ) ;
  assign w1182 = \pi104 | \pi232 ;
  assign w1183 = ( \pi105 & \pi233 ) | ( \pi105 & ~w1181 ) | ( \pi233 & ~w1181 ) ;
  assign w1184 = ( \pi105 & w1178 ) | ( \pi105 & ~w1183 ) | ( w1178 & ~w1183 ) ;
  assign w1185 = ~w1181 & w1184 ;
  assign w1186 = ( \pi104 & ~w1182 ) | ( \pi104 & w1185 ) | ( ~w1182 & w1185 ) ;
  assign w1187 = \pi104 & ~\pi232 ;
  assign w1188 = ( \pi105 & ~\pi233 ) | ( \pi105 & w1187 ) | ( ~\pi233 & w1187 ) ;
  assign w1189 = \pi107 | w1186 ;
  assign w1190 = ( \pi106 & ~\pi234 ) | ( \pi106 & w1188 ) | ( ~\pi234 & w1188 ) ;
  assign w1191 = \pi235 & ~w1186 ;
  assign w1192 = ( w1189 & w1190 ) | ( w1189 & ~w1191 ) | ( w1190 & ~w1191 ) ;
  assign w1193 = \pi108 | \pi236 ;
  assign w1194 = ~\pi109 & \pi237 ;
  assign w1195 = ( ~\pi108 & w1193 ) | ( ~\pi108 & w1194 ) | ( w1193 & w1194 ) ;
  assign w1196 = ( w890 & w1192 ) | ( w890 & ~w1195 ) | ( w1192 & ~w1195 ) ;
  assign w1197 = ( \pi110 & ~\pi238 ) | ( \pi110 & w1196 ) | ( ~\pi238 & w1196 ) ;
  assign w1198 = ~w890 & w1197 ;
  assign w1199 = w891 & ~w1198 ;
  assign w1200 = ( \pi108 & ~\pi236 ) | ( \pi108 & w1199 ) | ( ~\pi236 & w1199 ) ;
  assign w1201 = ( \pi109 & ~\pi237 ) | ( \pi109 & w1200 ) | ( ~\pi237 & w1200 ) ;
  assign w1202 = ( w1198 & ~w1199 ) | ( w1198 & w1201 ) | ( ~w1199 & w1201 ) ;
  assign w1203 = \pi111 | w1202 ;
  assign w1204 = ( ~\pi239 & w1202 ) | ( ~\pi239 & w1203 ) | ( w1202 & w1203 ) ;
  assign w1205 = ~\pi113 & \pi241 ;
  assign w1206 = w1204 & ~w1205 ;
  assign w1207 = \pi114 & \pi242 ;
  assign w1208 = \pi115 & \pi243 ;
  assign w1209 = ( ~\pi243 & w1206 ) | ( ~\pi243 & w1208 ) | ( w1206 & w1208 ) ;
  assign w1210 = ( ~\pi242 & w1207 ) | ( ~\pi242 & w1209 ) | ( w1207 & w1209 ) ;
  assign w1211 = \pi112 & ~\pi240 ;
  assign w1212 = ( \pi113 & ~\pi241 ) | ( \pi113 & w1211 ) | ( ~\pi241 & w1211 ) ;
  assign w1213 = ( \pi114 & ~\pi242 ) | ( \pi114 & w1212 ) | ( ~\pi242 & w1212 ) ;
  assign w1214 = ( \pi115 & ~\pi243 ) | ( \pi115 & w1213 ) | ( ~\pi243 & w1213 ) ;
  assign w1215 = \pi116 & \pi244 ;
  assign w1216 = \pi117 & \pi245 ;
  assign w1217 = ( \pi245 & w886 ) | ( \pi245 & ~w1216 ) | ( w886 & ~w1216 ) ;
  assign w1218 = ( \pi244 & ~w1215 ) | ( \pi244 & w1217 ) | ( ~w1215 & w1217 ) ;
  assign w1219 = w1214 & ~w1218 ;
  assign w1220 = ( w1210 & ~w1218 ) | ( w1210 & w1219 ) | ( ~w1218 & w1219 ) ;
  assign w1221 = ~\pi112 & \pi240 ;
  assign w1222 = ( w1219 & w1220 ) | ( w1219 & ~w1221 ) | ( w1220 & ~w1221 ) ;
  assign w1223 = \pi119 | w1222 ;
  assign w1224 = ( \pi118 & ~\pi246 ) | ( \pi118 & w888 ) | ( ~\pi246 & w888 ) ;
  assign w1225 = \pi247 & ~w1222 ;
  assign w1226 = ( w1223 & w1224 ) | ( w1223 & ~w1225 ) | ( w1224 & ~w1225 ) ;
  assign w1227 = \pi122 | \pi250 ;
  assign w1228 = ~\pi123 & \pi251 ;
  assign w1229 = ( ~\pi122 & w1227 ) | ( ~\pi122 & w1228 ) | ( w1227 & w1228 ) ;
  assign w1230 = \pi120 | \pi248 ;
  assign w1231 = ( \pi121 & \pi249 ) | ( \pi121 & ~w1229 ) | ( \pi249 & ~w1229 ) ;
  assign w1232 = ( \pi121 & w1226 ) | ( \pi121 & ~w1231 ) | ( w1226 & ~w1231 ) ;
  assign w1233 = ~w1229 & w1232 ;
  assign w1234 = ( \pi120 & ~w1230 ) | ( \pi120 & w1233 ) | ( ~w1230 & w1233 ) ;
  assign w1235 = \pi120 & ~\pi248 ;
  assign w1236 = ( \pi121 & ~\pi249 ) | ( \pi121 & w1235 ) | ( ~\pi249 & w1235 ) ;
  assign w1237 = \pi123 | w1234 ;
  assign w1238 = ( \pi122 & ~\pi250 ) | ( \pi122 & w1236 ) | ( ~\pi250 & w1236 ) ;
  assign w1239 = \pi251 & ~w1234 ;
  assign w1240 = ( w1237 & w1238 ) | ( w1237 & ~w1239 ) | ( w1238 & ~w1239 ) ;
  assign w1241 = \pi127 & ~\pi255 ;
  assign w1242 = \pi125 | \pi253 ;
  assign w1243 = ~\pi126 & \pi254 ;
  assign w1244 = ( ~\pi125 & w1242 ) | ( ~\pi125 & w1243 ) | ( w1242 & w1243 ) ;
  assign w1245 = \pi124 & ~\pi252 ;
  assign w1246 = ( \pi125 & ~\pi253 ) | ( \pi125 & w1245 ) | ( ~\pi253 & w1245 ) ;
  assign w1247 = ( \pi126 & ~\pi254 ) | ( \pi126 & w1246 ) | ( ~\pi254 & w1246 ) ;
  assign w1248 = ~w1241 & w1247 ;
  assign w1249 = ( \pi124 & \pi252 ) | ( \pi124 & w1248 ) | ( \pi252 & w1248 ) ;
  assign w1250 = ( ~\pi252 & w1240 ) | ( ~\pi252 & w1249 ) | ( w1240 & w1249 ) ;
  assign w1251 = ( w1241 & w1244 ) | ( w1241 & ~w1248 ) | ( w1244 & ~w1248 ) ;
  assign w1252 = ( w1248 & w1250 ) | ( w1248 & ~w1251 ) | ( w1250 & ~w1251 ) ;
  assign w1253 = ( \pi127 & \pi255 ) | ( \pi127 & w1252 ) | ( \pi255 & w1252 ) ;
  assign w1254 = \pi127 & w1253 ;
  assign w1255 = ( ~\pi127 & \pi255 ) | ( ~\pi127 & w1252 ) | ( \pi255 & w1252 ) ;
  assign w1256 = w1252 | w1255 ;
  assign w1257 = \pi247 ^ w1256 ;
  assign w1258 = ( \pi119 & \pi247 ) | ( \pi119 & w1257 ) | ( \pi247 & w1257 ) ;
  assign w1259 = ( ~\pi383 & \pi511 ) | ( ~\pi383 & w881 ) | ( \pi511 & w881 ) ;
  assign w1260 = w881 | w1259 ;
  assign w1261 = \pi503 ^ w1260 ;
  assign w1262 = ( \pi375 & \pi503 ) | ( \pi375 & w1261 ) | ( \pi503 & w1261 ) ;
  assign w1263 = \pi502 ^ w1260 ;
  assign w1264 = ( \pi374 & \pi502 ) | ( \pi374 & w1263 ) | ( \pi502 & w1263 ) ;
  assign w1265 = \pi246 ^ w1256 ;
  assign w1266 = ( \pi118 & \pi246 ) | ( \pi118 & w1265 ) | ( \pi246 & w1265 ) ;
  assign w1267 = \pi244 ^ w1256 ;
  assign w1268 = ( \pi116 & \pi244 ) | ( \pi116 & w1267 ) | ( \pi244 & w1267 ) ;
  assign w1269 = \pi245 ^ w1256 ;
  assign w1270 = ( \pi117 & \pi245 ) | ( \pi117 & w1269 ) | ( \pi245 & w1269 ) ;
  assign w1271 = \pi500 ^ w1260 ;
  assign w1272 = ( \pi372 & \pi500 ) | ( \pi372 & w1271 ) | ( \pi500 & w1271 ) ;
  assign w1273 = w1268 & ~w1272 ;
  assign w1274 = \pi501 ^ w1260 ;
  assign w1275 = ( \pi373 & \pi501 ) | ( \pi373 & w1274 ) | ( \pi501 & w1274 ) ;
  assign w1276 = ( w1270 & w1273 ) | ( w1270 & ~w1275 ) | ( w1273 & ~w1275 ) ;
  assign w1277 = \pi496 ^ w1260 ;
  assign w1278 = ( \pi368 & \pi496 ) | ( \pi368 & w1277 ) | ( \pi496 & w1277 ) ;
  assign w1279 = \pi240 ^ w1256 ;
  assign w1280 = ( \pi112 & \pi240 ) | ( \pi112 & w1279 ) | ( \pi240 & w1279 ) ;
  assign w1281 = \pi243 ^ w1256 ;
  assign w1282 = ( \pi115 & \pi243 ) | ( \pi115 & w1281 ) | ( \pi243 & w1281 ) ;
  assign w1283 = \pi499 ^ w1260 ;
  assign w1284 = ( \pi371 & \pi499 ) | ( \pi371 & w1283 ) | ( \pi499 & w1283 ) ;
  assign w1285 = \pi498 ^ w1260 ;
  assign w1286 = ( \pi370 & \pi498 ) | ( \pi370 & w1285 ) | ( \pi498 & w1285 ) ;
  assign w1287 = \pi242 ^ w1256 ;
  assign w1288 = ( \pi114 & \pi242 ) | ( \pi114 & w1287 ) | ( \pi242 & w1287 ) ;
  assign w1289 = w1286 | w1288 ;
  assign w1290 = ~w1282 & w1284 ;
  assign w1291 = ( ~w1288 & w1289 ) | ( ~w1288 & w1290 ) | ( w1289 & w1290 ) ;
  assign w1292 = \pi241 ^ w1256 ;
  assign w1293 = ( \pi113 & \pi241 ) | ( \pi113 & w1292 ) | ( \pi241 & w1292 ) ;
  assign w1294 = ( ~\pi369 & w1260 ) | ( ~\pi369 & w1293 ) | ( w1260 & w1293 ) ;
  assign w1295 = ( \pi497 & w1260 ) | ( \pi497 & ~w1293 ) | ( w1260 & ~w1293 ) ;
  assign w1296 = ~w1294 & w1295 ;
  assign w1297 = \pi239 ^ w1256 ;
  assign w1298 = ( \pi111 & \pi239 ) | ( \pi111 & w1297 ) | ( \pi239 & w1297 ) ;
  assign w1299 = \pi495 ^ w1260 ;
  assign w1300 = ( \pi367 & \pi495 ) | ( \pi367 & w1299 ) | ( \pi495 & w1299 ) ;
  assign w1301 = \pi494 ^ w1260 ;
  assign w1302 = ( \pi366 & \pi494 ) | ( \pi366 & w1301 ) | ( \pi494 & w1301 ) ;
  assign w1303 = \pi238 ^ w1256 ;
  assign w1304 = ( \pi110 & \pi238 ) | ( \pi110 & w1303 ) | ( \pi238 & w1303 ) ;
  assign w1305 = w1302 | w1304 ;
  assign w1306 = ~w1298 & w1300 ;
  assign w1307 = ( ~w1304 & w1305 ) | ( ~w1304 & w1306 ) | ( w1305 & w1306 ) ;
  assign w1308 = \pi237 ^ w1256 ;
  assign w1309 = ( \pi109 & \pi237 ) | ( \pi109 & w1308 ) | ( \pi237 & w1308 ) ;
  assign w1310 = \pi493 ^ w1260 ;
  assign w1311 = ( \pi365 & \pi493 ) | ( \pi365 & w1310 ) | ( \pi493 & w1310 ) ;
  assign w1312 = \pi236 ^ w1256 ;
  assign w1313 = ( \pi108 & \pi236 ) | ( \pi108 & w1312 ) | ( \pi236 & w1312 ) ;
  assign w1314 = \pi492 ^ w1260 ;
  assign w1315 = ( \pi364 & \pi492 ) | ( \pi364 & w1314 ) | ( \pi492 & w1314 ) ;
  assign w1316 = w1313 & ~w1315 ;
  assign w1317 = ( w1309 & ~w1311 ) | ( w1309 & w1316 ) | ( ~w1311 & w1316 ) ;
  assign w1318 = \pi231 ^ w1256 ;
  assign w1319 = ( \pi103 & \pi231 ) | ( \pi103 & w1318 ) | ( \pi231 & w1318 ) ;
  assign w1320 = \pi487 ^ w1260 ;
  assign w1321 = ( \pi359 & \pi487 ) | ( \pi359 & w1320 ) | ( \pi487 & w1320 ) ;
  assign w1322 = \pi486 ^ w1260 ;
  assign w1323 = ( \pi358 & \pi486 ) | ( \pi358 & w1322 ) | ( \pi486 & w1322 ) ;
  assign w1324 = \pi230 ^ w1256 ;
  assign w1325 = ( \pi102 & \pi230 ) | ( \pi102 & w1324 ) | ( \pi230 & w1324 ) ;
  assign w1326 = \pi229 ^ w1256 ;
  assign w1327 = ( \pi101 & \pi229 ) | ( \pi101 & w1326 ) | ( \pi229 & w1326 ) ;
  assign w1328 = \pi228 ^ w1256 ;
  assign w1329 = ( \pi100 & \pi228 ) | ( \pi100 & w1328 ) | ( \pi228 & w1328 ) ;
  assign w1330 = \pi484 ^ w1260 ;
  assign w1331 = ( \pi356 & \pi484 ) | ( \pi356 & w1330 ) | ( \pi484 & w1330 ) ;
  assign w1332 = w1329 & ~w1331 ;
  assign w1333 = \pi485 ^ w1260 ;
  assign w1334 = ( \pi357 & \pi485 ) | ( \pi357 & w1333 ) | ( \pi485 & w1333 ) ;
  assign w1335 = ( w1327 & w1332 ) | ( w1327 & ~w1334 ) | ( w1332 & ~w1334 ) ;
  assign w1336 = \pi480 ^ w1260 ;
  assign w1337 = ( \pi352 & \pi480 ) | ( \pi352 & w1336 ) | ( \pi480 & w1336 ) ;
  assign w1338 = \pi224 ^ w1256 ;
  assign w1339 = ( \pi096 & \pi224 ) | ( \pi096 & w1338 ) | ( \pi224 & w1338 ) ;
  assign w1340 = \pi227 ^ w1256 ;
  assign w1341 = ( \pi099 & \pi227 ) | ( \pi099 & w1340 ) | ( \pi227 & w1340 ) ;
  assign w1342 = \pi483 ^ w1260 ;
  assign w1343 = ( \pi355 & \pi483 ) | ( \pi355 & w1342 ) | ( \pi483 & w1342 ) ;
  assign w1344 = \pi482 ^ w1260 ;
  assign w1345 = ( \pi354 & \pi482 ) | ( \pi354 & w1344 ) | ( \pi482 & w1344 ) ;
  assign w1346 = \pi226 ^ w1256 ;
  assign w1347 = ( \pi098 & \pi226 ) | ( \pi098 & w1346 ) | ( \pi226 & w1346 ) ;
  assign w1348 = w1345 | w1347 ;
  assign w1349 = ~w1341 & w1343 ;
  assign w1350 = ( ~w1347 & w1348 ) | ( ~w1347 & w1349 ) | ( w1348 & w1349 ) ;
  assign w1351 = \pi225 ^ w1256 ;
  assign w1352 = ( \pi097 & \pi225 ) | ( \pi097 & w1351 ) | ( \pi225 & w1351 ) ;
  assign w1353 = ( ~\pi353 & w1260 ) | ( ~\pi353 & w1352 ) | ( w1260 & w1352 ) ;
  assign w1354 = ( \pi481 & w1260 ) | ( \pi481 & ~w1352 ) | ( w1260 & ~w1352 ) ;
  assign w1355 = ~w1353 & w1354 ;
  assign w1356 = \pi223 ^ w1256 ;
  assign w1357 = ( \pi095 & \pi223 ) | ( \pi095 & w1356 ) | ( \pi223 & w1356 ) ;
  assign w1358 = \pi479 ^ w1260 ;
  assign w1359 = ( \pi351 & \pi479 ) | ( \pi351 & w1358 ) | ( \pi479 & w1358 ) ;
  assign w1360 = \pi478 ^ w1260 ;
  assign w1361 = ( \pi350 & \pi478 ) | ( \pi350 & w1360 ) | ( \pi478 & w1360 ) ;
  assign w1362 = \pi222 ^ w1256 ;
  assign w1363 = ( \pi094 & \pi222 ) | ( \pi094 & w1362 ) | ( \pi222 & w1362 ) ;
  assign w1364 = w1361 | w1363 ;
  assign w1365 = ~w1357 & w1359 ;
  assign w1366 = ( ~w1363 & w1364 ) | ( ~w1363 & w1365 ) | ( w1364 & w1365 ) ;
  assign w1367 = \pi221 ^ w1256 ;
  assign w1368 = ( \pi093 & \pi221 ) | ( \pi093 & w1367 ) | ( \pi221 & w1367 ) ;
  assign w1369 = \pi477 ^ w1260 ;
  assign w1370 = ( \pi349 & \pi477 ) | ( \pi349 & w1369 ) | ( \pi477 & w1369 ) ;
  assign w1371 = \pi220 ^ w1256 ;
  assign w1372 = ( \pi092 & \pi220 ) | ( \pi092 & w1371 ) | ( \pi220 & w1371 ) ;
  assign w1373 = \pi476 ^ w1260 ;
  assign w1374 = ( \pi348 & \pi476 ) | ( \pi348 & w1373 ) | ( \pi476 & w1373 ) ;
  assign w1375 = w1372 & ~w1374 ;
  assign w1376 = ( w1368 & ~w1370 ) | ( w1368 & w1375 ) | ( ~w1370 & w1375 ) ;
  assign w1377 = \pi215 ^ w1256 ;
  assign w1378 = ( \pi087 & \pi215 ) | ( \pi087 & w1377 ) | ( \pi215 & w1377 ) ;
  assign w1379 = ( \pi343 & w1260 ) | ( \pi343 & ~w1378 ) | ( w1260 & ~w1378 ) ;
  assign w1380 = ( ~\pi471 & w1260 ) | ( ~\pi471 & w1378 ) | ( w1260 & w1378 ) ;
  assign w1381 = ~w1379 & w1380 ;
  assign w1382 = ( ~\pi343 & w1260 ) | ( ~\pi343 & w1378 ) | ( w1260 & w1378 ) ;
  assign w1383 = ( \pi471 & w1260 ) | ( \pi471 & ~w1378 ) | ( w1260 & ~w1378 ) ;
  assign w1384 = ~w1382 & w1383 ;
  assign w1385 = \pi470 ^ w1260 ;
  assign w1386 = ( \pi342 & \pi470 ) | ( \pi342 & w1385 ) | ( \pi470 & w1385 ) ;
  assign w1387 = \pi214 ^ w1256 ;
  assign w1388 = ( \pi086 & \pi214 ) | ( \pi086 & w1387 ) | ( \pi214 & w1387 ) ;
  assign w1389 = \pi213 ^ w1256 ;
  assign w1390 = ( \pi085 & \pi213 ) | ( \pi085 & w1389 ) | ( \pi213 & w1389 ) ;
  assign w1391 = \pi212 ^ w1256 ;
  assign w1392 = ( \pi084 & \pi212 ) | ( \pi084 & w1391 ) | ( \pi212 & w1391 ) ;
  assign w1393 = \pi468 ^ w1260 ;
  assign w1394 = ( \pi340 & \pi468 ) | ( \pi340 & w1393 ) | ( \pi468 & w1393 ) ;
  assign w1395 = w1392 & ~w1394 ;
  assign w1396 = \pi469 ^ w1260 ;
  assign w1397 = ( \pi341 & \pi469 ) | ( \pi341 & w1396 ) | ( \pi469 & w1396 ) ;
  assign w1398 = ( w1390 & w1395 ) | ( w1390 & ~w1397 ) | ( w1395 & ~w1397 ) ;
  assign w1399 = \pi464 ^ w1260 ;
  assign w1400 = ( \pi336 & \pi464 ) | ( \pi336 & w1399 ) | ( \pi464 & w1399 ) ;
  assign w1401 = \pi208 ^ w1256 ;
  assign w1402 = ( \pi080 & \pi208 ) | ( \pi080 & w1401 ) | ( \pi208 & w1401 ) ;
  assign w1403 = \pi211 ^ w1256 ;
  assign w1404 = ( \pi083 & \pi211 ) | ( \pi083 & w1403 ) | ( \pi211 & w1403 ) ;
  assign w1405 = \pi467 ^ w1260 ;
  assign w1406 = ( \pi339 & \pi467 ) | ( \pi339 & w1405 ) | ( \pi467 & w1405 ) ;
  assign w1407 = \pi466 ^ w1260 ;
  assign w1408 = ( \pi338 & \pi466 ) | ( \pi338 & w1407 ) | ( \pi466 & w1407 ) ;
  assign w1409 = \pi210 ^ w1256 ;
  assign w1410 = ( \pi082 & \pi210 ) | ( \pi082 & w1409 ) | ( \pi210 & w1409 ) ;
  assign w1411 = w1408 | w1410 ;
  assign w1412 = ~w1404 & w1406 ;
  assign w1413 = ( ~w1410 & w1411 ) | ( ~w1410 & w1412 ) | ( w1411 & w1412 ) ;
  assign w1414 = \pi209 ^ w1256 ;
  assign w1415 = ( \pi081 & \pi209 ) | ( \pi081 & w1414 ) | ( \pi209 & w1414 ) ;
  assign w1416 = ( ~\pi337 & w1260 ) | ( ~\pi337 & w1415 ) | ( w1260 & w1415 ) ;
  assign w1417 = ( \pi465 & w1260 ) | ( \pi465 & ~w1415 ) | ( w1260 & ~w1415 ) ;
  assign w1418 = ~w1416 & w1417 ;
  assign w1419 = \pi207 ^ w1256 ;
  assign w1420 = ( \pi079 & \pi207 ) | ( \pi079 & w1419 ) | ( \pi207 & w1419 ) ;
  assign w1421 = \pi463 ^ w1260 ;
  assign w1422 = ( \pi335 & \pi463 ) | ( \pi335 & w1421 ) | ( \pi463 & w1421 ) ;
  assign w1423 = \pi206 ^ w1256 ;
  assign w1424 = ( \pi078 & \pi206 ) | ( \pi078 & w1423 ) | ( \pi206 & w1423 ) ;
  assign w1425 = w1260 | w1424 ;
  assign w1426 = \pi462 | w1425 ;
  assign w1427 = ~w1420 & w1422 ;
  assign w1428 = ( ~\pi334 & w1424 ) | ( ~\pi334 & w1425 ) | ( w1424 & w1425 ) ;
  assign w1429 = ( w1426 & w1427 ) | ( w1426 & ~w1428 ) | ( w1427 & ~w1428 ) ;
  assign w1430 = \pi205 ^ w1256 ;
  assign w1431 = ( \pi077 & \pi205 ) | ( \pi077 & w1430 ) | ( \pi205 & w1430 ) ;
  assign w1432 = \pi204 ^ w1256 ;
  assign w1433 = ( \pi076 & \pi204 ) | ( \pi076 & w1432 ) | ( \pi204 & w1432 ) ;
  assign w1434 = \pi460 ^ w1260 ;
  assign w1435 = ( \pi332 & \pi460 ) | ( \pi332 & w1434 ) | ( \pi460 & w1434 ) ;
  assign w1436 = w1433 & ~w1435 ;
  assign w1437 = \pi461 ^ w1260 ;
  assign w1438 = ( \pi333 & \pi461 ) | ( \pi333 & w1437 ) | ( \pi461 & w1437 ) ;
  assign w1439 = ( w1431 & w1436 ) | ( w1431 & ~w1438 ) | ( w1436 & ~w1438 ) ;
  assign w1440 = ~w1422 & w1424 ;
  assign w1441 = ( w1420 & w1424 ) | ( w1420 & w1440 ) | ( w1424 & w1440 ) ;
  assign w1442 = \pi334 ^ w1260 ;
  assign w1443 = ( \pi334 & \pi462 ) | ( \pi334 & ~w1442 ) | ( \pi462 & ~w1442 ) ;
  assign w1444 = w1441 & ~w1443 ;
  assign w1445 = \pi199 ^ w1256 ;
  assign w1446 = ( \pi071 & \pi199 ) | ( \pi071 & w1445 ) | ( \pi199 & w1445 ) ;
  assign w1447 = \pi455 ^ w1260 ;
  assign w1448 = ( \pi327 & \pi455 ) | ( \pi327 & w1447 ) | ( \pi455 & w1447 ) ;
  assign w1449 = \pi454 ^ w1260 ;
  assign w1450 = ( \pi326 & \pi454 ) | ( \pi326 & w1449 ) | ( \pi454 & w1449 ) ;
  assign w1451 = \pi198 ^ w1256 ;
  assign w1452 = ( \pi070 & \pi198 ) | ( \pi070 & w1451 ) | ( \pi198 & w1451 ) ;
  assign w1453 = \pi197 ^ w1256 ;
  assign w1454 = ( \pi069 & \pi197 ) | ( \pi069 & w1453 ) | ( \pi197 & w1453 ) ;
  assign w1455 = \pi453 ^ w1260 ;
  assign w1456 = ( \pi325 & \pi453 ) | ( \pi325 & w1455 ) | ( \pi453 & w1455 ) ;
  assign w1457 = \pi196 ^ w1256 ;
  assign w1458 = ( \pi068 & \pi196 ) | ( \pi068 & w1457 ) | ( \pi196 & w1457 ) ;
  assign w1459 = \pi452 ^ w1260 ;
  assign w1460 = ( \pi324 & \pi452 ) | ( \pi324 & w1459 ) | ( \pi452 & w1459 ) ;
  assign w1461 = w1458 & ~w1460 ;
  assign w1462 = ( w1454 & ~w1456 ) | ( w1454 & w1461 ) | ( ~w1456 & w1461 ) ;
  assign w1463 = \pi195 ^ w1256 ;
  assign w1464 = ( \pi067 & \pi195 ) | ( \pi067 & w1463 ) | ( \pi195 & w1463 ) ;
  assign w1465 = \pi451 ^ w1260 ;
  assign w1466 = ( \pi323 & \pi451 ) | ( \pi323 & w1465 ) | ( \pi451 & w1465 ) ;
  assign w1467 = \pi450 ^ w1260 ;
  assign w1468 = ( \pi322 & \pi450 ) | ( \pi322 & w1467 ) | ( \pi450 & w1467 ) ;
  assign w1469 = \pi194 ^ w1256 ;
  assign w1470 = ( \pi066 & \pi194 ) | ( \pi066 & w1469 ) | ( \pi194 & w1469 ) ;
  assign w1471 = \pi448 ^ w1260 ;
  assign w1472 = ( \pi320 & \pi448 ) | ( \pi320 & w1471 ) | ( \pi448 & w1471 ) ;
  assign w1473 = \pi192 ^ w1256 ;
  assign w1474 = ( \pi064 & \pi192 ) | ( \pi064 & w1473 ) | ( \pi192 & w1473 ) ;
  assign w1475 = \pi193 ^ w1256 ;
  assign w1476 = ( \pi065 & \pi193 ) | ( \pi065 & w1475 ) | ( \pi193 & w1475 ) ;
  assign w1477 = \pi191 ^ w1256 ;
  assign w1478 = ( \pi063 & \pi191 ) | ( \pi063 & w1477 ) | ( \pi191 & w1477 ) ;
  assign w1479 = ( ~\pi319 & w1260 ) | ( ~\pi319 & w1478 ) | ( w1260 & w1478 ) ;
  assign w1480 = ( \pi447 & w1260 ) | ( \pi447 & ~w1478 ) | ( w1260 & ~w1478 ) ;
  assign w1481 = ~w1479 & w1480 ;
  assign w1482 = \pi446 ^ w1260 ;
  assign w1483 = ( \pi318 & \pi446 ) | ( \pi318 & w1482 ) | ( \pi446 & w1482 ) ;
  assign w1484 = \pi190 ^ w1256 ;
  assign w1485 = ( \pi062 & \pi190 ) | ( \pi062 & w1484 ) | ( \pi190 & w1484 ) ;
  assign w1486 = \pi188 ^ w1256 ;
  assign w1487 = ( \pi060 & \pi188 ) | ( \pi060 & w1486 ) | ( \pi188 & w1486 ) ;
  assign w1488 = \pi444 ^ w1260 ;
  assign w1489 = ( \pi316 & \pi444 ) | ( \pi316 & w1488 ) | ( \pi444 & w1488 ) ;
  assign w1490 = \pi189 ^ w1256 ;
  assign w1491 = ( \pi061 & \pi189 ) | ( \pi061 & w1490 ) | ( \pi189 & w1490 ) ;
  assign w1492 = w1260 | w1491 ;
  assign w1493 = \pi445 | w1492 ;
  assign w1494 = ~w1487 & w1489 ;
  assign w1495 = ( ~\pi317 & w1491 ) | ( ~\pi317 & w1492 ) | ( w1491 & w1492 ) ;
  assign w1496 = ( w1493 & w1494 ) | ( w1493 & ~w1495 ) | ( w1494 & ~w1495 ) ;
  assign w1497 = w1481 | w1496 ;
  assign w1498 = ( w1483 & ~w1485 ) | ( w1483 & w1496 ) | ( ~w1485 & w1496 ) ;
  assign w1499 = w1497 | w1498 ;
  assign w1500 = \pi187 ^ w1256 ;
  assign w1501 = ( \pi059 & \pi187 ) | ( \pi059 & w1500 ) | ( \pi187 & w1500 ) ;
  assign w1502 = \pi443 ^ w1260 ;
  assign w1503 = ( \pi315 & \pi443 ) | ( \pi315 & w1502 ) | ( \pi443 & w1502 ) ;
  assign w1504 = \pi186 ^ w1256 ;
  assign w1505 = ( \pi058 & \pi186 ) | ( \pi058 & w1504 ) | ( \pi186 & w1504 ) ;
  assign w1506 = \pi442 ^ w1260 ;
  assign w1507 = ( \pi314 & \pi442 ) | ( \pi314 & w1506 ) | ( \pi442 & w1506 ) ;
  assign w1508 = \pi185 ^ w1256 ;
  assign w1509 = ( \pi057 & \pi185 ) | ( \pi057 & w1508 ) | ( \pi185 & w1508 ) ;
  assign w1510 = \pi441 ^ w1260 ;
  assign w1511 = ( \pi313 & \pi441 ) | ( \pi313 & w1510 ) | ( \pi441 & w1510 ) ;
  assign w1512 = \pi184 ^ w1256 ;
  assign w1513 = ( \pi056 & \pi184 ) | ( \pi056 & w1512 ) | ( \pi184 & w1512 ) ;
  assign w1514 = \pi440 ^ w1260 ;
  assign w1515 = ( \pi312 & \pi440 ) | ( \pi312 & w1514 ) | ( \pi440 & w1514 ) ;
  assign w1516 = w1513 & ~w1515 ;
  assign w1517 = ( w1509 & ~w1511 ) | ( w1509 & w1516 ) | ( ~w1511 & w1516 ) ;
  assign w1518 = ~w1499 & w1501 ;
  assign w1519 = ( w1505 & ~w1507 ) | ( w1505 & w1517 ) | ( ~w1507 & w1517 ) ;
  assign w1520 = w1499 | w1503 ;
  assign w1521 = ( w1518 & w1519 ) | ( w1518 & ~w1520 ) | ( w1519 & ~w1520 ) ;
  assign w1522 = w1487 & ~w1489 ;
  assign w1523 = \pi445 ^ w1260 ;
  assign w1524 = ( \pi317 & \pi445 ) | ( \pi317 & w1523 ) | ( \pi445 & w1523 ) ;
  assign w1525 = ( w1491 & w1522 ) | ( w1491 & ~w1524 ) | ( w1522 & ~w1524 ) ;
  assign w1526 = \pi175 ^ w1256 ;
  assign w1527 = ( \pi047 & \pi175 ) | ( \pi047 & w1526 ) | ( \pi175 & w1526 ) ;
  assign w1528 = \pi431 ^ w1260 ;
  assign w1529 = ( \pi303 & \pi431 ) | ( \pi303 & w1528 ) | ( \pi431 & w1528 ) ;
  assign w1530 = ~w1527 & w1529 ;
  assign w1531 = \pi430 ^ w1260 ;
  assign w1532 = ( \pi302 & \pi430 ) | ( \pi302 & w1531 ) | ( \pi430 & w1531 ) ;
  assign w1533 = \pi174 ^ w1256 ;
  assign w1534 = ( \pi046 & \pi174 ) | ( \pi046 & w1533 ) | ( \pi174 & w1533 ) ;
  assign w1535 = \pi172 ^ w1256 ;
  assign w1536 = ( \pi044 & \pi172 ) | ( \pi044 & w1535 ) | ( \pi172 & w1535 ) ;
  assign w1537 = \pi428 ^ w1260 ;
  assign w1538 = ( \pi300 & \pi428 ) | ( \pi300 & w1537 ) | ( \pi428 & w1537 ) ;
  assign w1539 = \pi173 ^ w1256 ;
  assign w1540 = ( \pi045 & \pi173 ) | ( \pi045 & w1539 ) | ( \pi173 & w1539 ) ;
  assign w1541 = w1260 | w1540 ;
  assign w1542 = \pi429 | w1541 ;
  assign w1543 = ~w1536 & w1538 ;
  assign w1544 = ( ~\pi301 & w1540 ) | ( ~\pi301 & w1541 ) | ( w1540 & w1541 ) ;
  assign w1545 = ( w1542 & w1543 ) | ( w1542 & ~w1544 ) | ( w1543 & ~w1544 ) ;
  assign w1546 = w1530 | w1545 ;
  assign w1547 = ( w1532 & ~w1534 ) | ( w1532 & w1545 ) | ( ~w1534 & w1545 ) ;
  assign w1548 = w1546 | w1547 ;
  assign w1549 = \pi171 ^ w1256 ;
  assign w1550 = ( \pi043 & \pi171 ) | ( \pi043 & w1549 ) | ( \pi171 & w1549 ) ;
  assign w1551 = \pi427 ^ w1260 ;
  assign w1552 = ( \pi299 & \pi427 ) | ( \pi299 & w1551 ) | ( \pi427 & w1551 ) ;
  assign w1553 = \pi170 ^ w1256 ;
  assign w1554 = ( \pi042 & \pi170 ) | ( \pi042 & w1553 ) | ( \pi170 & w1553 ) ;
  assign w1555 = \pi426 ^ w1260 ;
  assign w1556 = ( \pi298 & \pi426 ) | ( \pi298 & w1555 ) | ( \pi426 & w1555 ) ;
  assign w1557 = w1554 & w1556 ;
  assign w1558 = ~w1550 & w1552 ;
  assign w1559 = ( w1556 & ~w1557 ) | ( w1556 & w1558 ) | ( ~w1557 & w1558 ) ;
  assign w1560 = \pi169 ^ w1256 ;
  assign w1561 = ( \pi041 & \pi169 ) | ( \pi041 & w1560 ) | ( \pi169 & w1560 ) ;
  assign w1562 = ( ~\pi297 & w1260 ) | ( ~\pi297 & w1561 ) | ( w1260 & w1561 ) ;
  assign w1563 = ( \pi425 & w1260 ) | ( \pi425 & ~w1561 ) | ( w1260 & ~w1561 ) ;
  assign w1564 = ~w1562 & w1563 ;
  assign w1565 = \pi168 ^ w1256 ;
  assign w1566 = ( \pi040 & \pi168 ) | ( \pi040 & w1565 ) | ( \pi168 & w1565 ) ;
  assign w1567 = \pi424 ^ w1260 ;
  assign w1568 = ( \pi296 & \pi424 ) | ( \pi296 & w1567 ) | ( \pi424 & w1567 ) ;
  assign w1569 = w1566 & ~w1568 ;
  assign w1570 = \pi425 ^ w1260 ;
  assign w1571 = ( \pi297 & \pi425 ) | ( \pi297 & w1570 ) | ( \pi425 & w1570 ) ;
  assign w1572 = ( w1561 & w1569 ) | ( w1561 & ~w1571 ) | ( w1569 & ~w1571 ) ;
  assign w1573 = ~w1548 & w1550 ;
  assign w1574 = ( w1554 & ~w1556 ) | ( w1554 & w1572 ) | ( ~w1556 & w1572 ) ;
  assign w1575 = w1548 | w1552 ;
  assign w1576 = ( w1573 & w1574 ) | ( w1573 & ~w1575 ) | ( w1574 & ~w1575 ) ;
  assign w1577 = w1536 & ~w1538 ;
  assign w1578 = \pi429 ^ w1260 ;
  assign w1579 = ( \pi301 & \pi429 ) | ( \pi301 & w1578 ) | ( \pi429 & w1578 ) ;
  assign w1580 = ( w1540 & w1577 ) | ( w1540 & ~w1579 ) | ( w1577 & ~w1579 ) ;
  assign w1581 = \pi160 ^ w1256 ;
  assign w1582 = ( \pi032 & \pi160 ) | ( \pi032 & w1581 ) | ( \pi160 & w1581 ) ;
  assign w1583 = ( ~\pi288 & w1260 ) | ( ~\pi288 & w1582 ) | ( w1260 & w1582 ) ;
  assign w1584 = ( \pi416 & w1260 ) | ( \pi416 & ~w1582 ) | ( w1260 & ~w1582 ) ;
  assign w1585 = ~w1583 & w1584 ;
  assign w1586 = \pi159 ^ w1256 ;
  assign w1587 = ( \pi031 & \pi159 ) | ( \pi031 & w1586 ) | ( \pi159 & w1586 ) ;
  assign w1588 = \pi158 ^ w1256 ;
  assign w1589 = ( \pi030 & \pi158 ) | ( \pi030 & w1588 ) | ( \pi158 & w1588 ) ;
  assign w1590 = \pi157 ^ w1256 ;
  assign w1591 = ( \pi029 & \pi157 ) | ( \pi029 & w1590 ) | ( \pi157 & w1590 ) ;
  assign w1592 = \pi156 ^ w1256 ;
  assign w1593 = ( \pi028 & \pi156 ) | ( \pi028 & w1592 ) | ( \pi156 & w1592 ) ;
  assign w1594 = \pi155 ^ w1256 ;
  assign w1595 = ( \pi027 & \pi155 ) | ( \pi027 & w1594 ) | ( \pi155 & w1594 ) ;
  assign w1596 = \pi154 ^ w1256 ;
  assign w1597 = ( \pi026 & \pi154 ) | ( \pi026 & w1596 ) | ( \pi154 & w1596 ) ;
  assign w1598 = \pi410 ^ w1260 ;
  assign w1599 = ( \pi282 & \pi410 ) | ( \pi282 & w1598 ) | ( \pi410 & w1598 ) ;
  assign w1600 = \pi409 ^ w1260 ;
  assign w1601 = ( \pi281 & \pi409 ) | ( \pi281 & w1600 ) | ( \pi409 & w1600 ) ;
  assign w1602 = \pi151 ^ w1256 ;
  assign w1603 = ( \pi023 & \pi151 ) | ( \pi023 & w1602 ) | ( \pi151 & w1602 ) ;
  assign w1604 = \pi150 ^ w1256 ;
  assign w1605 = ( \pi022 & \pi150 ) | ( \pi022 & w1604 ) | ( \pi150 & w1604 ) ;
  assign w1606 = \pi149 ^ w1256 ;
  assign w1607 = ( \pi021 & \pi149 ) | ( \pi021 & w1606 ) | ( \pi149 & w1606 ) ;
  assign w1608 = \pi148 ^ w1256 ;
  assign w1609 = ( \pi020 & \pi148 ) | ( \pi020 & w1608 ) | ( \pi148 & w1608 ) ;
  assign w1610 = \pi147 ^ w1256 ;
  assign w1611 = ( \pi019 & \pi147 ) | ( \pi019 & w1610 ) | ( \pi147 & w1610 ) ;
  assign w1612 = \pi146 ^ w1256 ;
  assign w1613 = ( \pi018 & \pi146 ) | ( \pi018 & w1612 ) | ( \pi146 & w1612 ) ;
  assign w1614 = \pi402 ^ w1260 ;
  assign w1615 = ( \pi274 & \pi402 ) | ( \pi274 & w1614 ) | ( \pi402 & w1614 ) ;
  assign w1616 = \pi401 ^ w1260 ;
  assign w1617 = ( \pi273 & \pi401 ) | ( \pi273 & w1616 ) | ( \pi401 & w1616 ) ;
  assign w1618 = \pi143 ^ w1256 ;
  assign w1619 = ( \pi015 & \pi143 ) | ( \pi015 & w1618 ) | ( \pi143 & w1618 ) ;
  assign w1620 = \pi142 ^ w1256 ;
  assign w1621 = ( \pi014 & \pi142 ) | ( \pi014 & w1620 ) | ( \pi142 & w1620 ) ;
  assign w1622 = \pi141 ^ w1256 ;
  assign w1623 = ( \pi013 & \pi141 ) | ( \pi013 & w1622 ) | ( \pi141 & w1622 ) ;
  assign w1624 = \pi140 ^ w1256 ;
  assign w1625 = ( \pi012 & \pi140 ) | ( \pi012 & w1624 ) | ( \pi140 & w1624 ) ;
  assign w1626 = \pi139 ^ w1256 ;
  assign w1627 = ( \pi011 & \pi139 ) | ( \pi011 & w1626 ) | ( \pi139 & w1626 ) ;
  assign w1628 = \pi138 ^ w1256 ;
  assign w1629 = ( \pi010 & \pi138 ) | ( \pi010 & w1628 ) | ( \pi138 & w1628 ) ;
  assign w1630 = \pi394 ^ w1260 ;
  assign w1631 = ( \pi266 & \pi394 ) | ( \pi266 & w1630 ) | ( \pi394 & w1630 ) ;
  assign w1632 = \pi393 ^ w1260 ;
  assign w1633 = ( \pi265 & \pi393 ) | ( \pi265 & w1632 ) | ( \pi393 & w1632 ) ;
  assign w1634 = \pi135 ^ w1256 ;
  assign w1635 = ( \pi007 & \pi135 ) | ( \pi007 & w1634 ) | ( \pi135 & w1634 ) ;
  assign w1636 = \pi134 ^ w1256 ;
  assign w1637 = ( \pi006 & \pi134 ) | ( \pi006 & w1636 ) | ( \pi134 & w1636 ) ;
  assign w1638 = \pi133 ^ w1256 ;
  assign w1639 = ( \pi005 & \pi133 ) | ( \pi005 & w1638 ) | ( \pi133 & w1638 ) ;
  assign w1640 = \pi132 ^ w1256 ;
  assign w1641 = ( \pi004 & \pi132 ) | ( \pi004 & w1640 ) | ( \pi132 & w1640 ) ;
  assign w1642 = \pi131 ^ w1256 ;
  assign w1643 = ( \pi003 & \pi131 ) | ( \pi003 & w1642 ) | ( \pi131 & w1642 ) ;
  assign w1644 = \pi385 ^ w1260 ;
  assign w1645 = ( \pi257 & \pi385 ) | ( \pi257 & w1644 ) | ( \pi385 & w1644 ) ;
  assign w1646 = \pi128 ^ w1256 ;
  assign w1647 = ( \pi000 & \pi128 ) | ( \pi000 & w1646 ) | ( \pi128 & w1646 ) ;
  assign w1648 = ( \pi256 & w1260 ) | ( \pi256 & ~w1647 ) | ( w1260 & ~w1647 ) ;
  assign w1649 = ( ~\pi384 & w1260 ) | ( ~\pi384 & w1647 ) | ( w1260 & w1647 ) ;
  assign w1650 = ~w1648 & w1649 ;
  assign w1651 = \pi129 ^ w1256 ;
  assign w1652 = ( \pi001 & \pi129 ) | ( \pi001 & w1651 ) | ( \pi129 & w1651 ) ;
  assign w1653 = \pi130 ^ w1256 ;
  assign w1654 = ( \pi002 & \pi130 ) | ( \pi002 & w1653 ) | ( \pi130 & w1653 ) ;
  assign w1655 = \pi386 ^ w1260 ;
  assign w1656 = ( \pi258 & \pi386 ) | ( \pi258 & w1655 ) | ( \pi386 & w1655 ) ;
  assign w1657 = ( ~w1645 & w1650 ) | ( ~w1645 & w1652 ) | ( w1650 & w1652 ) ;
  assign w1658 = ( w1654 & ~w1656 ) | ( w1654 & w1657 ) | ( ~w1656 & w1657 ) ;
  assign w1659 = \pi259 ^ w1260 ;
  assign w1660 = ( \pi259 & \pi387 ) | ( \pi259 & ~w1659 ) | ( \pi387 & ~w1659 ) ;
  assign w1661 = ( w1643 & w1658 ) | ( w1643 & ~w1660 ) | ( w1658 & ~w1660 ) ;
  assign w1662 = \pi260 ^ w1260 ;
  assign w1663 = ( \pi260 & \pi388 ) | ( \pi260 & ~w1662 ) | ( \pi388 & ~w1662 ) ;
  assign w1664 = ( w1641 & w1661 ) | ( w1641 & ~w1663 ) | ( w1661 & ~w1663 ) ;
  assign w1665 = \pi261 ^ w1260 ;
  assign w1666 = ( \pi261 & \pi389 ) | ( \pi261 & ~w1665 ) | ( \pi389 & ~w1665 ) ;
  assign w1667 = ( w1639 & w1664 ) | ( w1639 & ~w1666 ) | ( w1664 & ~w1666 ) ;
  assign w1668 = \pi262 ^ w1260 ;
  assign w1669 = ( \pi262 & \pi390 ) | ( \pi262 & ~w1668 ) | ( \pi390 & ~w1668 ) ;
  assign w1670 = ( w1637 & w1667 ) | ( w1637 & ~w1669 ) | ( w1667 & ~w1669 ) ;
  assign w1671 = \pi263 ^ w1260 ;
  assign w1672 = ( \pi263 & \pi391 ) | ( \pi263 & ~w1671 ) | ( \pi391 & ~w1671 ) ;
  assign w1673 = ( w1635 & w1670 ) | ( w1635 & ~w1672 ) | ( w1670 & ~w1672 ) ;
  assign w1674 = \pi136 ^ w1256 ;
  assign w1675 = ( \pi008 & \pi136 ) | ( \pi008 & w1674 ) | ( \pi136 & w1674 ) ;
  assign w1676 = \pi264 ^ w1260 ;
  assign w1677 = ( \pi264 & \pi392 ) | ( \pi264 & ~w1676 ) | ( \pi392 & ~w1676 ) ;
  assign w1678 = ( w1673 & w1675 ) | ( w1673 & ~w1677 ) | ( w1675 & ~w1677 ) ;
  assign w1679 = \pi137 ^ w1256 ;
  assign w1680 = ( \pi009 & \pi137 ) | ( \pi009 & w1679 ) | ( \pi137 & w1679 ) ;
  assign w1681 = ( ~w1633 & w1678 ) | ( ~w1633 & w1680 ) | ( w1678 & w1680 ) ;
  assign w1682 = ( w1629 & ~w1631 ) | ( w1629 & w1681 ) | ( ~w1631 & w1681 ) ;
  assign w1683 = \pi267 ^ w1260 ;
  assign w1684 = ( \pi267 & \pi395 ) | ( \pi267 & ~w1683 ) | ( \pi395 & ~w1683 ) ;
  assign w1685 = ( w1627 & w1682 ) | ( w1627 & ~w1684 ) | ( w1682 & ~w1684 ) ;
  assign w1686 = \pi268 ^ w1260 ;
  assign w1687 = ( \pi268 & \pi396 ) | ( \pi268 & ~w1686 ) | ( \pi396 & ~w1686 ) ;
  assign w1688 = ( w1625 & w1685 ) | ( w1625 & ~w1687 ) | ( w1685 & ~w1687 ) ;
  assign w1689 = \pi269 ^ w1260 ;
  assign w1690 = ( \pi269 & \pi397 ) | ( \pi269 & ~w1689 ) | ( \pi397 & ~w1689 ) ;
  assign w1691 = ( w1623 & w1688 ) | ( w1623 & ~w1690 ) | ( w1688 & ~w1690 ) ;
  assign w1692 = \pi270 ^ w1260 ;
  assign w1693 = ( \pi270 & \pi398 ) | ( \pi270 & ~w1692 ) | ( \pi398 & ~w1692 ) ;
  assign w1694 = ( w1621 & w1691 ) | ( w1621 & ~w1693 ) | ( w1691 & ~w1693 ) ;
  assign w1695 = \pi271 ^ w1260 ;
  assign w1696 = ( \pi271 & \pi399 ) | ( \pi271 & ~w1695 ) | ( \pi399 & ~w1695 ) ;
  assign w1697 = ( w1619 & w1694 ) | ( w1619 & ~w1696 ) | ( w1694 & ~w1696 ) ;
  assign w1698 = \pi144 ^ w1256 ;
  assign w1699 = ( \pi016 & \pi144 ) | ( \pi016 & w1698 ) | ( \pi144 & w1698 ) ;
  assign w1700 = \pi272 ^ w1260 ;
  assign w1701 = ( \pi272 & \pi400 ) | ( \pi272 & ~w1700 ) | ( \pi400 & ~w1700 ) ;
  assign w1702 = ( w1697 & w1699 ) | ( w1697 & ~w1701 ) | ( w1699 & ~w1701 ) ;
  assign w1703 = \pi145 ^ w1256 ;
  assign w1704 = ( \pi017 & \pi145 ) | ( \pi017 & w1703 ) | ( \pi145 & w1703 ) ;
  assign w1705 = ( ~w1617 & w1702 ) | ( ~w1617 & w1704 ) | ( w1702 & w1704 ) ;
  assign w1706 = ( w1613 & ~w1615 ) | ( w1613 & w1705 ) | ( ~w1615 & w1705 ) ;
  assign w1707 = \pi275 ^ w1260 ;
  assign w1708 = ( \pi275 & \pi403 ) | ( \pi275 & ~w1707 ) | ( \pi403 & ~w1707 ) ;
  assign w1709 = ( w1611 & w1706 ) | ( w1611 & ~w1708 ) | ( w1706 & ~w1708 ) ;
  assign w1710 = \pi276 ^ w1260 ;
  assign w1711 = ( \pi276 & \pi404 ) | ( \pi276 & ~w1710 ) | ( \pi404 & ~w1710 ) ;
  assign w1712 = ( w1609 & w1709 ) | ( w1609 & ~w1711 ) | ( w1709 & ~w1711 ) ;
  assign w1713 = \pi277 ^ w1260 ;
  assign w1714 = ( \pi277 & \pi405 ) | ( \pi277 & ~w1713 ) | ( \pi405 & ~w1713 ) ;
  assign w1715 = ( w1607 & w1712 ) | ( w1607 & ~w1714 ) | ( w1712 & ~w1714 ) ;
  assign w1716 = \pi278 ^ w1260 ;
  assign w1717 = ( \pi278 & \pi406 ) | ( \pi278 & ~w1716 ) | ( \pi406 & ~w1716 ) ;
  assign w1718 = ( w1605 & w1715 ) | ( w1605 & ~w1717 ) | ( w1715 & ~w1717 ) ;
  assign w1719 = \pi279 ^ w1260 ;
  assign w1720 = ( \pi279 & \pi407 ) | ( \pi279 & ~w1719 ) | ( \pi407 & ~w1719 ) ;
  assign w1721 = ( w1603 & w1718 ) | ( w1603 & ~w1720 ) | ( w1718 & ~w1720 ) ;
  assign w1722 = \pi152 ^ w1256 ;
  assign w1723 = ( \pi024 & \pi152 ) | ( \pi024 & w1722 ) | ( \pi152 & w1722 ) ;
  assign w1724 = \pi280 ^ w1260 ;
  assign w1725 = ( \pi280 & \pi408 ) | ( \pi280 & ~w1724 ) | ( \pi408 & ~w1724 ) ;
  assign w1726 = ( w1721 & w1723 ) | ( w1721 & ~w1725 ) | ( w1723 & ~w1725 ) ;
  assign w1727 = \pi153 ^ w1256 ;
  assign w1728 = ( \pi025 & \pi153 ) | ( \pi025 & w1727 ) | ( \pi153 & w1727 ) ;
  assign w1729 = ( ~w1601 & w1726 ) | ( ~w1601 & w1728 ) | ( w1726 & w1728 ) ;
  assign w1730 = ( w1597 & ~w1599 ) | ( w1597 & w1729 ) | ( ~w1599 & w1729 ) ;
  assign w1731 = \pi283 ^ w1260 ;
  assign w1732 = ( \pi283 & \pi411 ) | ( \pi283 & ~w1731 ) | ( \pi411 & ~w1731 ) ;
  assign w1733 = ( w1595 & w1730 ) | ( w1595 & ~w1732 ) | ( w1730 & ~w1732 ) ;
  assign w1734 = \pi284 ^ w1260 ;
  assign w1735 = ( \pi284 & \pi412 ) | ( \pi284 & ~w1734 ) | ( \pi412 & ~w1734 ) ;
  assign w1736 = ( w1593 & w1733 ) | ( w1593 & ~w1735 ) | ( w1733 & ~w1735 ) ;
  assign w1737 = \pi285 ^ w1260 ;
  assign w1738 = ( \pi285 & \pi413 ) | ( \pi285 & ~w1737 ) | ( \pi413 & ~w1737 ) ;
  assign w1739 = ( w1591 & w1736 ) | ( w1591 & ~w1738 ) | ( w1736 & ~w1738 ) ;
  assign w1740 = \pi286 ^ w1260 ;
  assign w1741 = ( \pi286 & \pi414 ) | ( \pi286 & ~w1740 ) | ( \pi414 & ~w1740 ) ;
  assign w1742 = ( w1589 & w1739 ) | ( w1589 & ~w1741 ) | ( w1739 & ~w1741 ) ;
  assign w1743 = \pi287 ^ w1260 ;
  assign w1744 = ( \pi287 & \pi415 ) | ( \pi287 & ~w1743 ) | ( \pi415 & ~w1743 ) ;
  assign w1745 = ( w1587 & w1742 ) | ( w1587 & ~w1744 ) | ( w1742 & ~w1744 ) ;
  assign w1746 = \pi167 ^ w1256 ;
  assign w1747 = ( \pi039 & \pi167 ) | ( \pi039 & w1746 ) | ( \pi167 & w1746 ) ;
  assign w1748 = \pi423 ^ w1260 ;
  assign w1749 = ( \pi295 & \pi423 ) | ( \pi295 & w1748 ) | ( \pi423 & w1748 ) ;
  assign w1750 = \pi422 ^ w1260 ;
  assign w1751 = ( \pi294 & \pi422 ) | ( \pi294 & w1750 ) | ( \pi422 & w1750 ) ;
  assign w1752 = \pi166 ^ w1256 ;
  assign w1753 = ( \pi038 & \pi166 ) | ( \pi038 & w1752 ) | ( \pi166 & w1752 ) ;
  assign w1754 = \pi164 ^ w1256 ;
  assign w1755 = ( \pi036 & \pi164 ) | ( \pi036 & w1754 ) | ( \pi164 & w1754 ) ;
  assign w1756 = \pi420 ^ w1260 ;
  assign w1757 = ( \pi292 & \pi420 ) | ( \pi292 & w1756 ) | ( \pi420 & w1756 ) ;
  assign w1758 = \pi165 ^ w1256 ;
  assign w1759 = ( \pi037 & \pi165 ) | ( \pi037 & w1758 ) | ( \pi165 & w1758 ) ;
  assign w1760 = w1260 | w1759 ;
  assign w1761 = \pi421 | w1760 ;
  assign w1762 = ~w1755 & w1757 ;
  assign w1763 = ( ~\pi293 & w1759 ) | ( ~\pi293 & w1760 ) | ( w1759 & w1760 ) ;
  assign w1764 = ( w1761 & w1762 ) | ( w1761 & ~w1763 ) | ( w1762 & ~w1763 ) ;
  assign w1765 = w1747 & w1749 ;
  assign w1766 = w1751 & w1753 ;
  assign w1767 = ( w1751 & w1764 ) | ( w1751 & ~w1766 ) | ( w1764 & ~w1766 ) ;
  assign w1768 = ( w1749 & ~w1765 ) | ( w1749 & w1767 ) | ( ~w1765 & w1767 ) ;
  assign w1769 = \pi161 ^ w1256 ;
  assign w1770 = ( \pi033 & \pi161 ) | ( \pi033 & w1769 ) | ( \pi161 & w1769 ) ;
  assign w1771 = \pi417 ^ w1260 ;
  assign w1772 = ( \pi289 & \pi417 ) | ( \pi289 & w1771 ) | ( \pi417 & w1771 ) ;
  assign w1773 = \pi163 ^ w1256 ;
  assign w1774 = ( \pi035 & \pi163 ) | ( \pi035 & w1773 ) | ( \pi163 & w1773 ) ;
  assign w1775 = ( ~\pi291 & w1260 ) | ( ~\pi291 & w1774 ) | ( w1260 & w1774 ) ;
  assign w1776 = ( \pi419 & w1260 ) | ( \pi419 & ~w1774 ) | ( w1260 & ~w1774 ) ;
  assign w1777 = ~w1775 & w1776 ;
  assign w1778 = \pi418 ^ w1260 ;
  assign w1779 = ( \pi290 & \pi418 ) | ( \pi290 & w1778 ) | ( \pi418 & w1778 ) ;
  assign w1780 = \pi162 ^ w1256 ;
  assign w1781 = ( \pi034 & \pi162 ) | ( \pi034 & w1780 ) | ( \pi162 & w1780 ) ;
  assign w1782 = w1770 & w1772 ;
  assign w1783 = w1779 & w1781 ;
  assign w1784 = ( w1777 & w1779 ) | ( w1777 & ~w1783 ) | ( w1779 & ~w1783 ) ;
  assign w1785 = ( w1772 & ~w1782 ) | ( w1772 & w1784 ) | ( ~w1782 & w1784 ) ;
  assign w1786 = w1755 & ~w1757 ;
  assign w1787 = \pi421 ^ w1260 ;
  assign w1788 = ( \pi293 & \pi421 ) | ( \pi293 & w1787 ) | ( \pi421 & w1787 ) ;
  assign w1789 = ( w1759 & w1786 ) | ( w1759 & ~w1788 ) | ( w1786 & ~w1788 ) ;
  assign w1790 = ~w1260 & w1582 ;
  assign w1791 = \pi416 & w1790 ;
  assign w1792 = w1770 & ~w1772 ;
  assign w1793 = ( ~\pi288 & w1582 ) | ( ~\pi288 & w1790 ) | ( w1582 & w1790 ) ;
  assign w1794 = ( ~w1791 & w1792 ) | ( ~w1791 & w1793 ) | ( w1792 & w1793 ) ;
  assign w1795 = w1785 & w1794 ;
  assign w1796 = ~w1779 & w1781 ;
  assign w1797 = ~w1777 & w1796 ;
  assign w1798 = ( w1794 & ~w1795 ) | ( w1794 & w1797 ) | ( ~w1795 & w1797 ) ;
  assign w1799 = w1774 & ~w1798 ;
  assign w1800 = ( \pi291 & w1260 ) | ( \pi291 & ~w1799 ) | ( w1260 & ~w1799 ) ;
  assign w1801 = ( ~\pi419 & w1260 ) | ( ~\pi419 & w1799 ) | ( w1260 & w1799 ) ;
  assign w1802 = ~w1800 & w1801 ;
  assign w1803 = ( ~w1768 & w1798 ) | ( ~w1768 & w1802 ) | ( w1798 & w1802 ) ;
  assign w1804 = w1747 | w1803 ;
  assign w1805 = ( ~w1751 & w1753 ) | ( ~w1751 & w1789 ) | ( w1753 & w1789 ) ;
  assign w1806 = w1749 & ~w1803 ;
  assign w1807 = ( w1804 & w1805 ) | ( w1804 & ~w1806 ) | ( w1805 & ~w1806 ) ;
  assign w1808 = w1745 & ~w1768 ;
  assign w1809 = w1585 | w1785 ;
  assign w1810 = w1808 & ~w1809 ;
  assign w1811 = w1807 | w1810 ;
  assign w1812 = w1548 | w1559 ;
  assign w1813 = ( ~w1566 & w1568 ) | ( ~w1566 & w1812 ) | ( w1568 & w1812 ) ;
  assign w1814 = ( w1564 & ~w1812 ) | ( w1564 & w1813 ) | ( ~w1812 & w1813 ) ;
  assign w1815 = w1812 | w1814 ;
  assign w1816 = w1811 & ~w1815 ;
  assign w1817 = ~w1530 & w1580 ;
  assign w1818 = ( w1530 & w1532 ) | ( w1530 & ~w1816 ) | ( w1532 & ~w1816 ) ;
  assign w1819 = ( w1534 & w1817 ) | ( w1534 & ~w1818 ) | ( w1817 & ~w1818 ) ;
  assign w1820 = w1816 | w1819 ;
  assign w1821 = \pi176 ^ w1256 ;
  assign w1822 = ( \pi048 & \pi176 ) | ( \pi048 & w1821 ) | ( \pi176 & w1821 ) ;
  assign w1823 = \pi183 ^ w1256 ;
  assign w1824 = ( \pi055 & \pi183 ) | ( \pi055 & w1823 ) | ( \pi183 & w1823 ) ;
  assign w1825 = \pi439 ^ w1260 ;
  assign w1826 = ( \pi311 & \pi439 ) | ( \pi311 & w1825 ) | ( \pi439 & w1825 ) ;
  assign w1827 = \pi438 ^ w1260 ;
  assign w1828 = ( \pi310 & \pi438 ) | ( \pi310 & w1827 ) | ( \pi438 & w1827 ) ;
  assign w1829 = \pi182 ^ w1256 ;
  assign w1830 = ( \pi054 & \pi182 ) | ( \pi054 & w1829 ) | ( \pi182 & w1829 ) ;
  assign w1831 = \pi181 ^ w1256 ;
  assign w1832 = ( \pi053 & \pi181 ) | ( \pi053 & w1831 ) | ( \pi181 & w1831 ) ;
  assign w1833 = \pi436 ^ w1260 ;
  assign w1834 = ( \pi308 & \pi436 ) | ( \pi308 & w1833 ) | ( \pi436 & w1833 ) ;
  assign w1835 = \pi180 ^ w1256 ;
  assign w1836 = ( \pi052 & \pi180 ) | ( \pi052 & w1835 ) | ( \pi180 & w1835 ) ;
  assign w1837 = w1260 | w1832 ;
  assign w1838 = \pi437 | w1837 ;
  assign w1839 = w1834 & ~w1836 ;
  assign w1840 = ( ~\pi309 & w1832 ) | ( ~\pi309 & w1837 ) | ( w1832 & w1837 ) ;
  assign w1841 = ( w1838 & w1839 ) | ( w1838 & ~w1840 ) | ( w1839 & ~w1840 ) ;
  assign w1842 = w1824 & w1826 ;
  assign w1843 = w1828 & w1830 ;
  assign w1844 = ( w1828 & w1841 ) | ( w1828 & ~w1843 ) | ( w1841 & ~w1843 ) ;
  assign w1845 = ( w1826 & ~w1842 ) | ( w1826 & w1844 ) | ( ~w1842 & w1844 ) ;
  assign w1846 = \pi177 ^ w1256 ;
  assign w1847 = ( \pi049 & \pi177 ) | ( \pi049 & w1846 ) | ( \pi177 & w1846 ) ;
  assign w1848 = \pi433 ^ w1260 ;
  assign w1849 = ( \pi305 & \pi433 ) | ( \pi305 & w1848 ) | ( \pi433 & w1848 ) ;
  assign w1850 = \pi179 ^ w1256 ;
  assign w1851 = ( \pi051 & \pi179 ) | ( \pi051 & w1850 ) | ( \pi179 & w1850 ) ;
  assign w1852 = ( ~\pi307 & w1260 ) | ( ~\pi307 & w1851 ) | ( w1260 & w1851 ) ;
  assign w1853 = ( \pi435 & w1260 ) | ( \pi435 & ~w1851 ) | ( w1260 & ~w1851 ) ;
  assign w1854 = ~w1852 & w1853 ;
  assign w1855 = \pi434 ^ w1260 ;
  assign w1856 = ( \pi306 & \pi434 ) | ( \pi306 & w1855 ) | ( \pi434 & w1855 ) ;
  assign w1857 = \pi178 ^ w1256 ;
  assign w1858 = ( \pi050 & \pi178 ) | ( \pi050 & w1857 ) | ( \pi178 & w1857 ) ;
  assign w1859 = w1847 | w1849 ;
  assign w1860 = ( ~w1845 & w1856 ) | ( ~w1845 & w1858 ) | ( w1856 & w1858 ) ;
  assign w1861 = ( w1854 & ~w1858 ) | ( w1854 & w1860 ) | ( ~w1858 & w1860 ) ;
  assign w1862 = w1845 | w1861 ;
  assign w1863 = ( ~w1847 & w1859 ) | ( ~w1847 & w1862 ) | ( w1859 & w1862 ) ;
  assign w1864 = ~\pi304 & w1260 ;
  assign w1865 = \pi432 | w1260 ;
  assign w1866 = ( ~w1822 & w1863 ) | ( ~w1822 & w1865 ) | ( w1863 & w1865 ) ;
  assign w1867 = ( w1863 & ~w1864 ) | ( w1863 & w1866 ) | ( ~w1864 & w1866 ) ;
  assign w1868 = ( \pi304 & w1260 ) | ( \pi304 & ~w1822 ) | ( w1260 & ~w1822 ) ;
  assign w1869 = ( ~\pi432 & w1260 ) | ( ~\pi432 & w1822 ) | ( w1260 & w1822 ) ;
  assign w1870 = ~w1868 & w1869 ;
  assign w1871 = w1854 | w1856 ;
  assign w1872 = ( w1847 & ~w1849 ) | ( w1847 & w1870 ) | ( ~w1849 & w1870 ) ;
  assign w1873 = ~w1854 & w1858 ;
  assign w1874 = ( ~w1871 & w1872 ) | ( ~w1871 & w1873 ) | ( w1872 & w1873 ) ;
  assign w1875 = w1851 & ~w1874 ;
  assign w1876 = ( \pi307 & w1260 ) | ( \pi307 & ~w1875 ) | ( w1260 & ~w1875 ) ;
  assign w1877 = ( ~\pi435 & w1260 ) | ( ~\pi435 & w1875 ) | ( w1260 & w1875 ) ;
  assign w1878 = ~w1876 & w1877 ;
  assign w1879 = ( ~w1845 & w1874 ) | ( ~w1845 & w1878 ) | ( w1874 & w1878 ) ;
  assign w1880 = ~w1834 & w1836 ;
  assign w1881 = \pi437 ^ w1260 ;
  assign w1882 = ( \pi309 & \pi437 ) | ( \pi309 & w1881 ) | ( \pi437 & w1881 ) ;
  assign w1883 = ( w1832 & w1880 ) | ( w1832 & ~w1882 ) | ( w1880 & ~w1882 ) ;
  assign w1884 = w1824 | w1879 ;
  assign w1885 = ( ~w1828 & w1830 ) | ( ~w1828 & w1883 ) | ( w1830 & w1883 ) ;
  assign w1886 = w1826 & ~w1879 ;
  assign w1887 = ( w1884 & w1885 ) | ( w1884 & ~w1886 ) | ( w1885 & ~w1886 ) ;
  assign w1888 = w1867 & ~w1887 ;
  assign w1889 = ( w1527 & w1529 ) | ( w1527 & ~w1888 ) | ( w1529 & ~w1888 ) ;
  assign w1890 = ( ~w1529 & w1820 ) | ( ~w1529 & w1889 ) | ( w1820 & w1889 ) ;
  assign w1891 = ( w1576 & w1887 ) | ( w1576 & ~w1888 ) | ( w1887 & ~w1888 ) ;
  assign w1892 = ( ~w1888 & w1890 ) | ( ~w1888 & w1891 ) | ( w1890 & w1891 ) ;
  assign w1893 = w1509 & w1511 ;
  assign w1894 = w1513 | w1515 ;
  assign w1895 = ( w1499 & ~w1513 ) | ( w1499 & w1894 ) | ( ~w1513 & w1894 ) ;
  assign w1896 = ( w1511 & ~w1893 ) | ( w1511 & w1895 ) | ( ~w1893 & w1895 ) ;
  assign w1897 = w1501 | w1503 ;
  assign w1898 = ( w1505 & w1507 ) | ( w1505 & ~w1892 ) | ( w1507 & ~w1892 ) ;
  assign w1899 = ( w1507 & w1896 ) | ( w1507 & ~w1898 ) | ( w1896 & ~w1898 ) ;
  assign w1900 = w1892 & ~w1899 ;
  assign w1901 = ( w1501 & ~w1897 ) | ( w1501 & w1900 ) | ( ~w1897 & w1900 ) ;
  assign w1902 = w1481 & ~w1521 ;
  assign w1903 = ( ~w1483 & w1485 ) | ( ~w1483 & w1525 ) | ( w1485 & w1525 ) ;
  assign w1904 = ( w1521 & ~w1902 ) | ( w1521 & w1903 ) | ( ~w1902 & w1903 ) ;
  assign w1905 = w1901 | w1904 ;
  assign w1906 = \pi319 & w1260 ;
  assign w1907 = \pi447 & ~w1260 ;
  assign w1908 = ( w1478 & w1905 ) | ( w1478 & ~w1907 ) | ( w1905 & ~w1907 ) ;
  assign w1909 = ( w1905 & ~w1906 ) | ( w1905 & w1908 ) | ( ~w1906 & w1908 ) ;
  assign w1910 = ~\pi321 & w1260 ;
  assign w1911 = \pi449 | w1260 ;
  assign w1912 = ( w1476 & w1909 ) | ( w1476 & ~w1911 ) | ( w1909 & ~w1911 ) ;
  assign w1913 = ( w1909 & w1910 ) | ( w1909 & w1912 ) | ( w1910 & w1912 ) ;
  assign w1914 = ( ~w1472 & w1474 ) | ( ~w1472 & w1913 ) | ( w1474 & w1913 ) ;
  assign w1915 = w1913 & w1914 ;
  assign w1916 = ~w1472 & w1474 ;
  assign w1917 = \pi449 ^ w1260 ;
  assign w1918 = ( \pi321 & \pi449 ) | ( \pi321 & w1917 ) | ( \pi449 & w1917 ) ;
  assign w1919 = ( w1476 & w1916 ) | ( w1476 & ~w1918 ) | ( w1916 & ~w1918 ) ;
  assign w1920 = w1915 | w1919 ;
  assign w1921 = ( ~w1468 & w1470 ) | ( ~w1468 & w1920 ) | ( w1470 & w1920 ) ;
  assign w1922 = ( w1464 & ~w1466 ) | ( w1464 & w1921 ) | ( ~w1466 & w1921 ) ;
  assign w1923 = w1458 & w1460 ;
  assign w1924 = ~w1454 & w1456 ;
  assign w1925 = ( w1460 & ~w1923 ) | ( w1460 & w1924 ) | ( ~w1923 & w1924 ) ;
  assign w1926 = ~w1446 & w1448 ;
  assign w1927 = ( w1922 & ~w1925 ) | ( w1922 & w1926 ) | ( ~w1925 & w1926 ) ;
  assign w1928 = ( ~w1450 & w1452 ) | ( ~w1450 & w1927 ) | ( w1452 & w1927 ) ;
  assign w1929 = ~w1926 & w1928 ;
  assign w1930 = ( ~w1450 & w1452 ) | ( ~w1450 & w1462 ) | ( w1452 & w1462 ) ;
  assign w1931 = ( w1462 & w1929 ) | ( w1462 & w1930 ) | ( w1929 & w1930 ) ;
  assign w1932 = ( w1446 & ~w1448 ) | ( w1446 & w1931 ) | ( ~w1448 & w1931 ) ;
  assign w1933 = w1929 | w1932 ;
  assign w1934 = \pi203 ^ w1256 ;
  assign w1935 = ( \pi075 & \pi203 ) | ( \pi075 & w1934 ) | ( \pi203 & w1934 ) ;
  assign w1936 = \pi459 ^ w1260 ;
  assign w1937 = ( \pi331 & \pi459 ) | ( \pi331 & w1936 ) | ( \pi459 & w1936 ) ;
  assign w1938 = \pi458 ^ w1260 ;
  assign w1939 = ( \pi330 & \pi458 ) | ( \pi330 & w1938 ) | ( \pi458 & w1938 ) ;
  assign w1940 = \pi202 ^ w1256 ;
  assign w1941 = ( \pi074 & \pi202 ) | ( \pi074 & w1940 ) | ( \pi202 & w1940 ) ;
  assign w1942 = w1939 | w1941 ;
  assign w1943 = ~w1935 & w1937 ;
  assign w1944 = ( ~w1941 & w1942 ) | ( ~w1941 & w1943 ) | ( w1942 & w1943 ) ;
  assign w1945 = \pi201 ^ w1256 ;
  assign w1946 = ( \pi073 & \pi201 ) | ( \pi073 & w1945 ) | ( \pi201 & w1945 ) ;
  assign w1947 = ( ~\pi329 & w1260 ) | ( ~\pi329 & w1946 ) | ( w1260 & w1946 ) ;
  assign w1948 = ( \pi457 & w1260 ) | ( \pi457 & ~w1946 ) | ( w1260 & ~w1946 ) ;
  assign w1949 = ~w1947 & w1948 ;
  assign w1950 = \pi456 ^ w1260 ;
  assign w1951 = ( \pi328 & \pi456 ) | ( \pi328 & w1950 ) | ( \pi456 & w1950 ) ;
  assign w1952 = \pi200 ^ w1256 ;
  assign w1953 = ( \pi072 & \pi200 ) | ( \pi072 & w1952 ) | ( \pi200 & w1952 ) ;
  assign w1954 = w1933 & ~w1944 ;
  assign w1955 = ( ~w1951 & w1953 ) | ( ~w1951 & w1954 ) | ( w1953 & w1954 ) ;
  assign w1956 = ( w1949 & w1954 ) | ( w1949 & ~w1955 ) | ( w1954 & ~w1955 ) ;
  assign w1957 = w1954 & ~w1956 ;
  assign w1958 = ~w1951 & w1953 ;
  assign w1959 = \pi457 ^ w1260 ;
  assign w1960 = ( \pi329 & \pi457 ) | ( \pi329 & w1959 ) | ( \pi457 & w1959 ) ;
  assign w1961 = ( w1946 & w1958 ) | ( w1946 & ~w1960 ) | ( w1958 & ~w1960 ) ;
  assign w1962 = ( ~w1939 & w1941 ) | ( ~w1939 & w1961 ) | ( w1941 & w1961 ) ;
  assign w1963 = ( w1935 & ~w1937 ) | ( w1935 & w1962 ) | ( ~w1937 & w1962 ) ;
  assign w1964 = w1260 | w1431 ;
  assign w1965 = \pi461 | w1964 ;
  assign w1966 = ~w1433 & w1435 ;
  assign w1967 = ( ~\pi333 & w1431 ) | ( ~\pi333 & w1964 ) | ( w1431 & w1964 ) ;
  assign w1968 = ( w1965 & w1966 ) | ( w1965 & ~w1967 ) | ( w1966 & ~w1967 ) ;
  assign w1969 = w1429 & ~w1444 ;
  assign w1970 = w1957 | w1963 ;
  assign w1971 = ( w1439 & ~w1968 ) | ( w1439 & w1970 ) | ( ~w1968 & w1970 ) ;
  assign w1972 = ( w1439 & w1444 ) | ( w1439 & ~w1969 ) | ( w1444 & ~w1969 ) ;
  assign w1973 = ( ~w1969 & w1971 ) | ( ~w1969 & w1972 ) | ( w1971 & w1972 ) ;
  assign w1974 = w1413 | w1418 ;
  assign w1975 = ( w1420 & ~w1422 ) | ( w1420 & w1973 ) | ( ~w1422 & w1973 ) ;
  assign w1976 = ( w1973 & ~w1974 ) | ( w1973 & w1975 ) | ( ~w1974 & w1975 ) ;
  assign w1977 = ~w1974 & w1976 ;
  assign w1978 = ~w1400 & w1402 ;
  assign w1979 = \pi465 ^ w1260 ;
  assign w1980 = ( \pi337 & \pi465 ) | ( \pi337 & w1979 ) | ( \pi465 & w1979 ) ;
  assign w1981 = ( w1415 & w1978 ) | ( w1415 & ~w1980 ) | ( w1978 & ~w1980 ) ;
  assign w1982 = ( ~w1408 & w1410 ) | ( ~w1408 & w1981 ) | ( w1410 & w1981 ) ;
  assign w1983 = ( w1404 & ~w1406 ) | ( w1404 & w1982 ) | ( ~w1406 & w1982 ) ;
  assign w1984 = w1400 & ~w1402 ;
  assign w1985 = w1977 | w1984 ;
  assign w1986 = ( w1983 & ~w1984 ) | ( w1983 & w1985 ) | ( ~w1984 & w1985 ) ;
  assign w1987 = w1260 | w1390 ;
  assign w1988 = \pi469 | w1987 ;
  assign w1989 = ~w1392 & w1394 ;
  assign w1990 = ( ~\pi341 & w1390 ) | ( ~\pi341 & w1987 ) | ( w1390 & w1987 ) ;
  assign w1991 = ( w1988 & w1989 ) | ( w1988 & ~w1990 ) | ( w1989 & ~w1990 ) ;
  assign w1992 = ( w1398 & w1986 ) | ( w1398 & ~w1991 ) | ( w1986 & ~w1991 ) ;
  assign w1993 = ( ~w1384 & w1398 ) | ( ~w1384 & w1992 ) | ( w1398 & w1992 ) ;
  assign w1994 = ( ~w1386 & w1388 ) | ( ~w1386 & w1993 ) | ( w1388 & w1993 ) ;
  assign w1995 = ~w1384 & w1994 ;
  assign w1996 = \pi219 ^ w1256 ;
  assign w1997 = ( \pi091 & \pi219 ) | ( \pi091 & w1996 ) | ( \pi219 & w1996 ) ;
  assign w1998 = \pi475 ^ w1260 ;
  assign w1999 = ( \pi347 & \pi475 ) | ( \pi347 & w1998 ) | ( \pi475 & w1998 ) ;
  assign w2000 = \pi474 ^ w1260 ;
  assign w2001 = ( \pi346 & \pi474 ) | ( \pi346 & w2000 ) | ( \pi474 & w2000 ) ;
  assign w2002 = \pi218 ^ w1256 ;
  assign w2003 = ( \pi090 & \pi218 ) | ( \pi090 & w2002 ) | ( \pi218 & w2002 ) ;
  assign w2004 = \pi217 ^ w1256 ;
  assign w2005 = ( \pi089 & \pi217 ) | ( \pi089 & w2004 ) | ( \pi217 & w2004 ) ;
  assign w2006 = \pi472 ^ w1260 ;
  assign w2007 = ( \pi344 & \pi472 ) | ( \pi344 & w2006 ) | ( \pi472 & w2006 ) ;
  assign w2008 = \pi216 ^ w1256 ;
  assign w2009 = ( \pi088 & \pi216 ) | ( \pi088 & w2008 ) | ( \pi216 & w2008 ) ;
  assign w2010 = w1260 | w2005 ;
  assign w2011 = \pi473 | w2010 ;
  assign w2012 = w2007 & ~w2009 ;
  assign w2013 = ( ~\pi345 & w2005 ) | ( ~\pi345 & w2010 ) | ( w2005 & w2010 ) ;
  assign w2014 = ( w2011 & w2012 ) | ( w2011 & ~w2013 ) | ( w2012 & ~w2013 ) ;
  assign w2015 = w1997 & w1999 ;
  assign w2016 = w2001 & w2003 ;
  assign w2017 = ( w2001 & w2014 ) | ( w2001 & ~w2016 ) | ( w2014 & ~w2016 ) ;
  assign w2018 = ( w1999 & ~w2015 ) | ( w1999 & w2017 ) | ( ~w2015 & w2017 ) ;
  assign w2019 = ~w2007 & w2009 ;
  assign w2020 = \pi473 ^ w1260 ;
  assign w2021 = ( \pi345 & \pi473 ) | ( \pi345 & w2020 ) | ( \pi473 & w2020 ) ;
  assign w2022 = ( w2005 & w2019 ) | ( w2005 & ~w2021 ) | ( w2019 & ~w2021 ) ;
  assign w2023 = ( ~w2001 & w2003 ) | ( ~w2001 & w2022 ) | ( w2003 & w2022 ) ;
  assign w2024 = ( w1997 & ~w1999 ) | ( w1997 & w2023 ) | ( ~w1999 & w2023 ) ;
  assign w2025 = w1368 & w1370 ;
  assign w2026 = w1372 | w1374 ;
  assign w2027 = ( w1366 & ~w1372 ) | ( w1366 & w2026 ) | ( ~w1372 & w2026 ) ;
  assign w2028 = ( w1370 & ~w2025 ) | ( w1370 & w2027 ) | ( ~w2025 & w2027 ) ;
  assign w2029 = w2024 & ~w2028 ;
  assign w2030 = ( w2018 & w2028 ) | ( w2018 & ~w2029 ) | ( w2028 & ~w2029 ) ;
  assign w2031 = w1381 | w1995 ;
  assign w2032 = ( w2029 & ~w2030 ) | ( w2029 & w2031 ) | ( ~w2030 & w2031 ) ;
  assign w2033 = ( ~w1357 & w1359 ) | ( ~w1357 & w2032 ) | ( w1359 & w2032 ) ;
  assign w2034 = ~w2032 & w2033 ;
  assign w2035 = ( ~w1361 & w1363 ) | ( ~w1361 & w1376 ) | ( w1363 & w1376 ) ;
  assign w2036 = ( w2032 & ~w2034 ) | ( w2032 & w2035 ) | ( ~w2034 & w2035 ) ;
  assign w2037 = w1357 & ~w1359 ;
  assign w2038 = w2036 & ~w2037 ;
  assign w2039 = ( ~w1355 & w2037 ) | ( ~w1355 & w2038 ) | ( w2037 & w2038 ) ;
  assign w2040 = ~w1337 & w1339 ;
  assign w2041 = \pi481 ^ w1260 ;
  assign w2042 = ( \pi353 & \pi481 ) | ( \pi353 & w2041 ) | ( \pi481 & w2041 ) ;
  assign w2043 = ( w1352 & w2040 ) | ( w1352 & ~w2042 ) | ( w2040 & ~w2042 ) ;
  assign w2044 = ( ~w1345 & w1347 ) | ( ~w1345 & w2043 ) | ( w1347 & w2043 ) ;
  assign w2045 = ( w1341 & ~w1343 ) | ( w1341 & w2044 ) | ( ~w1343 & w2044 ) ;
  assign w2046 = w1260 | w1327 ;
  assign w2047 = \pi485 | w2046 ;
  assign w2048 = ~w1329 & w1331 ;
  assign w2049 = ( ~\pi357 & w1327 ) | ( ~\pi357 & w2046 ) | ( w1327 & w2046 ) ;
  assign w2050 = ( w2047 & w2048 ) | ( w2047 & ~w2049 ) | ( w2048 & ~w2049 ) ;
  assign w2051 = w1319 & w1321 ;
  assign w2052 = w1323 & w1325 ;
  assign w2053 = ( w1323 & w2050 ) | ( w1323 & ~w2052 ) | ( w2050 & ~w2052 ) ;
  assign w2054 = ( w1321 & ~w2051 ) | ( w1321 & w2053 ) | ( ~w2051 & w2053 ) ;
  assign w2055 = w2045 & ~w2054 ;
  assign w2056 = ( w1337 & w1339 ) | ( w1337 & ~w2055 ) | ( w1339 & ~w2055 ) ;
  assign w2057 = ( w1339 & w2039 ) | ( w1339 & ~w2056 ) | ( w2039 & ~w2056 ) ;
  assign w2058 = ( w1350 & w2054 ) | ( w1350 & ~w2055 ) | ( w2054 & ~w2055 ) ;
  assign w2059 = ( w2055 & w2057 ) | ( w2055 & ~w2058 ) | ( w2057 & ~w2058 ) ;
  assign w2060 = w1319 | w2059 ;
  assign w2061 = ( ~w1323 & w1325 ) | ( ~w1323 & w1335 ) | ( w1325 & w1335 ) ;
  assign w2062 = w1321 & ~w2059 ;
  assign w2063 = ( w2060 & w2061 ) | ( w2060 & ~w2062 ) | ( w2061 & ~w2062 ) ;
  assign w2064 = \pi235 ^ w1256 ;
  assign w2065 = ( \pi107 & \pi235 ) | ( \pi107 & w2064 ) | ( \pi235 & w2064 ) ;
  assign w2066 = \pi491 ^ w1260 ;
  assign w2067 = ( \pi363 & \pi491 ) | ( \pi363 & w2066 ) | ( \pi491 & w2066 ) ;
  assign w2068 = \pi490 ^ w1260 ;
  assign w2069 = ( \pi362 & \pi490 ) | ( \pi362 & w2068 ) | ( \pi490 & w2068 ) ;
  assign w2070 = \pi234 ^ w1256 ;
  assign w2071 = ( \pi106 & \pi234 ) | ( \pi106 & w2070 ) | ( \pi234 & w2070 ) ;
  assign w2072 = \pi233 ^ w1256 ;
  assign w2073 = ( \pi105 & \pi233 ) | ( \pi105 & w2072 ) | ( \pi233 & w2072 ) ;
  assign w2074 = \pi488 ^ w1260 ;
  assign w2075 = ( \pi360 & \pi488 ) | ( \pi360 & w2074 ) | ( \pi488 & w2074 ) ;
  assign w2076 = \pi232 ^ w1256 ;
  assign w2077 = ( \pi104 & \pi232 ) | ( \pi104 & w2076 ) | ( \pi232 & w2076 ) ;
  assign w2078 = w1260 | w2073 ;
  assign w2079 = \pi489 | w2078 ;
  assign w2080 = w2075 & ~w2077 ;
  assign w2081 = ( ~\pi361 & w2073 ) | ( ~\pi361 & w2078 ) | ( w2073 & w2078 ) ;
  assign w2082 = ( w2079 & w2080 ) | ( w2079 & ~w2081 ) | ( w2080 & ~w2081 ) ;
  assign w2083 = w2065 | w2067 ;
  assign w2084 = ( w2063 & w2069 ) | ( w2063 & w2071 ) | ( w2069 & w2071 ) ;
  assign w2085 = ( ~w2071 & w2082 ) | ( ~w2071 & w2084 ) | ( w2082 & w2084 ) ;
  assign w2086 = w2063 & ~w2085 ;
  assign w2087 = ( w2065 & ~w2083 ) | ( w2065 & w2086 ) | ( ~w2083 & w2086 ) ;
  assign w2088 = ~w2075 & w2077 ;
  assign w2089 = \pi489 ^ w1260 ;
  assign w2090 = ( \pi361 & \pi489 ) | ( \pi361 & w2089 ) | ( \pi489 & w2089 ) ;
  assign w2091 = ( w2073 & w2088 ) | ( w2073 & ~w2090 ) | ( w2088 & ~w2090 ) ;
  assign w2092 = ( ~w2069 & w2071 ) | ( ~w2069 & w2091 ) | ( w2071 & w2091 ) ;
  assign w2093 = ( w2065 & ~w2067 ) | ( w2065 & w2092 ) | ( ~w2067 & w2092 ) ;
  assign w2094 = w1309 & w1311 ;
  assign w2095 = w1313 | w1315 ;
  assign w2096 = ( w1307 & ~w1313 ) | ( w1307 & w2095 ) | ( ~w1313 & w2095 ) ;
  assign w2097 = ( w1311 & ~w2094 ) | ( w1311 & w2096 ) | ( ~w2094 & w2096 ) ;
  assign w2098 = ( w2087 & w2093 ) | ( w2087 & ~w2097 ) | ( w2093 & ~w2097 ) ;
  assign w2099 = ~w2097 & w2098 ;
  assign w2100 = ( ~w1298 & w1300 ) | ( ~w1298 & w2099 ) | ( w1300 & w2099 ) ;
  assign w2101 = ~w2099 & w2100 ;
  assign w2102 = ( ~w1302 & w1304 ) | ( ~w1302 & w1317 ) | ( w1304 & w1317 ) ;
  assign w2103 = ( w2099 & ~w2101 ) | ( w2099 & w2102 ) | ( ~w2101 & w2102 ) ;
  assign w2104 = w1298 & ~w1300 ;
  assign w2105 = w2103 & ~w2104 ;
  assign w2106 = ( ~w1296 & w2104 ) | ( ~w1296 & w2105 ) | ( w2104 & w2105 ) ;
  assign w2107 = ~w1278 & w1280 ;
  assign w2108 = \pi497 ^ w1260 ;
  assign w2109 = ( \pi369 & \pi497 ) | ( \pi369 & w2108 ) | ( \pi497 & w2108 ) ;
  assign w2110 = ( w1293 & w2107 ) | ( w1293 & ~w2109 ) | ( w2107 & ~w2109 ) ;
  assign w2111 = ( ~w1286 & w1288 ) | ( ~w1286 & w2110 ) | ( w1288 & w2110 ) ;
  assign w2112 = ( w1282 & ~w1284 ) | ( w1282 & w2111 ) | ( ~w1284 & w2111 ) ;
  assign w2113 = w1260 | w1270 ;
  assign w2114 = \pi501 | w2113 ;
  assign w2115 = ~w1268 & w1272 ;
  assign w2116 = ( ~\pi373 & w1270 ) | ( ~\pi373 & w2113 ) | ( w1270 & w2113 ) ;
  assign w2117 = ( w2114 & w2115 ) | ( w2114 & ~w2116 ) | ( w2115 & ~w2116 ) ;
  assign w2118 = w1258 & w1262 ;
  assign w2119 = w1264 & w1266 ;
  assign w2120 = ( w1264 & w2117 ) | ( w1264 & ~w2119 ) | ( w2117 & ~w2119 ) ;
  assign w2121 = ( w1262 & ~w2118 ) | ( w1262 & w2120 ) | ( ~w2118 & w2120 ) ;
  assign w2122 = w2112 & ~w2121 ;
  assign w2123 = ( w1278 & w1280 ) | ( w1278 & ~w2122 ) | ( w1280 & ~w2122 ) ;
  assign w2124 = ( w1280 & w2106 ) | ( w1280 & ~w2123 ) | ( w2106 & ~w2123 ) ;
  assign w2125 = ( w1291 & w2121 ) | ( w1291 & ~w2122 ) | ( w2121 & ~w2122 ) ;
  assign w2126 = ( w2122 & w2124 ) | ( w2122 & ~w2125 ) | ( w2124 & ~w2125 ) ;
  assign w2127 = w1258 | w2126 ;
  assign w2128 = ( ~w1264 & w1266 ) | ( ~w1264 & w1276 ) | ( w1266 & w1276 ) ;
  assign w2129 = w1262 & ~w2126 ;
  assign w2130 = ( w2127 & w2128 ) | ( w2127 & ~w2129 ) | ( w2128 & ~w2129 ) ;
  assign w2131 = \pi251 ^ w1256 ;
  assign w2132 = ( \pi123 & \pi251 ) | ( \pi123 & w2131 ) | ( \pi251 & w2131 ) ;
  assign w2133 = \pi507 ^ w1260 ;
  assign w2134 = ( \pi379 & \pi507 ) | ( \pi379 & w2133 ) | ( \pi507 & w2133 ) ;
  assign w2135 = \pi506 ^ w1260 ;
  assign w2136 = ( \pi378 & \pi506 ) | ( \pi378 & w2135 ) | ( \pi506 & w2135 ) ;
  assign w2137 = \pi250 ^ w1256 ;
  assign w2138 = ( \pi122 & \pi250 ) | ( \pi122 & w2137 ) | ( \pi250 & w2137 ) ;
  assign w2139 = \pi249 ^ w1256 ;
  assign w2140 = ( \pi121 & \pi249 ) | ( \pi121 & w2139 ) | ( \pi249 & w2139 ) ;
  assign w2141 = \pi504 ^ w1260 ;
  assign w2142 = ( \pi376 & \pi504 ) | ( \pi376 & w2141 ) | ( \pi504 & w2141 ) ;
  assign w2143 = \pi248 ^ w1256 ;
  assign w2144 = ( \pi120 & \pi248 ) | ( \pi120 & w2143 ) | ( \pi248 & w2143 ) ;
  assign w2145 = w1260 | w2140 ;
  assign w2146 = \pi505 | w2145 ;
  assign w2147 = w2142 & ~w2144 ;
  assign w2148 = ( ~\pi377 & w2140 ) | ( ~\pi377 & w2145 ) | ( w2140 & w2145 ) ;
  assign w2149 = ( w2146 & w2147 ) | ( w2146 & ~w2148 ) | ( w2147 & ~w2148 ) ;
  assign w2150 = w2132 | w2134 ;
  assign w2151 = ( w2130 & w2136 ) | ( w2130 & w2138 ) | ( w2136 & w2138 ) ;
  assign w2152 = ( ~w2138 & w2149 ) | ( ~w2138 & w2151 ) | ( w2149 & w2151 ) ;
  assign w2153 = w2130 & ~w2152 ;
  assign w2154 = ( w2132 & ~w2150 ) | ( w2132 & w2153 ) | ( ~w2150 & w2153 ) ;
  assign w2155 = ~w2142 & w2144 ;
  assign w2156 = \pi505 ^ w1260 ;
  assign w2157 = ( \pi377 & \pi505 ) | ( \pi377 & w2156 ) | ( \pi505 & w2156 ) ;
  assign w2158 = ( w2140 & w2155 ) | ( w2140 & ~w2157 ) | ( w2155 & ~w2157 ) ;
  assign w2159 = w2132 | w2154 ;
  assign w2160 = ( ~w2136 & w2138 ) | ( ~w2136 & w2158 ) | ( w2138 & w2158 ) ;
  assign w2161 = w2134 & ~w2154 ;
  assign w2162 = ( w2159 & w2160 ) | ( w2159 & ~w2161 ) | ( w2160 & ~w2161 ) ;
  assign w2163 = \pi252 ^ w1256 ;
  assign w2164 = ( \pi124 & \pi252 ) | ( \pi124 & w2163 ) | ( \pi252 & w2163 ) ;
  assign w2165 = \pi508 ^ w1260 ;
  assign w2166 = ( \pi380 & \pi508 ) | ( \pi380 & w2165 ) | ( \pi508 & w2165 ) ;
  assign w2167 = ~w2164 & w2166 ;
  assign w2168 = \pi254 ^ w1256 ;
  assign w2169 = ( \pi126 & \pi254 ) | ( \pi126 & w2168 ) | ( \pi254 & w2168 ) ;
  assign w2170 = \pi510 ^ w1260 ;
  assign w2171 = ( \pi382 & \pi510 ) | ( \pi382 & w2170 ) | ( \pi510 & w2170 ) ;
  assign w2172 = \pi253 ^ w1256 ;
  assign w2173 = ( \pi125 & \pi253 ) | ( \pi125 & w2172 ) | ( \pi253 & w2172 ) ;
  assign w2174 = \pi509 ^ w1260 ;
  assign w2175 = ( \pi381 & \pi509 ) | ( \pi381 & w2174 ) | ( \pi509 & w2174 ) ;
  assign w2176 = w2173 & w2175 ;
  assign w2177 = ~w2169 & w2171 ;
  assign w2178 = ( w2175 & ~w2176 ) | ( w2175 & w2177 ) | ( ~w2176 & w2177 ) ;
  assign w2179 = w2164 & ~w2166 ;
  assign w2180 = ( w2173 & ~w2175 ) | ( w2173 & w2179 ) | ( ~w2175 & w2179 ) ;
  assign w2181 = ( w2169 & ~w2171 ) | ( w2169 & w2180 ) | ( ~w2171 & w2180 ) ;
  assign w2182 = ~w883 & w1254 ;
  assign w2183 = ( w2162 & w2167 ) | ( w2162 & w2181 ) | ( w2167 & w2181 ) ;
  assign w2184 = ( w2162 & ~w2178 ) | ( w2162 & w2183 ) | ( ~w2178 & w2183 ) ;
  assign w2185 = ~w2183 & w2184 ;
  assign w2186 = ( w2181 & ~w2182 ) | ( w2181 & w2185 ) | ( ~w2182 & w2185 ) ;
  assign w2187 = ( w883 & ~w1254 ) | ( w883 & w2186 ) | ( ~w1254 & w2186 ) ;
  assign w2188 = w2186 | w2187 ;
  assign w2189 = w1647 ^ w2188 ;
  assign w2190 = \pi256 ^ w1260 ;
  assign w2191 = ( \pi256 & \pi384 ) | ( \pi256 & ~w2190 ) | ( \pi384 & ~w2190 ) ;
  assign w2192 = ( w1647 & ~w2189 ) | ( w1647 & w2191 ) | ( ~w2189 & w2191 ) ;
  assign w2193 = w1645 ^ w2188 ;
  assign w2194 = ( w1645 & w1652 ) | ( w1645 & w2193 ) | ( w1652 & w2193 ) ;
  assign w2195 = w1656 ^ w2188 ;
  assign w2196 = ( w1654 & w1656 ) | ( w1654 & w2195 ) | ( w1656 & w2195 ) ;
  assign w2197 = w1643 ^ w2188 ;
  assign w2198 = ( w1643 & w1660 ) | ( w1643 & ~w2197 ) | ( w1660 & ~w2197 ) ;
  assign w2199 = w1641 ^ w2188 ;
  assign w2200 = ( w1641 & w1663 ) | ( w1641 & ~w2199 ) | ( w1663 & ~w2199 ) ;
  assign w2201 = w1639 ^ w2188 ;
  assign w2202 = ( w1639 & w1666 ) | ( w1639 & ~w2201 ) | ( w1666 & ~w2201 ) ;
  assign w2203 = w1637 ^ w2188 ;
  assign w2204 = ( w1637 & w1669 ) | ( w1637 & ~w2203 ) | ( w1669 & ~w2203 ) ;
  assign w2205 = w1635 ^ w2188 ;
  assign w2206 = ( w1635 & w1672 ) | ( w1635 & ~w2205 ) | ( w1672 & ~w2205 ) ;
  assign w2207 = w1675 ^ w2188 ;
  assign w2208 = ( w1675 & w1677 ) | ( w1675 & ~w2207 ) | ( w1677 & ~w2207 ) ;
  assign w2209 = w1633 ^ w2188 ;
  assign w2210 = ( w1633 & w1680 ) | ( w1633 & w2209 ) | ( w1680 & w2209 ) ;
  assign w2211 = w1631 ^ w2188 ;
  assign w2212 = ( w1629 & w1631 ) | ( w1629 & w2211 ) | ( w1631 & w2211 ) ;
  assign w2213 = w1627 ^ w2188 ;
  assign w2214 = ( w1627 & w1684 ) | ( w1627 & ~w2213 ) | ( w1684 & ~w2213 ) ;
  assign w2215 = w1625 ^ w2188 ;
  assign w2216 = ( w1625 & w1687 ) | ( w1625 & ~w2215 ) | ( w1687 & ~w2215 ) ;
  assign w2217 = w1623 ^ w2188 ;
  assign w2218 = ( w1623 & w1690 ) | ( w1623 & ~w2217 ) | ( w1690 & ~w2217 ) ;
  assign w2219 = w1621 ^ w2188 ;
  assign w2220 = ( w1621 & w1693 ) | ( w1621 & ~w2219 ) | ( w1693 & ~w2219 ) ;
  assign w2221 = w1619 ^ w2188 ;
  assign w2222 = ( w1619 & w1696 ) | ( w1619 & ~w2221 ) | ( w1696 & ~w2221 ) ;
  assign w2223 = w1699 ^ w2188 ;
  assign w2224 = ( w1699 & w1701 ) | ( w1699 & ~w2223 ) | ( w1701 & ~w2223 ) ;
  assign w2225 = w1617 ^ w2188 ;
  assign w2226 = ( w1617 & w1704 ) | ( w1617 & w2225 ) | ( w1704 & w2225 ) ;
  assign w2227 = w1615 ^ w2188 ;
  assign w2228 = ( w1613 & w1615 ) | ( w1613 & w2227 ) | ( w1615 & w2227 ) ;
  assign w2229 = w1611 ^ w2188 ;
  assign w2230 = ( w1611 & w1708 ) | ( w1611 & ~w2229 ) | ( w1708 & ~w2229 ) ;
  assign w2231 = w1609 ^ w2188 ;
  assign w2232 = ( w1609 & w1711 ) | ( w1609 & ~w2231 ) | ( w1711 & ~w2231 ) ;
  assign w2233 = w1607 ^ w2188 ;
  assign w2234 = ( w1607 & w1714 ) | ( w1607 & ~w2233 ) | ( w1714 & ~w2233 ) ;
  assign w2235 = w1605 ^ w2188 ;
  assign w2236 = ( w1605 & w1717 ) | ( w1605 & ~w2235 ) | ( w1717 & ~w2235 ) ;
  assign w2237 = w1603 ^ w2188 ;
  assign w2238 = ( w1603 & w1720 ) | ( w1603 & ~w2237 ) | ( w1720 & ~w2237 ) ;
  assign w2239 = w1723 ^ w2188 ;
  assign w2240 = ( w1723 & w1725 ) | ( w1723 & ~w2239 ) | ( w1725 & ~w2239 ) ;
  assign w2241 = w1601 ^ w2188 ;
  assign w2242 = ( w1601 & w1728 ) | ( w1601 & w2241 ) | ( w1728 & w2241 ) ;
  assign w2243 = w1599 ^ w2188 ;
  assign w2244 = ( w1597 & w1599 ) | ( w1597 & w2243 ) | ( w1599 & w2243 ) ;
  assign w2245 = w1595 ^ w2188 ;
  assign w2246 = ( w1595 & w1732 ) | ( w1595 & ~w2245 ) | ( w1732 & ~w2245 ) ;
  assign w2247 = w1593 ^ w2188 ;
  assign w2248 = ( w1593 & w1735 ) | ( w1593 & ~w2247 ) | ( w1735 & ~w2247 ) ;
  assign w2249 = w1591 ^ w2188 ;
  assign w2250 = ( w1591 & w1738 ) | ( w1591 & ~w2249 ) | ( w1738 & ~w2249 ) ;
  assign w2251 = w1589 ^ w2188 ;
  assign w2252 = ( w1589 & w1741 ) | ( w1589 & ~w2251 ) | ( w1741 & ~w2251 ) ;
  assign w2253 = w1587 ^ w2188 ;
  assign w2254 = ( w1587 & w1744 ) | ( w1587 & ~w2253 ) | ( w1744 & ~w2253 ) ;
  assign w2255 = w1582 ^ w2188 ;
  assign w2256 = \pi288 ^ w1260 ;
  assign w2257 = ( \pi288 & \pi416 ) | ( \pi288 & ~w2256 ) | ( \pi416 & ~w2256 ) ;
  assign w2258 = ( w1582 & ~w2255 ) | ( w1582 & w2257 ) | ( ~w2255 & w2257 ) ;
  assign w2259 = w1772 ^ w2188 ;
  assign w2260 = ( w1770 & w1772 ) | ( w1770 & w2259 ) | ( w1772 & w2259 ) ;
  assign w2261 = w1779 ^ w2188 ;
  assign w2262 = ( w1779 & w1781 ) | ( w1779 & w2261 ) | ( w1781 & w2261 ) ;
  assign w2263 = w1774 ^ w2188 ;
  assign w2264 = \pi291 ^ w1260 ;
  assign w2265 = ( \pi291 & \pi419 ) | ( \pi291 & ~w2264 ) | ( \pi419 & ~w2264 ) ;
  assign w2266 = ( w1774 & ~w2263 ) | ( w1774 & w2265 ) | ( ~w2263 & w2265 ) ;
  assign w2267 = w1757 ^ w2188 ;
  assign w2268 = ( w1755 & w1757 ) | ( w1755 & w2267 ) | ( w1757 & w2267 ) ;
  assign w2269 = w1759 ^ w2188 ;
  assign w2270 = \pi293 ^ w1260 ;
  assign w2271 = ( \pi293 & \pi421 ) | ( \pi293 & ~w2270 ) | ( \pi421 & ~w2270 ) ;
  assign w2272 = ( w1759 & ~w2269 ) | ( w1759 & w2271 ) | ( ~w2269 & w2271 ) ;
  assign w2273 = w1751 ^ w2188 ;
  assign w2274 = ( w1751 & w1753 ) | ( w1751 & w2273 ) | ( w1753 & w2273 ) ;
  assign w2275 = w1749 ^ w2188 ;
  assign w2276 = ( w1747 & w1749 ) | ( w1747 & w2275 ) | ( w1749 & w2275 ) ;
  assign w2277 = w1568 ^ w2188 ;
  assign w2278 = ( w1566 & w1568 ) | ( w1566 & w2277 ) | ( w1568 & w2277 ) ;
  assign w2279 = w1561 ^ w2188 ;
  assign w2280 = \pi297 ^ w1260 ;
  assign w2281 = ( \pi297 & \pi425 ) | ( \pi297 & ~w2280 ) | ( \pi425 & ~w2280 ) ;
  assign w2282 = ( w1561 & ~w2279 ) | ( w1561 & w2281 ) | ( ~w2279 & w2281 ) ;
  assign w2283 = w1556 ^ w2188 ;
  assign w2284 = ( w1554 & w1556 ) | ( w1554 & w2283 ) | ( w1556 & w2283 ) ;
  assign w2285 = w1552 ^ w2188 ;
  assign w2286 = ( w1550 & w1552 ) | ( w1550 & w2285 ) | ( w1552 & w2285 ) ;
  assign w2287 = w1538 ^ w2188 ;
  assign w2288 = ( w1536 & w1538 ) | ( w1536 & w2287 ) | ( w1538 & w2287 ) ;
  assign w2289 = w1540 ^ w2188 ;
  assign w2290 = \pi301 ^ w1260 ;
  assign w2291 = ( \pi301 & \pi429 ) | ( \pi301 & ~w2290 ) | ( \pi429 & ~w2290 ) ;
  assign w2292 = ( w1540 & ~w2289 ) | ( w1540 & w2291 ) | ( ~w2289 & w2291 ) ;
  assign w2293 = w1532 ^ w2188 ;
  assign w2294 = ( w1532 & w1534 ) | ( w1532 & w2293 ) | ( w1534 & w2293 ) ;
  assign w2295 = w1529 ^ w2188 ;
  assign w2296 = ( w1527 & w1529 ) | ( w1527 & w2295 ) | ( w1529 & w2295 ) ;
  assign w2297 = w1822 ^ w2188 ;
  assign w2298 = \pi304 ^ w1260 ;
  assign w2299 = ( \pi304 & \pi432 ) | ( \pi304 & ~w2298 ) | ( \pi432 & ~w2298 ) ;
  assign w2300 = ( w1822 & ~w2297 ) | ( w1822 & w2299 ) | ( ~w2297 & w2299 ) ;
  assign w2301 = w1849 ^ w2188 ;
  assign w2302 = ( w1847 & w1849 ) | ( w1847 & w2301 ) | ( w1849 & w2301 ) ;
  assign w2303 = w1856 ^ w2188 ;
  assign w2304 = ( w1856 & w1858 ) | ( w1856 & w2303 ) | ( w1858 & w2303 ) ;
  assign w2305 = w1851 ^ w2188 ;
  assign w2306 = \pi307 ^ w1260 ;
  assign w2307 = ( \pi307 & \pi435 ) | ( \pi307 & ~w2306 ) | ( \pi435 & ~w2306 ) ;
  assign w2308 = ( w1851 & ~w2305 ) | ( w1851 & w2307 ) | ( ~w2305 & w2307 ) ;
  assign w2309 = w1834 ^ w2188 ;
  assign w2310 = ( w1834 & w1836 ) | ( w1834 & w2309 ) | ( w1836 & w2309 ) ;
  assign w2311 = w1832 ^ w2188 ;
  assign w2312 = \pi309 ^ w1260 ;
  assign w2313 = ( \pi309 & \pi437 ) | ( \pi309 & ~w2312 ) | ( \pi437 & ~w2312 ) ;
  assign w2314 = ( w1832 & ~w2311 ) | ( w1832 & w2313 ) | ( ~w2311 & w2313 ) ;
  assign w2315 = w1828 ^ w2188 ;
  assign w2316 = ( w1828 & w1830 ) | ( w1828 & w2315 ) | ( w1830 & w2315 ) ;
  assign w2317 = w1826 ^ w2188 ;
  assign w2318 = ( w1824 & w1826 ) | ( w1824 & w2317 ) | ( w1826 & w2317 ) ;
  assign w2319 = w1515 ^ w2188 ;
  assign w2320 = ( w1513 & w1515 ) | ( w1513 & w2319 ) | ( w1515 & w2319 ) ;
  assign w2321 = w1511 ^ w2188 ;
  assign w2322 = ( w1509 & w1511 ) | ( w1509 & w2321 ) | ( w1511 & w2321 ) ;
  assign w2323 = w1507 ^ w2188 ;
  assign w2324 = ( w1505 & w1507 ) | ( w1505 & w2323 ) | ( w1507 & w2323 ) ;
  assign w2325 = w1503 ^ w2188 ;
  assign w2326 = ( w1501 & w1503 ) | ( w1501 & w2325 ) | ( w1503 & w2325 ) ;
  assign w2327 = w1489 ^ w2188 ;
  assign w2328 = ( w1487 & w1489 ) | ( w1487 & w2327 ) | ( w1489 & w2327 ) ;
  assign w2329 = w1491 ^ w2188 ;
  assign w2330 = \pi317 ^ w1260 ;
  assign w2331 = ( \pi317 & \pi445 ) | ( \pi317 & ~w2330 ) | ( \pi445 & ~w2330 ) ;
  assign w2332 = ( w1491 & ~w2329 ) | ( w1491 & w2331 ) | ( ~w2329 & w2331 ) ;
  assign w2333 = w1483 ^ w2188 ;
  assign w2334 = ( w1483 & w1485 ) | ( w1483 & w2333 ) | ( w1485 & w2333 ) ;
  assign w2335 = w1478 ^ w2188 ;
  assign w2336 = \pi319 ^ w1260 ;
  assign w2337 = ( \pi319 & \pi447 ) | ( \pi319 & ~w2336 ) | ( \pi447 & ~w2336 ) ;
  assign w2338 = ( w1478 & ~w2335 ) | ( w1478 & w2337 ) | ( ~w2335 & w2337 ) ;
  assign w2339 = w1472 ^ w2188 ;
  assign w2340 = ( w1472 & w1474 ) | ( w1472 & w2339 ) | ( w1474 & w2339 ) ;
  assign w2341 = w1476 ^ w2188 ;
  assign w2342 = \pi321 ^ w1260 ;
  assign w2343 = ( \pi321 & \pi449 ) | ( \pi321 & ~w2342 ) | ( \pi449 & ~w2342 ) ;
  assign w2344 = ( w1476 & ~w2341 ) | ( w1476 & w2343 ) | ( ~w2341 & w2343 ) ;
  assign w2345 = w1468 ^ w2188 ;
  assign w2346 = ( w1468 & w1470 ) | ( w1468 & w2345 ) | ( w1470 & w2345 ) ;
  assign w2347 = w1466 ^ w2188 ;
  assign w2348 = ( w1464 & w1466 ) | ( w1464 & w2347 ) | ( w1466 & w2347 ) ;
  assign w2349 = w1460 ^ w2188 ;
  assign w2350 = ( w1458 & w1460 ) | ( w1458 & w2349 ) | ( w1460 & w2349 ) ;
  assign w2351 = w1456 ^ w2188 ;
  assign w2352 = ( w1454 & w1456 ) | ( w1454 & w2351 ) | ( w1456 & w2351 ) ;
  assign w2353 = w1450 ^ w2188 ;
  assign w2354 = ( w1450 & w1452 ) | ( w1450 & w2353 ) | ( w1452 & w2353 ) ;
  assign w2355 = w1448 ^ w2188 ;
  assign w2356 = ( w1446 & w1448 ) | ( w1446 & w2355 ) | ( w1448 & w2355 ) ;
  assign w2357 = w1951 ^ w2188 ;
  assign w2358 = ( w1951 & w1953 ) | ( w1951 & w2357 ) | ( w1953 & w2357 ) ;
  assign w2359 = w1946 ^ w2188 ;
  assign w2360 = \pi329 ^ w1260 ;
  assign w2361 = ( \pi329 & \pi457 ) | ( \pi329 & ~w2360 ) | ( \pi457 & ~w2360 ) ;
  assign w2362 = ( w1946 & ~w2359 ) | ( w1946 & w2361 ) | ( ~w2359 & w2361 ) ;
  assign w2363 = w1939 ^ w2188 ;
  assign w2364 = ( w1939 & w1941 ) | ( w1939 & w2363 ) | ( w1941 & w2363 ) ;
  assign w2365 = w1937 ^ w2188 ;
  assign w2366 = ( w1935 & w1937 ) | ( w1935 & w2365 ) | ( w1937 & w2365 ) ;
  assign w2367 = w1435 ^ w2188 ;
  assign w2368 = ( w1433 & w1435 ) | ( w1433 & w2367 ) | ( w1435 & w2367 ) ;
  assign w2369 = w1431 ^ w2188 ;
  assign w2370 = \pi333 ^ w1260 ;
  assign w2371 = ( \pi333 & \pi461 ) | ( \pi333 & ~w2370 ) | ( \pi461 & ~w2370 ) ;
  assign w2372 = ( w1431 & ~w2369 ) | ( w1431 & w2371 ) | ( ~w2369 & w2371 ) ;
  assign w2373 = w1424 ^ w2188 ;
  assign w2374 = ( w1424 & w1443 ) | ( w1424 & ~w2373 ) | ( w1443 & ~w2373 ) ;
  assign w2375 = w1422 ^ w2188 ;
  assign w2376 = ( w1420 & w1422 ) | ( w1420 & w2375 ) | ( w1422 & w2375 ) ;
  assign w2377 = w1400 ^ w2188 ;
  assign w2378 = ( w1400 & w1402 ) | ( w1400 & w2377 ) | ( w1402 & w2377 ) ;
  assign w2379 = w1415 ^ w2188 ;
  assign w2380 = \pi337 ^ w1260 ;
  assign w2381 = ( \pi337 & \pi465 ) | ( \pi337 & ~w2380 ) | ( \pi465 & ~w2380 ) ;
  assign w2382 = ( w1415 & ~w2379 ) | ( w1415 & w2381 ) | ( ~w2379 & w2381 ) ;
  assign w2383 = w1408 ^ w2188 ;
  assign w2384 = ( w1408 & w1410 ) | ( w1408 & w2383 ) | ( w1410 & w2383 ) ;
  assign w2385 = w1406 ^ w2188 ;
  assign w2386 = ( w1404 & w1406 ) | ( w1404 & w2385 ) | ( w1406 & w2385 ) ;
  assign w2387 = w1394 ^ w2188 ;
  assign w2388 = ( w1392 & w1394 ) | ( w1392 & w2387 ) | ( w1394 & w2387 ) ;
  assign w2389 = w1390 ^ w2188 ;
  assign w2390 = \pi341 ^ w1260 ;
  assign w2391 = ( \pi341 & \pi469 ) | ( \pi341 & ~w2390 ) | ( \pi469 & ~w2390 ) ;
  assign w2392 = ( w1390 & ~w2389 ) | ( w1390 & w2391 ) | ( ~w2389 & w2391 ) ;
  assign w2393 = w1386 ^ w2188 ;
  assign w2394 = ( w1386 & w1388 ) | ( w1386 & w2393 ) | ( w1388 & w2393 ) ;
  assign w2395 = w1378 ^ w2188 ;
  assign w2396 = \pi343 ^ w1260 ;
  assign w2397 = ( \pi343 & \pi471 ) | ( \pi343 & ~w2396 ) | ( \pi471 & ~w2396 ) ;
  assign w2398 = ( w1378 & ~w2395 ) | ( w1378 & w2397 ) | ( ~w2395 & w2397 ) ;
  assign w2399 = w2007 ^ w2188 ;
  assign w2400 = ( w2007 & w2009 ) | ( w2007 & w2399 ) | ( w2009 & w2399 ) ;
  assign w2401 = w2005 ^ w2188 ;
  assign w2402 = \pi345 ^ w1260 ;
  assign w2403 = ( \pi345 & \pi473 ) | ( \pi345 & ~w2402 ) | ( \pi473 & ~w2402 ) ;
  assign w2404 = ( w2005 & ~w2401 ) | ( w2005 & w2403 ) | ( ~w2401 & w2403 ) ;
  assign w2405 = w2001 ^ w2188 ;
  assign w2406 = ( w2001 & w2003 ) | ( w2001 & w2405 ) | ( w2003 & w2405 ) ;
  assign w2407 = w1999 ^ w2188 ;
  assign w2408 = ( w1997 & w1999 ) | ( w1997 & w2407 ) | ( w1999 & w2407 ) ;
  assign w2409 = w1374 ^ w2188 ;
  assign w2410 = ( w1372 & w1374 ) | ( w1372 & w2409 ) | ( w1374 & w2409 ) ;
  assign w2411 = w1370 ^ w2188 ;
  assign w2412 = ( w1368 & w1370 ) | ( w1368 & w2411 ) | ( w1370 & w2411 ) ;
  assign w2413 = w1361 ^ w2188 ;
  assign w2414 = ( w1361 & w1363 ) | ( w1361 & w2413 ) | ( w1363 & w2413 ) ;
  assign w2415 = w1359 ^ w2188 ;
  assign w2416 = ( w1357 & w1359 ) | ( w1357 & w2415 ) | ( w1359 & w2415 ) ;
  assign w2417 = w1337 ^ w2188 ;
  assign w2418 = ( w1337 & w1339 ) | ( w1337 & w2417 ) | ( w1339 & w2417 ) ;
  assign w2419 = w1352 ^ w2188 ;
  assign w2420 = \pi353 ^ w1260 ;
  assign w2421 = ( \pi353 & \pi481 ) | ( \pi353 & ~w2420 ) | ( \pi481 & ~w2420 ) ;
  assign w2422 = ( w1352 & ~w2419 ) | ( w1352 & w2421 ) | ( ~w2419 & w2421 ) ;
  assign w2423 = w1345 ^ w2188 ;
  assign w2424 = ( w1345 & w1347 ) | ( w1345 & w2423 ) | ( w1347 & w2423 ) ;
  assign w2425 = w1343 ^ w2188 ;
  assign w2426 = ( w1341 & w1343 ) | ( w1341 & w2425 ) | ( w1343 & w2425 ) ;
  assign w2427 = w1331 ^ w2188 ;
  assign w2428 = ( w1329 & w1331 ) | ( w1329 & w2427 ) | ( w1331 & w2427 ) ;
  assign w2429 = w1327 ^ w2188 ;
  assign w2430 = \pi357 ^ w1260 ;
  assign w2431 = ( \pi357 & \pi485 ) | ( \pi357 & ~w2430 ) | ( \pi485 & ~w2430 ) ;
  assign w2432 = ( w1327 & ~w2429 ) | ( w1327 & w2431 ) | ( ~w2429 & w2431 ) ;
  assign w2433 = w1323 ^ w2188 ;
  assign w2434 = ( w1323 & w1325 ) | ( w1323 & w2433 ) | ( w1325 & w2433 ) ;
  assign w2435 = w1321 ^ w2188 ;
  assign w2436 = ( w1319 & w1321 ) | ( w1319 & w2435 ) | ( w1321 & w2435 ) ;
  assign w2437 = w2075 ^ w2188 ;
  assign w2438 = ( w2075 & w2077 ) | ( w2075 & w2437 ) | ( w2077 & w2437 ) ;
  assign w2439 = w2073 ^ w2188 ;
  assign w2440 = \pi361 ^ w1260 ;
  assign w2441 = ( \pi361 & \pi489 ) | ( \pi361 & ~w2440 ) | ( \pi489 & ~w2440 ) ;
  assign w2442 = ( w2073 & ~w2439 ) | ( w2073 & w2441 ) | ( ~w2439 & w2441 ) ;
  assign w2443 = w2069 ^ w2188 ;
  assign w2444 = ( w2069 & w2071 ) | ( w2069 & w2443 ) | ( w2071 & w2443 ) ;
  assign w2445 = w2067 ^ w2188 ;
  assign w2446 = ( w2065 & w2067 ) | ( w2065 & w2445 ) | ( w2067 & w2445 ) ;
  assign w2447 = w1315 ^ w2188 ;
  assign w2448 = ( w1313 & w1315 ) | ( w1313 & w2447 ) | ( w1315 & w2447 ) ;
  assign w2449 = w1311 ^ w2188 ;
  assign w2450 = ( w1309 & w1311 ) | ( w1309 & w2449 ) | ( w1311 & w2449 ) ;
  assign w2451 = w1302 ^ w2188 ;
  assign w2452 = ( w1302 & w1304 ) | ( w1302 & w2451 ) | ( w1304 & w2451 ) ;
  assign w2453 = w1300 ^ w2188 ;
  assign w2454 = ( w1298 & w1300 ) | ( w1298 & w2453 ) | ( w1300 & w2453 ) ;
  assign w2455 = w1278 ^ w2188 ;
  assign w2456 = ( w1278 & w1280 ) | ( w1278 & w2455 ) | ( w1280 & w2455 ) ;
  assign w2457 = w1293 ^ w2188 ;
  assign w2458 = \pi369 ^ w1260 ;
  assign w2459 = ( \pi369 & \pi497 ) | ( \pi369 & ~w2458 ) | ( \pi497 & ~w2458 ) ;
  assign w2460 = ( w1293 & ~w2457 ) | ( w1293 & w2459 ) | ( ~w2457 & w2459 ) ;
  assign w2461 = w1286 ^ w2188 ;
  assign w2462 = ( w1286 & w1288 ) | ( w1286 & w2461 ) | ( w1288 & w2461 ) ;
  assign w2463 = w1284 ^ w2188 ;
  assign w2464 = ( w1282 & w1284 ) | ( w1282 & w2463 ) | ( w1284 & w2463 ) ;
  assign w2465 = w1272 ^ w2188 ;
  assign w2466 = ( w1268 & w1272 ) | ( w1268 & w2465 ) | ( w1272 & w2465 ) ;
  assign w2467 = w1270 ^ w2188 ;
  assign w2468 = \pi373 ^ w1260 ;
  assign w2469 = ( \pi373 & \pi501 ) | ( \pi373 & ~w2468 ) | ( \pi501 & ~w2468 ) ;
  assign w2470 = ( w1270 & ~w2467 ) | ( w1270 & w2469 ) | ( ~w2467 & w2469 ) ;
  assign w2471 = w1264 ^ w2188 ;
  assign w2472 = ( w1264 & w1266 ) | ( w1264 & w2471 ) | ( w1266 & w2471 ) ;
  assign w2473 = w1262 ^ w2188 ;
  assign w2474 = ( w1258 & w1262 ) | ( w1258 & w2473 ) | ( w1262 & w2473 ) ;
  assign w2475 = w2142 ^ w2188 ;
  assign w2476 = ( w2142 & w2144 ) | ( w2142 & w2475 ) | ( w2144 & w2475 ) ;
  assign w2477 = w2140 ^ w2188 ;
  assign w2478 = \pi377 ^ w1260 ;
  assign w2479 = ( \pi377 & \pi505 ) | ( \pi377 & ~w2478 ) | ( \pi505 & ~w2478 ) ;
  assign w2480 = ( w2140 & ~w2477 ) | ( w2140 & w2479 ) | ( ~w2477 & w2479 ) ;
  assign w2481 = w2136 ^ w2188 ;
  assign w2482 = ( w2136 & w2138 ) | ( w2136 & w2481 ) | ( w2138 & w2481 ) ;
  assign w2483 = w2134 ^ w2188 ;
  assign w2484 = ( w2132 & w2134 ) | ( w2132 & w2483 ) | ( w2134 & w2483 ) ;
  assign w2485 = w2166 ^ w2188 ;
  assign w2486 = ( w2164 & w2166 ) | ( w2164 & w2485 ) | ( w2166 & w2485 ) ;
  assign w2487 = w2175 ^ w2188 ;
  assign w2488 = ( w2173 & w2175 ) | ( w2173 & w2487 ) | ( w2175 & w2487 ) ;
  assign w2489 = w2171 ^ w2188 ;
  assign w2490 = ( w2169 & w2171 ) | ( w2169 & w2489 ) | ( w2171 & w2489 ) ;
  assign w2491 = ( w883 & w1254 ) | ( w883 & w2186 ) | ( w1254 & w2186 ) ;
  assign w2492 = w1254 & w2491 ;
  assign w2493 = w1260 ^ w2188 ;
  assign w2494 = ( w1256 & w1260 ) | ( w1256 & w2493 ) | ( w1260 & w2493 ) ;
  assign \po000 = w2192 ;
  assign \po001 = w2194 ;
  assign \po002 = w2196 ;
  assign \po003 = w2198 ;
  assign \po004 = w2200 ;
  assign \po005 = w2202 ;
  assign \po006 = w2204 ;
  assign \po007 = w2206 ;
  assign \po008 = w2208 ;
  assign \po009 = w2210 ;
  assign \po010 = w2212 ;
  assign \po011 = w2214 ;
  assign \po012 = w2216 ;
  assign \po013 = w2218 ;
  assign \po014 = w2220 ;
  assign \po015 = w2222 ;
  assign \po016 = w2224 ;
  assign \po017 = w2226 ;
  assign \po018 = w2228 ;
  assign \po019 = w2230 ;
  assign \po020 = w2232 ;
  assign \po021 = w2234 ;
  assign \po022 = w2236 ;
  assign \po023 = w2238 ;
  assign \po024 = w2240 ;
  assign \po025 = w2242 ;
  assign \po026 = w2244 ;
  assign \po027 = w2246 ;
  assign \po028 = w2248 ;
  assign \po029 = w2250 ;
  assign \po030 = w2252 ;
  assign \po031 = w2254 ;
  assign \po032 = w2258 ;
  assign \po033 = w2260 ;
  assign \po034 = w2262 ;
  assign \po035 = w2266 ;
  assign \po036 = w2268 ;
  assign \po037 = w2272 ;
  assign \po038 = w2274 ;
  assign \po039 = w2276 ;
  assign \po040 = w2278 ;
  assign \po041 = w2282 ;
  assign \po042 = w2284 ;
  assign \po043 = w2286 ;
  assign \po044 = w2288 ;
  assign \po045 = w2292 ;
  assign \po046 = w2294 ;
  assign \po047 = w2296 ;
  assign \po048 = w2300 ;
  assign \po049 = w2302 ;
  assign \po050 = w2304 ;
  assign \po051 = w2308 ;
  assign \po052 = w2310 ;
  assign \po053 = w2314 ;
  assign \po054 = w2316 ;
  assign \po055 = w2318 ;
  assign \po056 = w2320 ;
  assign \po057 = w2322 ;
  assign \po058 = w2324 ;
  assign \po059 = w2326 ;
  assign \po060 = w2328 ;
  assign \po061 = w2332 ;
  assign \po062 = w2334 ;
  assign \po063 = w2338 ;
  assign \po064 = w2340 ;
  assign \po065 = w2344 ;
  assign \po066 = w2346 ;
  assign \po067 = w2348 ;
  assign \po068 = w2350 ;
  assign \po069 = w2352 ;
  assign \po070 = w2354 ;
  assign \po071 = w2356 ;
  assign \po072 = w2358 ;
  assign \po073 = w2362 ;
  assign \po074 = w2364 ;
  assign \po075 = w2366 ;
  assign \po076 = w2368 ;
  assign \po077 = w2372 ;
  assign \po078 = w2374 ;
  assign \po079 = w2376 ;
  assign \po080 = w2378 ;
  assign \po081 = w2382 ;
  assign \po082 = w2384 ;
  assign \po083 = w2386 ;
  assign \po084 = w2388 ;
  assign \po085 = w2392 ;
  assign \po086 = w2394 ;
  assign \po087 = w2398 ;
  assign \po088 = w2400 ;
  assign \po089 = w2404 ;
  assign \po090 = w2406 ;
  assign \po091 = w2408 ;
  assign \po092 = w2410 ;
  assign \po093 = w2412 ;
  assign \po094 = w2414 ;
  assign \po095 = w2416 ;
  assign \po096 = w2418 ;
  assign \po097 = w2422 ;
  assign \po098 = w2424 ;
  assign \po099 = w2426 ;
  assign \po100 = w2428 ;
  assign \po101 = w2432 ;
  assign \po102 = w2434 ;
  assign \po103 = w2436 ;
  assign \po104 = w2438 ;
  assign \po105 = w2442 ;
  assign \po106 = w2444 ;
  assign \po107 = w2446 ;
  assign \po108 = w2448 ;
  assign \po109 = w2450 ;
  assign \po110 = w2452 ;
  assign \po111 = w2454 ;
  assign \po112 = w2456 ;
  assign \po113 = w2460 ;
  assign \po114 = w2462 ;
  assign \po115 = w2464 ;
  assign \po116 = w2466 ;
  assign \po117 = w2470 ;
  assign \po118 = w2472 ;
  assign \po119 = w2474 ;
  assign \po120 = w2476 ;
  assign \po121 = w2480 ;
  assign \po122 = w2482 ;
  assign \po123 = w2484 ;
  assign \po124 = w2486 ;
  assign \po125 = w2488 ;
  assign \po126 = w2490 ;
  assign \po127 = w2492 ;
  assign \po128 = ~w2494 ;
  assign \po129 = ~w2188 ;
endmodule
