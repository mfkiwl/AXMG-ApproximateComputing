module adder( \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 , \pi135 , \pi136 , \pi137 , \pi138 , \pi139 , \pi140 , \pi141 , \pi142 , \pi143 , \pi144 , \pi145 , \pi146 , \pi147 , \pi148 , \pi149 , \pi150 , \pi151 , \pi152 , \pi153 , \pi154 , \pi155 , \pi156 , \pi157 , \pi158 , \pi159 , \pi160 , \pi161 , \pi162 , \pi163 , \pi164 , \pi165 , \pi166 , \pi167 , \pi168 , \pi169 , \pi170 , \pi171 , \pi172 , \pi173 , \pi174 , \pi175 , \pi176 , \pi177 , \pi178 , \pi179 , \pi180 , \pi181 , \pi182 , \pi183 , \pi184 , \pi185 , \pi186 , \pi187 , \pi188 , \pi189 , \pi190 , \pi191 , \pi192 , \pi193 , \pi194 , \pi195 , \pi196 , \pi197 , \pi198 , \pi199 , \pi200 , \pi201 , \pi202 , \pi203 , \pi204 , \pi205 , \pi206 , \pi207 , \pi208 , \pi209 , \pi210 , \pi211 , \pi212 , \pi213 , \pi214 , \pi215 , \pi216 , \pi217 , \pi218 , \pi219 , \pi220 , \pi221 , \pi222 , \pi223 , \pi224 , \pi225 , \pi226 , \pi227 , \pi228 , \pi229 , \pi230 , \pi231 , \pi232 , \pi233 , \pi234 , \pi235 , \pi236 , \pi237 , \pi238 , \pi239 , \pi240 , \pi241 , \pi242 , \pi243 , \pi244 , \pi245 , \pi246 , \pi247 , \pi248 , \pi249 , \pi250 , \pi251 , \pi252 , \pi253 , \pi254 , \pi255 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 , \po128 );
  input \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \pi128 , \pi129 , \pi130 , \pi131 , \pi132 , \pi133 , \pi134 , \pi135 , \pi136 , \pi137 , \pi138 , \pi139 , \pi140 , \pi141 , \pi142 , \pi143 , \pi144 , \pi145 , \pi146 , \pi147 , \pi148 , \pi149 , \pi150 , \pi151 , \pi152 , \pi153 , \pi154 , \pi155 , \pi156 , \pi157 , \pi158 , \pi159 , \pi160 , \pi161 , \pi162 , \pi163 , \pi164 , \pi165 , \pi166 , \pi167 , \pi168 , \pi169 , \pi170 , \pi171 , \pi172 , \pi173 , \pi174 , \pi175 , \pi176 , \pi177 , \pi178 , \pi179 , \pi180 , \pi181 , \pi182 , \pi183 , \pi184 , \pi185 , \pi186 , \pi187 , \pi188 , \pi189 , \pi190 , \pi191 , \pi192 , \pi193 , \pi194 , \pi195 , \pi196 , \pi197 , \pi198 , \pi199 , \pi200 , \pi201 , \pi202 , \pi203 , \pi204 , \pi205 , \pi206 , \pi207 , \pi208 , \pi209 , \pi210 , \pi211 , \pi212 , \pi213 , \pi214 , \pi215 , \pi216 , \pi217 , \pi218 , \pi219 , \pi220 , \pi221 , \pi222 , \pi223 , \pi224 , \pi225 , \pi226 , \pi227 , \pi228 , \pi229 , \pi230 , \pi231 , \pi232 , \pi233 , \pi234 , \pi235 , \pi236 , \pi237 , \pi238 , \pi239 , \pi240 , \pi241 , \pi242 , \pi243 , \pi244 , \pi245 , \pi246 , \pi247 , \pi248 , \pi249 , \pi250 , \pi251 , \pi252 , \pi253 , \pi254 , \pi255 ;
  output \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 , \po128 ;
  wire zero , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 ;
  assign zero = 0;
  assign w257 = \pi000 ^ \pi128 ;
  assign w258 = \pi000 & \pi128 ;
  assign w259 = \pi129 ^ w258 ;
  assign w260 = \pi001 ^ w259 ;
  assign w261 = ( \pi001 & \pi129 ) | ( \pi001 & w258 ) | ( \pi129 & w258 ) ;
  assign w262 = \pi002 ^ w261 ;
  assign w263 = \pi130 ^ w262 ;
  assign w264 = ( \pi002 & \pi130 ) | ( \pi002 & w261 ) | ( \pi130 & w261 ) ;
  assign w265 = \pi003 ^ w264 ;
  assign w266 = \pi131 ^ w265 ;
  assign w267 = ( \pi003 & \pi131 ) | ( \pi003 & w264 ) | ( \pi131 & w264 ) ;
  assign w268 = \pi004 ^ \pi132 ;
  assign w269 = w267 ^ w268 ;
  assign w270 = ( \pi004 & \pi132 ) | ( \pi004 & w267 ) | ( \pi132 & w267 ) ;
  assign w271 = \pi005 ^ w270 ;
  assign w272 = \pi133 ^ w271 ;
  assign w273 = ( \pi005 & \pi133 ) | ( \pi005 & w270 ) | ( \pi133 & w270 ) ;
  assign w274 = \pi006 ^ \pi134 ;
  assign w275 = w273 ^ w274 ;
  assign w276 = ( \pi006 & \pi134 ) | ( \pi006 & w273 ) | ( \pi134 & w273 ) ;
  assign w277 = \pi007 ^ w276 ;
  assign w278 = \pi135 ^ w277 ;
  assign w279 = ( \pi007 & \pi135 ) | ( \pi007 & w276 ) | ( \pi135 & w276 ) ;
  assign w280 = \pi008 ^ \pi136 ;
  assign w281 = w279 ^ w280 ;
  assign w282 = ( \pi008 & \pi136 ) | ( \pi008 & w279 ) | ( \pi136 & w279 ) ;
  assign w283 = \pi009 ^ w282 ;
  assign w284 = \pi137 ^ w283 ;
  assign w285 = ( \pi009 & \pi137 ) | ( \pi009 & w282 ) | ( \pi137 & w282 ) ;
  assign w286 = \pi010 ^ \pi138 ;
  assign w287 = w285 ^ w286 ;
  assign w288 = ( \pi010 & \pi138 ) | ( \pi010 & w285 ) | ( \pi138 & w285 ) ;
  assign w289 = \pi011 ^ w288 ;
  assign w290 = \pi139 ^ w289 ;
  assign w291 = ( \pi011 & \pi139 ) | ( \pi011 & w288 ) | ( \pi139 & w288 ) ;
  assign w292 = \pi012 ^ \pi140 ;
  assign w293 = w291 ^ w292 ;
  assign w294 = ( \pi012 & \pi140 ) | ( \pi012 & w291 ) | ( \pi140 & w291 ) ;
  assign w295 = \pi013 ^ w294 ;
  assign w296 = \pi141 ^ w295 ;
  assign w297 = ( \pi013 & \pi141 ) | ( \pi013 & w294 ) | ( \pi141 & w294 ) ;
  assign w298 = \pi014 ^ w297 ;
  assign w299 = \pi142 ^ w298 ;
  assign w300 = ( \pi014 & \pi142 ) | ( \pi014 & w297 ) | ( \pi142 & w297 ) ;
  assign w301 = \pi015 ^ w300 ;
  assign w302 = \pi143 ^ w301 ;
  assign w303 = ( \pi015 & \pi143 ) | ( \pi015 & w300 ) | ( \pi143 & w300 ) ;
  assign w304 = \pi016 ^ w303 ;
  assign w305 = \pi144 ^ w304 ;
  assign w306 = ( \pi016 & \pi144 ) | ( \pi016 & w303 ) | ( \pi144 & w303 ) ;
  assign w307 = \pi017 ^ w306 ;
  assign w308 = \pi145 ^ w307 ;
  assign w309 = ( \pi017 & \pi145 ) | ( \pi017 & w306 ) | ( \pi145 & w306 ) ;
  assign w310 = \pi018 ^ w309 ;
  assign w311 = \pi146 ^ w310 ;
  assign w312 = ( \pi018 & \pi146 ) | ( \pi018 & w309 ) | ( \pi146 & w309 ) ;
  assign w313 = \pi019 ^ w312 ;
  assign w314 = \pi147 ^ w313 ;
  assign w315 = ( \pi019 & \pi147 ) | ( \pi019 & w312 ) | ( \pi147 & w312 ) ;
  assign w316 = \pi020 ^ w315 ;
  assign w317 = \pi148 ^ w316 ;
  assign w318 = ( \pi020 & \pi148 ) | ( \pi020 & w315 ) | ( \pi148 & w315 ) ;
  assign w319 = \pi021 ^ w318 ;
  assign w320 = \pi149 ^ w319 ;
  assign w321 = ( \pi021 & \pi149 ) | ( \pi021 & w318 ) | ( \pi149 & w318 ) ;
  assign w322 = \pi022 ^ w321 ;
  assign w323 = \pi150 ^ w322 ;
  assign w324 = ( \pi022 & \pi150 ) | ( \pi022 & w321 ) | ( \pi150 & w321 ) ;
  assign w325 = \pi023 ^ w324 ;
  assign w326 = \pi151 ^ w325 ;
  assign w327 = ( \pi023 & \pi151 ) | ( \pi023 & w324 ) | ( \pi151 & w324 ) ;
  assign w328 = \pi024 ^ w327 ;
  assign w329 = \pi152 ^ w328 ;
  assign w330 = ( \pi024 & \pi152 ) | ( \pi024 & w327 ) | ( \pi152 & w327 ) ;
  assign w331 = \pi025 ^ w330 ;
  assign w332 = \pi153 ^ w331 ;
  assign w333 = ( \pi025 & \pi153 ) | ( \pi025 & w330 ) | ( \pi153 & w330 ) ;
  assign w334 = \pi026 ^ w333 ;
  assign w335 = \pi154 ^ w334 ;
  assign w336 = ( \pi026 & \pi154 ) | ( \pi026 & w333 ) | ( \pi154 & w333 ) ;
  assign w337 = \pi027 ^ w336 ;
  assign w338 = \pi155 ^ w337 ;
  assign w339 = ( \pi027 & \pi155 ) | ( \pi027 & w336 ) | ( \pi155 & w336 ) ;
  assign w340 = \pi028 ^ w339 ;
  assign w341 = \pi156 ^ w340 ;
  assign w342 = ( \pi028 & \pi156 ) | ( \pi028 & w339 ) | ( \pi156 & w339 ) ;
  assign w343 = \pi029 ^ w342 ;
  assign w344 = \pi157 ^ w343 ;
  assign w345 = ( \pi029 & \pi157 ) | ( \pi029 & w342 ) | ( \pi157 & w342 ) ;
  assign w346 = \pi030 ^ w345 ;
  assign w347 = \pi158 ^ w346 ;
  assign w348 = ( \pi030 & \pi158 ) | ( \pi030 & w345 ) | ( \pi158 & w345 ) ;
  assign w349 = \pi031 ^ w348 ;
  assign w350 = \pi159 ^ w349 ;
  assign w351 = ( \pi031 & \pi159 ) | ( \pi031 & w348 ) | ( \pi159 & w348 ) ;
  assign w352 = \pi032 ^ w351 ;
  assign w353 = \pi160 ^ w352 ;
  assign w354 = ( \pi032 & \pi160 ) | ( \pi032 & w351 ) | ( \pi160 & w351 ) ;
  assign w355 = \pi033 ^ w354 ;
  assign w356 = \pi161 ^ w355 ;
  assign w357 = ( \pi033 & \pi161 ) | ( \pi033 & w354 ) | ( \pi161 & w354 ) ;
  assign w358 = \pi034 ^ w357 ;
  assign w359 = \pi162 ^ w358 ;
  assign w360 = ( \pi034 & \pi162 ) | ( \pi034 & w357 ) | ( \pi162 & w357 ) ;
  assign w361 = \pi035 ^ w360 ;
  assign w362 = \pi163 ^ w361 ;
  assign w363 = ( \pi035 & \pi163 ) | ( \pi035 & w360 ) | ( \pi163 & w360 ) ;
  assign w364 = \pi036 ^ w363 ;
  assign w365 = \pi164 ^ w364 ;
  assign w366 = ( \pi036 & \pi164 ) | ( \pi036 & w363 ) | ( \pi164 & w363 ) ;
  assign w367 = \pi037 ^ w366 ;
  assign w368 = \pi165 ^ w367 ;
  assign w369 = ( \pi037 & \pi165 ) | ( \pi037 & w366 ) | ( \pi165 & w366 ) ;
  assign w370 = \pi038 ^ w369 ;
  assign w371 = \pi166 ^ w370 ;
  assign w372 = ( \pi038 & \pi166 ) | ( \pi038 & w369 ) | ( \pi166 & w369 ) ;
  assign w373 = \pi039 ^ w372 ;
  assign w374 = \pi167 ^ w373 ;
  assign w375 = ( \pi039 & \pi167 ) | ( \pi039 & w372 ) | ( \pi167 & w372 ) ;
  assign w376 = \pi040 ^ w375 ;
  assign w377 = \pi168 ^ w376 ;
  assign w378 = ( \pi040 & \pi168 ) | ( \pi040 & w375 ) | ( \pi168 & w375 ) ;
  assign w379 = \pi041 ^ w378 ;
  assign w380 = \pi169 ^ w379 ;
  assign w381 = ( \pi041 & \pi169 ) | ( \pi041 & w378 ) | ( \pi169 & w378 ) ;
  assign w382 = \pi042 ^ w381 ;
  assign w383 = \pi170 ^ w382 ;
  assign w384 = ( \pi042 & \pi170 ) | ( \pi042 & w381 ) | ( \pi170 & w381 ) ;
  assign w385 = \pi043 ^ w384 ;
  assign w386 = \pi171 ^ w385 ;
  assign w387 = ( \pi043 & \pi171 ) | ( \pi043 & w384 ) | ( \pi171 & w384 ) ;
  assign w388 = \pi044 ^ w387 ;
  assign w389 = \pi172 ^ w388 ;
  assign w390 = ( \pi044 & \pi172 ) | ( \pi044 & w387 ) | ( \pi172 & w387 ) ;
  assign w391 = \pi045 ^ w390 ;
  assign w392 = \pi173 ^ w391 ;
  assign w393 = ( \pi045 & \pi173 ) | ( \pi045 & w390 ) | ( \pi173 & w390 ) ;
  assign w394 = \pi046 ^ w393 ;
  assign w395 = \pi174 ^ w394 ;
  assign w396 = ( \pi046 & \pi174 ) | ( \pi046 & w393 ) | ( \pi174 & w393 ) ;
  assign w397 = \pi047 ^ w396 ;
  assign w398 = \pi175 ^ w397 ;
  assign w399 = ( \pi047 & \pi175 ) | ( \pi047 & w396 ) | ( \pi175 & w396 ) ;
  assign w400 = \pi048 ^ w399 ;
  assign w401 = \pi176 ^ w400 ;
  assign w402 = ( \pi048 & \pi176 ) | ( \pi048 & w399 ) | ( \pi176 & w399 ) ;
  assign w403 = \pi049 ^ w402 ;
  assign w404 = \pi177 ^ w403 ;
  assign w405 = ( \pi049 & \pi177 ) | ( \pi049 & w402 ) | ( \pi177 & w402 ) ;
  assign w406 = \pi050 ^ w405 ;
  assign w407 = \pi178 ^ w406 ;
  assign w408 = ( \pi050 & \pi178 ) | ( \pi050 & w405 ) | ( \pi178 & w405 ) ;
  assign w409 = \pi051 ^ w408 ;
  assign w410 = \pi179 ^ w409 ;
  assign w411 = ( \pi051 & \pi179 ) | ( \pi051 & w408 ) | ( \pi179 & w408 ) ;
  assign w412 = \pi052 ^ w411 ;
  assign w413 = \pi180 ^ w412 ;
  assign w414 = ( \pi052 & \pi180 ) | ( \pi052 & w411 ) | ( \pi180 & w411 ) ;
  assign w415 = \pi053 ^ w414 ;
  assign w416 = \pi181 ^ w415 ;
  assign w417 = ( \pi053 & \pi181 ) | ( \pi053 & w414 ) | ( \pi181 & w414 ) ;
  assign w418 = \pi054 ^ w417 ;
  assign w419 = \pi182 ^ w418 ;
  assign w420 = ( \pi054 & \pi182 ) | ( \pi054 & w417 ) | ( \pi182 & w417 ) ;
  assign w421 = \pi055 ^ w420 ;
  assign w422 = \pi183 ^ w421 ;
  assign w423 = ( \pi055 & \pi183 ) | ( \pi055 & w420 ) | ( \pi183 & w420 ) ;
  assign w424 = \pi056 ^ w423 ;
  assign w425 = \pi184 ^ w424 ;
  assign w426 = ( \pi056 & \pi184 ) | ( \pi056 & w423 ) | ( \pi184 & w423 ) ;
  assign w427 = \pi057 ^ w426 ;
  assign w428 = \pi185 ^ w427 ;
  assign w429 = ( \pi057 & \pi185 ) | ( \pi057 & w426 ) | ( \pi185 & w426 ) ;
  assign w430 = \pi058 ^ w429 ;
  assign w431 = \pi186 ^ w430 ;
  assign w432 = ( \pi058 & \pi186 ) | ( \pi058 & w429 ) | ( \pi186 & w429 ) ;
  assign w433 = \pi059 ^ w432 ;
  assign w434 = \pi187 ^ w433 ;
  assign w435 = ( \pi059 & \pi187 ) | ( \pi059 & w432 ) | ( \pi187 & w432 ) ;
  assign w436 = \pi060 ^ w435 ;
  assign w437 = \pi188 ^ w436 ;
  assign w438 = ( \pi060 & \pi188 ) | ( \pi060 & w435 ) | ( \pi188 & w435 ) ;
  assign w439 = \pi061 ^ w438 ;
  assign w440 = \pi189 ^ w439 ;
  assign w441 = ( \pi061 & \pi189 ) | ( \pi061 & w438 ) | ( \pi189 & w438 ) ;
  assign w442 = \pi062 ^ w441 ;
  assign w443 = \pi190 ^ w442 ;
  assign w444 = ( \pi062 & \pi190 ) | ( \pi062 & w441 ) | ( \pi190 & w441 ) ;
  assign w445 = \pi063 ^ w444 ;
  assign w446 = \pi191 ^ w445 ;
  assign w447 = ( \pi063 & \pi191 ) | ( \pi063 & w444 ) | ( \pi191 & w444 ) ;
  assign w448 = \pi064 ^ w447 ;
  assign w449 = \pi192 ^ w448 ;
  assign w450 = ( \pi064 & \pi192 ) | ( \pi064 & w447 ) | ( \pi192 & w447 ) ;
  assign w451 = \pi065 ^ w450 ;
  assign w452 = \pi193 ^ w451 ;
  assign w453 = ( \pi065 & \pi193 ) | ( \pi065 & w450 ) | ( \pi193 & w450 ) ;
  assign w454 = \pi066 ^ w453 ;
  assign w455 = \pi194 ^ w454 ;
  assign w456 = ( \pi066 & \pi194 ) | ( \pi066 & w453 ) | ( \pi194 & w453 ) ;
  assign w457 = \pi067 ^ w456 ;
  assign w458 = \pi195 ^ w457 ;
  assign w459 = ( \pi067 & \pi195 ) | ( \pi067 & w456 ) | ( \pi195 & w456 ) ;
  assign w460 = \pi068 ^ w459 ;
  assign w461 = \pi196 ^ w460 ;
  assign w462 = ( \pi068 & \pi196 ) | ( \pi068 & w459 ) | ( \pi196 & w459 ) ;
  assign w463 = \pi069 ^ w462 ;
  assign w464 = \pi197 ^ w463 ;
  assign w465 = ( \pi069 & \pi197 ) | ( \pi069 & w462 ) | ( \pi197 & w462 ) ;
  assign w466 = \pi070 ^ w465 ;
  assign w467 = \pi198 ^ w466 ;
  assign w468 = ( \pi070 & \pi198 ) | ( \pi070 & w465 ) | ( \pi198 & w465 ) ;
  assign w469 = \pi071 ^ w468 ;
  assign w470 = \pi199 ^ w469 ;
  assign w471 = ( \pi071 & \pi199 ) | ( \pi071 & w468 ) | ( \pi199 & w468 ) ;
  assign w472 = \pi072 ^ w471 ;
  assign w473 = \pi200 ^ w472 ;
  assign w474 = ( \pi072 & \pi200 ) | ( \pi072 & w471 ) | ( \pi200 & w471 ) ;
  assign w475 = \pi073 ^ w474 ;
  assign w476 = \pi201 ^ w475 ;
  assign w477 = ( \pi073 & \pi201 ) | ( \pi073 & w474 ) | ( \pi201 & w474 ) ;
  assign w478 = \pi074 ^ w477 ;
  assign w479 = \pi202 ^ w478 ;
  assign w480 = ( \pi074 & \pi202 ) | ( \pi074 & w477 ) | ( \pi202 & w477 ) ;
  assign w481 = \pi075 ^ w480 ;
  assign w482 = \pi203 ^ w481 ;
  assign w483 = ( \pi075 & \pi203 ) | ( \pi075 & w480 ) | ( \pi203 & w480 ) ;
  assign w484 = \pi076 ^ w483 ;
  assign w485 = \pi204 ^ w484 ;
  assign w486 = ( \pi076 & \pi204 ) | ( \pi076 & w483 ) | ( \pi204 & w483 ) ;
  assign w487 = \pi077 ^ w486 ;
  assign w488 = \pi205 ^ w487 ;
  assign w489 = ( \pi077 & \pi205 ) | ( \pi077 & w486 ) | ( \pi205 & w486 ) ;
  assign w490 = \pi078 ^ w489 ;
  assign w491 = \pi206 ^ w490 ;
  assign w492 = ( \pi078 & \pi206 ) | ( \pi078 & w489 ) | ( \pi206 & w489 ) ;
  assign w493 = \pi079 ^ w492 ;
  assign w494 = \pi207 ^ w493 ;
  assign w495 = ( \pi079 & \pi207 ) | ( \pi079 & w492 ) | ( \pi207 & w492 ) ;
  assign w496 = \pi080 ^ w495 ;
  assign w497 = \pi208 ^ w496 ;
  assign w498 = ( \pi080 & \pi208 ) | ( \pi080 & w495 ) | ( \pi208 & w495 ) ;
  assign w499 = \pi081 ^ w498 ;
  assign w500 = \pi209 ^ w499 ;
  assign w501 = ( \pi081 & \pi209 ) | ( \pi081 & w498 ) | ( \pi209 & w498 ) ;
  assign w502 = \pi082 ^ w501 ;
  assign w503 = \pi210 ^ w502 ;
  assign w504 = ( \pi082 & \pi210 ) | ( \pi082 & w501 ) | ( \pi210 & w501 ) ;
  assign w505 = \pi083 ^ w504 ;
  assign w506 = \pi211 ^ w505 ;
  assign w507 = ( \pi083 & \pi211 ) | ( \pi083 & w504 ) | ( \pi211 & w504 ) ;
  assign w508 = \pi084 ^ w507 ;
  assign w509 = \pi212 ^ w508 ;
  assign w510 = ( \pi084 & \pi212 ) | ( \pi084 & w507 ) | ( \pi212 & w507 ) ;
  assign w511 = \pi085 ^ w510 ;
  assign w512 = \pi213 ^ w511 ;
  assign w513 = ( \pi085 & \pi213 ) | ( \pi085 & w510 ) | ( \pi213 & w510 ) ;
  assign w514 = \pi086 ^ w513 ;
  assign w515 = \pi214 ^ w514 ;
  assign w516 = ( \pi086 & \pi214 ) | ( \pi086 & w513 ) | ( \pi214 & w513 ) ;
  assign w517 = \pi087 ^ w516 ;
  assign w518 = \pi215 ^ w517 ;
  assign w519 = ( \pi087 & \pi215 ) | ( \pi087 & w516 ) | ( \pi215 & w516 ) ;
  assign w520 = \pi088 ^ w519 ;
  assign w521 = \pi216 ^ w520 ;
  assign w522 = ( \pi088 & \pi216 ) | ( \pi088 & w519 ) | ( \pi216 & w519 ) ;
  assign w523 = \pi089 ^ w522 ;
  assign w524 = \pi217 ^ w523 ;
  assign w525 = ( \pi089 & \pi217 ) | ( \pi089 & w522 ) | ( \pi217 & w522 ) ;
  assign w526 = \pi090 ^ w525 ;
  assign w527 = \pi218 ^ w526 ;
  assign w528 = ( \pi090 & \pi218 ) | ( \pi090 & w525 ) | ( \pi218 & w525 ) ;
  assign w529 = \pi091 ^ w528 ;
  assign w530 = \pi219 ^ w529 ;
  assign w531 = ( \pi091 & \pi219 ) | ( \pi091 & w528 ) | ( \pi219 & w528 ) ;
  assign w532 = \pi092 ^ w531 ;
  assign w533 = \pi220 ^ w532 ;
  assign w534 = ( \pi092 & \pi220 ) | ( \pi092 & w531 ) | ( \pi220 & w531 ) ;
  assign w535 = \pi093 ^ w534 ;
  assign w536 = \pi221 ^ w535 ;
  assign w537 = ( \pi093 & \pi221 ) | ( \pi093 & w534 ) | ( \pi221 & w534 ) ;
  assign w538 = \pi094 ^ w537 ;
  assign w539 = \pi222 ^ w538 ;
  assign w540 = ( \pi094 & \pi222 ) | ( \pi094 & w537 ) | ( \pi222 & w537 ) ;
  assign w541 = \pi095 ^ w540 ;
  assign w542 = \pi223 ^ w541 ;
  assign w543 = ( \pi095 & \pi223 ) | ( \pi095 & w540 ) | ( \pi223 & w540 ) ;
  assign w544 = \pi096 ^ w543 ;
  assign w545 = \pi224 ^ w544 ;
  assign w546 = ( \pi096 & \pi224 ) | ( \pi096 & w543 ) | ( \pi224 & w543 ) ;
  assign w547 = \pi097 ^ w546 ;
  assign w548 = \pi225 ^ w547 ;
  assign w549 = ( \pi097 & \pi225 ) | ( \pi097 & w546 ) | ( \pi225 & w546 ) ;
  assign w550 = \pi098 ^ w549 ;
  assign w551 = \pi226 ^ w550 ;
  assign w552 = ( \pi098 & \pi226 ) | ( \pi098 & w549 ) | ( \pi226 & w549 ) ;
  assign w553 = \pi099 ^ w552 ;
  assign w554 = \pi227 ^ w553 ;
  assign w555 = ( \pi099 & \pi227 ) | ( \pi099 & w552 ) | ( \pi227 & w552 ) ;
  assign w556 = \pi100 ^ w555 ;
  assign w557 = \pi228 ^ w556 ;
  assign w558 = ( \pi100 & \pi228 ) | ( \pi100 & w555 ) | ( \pi228 & w555 ) ;
  assign w559 = \pi101 ^ w558 ;
  assign w560 = \pi229 ^ w559 ;
  assign w561 = ( \pi101 & \pi229 ) | ( \pi101 & w558 ) | ( \pi229 & w558 ) ;
  assign w562 = \pi102 ^ w561 ;
  assign w563 = \pi230 ^ w562 ;
  assign w564 = ( \pi102 & \pi230 ) | ( \pi102 & w561 ) | ( \pi230 & w561 ) ;
  assign w565 = \pi103 ^ w564 ;
  assign w566 = \pi231 ^ w565 ;
  assign w567 = ( \pi103 & \pi231 ) | ( \pi103 & w564 ) | ( \pi231 & w564 ) ;
  assign w568 = \pi104 ^ w567 ;
  assign w569 = \pi232 ^ w568 ;
  assign w570 = ( \pi104 & \pi232 ) | ( \pi104 & w567 ) | ( \pi232 & w567 ) ;
  assign w571 = \pi105 ^ w570 ;
  assign w572 = \pi233 ^ w571 ;
  assign w573 = ( \pi105 & \pi233 ) | ( \pi105 & w570 ) | ( \pi233 & w570 ) ;
  assign w574 = \pi106 ^ w573 ;
  assign w575 = \pi234 ^ w574 ;
  assign w576 = ( \pi106 & \pi234 ) | ( \pi106 & w573 ) | ( \pi234 & w573 ) ;
  assign w577 = \pi107 ^ w576 ;
  assign w578 = \pi235 ^ w577 ;
  assign w579 = ( \pi107 & \pi235 ) | ( \pi107 & w576 ) | ( \pi235 & w576 ) ;
  assign w580 = \pi108 ^ w579 ;
  assign w581 = \pi236 ^ w580 ;
  assign w582 = ( \pi108 & \pi236 ) | ( \pi108 & w579 ) | ( \pi236 & w579 ) ;
  assign w583 = \pi109 ^ w582 ;
  assign w584 = \pi237 ^ w583 ;
  assign w585 = ( \pi109 & \pi237 ) | ( \pi109 & w582 ) | ( \pi237 & w582 ) ;
  assign w586 = \pi110 ^ w585 ;
  assign w587 = \pi238 ^ w586 ;
  assign w588 = ( \pi110 & \pi238 ) | ( \pi110 & w585 ) | ( \pi238 & w585 ) ;
  assign w589 = \pi111 ^ w588 ;
  assign w590 = \pi239 ^ w589 ;
  assign w591 = ( \pi111 & \pi239 ) | ( \pi111 & w588 ) | ( \pi239 & w588 ) ;
  assign w592 = \pi112 ^ w591 ;
  assign w593 = \pi240 ^ w592 ;
  assign w594 = ( \pi112 & \pi240 ) | ( \pi112 & w591 ) | ( \pi240 & w591 ) ;
  assign w595 = \pi113 ^ w594 ;
  assign w596 = \pi241 ^ w595 ;
  assign w597 = ( \pi113 & \pi241 ) | ( \pi113 & w594 ) | ( \pi241 & w594 ) ;
  assign w598 = \pi114 ^ w597 ;
  assign w599 = \pi242 ^ w598 ;
  assign w600 = ( \pi114 & \pi242 ) | ( \pi114 & w597 ) | ( \pi242 & w597 ) ;
  assign w601 = \pi115 ^ w600 ;
  assign w602 = \pi243 ^ w601 ;
  assign w603 = ( \pi115 & \pi243 ) | ( \pi115 & w600 ) | ( \pi243 & w600 ) ;
  assign w604 = \pi116 ^ w603 ;
  assign w605 = \pi244 ^ w604 ;
  assign w606 = ( \pi116 & \pi244 ) | ( \pi116 & w603 ) | ( \pi244 & w603 ) ;
  assign w607 = \pi117 ^ w606 ;
  assign w608 = \pi245 ^ w607 ;
  assign w609 = ( \pi117 & \pi245 ) | ( \pi117 & w606 ) | ( \pi245 & w606 ) ;
  assign w610 = \pi118 ^ w609 ;
  assign w611 = \pi246 ^ w610 ;
  assign w612 = ( \pi118 & \pi246 ) | ( \pi118 & w609 ) | ( \pi246 & w609 ) ;
  assign w613 = \pi119 ^ w612 ;
  assign w614 = \pi247 ^ w613 ;
  assign w615 = ( \pi119 & \pi247 ) | ( \pi119 & w612 ) | ( \pi247 & w612 ) ;
  assign w616 = \pi120 ^ w615 ;
  assign w617 = \pi248 ^ w616 ;
  assign w618 = ( \pi120 & \pi248 ) | ( \pi120 & w615 ) | ( \pi248 & w615 ) ;
  assign w619 = \pi121 ^ w618 ;
  assign w620 = \pi249 ^ w619 ;
  assign w621 = ( \pi121 & \pi249 ) | ( \pi121 & w618 ) | ( \pi249 & w618 ) ;
  assign w622 = \pi122 ^ w621 ;
  assign w623 = \pi250 ^ w622 ;
  assign w624 = ( \pi122 & \pi250 ) | ( \pi122 & w621 ) | ( \pi250 & w621 ) ;
  assign w625 = \pi123 ^ w624 ;
  assign w626 = \pi251 ^ w625 ;
  assign w627 = ( \pi123 & \pi251 ) | ( \pi123 & w624 ) | ( \pi251 & w624 ) ;
  assign w628 = \pi124 ^ w627 ;
  assign w629 = \pi252 ^ w628 ;
  assign w630 = ( \pi124 & \pi252 ) | ( \pi124 & w627 ) | ( \pi252 & w627 ) ;
  assign w631 = \pi125 ^ w630 ;
  assign w632 = \pi253 ^ w631 ;
  assign w633 = ( \pi125 & \pi253 ) | ( \pi125 & w630 ) | ( \pi253 & w630 ) ;
  assign w634 = \pi126 ^ w633 ;
  assign w635 = \pi254 ^ w634 ;
  assign w636 = ( \pi126 & \pi254 ) | ( \pi126 & w633 ) | ( \pi254 & w633 ) ;
  assign w637 = \pi127 ^ w636 ;
  assign w638 = \pi255 ^ w637 ;
  assign w639 = ( \pi127 & \pi255 ) | ( \pi127 & w636 ) | ( \pi255 & w636 ) ;
  assign \po000 = w257 ;
  assign \po001 = w260 ;
  assign \po002 = w263 ;
  assign \po003 = w266 ;
  assign \po004 = w269 ;
  assign \po005 = w272 ;
  assign \po006 = w275 ;
  assign \po007 = w278 ;
  assign \po008 = w281 ;
  assign \po009 = w284 ;
  assign \po010 = w287 ;
  assign \po011 = w290 ;
  assign \po012 = w293 ;
  assign \po013 = w296 ;
  assign \po014 = w299 ;
  assign \po015 = w302 ;
  assign \po016 = w305 ;
  assign \po017 = w308 ;
  assign \po018 = w311 ;
  assign \po019 = w314 ;
  assign \po020 = w317 ;
  assign \po021 = w320 ;
  assign \po022 = w323 ;
  assign \po023 = w326 ;
  assign \po024 = w329 ;
  assign \po025 = w332 ;
  assign \po026 = w335 ;
  assign \po027 = w338 ;
  assign \po028 = w341 ;
  assign \po029 = w344 ;
  assign \po030 = w347 ;
  assign \po031 = w350 ;
  assign \po032 = w353 ;
  assign \po033 = w356 ;
  assign \po034 = w359 ;
  assign \po035 = w362 ;
  assign \po036 = w365 ;
  assign \po037 = w368 ;
  assign \po038 = w371 ;
  assign \po039 = w374 ;
  assign \po040 = w377 ;
  assign \po041 = w380 ;
  assign \po042 = w383 ;
  assign \po043 = w386 ;
  assign \po044 = w389 ;
  assign \po045 = w392 ;
  assign \po046 = w395 ;
  assign \po047 = w398 ;
  assign \po048 = w401 ;
  assign \po049 = w404 ;
  assign \po050 = w407 ;
  assign \po051 = w410 ;
  assign \po052 = w413 ;
  assign \po053 = w416 ;
  assign \po054 = w419 ;
  assign \po055 = w422 ;
  assign \po056 = w425 ;
  assign \po057 = w428 ;
  assign \po058 = w431 ;
  assign \po059 = w434 ;
  assign \po060 = w437 ;
  assign \po061 = w440 ;
  assign \po062 = w443 ;
  assign \po063 = w446 ;
  assign \po064 = w449 ;
  assign \po065 = w452 ;
  assign \po066 = w455 ;
  assign \po067 = w458 ;
  assign \po068 = w461 ;
  assign \po069 = w464 ;
  assign \po070 = w467 ;
  assign \po071 = w470 ;
  assign \po072 = w473 ;
  assign \po073 = w476 ;
  assign \po074 = w479 ;
  assign \po075 = w482 ;
  assign \po076 = w485 ;
  assign \po077 = w488 ;
  assign \po078 = w491 ;
  assign \po079 = w494 ;
  assign \po080 = w497 ;
  assign \po081 = w500 ;
  assign \po082 = w503 ;
  assign \po083 = w506 ;
  assign \po084 = w509 ;
  assign \po085 = w512 ;
  assign \po086 = w515 ;
  assign \po087 = w518 ;
  assign \po088 = w521 ;
  assign \po089 = w524 ;
  assign \po090 = w527 ;
  assign \po091 = w530 ;
  assign \po092 = w533 ;
  assign \po093 = w536 ;
  assign \po094 = w539 ;
  assign \po095 = w542 ;
  assign \po096 = w545 ;
  assign \po097 = w548 ;
  assign \po098 = w551 ;
  assign \po099 = w554 ;
  assign \po100 = w557 ;
  assign \po101 = w560 ;
  assign \po102 = w563 ;
  assign \po103 = w566 ;
  assign \po104 = w569 ;
  assign \po105 = w572 ;
  assign \po106 = w575 ;
  assign \po107 = w578 ;
  assign \po108 = w581 ;
  assign \po109 = w584 ;
  assign \po110 = w587 ;
  assign \po111 = w590 ;
  assign \po112 = w593 ;
  assign \po113 = w596 ;
  assign \po114 = w599 ;
  assign \po115 = w602 ;
  assign \po116 = w605 ;
  assign \po117 = w608 ;
  assign \po118 = w611 ;
  assign \po119 = w614 ;
  assign \po120 = w617 ;
  assign \po121 = w620 ;
  assign \po122 = w623 ;
  assign \po123 = w626 ;
  assign \po124 = w629 ;
  assign \po125 = w632 ;
  assign \po126 = w635 ;
  assign \po127 = w638 ;
  assign \po128 = w639 ;
endmodule
