module sqrt( \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po23 , \po24 , \po25 , \po26 , \po27 , \po28 , \po29 , \po30 , \po31 , \po32 , \po33 , \po34 , \po35 , \po36 , \po37 , \po38 , \po39 , \po40 , \po41 , \po42 , \po43 , \po44 , \po45 , \po46 , \po47 , \po48 , \po49 , \po50 , \po51 , \po52 , \po53 , \po54 , \po55 , \po56 , \po57 , \po58 , \po59 , \po60 , \po61 , \po62 , \po63 );
  input \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 ;
  output \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po23 , \po24 , \po25 , \po26 , \po27 , \po28 , \po29 , \po30 , \po31 , \po32 , \po33 , \po34 , \po35 , \po36 , \po37 , \po38 , \po39 , \po40 , \po41 , \po42 , \po43 , \po44 , \po45 , \po46 , \po47 , \po48 , \po49 , \po50 , \po51 , \po52 , \po53 , \po54 , \po55 , \po56 , \po57 , \po58 , \po59 , \po60 , \po61 , \po62 , \po63 ;
  wire zero , w129 , w130 , w131 , w132 , w133 , w134 , w135 , w136 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w146 , w147 , w148 , w149 , w150 , w151 , w152 , w153 , w154 , w155 , w156 , w157 , w158 , w159 , w160 , w161 , w162 , w163 , w164 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w174 , w175 , w176 , w177 , w178 , w179 , w180 , w181 , w182 , w183 , w184 , w185 , w186 , w187 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w203 , w204 , w205 , w206 , w207 , w208 , w209 , w210 , w211 , w212 , w213 , w214 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w224 , w225 , w226 , w227 , w228 , w229 , w230 , w231 , w232 , w233 , w234 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w250 , w251 , w252 , w253 , w254 , w255 , w256 , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 , w2495 , w2496 , w2497 , w2498 , w2499 , w2500 , w2501 , w2502 , w2503 , w2504 , w2505 , w2506 , w2507 , w2508 , w2509 , w2510 , w2511 , w2512 , w2513 , w2514 , w2515 , w2516 , w2517 , w2518 , w2519 , w2520 , w2521 , w2522 , w2523 , w2524 , w2525 , w2526 , w2527 , w2528 , w2529 , w2530 , w2531 , w2532 , w2533 , w2534 , w2535 , w2536 , w2537 , w2538 , w2539 , w2540 , w2541 , w2542 , w2543 , w2544 , w2545 , w2546 , w2547 , w2548 , w2549 , w2550 , w2551 , w2552 , w2553 , w2554 , w2555 , w2556 , w2557 , w2558 , w2559 , w2560 , w2561 , w2562 , w2563 , w2564 , w2565 , w2566 , w2567 , w2568 , w2569 , w2570 , w2571 , w2572 , w2573 , w2574 , w2575 , w2576 , w2577 , w2578 , w2579 , w2580 , w2581 , w2582 , w2583 , w2584 , w2585 , w2586 , w2587 , w2588 , w2589 , w2590 , w2591 , w2592 , w2593 , w2594 , w2595 , w2596 , w2597 , w2598 , w2599 , w2600 , w2601 , w2602 , w2603 , w2604 , w2605 , w2606 , w2607 , w2608 , w2609 , w2610 , w2611 , w2612 , w2613 , w2614 , w2615 , w2616 , w2617 , w2618 , w2619 , w2620 , w2621 , w2622 , w2623 , w2624 , w2625 , w2626 , w2627 , w2628 , w2629 , w2630 , w2631 , w2632 , w2633 , w2634 , w2635 , w2636 , w2637 , w2638 , w2639 , w2640 , w2641 , w2642 , w2643 , w2644 , w2645 , w2646 , w2647 , w2648 , w2649 , w2650 , w2651 , w2652 , w2653 , w2654 , w2655 , w2656 , w2657 , w2658 , w2659 , w2660 , w2661 , w2662 , w2663 , w2664 , w2665 , w2666 , w2667 , w2668 , w2669 , w2670 , w2671 , w2672 , w2673 , w2674 , w2675 , w2676 , w2677 , w2678 , w2679 , w2680 , w2681 , w2682 , w2683 , w2684 , w2685 , w2686 , w2687 , w2688 , w2689 , w2690 , w2691 , w2692 , w2693 , w2694 , w2695 , w2696 , w2697 , w2698 , w2699 , w2700 , w2701 , w2702 , w2703 , w2704 , w2705 , w2706 , w2707 , w2708 , w2709 , w2710 , w2711 , w2712 , w2713 , w2714 , w2715 , w2716 , w2717 , w2718 , w2719 , w2720 , w2721 , w2722 , w2723 , w2724 , w2725 , w2726 , w2727 , w2728 , w2729 , w2730 , w2731 , w2732 , w2733 , w2734 , w2735 , w2736 , w2737 , w2738 , w2739 , w2740 , w2741 , w2742 , w2743 , w2744 , w2745 , w2746 , w2747 , w2748 , w2749 , w2750 , w2751 , w2752 , w2753 , w2754 , w2755 , w2756 , w2757 , w2758 , w2759 , w2760 , w2761 , w2762 , w2763 , w2764 , w2765 , w2766 , w2767 , w2768 , w2769 , w2770 , w2771 , w2772 , w2773 , w2774 , w2775 , w2776 , w2777 , w2778 , w2779 , w2780 , w2781 , w2782 , w2783 , w2784 , w2785 , w2786 , w2787 , w2788 , w2789 , w2790 , w2791 , w2792 , w2793 , w2794 , w2795 , w2796 , w2797 , w2798 , w2799 , w2800 , w2801 , w2802 , w2803 , w2804 , w2805 , w2806 , w2807 , w2808 , w2809 , w2810 , w2811 , w2812 , w2813 , w2814 , w2815 , w2816 , w2817 , w2818 , w2819 , w2820 , w2821 , w2822 , w2823 , w2824 , w2825 , w2826 , w2827 , w2828 , w2829 , w2830 , w2831 , w2832 , w2833 , w2834 , w2835 , w2836 , w2837 , w2838 , w2839 , w2840 , w2841 , w2842 , w2843 , w2844 , w2845 , w2846 , w2847 , w2848 , w2849 , w2850 , w2851 , w2852 , w2853 , w2854 , w2855 , w2856 , w2857 , w2858 , w2859 , w2860 , w2861 , w2862 , w2863 , w2864 , w2865 , w2866 , w2867 , w2868 , w2869 , w2870 , w2871 , w2872 , w2873 , w2874 , w2875 , w2876 , w2877 , w2878 , w2879 , w2880 , w2881 , w2882 , w2883 , w2884 , w2885 , w2886 , w2887 , w2888 , w2889 , w2890 , w2891 , w2892 , w2893 , w2894 , w2895 , w2896 , w2897 , w2898 , w2899 , w2900 , w2901 , w2902 , w2903 , w2904 , w2905 , w2906 , w2907 , w2908 , w2909 , w2910 , w2911 , w2912 , w2913 , w2914 , w2915 , w2916 , w2917 , w2918 , w2919 , w2920 , w2921 , w2922 , w2923 , w2924 , w2925 , w2926 , w2927 , w2928 , w2929 , w2930 , w2931 , w2932 , w2933 , w2934 , w2935 , w2936 , w2937 , w2938 , w2939 , w2940 , w2941 , w2942 , w2943 , w2944 , w2945 , w2946 , w2947 , w2948 , w2949 , w2950 , w2951 , w2952 , w2953 , w2954 , w2955 , w2956 , w2957 , w2958 , w2959 , w2960 , w2961 , w2962 , w2963 , w2964 , w2965 , w2966 , w2967 , w2968 , w2969 , w2970 , w2971 , w2972 , w2973 , w2974 , w2975 , w2976 , w2977 , w2978 , w2979 , w2980 , w2981 , w2982 , w2983 , w2984 , w2985 , w2986 , w2987 , w2988 , w2989 , w2990 , w2991 , w2992 , w2993 , w2994 , w2995 , w2996 , w2997 , w2998 , w2999 , w3000 , w3001 , w3002 , w3003 , w3004 , w3005 , w3006 , w3007 , w3008 , w3009 , w3010 , w3011 , w3012 , w3013 , w3014 , w3015 , w3016 , w3017 , w3018 , w3019 , w3020 , w3021 , w3022 , w3023 , w3024 , w3025 , w3026 , w3027 , w3028 , w3029 , w3030 , w3031 , w3032 , w3033 , w3034 , w3035 , w3036 , w3037 , w3038 , w3039 , w3040 , w3041 , w3042 , w3043 , w3044 , w3045 , w3046 , w3047 , w3048 , w3049 , w3050 , w3051 , w3052 , w3053 , w3054 , w3055 , w3056 , w3057 , w3058 , w3059 , w3060 , w3061 , w3062 , w3063 , w3064 , w3065 , w3066 , w3067 , w3068 , w3069 , w3070 , w3071 , w3072 , w3073 , w3074 , w3075 , w3076 , w3077 , w3078 , w3079 , w3080 , w3081 , w3082 , w3083 , w3084 , w3085 , w3086 , w3087 , w3088 , w3089 , w3090 , w3091 , w3092 , w3093 , w3094 , w3095 , w3096 , w3097 , w3098 , w3099 , w3100 , w3101 , w3102 , w3103 , w3104 , w3105 , w3106 , w3107 , w3108 , w3109 , w3110 , w3111 , w3112 , w3113 , w3114 , w3115 , w3116 , w3117 , w3118 , w3119 , w3120 , w3121 , w3122 , w3123 , w3124 , w3125 , w3126 , w3127 , w3128 , w3129 , w3130 , w3131 , w3132 , w3133 , w3134 , w3135 , w3136 , w3137 , w3138 , w3139 , w3140 , w3141 , w3142 , w3143 , w3144 , w3145 , w3146 , w3147 , w3148 , w3149 , w3150 , w3151 , w3152 , w3153 , w3154 , w3155 , w3156 , w3157 , w3158 , w3159 , w3160 , w3161 , w3162 , w3163 , w3164 , w3165 , w3166 , w3167 , w3168 , w3169 , w3170 , w3171 , w3172 , w3173 , w3174 , w3175 , w3176 , w3177 , w3178 , w3179 , w3180 , w3181 , w3182 , w3183 , w3184 , w3185 , w3186 , w3187 , w3188 , w3189 , w3190 , w3191 , w3192 , w3193 , w3194 , w3195 , w3196 , w3197 , w3198 , w3199 , w3200 , w3201 , w3202 , w3203 , w3204 , w3205 , w3206 , w3207 , w3208 , w3209 , w3210 , w3211 , w3212 , w3213 , w3214 , w3215 , w3216 , w3217 , w3218 , w3219 , w3220 , w3221 , w3222 , w3223 , w3224 , w3225 , w3226 , w3227 , w3228 , w3229 , w3230 , w3231 , w3232 , w3233 , w3234 , w3235 , w3236 , w3237 , w3238 , w3239 , w3240 , w3241 , w3242 , w3243 , w3244 , w3245 , w3246 , w3247 , w3248 , w3249 , w3250 , w3251 , w3252 , w3253 , w3254 , w3255 , w3256 , w3257 , w3258 , w3259 , w3260 , w3261 , w3262 , w3263 , w3264 , w3265 , w3266 , w3267 , w3268 , w3269 , w3270 , w3271 , w3272 , w3273 , w3274 , w3275 , w3276 , w3277 , w3278 , w3279 , w3280 , w3281 , w3282 , w3283 , w3284 , w3285 , w3286 , w3287 , w3288 , w3289 , w3290 , w3291 , w3292 , w3293 , w3294 , w3295 , w3296 , w3297 , w3298 , w3299 , w3300 , w3301 , w3302 , w3303 , w3304 , w3305 , w3306 , w3307 , w3308 , w3309 , w3310 , w3311 , w3312 , w3313 , w3314 , w3315 , w3316 , w3317 , w3318 , w3319 , w3320 , w3321 , w3322 , w3323 , w3324 , w3325 , w3326 , w3327 , w3328 , w3329 , w3330 , w3331 , w3332 , w3333 , w3334 , w3335 , w3336 , w3337 , w3338 , w3339 , w3340 , w3341 , w3342 , w3343 , w3344 , w3345 , w3346 , w3347 , w3348 , w3349 , w3350 , w3351 , w3352 , w3353 , w3354 , w3355 , w3356 , w3357 , w3358 , w3359 , w3360 , w3361 , w3362 , w3363 , w3364 , w3365 , w3366 , w3367 , w3368 , w3369 , w3370 , w3371 , w3372 , w3373 , w3374 , w3375 , w3376 , w3377 , w3378 , w3379 , w3380 , w3381 , w3382 , w3383 , w3384 , w3385 , w3386 , w3387 , w3388 , w3389 , w3390 , w3391 , w3392 , w3393 , w3394 , w3395 , w3396 , w3397 , w3398 , w3399 , w3400 , w3401 , w3402 , w3403 , w3404 , w3405 , w3406 , w3407 , w3408 , w3409 , w3410 , w3411 , w3412 , w3413 , w3414 , w3415 , w3416 , w3417 , w3418 , w3419 , w3420 , w3421 , w3422 , w3423 , w3424 , w3425 , w3426 , w3427 , w3428 , w3429 , w3430 , w3431 , w3432 , w3433 , w3434 , w3435 , w3436 , w3437 , w3438 , w3439 , w3440 , w3441 , w3442 , w3443 , w3444 , w3445 , w3446 , w3447 , w3448 , w3449 , w3450 , w3451 , w3452 , w3453 , w3454 , w3455 , w3456 , w3457 , w3458 , w3459 , w3460 , w3461 , w3462 , w3463 , w3464 , w3465 , w3466 , w3467 , w3468 , w3469 , w3470 , w3471 , w3472 , w3473 , w3474 , w3475 , w3476 , w3477 , w3478 , w3479 , w3480 , w3481 , w3482 , w3483 , w3484 , w3485 , w3486 , w3487 , w3488 , w3489 , w3490 , w3491 , w3492 , w3493 , w3494 , w3495 , w3496 , w3497 , w3498 , w3499 , w3500 , w3501 , w3502 , w3503 , w3504 , w3505 , w3506 , w3507 , w3508 , w3509 , w3510 , w3511 , w3512 , w3513 , w3514 , w3515 , w3516 , w3517 , w3518 , w3519 , w3520 , w3521 , w3522 , w3523 , w3524 , w3525 , w3526 , w3527 , w3528 , w3529 , w3530 , w3531 , w3532 , w3533 , w3534 , w3535 , w3536 , w3537 , w3538 , w3539 , w3540 , w3541 , w3542 , w3543 , w3544 , w3545 , w3546 , w3547 , w3548 , w3549 , w3550 , w3551 , w3552 , w3553 , w3554 , w3555 , w3556 , w3557 , w3558 , w3559 , w3560 , w3561 , w3562 , w3563 , w3564 , w3565 , w3566 , w3567 , w3568 , w3569 , w3570 , w3571 , w3572 , w3573 , w3574 , w3575 , w3576 , w3577 , w3578 , w3579 , w3580 , w3581 , w3582 , w3583 , w3584 , w3585 , w3586 , w3587 , w3588 , w3589 , w3590 , w3591 , w3592 , w3593 , w3594 , w3595 , w3596 , w3597 , w3598 , w3599 , w3600 , w3601 , w3602 , w3603 , w3604 , w3605 , w3606 , w3607 , w3608 , w3609 , w3610 , w3611 , w3612 , w3613 , w3614 , w3615 , w3616 , w3617 , w3618 , w3619 , w3620 , w3621 , w3622 , w3623 , w3624 , w3625 , w3626 , w3627 , w3628 , w3629 , w3630 , w3631 , w3632 , w3633 , w3634 , w3635 , w3636 , w3637 , w3638 , w3639 , w3640 , w3641 , w3642 , w3643 , w3644 , w3645 , w3646 , w3647 , w3648 , w3649 , w3650 , w3651 , w3652 , w3653 , w3654 , w3655 , w3656 , w3657 , w3658 , w3659 , w3660 , w3661 , w3662 , w3663 , w3664 , w3665 , w3666 , w3667 , w3668 , w3669 , w3670 , w3671 , w3672 , w3673 , w3674 , w3675 , w3676 , w3677 , w3678 , w3679 , w3680 , w3681 , w3682 , w3683 , w3684 , w3685 , w3686 , w3687 , w3688 , w3689 , w3690 , w3691 , w3692 , w3693 , w3694 , w3695 , w3696 , w3697 , w3698 , w3699 , w3700 , w3701 , w3702 , w3703 , w3704 , w3705 , w3706 , w3707 , w3708 , w3709 , w3710 , w3711 , w3712 , w3713 , w3714 , w3715 , w3716 , w3717 , w3718 , w3719 , w3720 , w3721 , w3722 , w3723 , w3724 , w3725 , w3726 , w3727 , w3728 , w3729 , w3730 , w3731 , w3732 , w3733 , w3734 , w3735 , w3736 , w3737 , w3738 , w3739 , w3740 , w3741 , w3742 , w3743 , w3744 , w3745 , w3746 , w3747 , w3748 , w3749 , w3750 , w3751 , w3752 , w3753 , w3754 , w3755 , w3756 , w3757 , w3758 , w3759 , w3760 , w3761 , w3762 , w3763 , w3764 , w3765 , w3766 , w3767 , w3768 , w3769 , w3770 , w3771 , w3772 , w3773 , w3774 , w3775 , w3776 , w3777 , w3778 , w3779 , w3780 , w3781 , w3782 , w3783 , w3784 , w3785 , w3786 , w3787 , w3788 , w3789 , w3790 , w3791 , w3792 , w3793 , w3794 , w3795 , w3796 , w3797 , w3798 , w3799 , w3800 , w3801 , w3802 , w3803 , w3804 , w3805 , w3806 , w3807 , w3808 , w3809 , w3810 , w3811 , w3812 , w3813 , w3814 , w3815 , w3816 , w3817 , w3818 , w3819 , w3820 , w3821 , w3822 , w3823 , w3824 , w3825 , w3826 , w3827 , w3828 , w3829 , w3830 , w3831 , w3832 , w3833 , w3834 , w3835 , w3836 , w3837 , w3838 , w3839 , w3840 , w3841 , w3842 , w3843 , w3844 , w3845 , w3846 , w3847 , w3848 , w3849 , w3850 , w3851 , w3852 , w3853 , w3854 , w3855 , w3856 , w3857 , w3858 , w3859 , w3860 , w3861 , w3862 , w3863 , w3864 , w3865 , w3866 , w3867 , w3868 , w3869 , w3870 , w3871 , w3872 , w3873 , w3874 , w3875 , w3876 , w3877 , w3878 , w3879 , w3880 , w3881 , w3882 , w3883 , w3884 , w3885 , w3886 , w3887 , w3888 , w3889 , w3890 , w3891 , w3892 , w3893 , w3894 , w3895 , w3896 , w3897 , w3898 , w3899 , w3900 , w3901 , w3902 , w3903 , w3904 , w3905 , w3906 , w3907 , w3908 , w3909 , w3910 , w3911 , w3912 , w3913 , w3914 , w3915 , w3916 , w3917 , w3918 , w3919 , w3920 , w3921 , w3922 , w3923 , w3924 , w3925 , w3926 , w3927 , w3928 , w3929 , w3930 , w3931 , w3932 , w3933 , w3934 , w3935 , w3936 , w3937 , w3938 , w3939 , w3940 , w3941 , w3942 , w3943 , w3944 , w3945 , w3946 , w3947 , w3948 , w3949 , w3950 , w3951 , w3952 , w3953 , w3954 , w3955 , w3956 , w3957 , w3958 , w3959 , w3960 , w3961 , w3962 , w3963 , w3964 , w3965 , w3966 , w3967 , w3968 , w3969 , w3970 , w3971 , w3972 , w3973 , w3974 , w3975 , w3976 , w3977 , w3978 , w3979 , w3980 , w3981 , w3982 , w3983 , w3984 , w3985 , w3986 , w3987 , w3988 , w3989 , w3990 , w3991 , w3992 , w3993 , w3994 , w3995 , w3996 , w3997 , w3998 , w3999 , w4000 , w4001 , w4002 , w4003 , w4004 , w4005 , w4006 , w4007 , w4008 , w4009 , w4010 , w4011 , w4012 , w4013 , w4014 , w4015 , w4016 , w4017 , w4018 , w4019 , w4020 , w4021 , w4022 , w4023 , w4024 , w4025 , w4026 , w4027 , w4028 , w4029 , w4030 , w4031 , w4032 , w4033 , w4034 , w4035 , w4036 , w4037 , w4038 , w4039 , w4040 , w4041 , w4042 , w4043 , w4044 , w4045 , w4046 , w4047 , w4048 , w4049 , w4050 , w4051 , w4052 , w4053 , w4054 , w4055 , w4056 , w4057 , w4058 , w4059 , w4060 , w4061 , w4062 , w4063 , w4064 , w4065 , w4066 , w4067 , w4068 , w4069 , w4070 , w4071 , w4072 , w4073 , w4074 , w4075 , w4076 , w4077 , w4078 , w4079 , w4080 , w4081 , w4082 , w4083 , w4084 , w4085 , w4086 , w4087 , w4088 , w4089 , w4090 , w4091 , w4092 , w4093 , w4094 , w4095 , w4096 , w4097 , w4098 , w4099 , w4100 , w4101 , w4102 , w4103 , w4104 , w4105 , w4106 , w4107 , w4108 , w4109 , w4110 , w4111 , w4112 , w4113 , w4114 , w4115 , w4116 , w4117 , w4118 , w4119 , w4120 , w4121 , w4122 , w4123 , w4124 , w4125 , w4126 , w4127 , w4128 , w4129 , w4130 , w4131 , w4132 , w4133 , w4134 , w4135 , w4136 , w4137 , w4138 , w4139 , w4140 , w4141 , w4142 , w4143 , w4144 , w4145 , w4146 , w4147 , w4148 , w4149 , w4150 , w4151 , w4152 , w4153 , w4154 , w4155 , w4156 , w4157 , w4158 , w4159 , w4160 , w4161 , w4162 , w4163 , w4164 , w4165 , w4166 , w4167 , w4168 , w4169 , w4170 , w4171 , w4172 , w4173 , w4174 , w4175 , w4176 , w4177 , w4178 , w4179 , w4180 , w4181 , w4182 , w4183 , w4184 , w4185 , w4186 , w4187 , w4188 , w4189 , w4190 , w4191 , w4192 , w4193 , w4194 , w4195 , w4196 , w4197 , w4198 , w4199 , w4200 , w4201 , w4202 , w4203 , w4204 , w4205 , w4206 , w4207 , w4208 , w4209 , w4210 , w4211 , w4212 , w4213 , w4214 , w4215 , w4216 , w4217 , w4218 , w4219 , w4220 , w4221 , w4222 , w4223 , w4224 , w4225 , w4226 , w4227 , w4228 , w4229 , w4230 , w4231 , w4232 , w4233 , w4234 , w4235 , w4236 , w4237 , w4238 , w4239 , w4240 , w4241 , w4242 , w4243 , w4244 , w4245 , w4246 , w4247 , w4248 , w4249 , w4250 , w4251 , w4252 , w4253 , w4254 , w4255 , w4256 , w4257 , w4258 , w4259 , w4260 , w4261 , w4262 , w4263 , w4264 , w4265 , w4266 , w4267 , w4268 , w4269 , w4270 , w4271 , w4272 , w4273 , w4274 , w4275 , w4276 , w4277 , w4278 , w4279 , w4280 , w4281 , w4282 , w4283 , w4284 , w4285 , w4286 , w4287 , w4288 , w4289 , w4290 , w4291 , w4292 , w4293 , w4294 , w4295 , w4296 , w4297 , w4298 , w4299 , w4300 , w4301 , w4302 , w4303 , w4304 , w4305 , w4306 , w4307 , w4308 , w4309 , w4310 , w4311 , w4312 , w4313 , w4314 , w4315 , w4316 , w4317 , w4318 , w4319 , w4320 , w4321 , w4322 , w4323 , w4324 , w4325 , w4326 , w4327 , w4328 , w4329 , w4330 , w4331 , w4332 , w4333 , w4334 , w4335 , w4336 , w4337 , w4338 , w4339 , w4340 , w4341 , w4342 , w4343 , w4344 , w4345 , w4346 , w4347 , w4348 , w4349 , w4350 , w4351 , w4352 , w4353 , w4354 , w4355 , w4356 , w4357 , w4358 , w4359 , w4360 , w4361 , w4362 , w4363 , w4364 , w4365 , w4366 , w4367 , w4368 , w4369 , w4370 , w4371 , w4372 , w4373 , w4374 , w4375 , w4376 , w4377 , w4378 , w4379 , w4380 , w4381 , w4382 , w4383 , w4384 , w4385 , w4386 , w4387 , w4388 , w4389 , w4390 , w4391 , w4392 , w4393 , w4394 , w4395 , w4396 , w4397 , w4398 , w4399 , w4400 , w4401 , w4402 , w4403 , w4404 , w4405 , w4406 , w4407 , w4408 , w4409 , w4410 , w4411 , w4412 , w4413 , w4414 , w4415 , w4416 , w4417 , w4418 , w4419 , w4420 , w4421 , w4422 , w4423 , w4424 , w4425 , w4426 , w4427 , w4428 , w4429 , w4430 , w4431 , w4432 , w4433 , w4434 , w4435 , w4436 , w4437 , w4438 , w4439 , w4440 , w4441 , w4442 , w4443 , w4444 , w4445 , w4446 , w4447 , w4448 , w4449 , w4450 , w4451 , w4452 , w4453 , w4454 , w4455 , w4456 , w4457 , w4458 , w4459 , w4460 , w4461 , w4462 , w4463 , w4464 , w4465 , w4466 , w4467 , w4468 , w4469 , w4470 , w4471 , w4472 , w4473 , w4474 , w4475 , w4476 , w4477 , w4478 , w4479 , w4480 , w4481 , w4482 , w4483 , w4484 , w4485 , w4486 , w4487 , w4488 , w4489 , w4490 , w4491 , w4492 , w4493 , w4494 , w4495 , w4496 , w4497 , w4498 , w4499 , w4500 , w4501 , w4502 , w4503 , w4504 , w4505 , w4506 , w4507 , w4508 , w4509 , w4510 , w4511 , w4512 , w4513 , w4514 , w4515 , w4516 , w4517 , w4518 , w4519 , w4520 , w4521 , w4522 , w4523 , w4524 , w4525 , w4526 , w4527 , w4528 , w4529 , w4530 , w4531 , w4532 , w4533 , w4534 , w4535 , w4536 , w4537 , w4538 , w4539 , w4540 , w4541 , w4542 , w4543 , w4544 , w4545 , w4546 , w4547 , w4548 , w4549 , w4550 , w4551 , w4552 , w4553 , w4554 , w4555 , w4556 , w4557 , w4558 , w4559 , w4560 , w4561 , w4562 , w4563 , w4564 , w4565 , w4566 , w4567 , w4568 , w4569 , w4570 , w4571 , w4572 , w4573 , w4574 , w4575 , w4576 , w4577 , w4578 , w4579 , w4580 , w4581 , w4582 , w4583 , w4584 , w4585 , w4586 , w4587 , w4588 , w4589 , w4590 , w4591 , w4592 , w4593 , w4594 , w4595 , w4596 , w4597 , w4598 , w4599 , w4600 , w4601 , w4602 , w4603 , w4604 , w4605 , w4606 , w4607 , w4608 , w4609 , w4610 , w4611 , w4612 , w4613 , w4614 , w4615 , w4616 , w4617 , w4618 , w4619 , w4620 , w4621 , w4622 , w4623 , w4624 , w4625 , w4626 , w4627 , w4628 , w4629 , w4630 , w4631 , w4632 , w4633 , w4634 , w4635 , w4636 , w4637 , w4638 , w4639 , w4640 , w4641 , w4642 , w4643 , w4644 , w4645 , w4646 , w4647 , w4648 , w4649 , w4650 , w4651 , w4652 , w4653 , w4654 , w4655 , w4656 , w4657 , w4658 , w4659 , w4660 , w4661 , w4662 , w4663 , w4664 , w4665 , w4666 , w4667 , w4668 , w4669 , w4670 , w4671 , w4672 , w4673 , w4674 , w4675 , w4676 , w4677 , w4678 , w4679 , w4680 , w4681 , w4682 , w4683 , w4684 , w4685 , w4686 , w4687 , w4688 , w4689 , w4690 , w4691 , w4692 , w4693 , w4694 , w4695 , w4696 , w4697 , w4698 , w4699 , w4700 , w4701 , w4702 , w4703 , w4704 , w4705 , w4706 , w4707 , w4708 , w4709 , w4710 , w4711 , w4712 , w4713 , w4714 , w4715 , w4716 , w4717 , w4718 , w4719 , w4720 , w4721 , w4722 , w4723 , w4724 , w4725 , w4726 , w4727 , w4728 , w4729 , w4730 , w4731 , w4732 , w4733 , w4734 , w4735 , w4736 , w4737 , w4738 , w4739 , w4740 , w4741 , w4742 , w4743 , w4744 , w4745 , w4746 , w4747 , w4748 , w4749 , w4750 , w4751 , w4752 , w4753 , w4754 , w4755 , w4756 , w4757 , w4758 , w4759 , w4760 , w4761 , w4762 , w4763 , w4764 , w4765 , w4766 , w4767 , w4768 , w4769 , w4770 , w4771 , w4772 , w4773 , w4774 , w4775 , w4776 , w4777 , w4778 , w4779 , w4780 , w4781 , w4782 , w4783 , w4784 , w4785 , w4786 , w4787 , w4788 , w4789 , w4790 , w4791 , w4792 , w4793 , w4794 , w4795 , w4796 , w4797 , w4798 , w4799 , w4800 , w4801 , w4802 , w4803 , w4804 , w4805 , w4806 , w4807 , w4808 , w4809 , w4810 , w4811 , w4812 , w4813 , w4814 , w4815 , w4816 , w4817 , w4818 , w4819 , w4820 , w4821 , w4822 , w4823 , w4824 , w4825 , w4826 , w4827 , w4828 , w4829 , w4830 , w4831 , w4832 , w4833 , w4834 , w4835 , w4836 , w4837 , w4838 , w4839 , w4840 , w4841 , w4842 , w4843 , w4844 , w4845 , w4846 , w4847 , w4848 , w4849 , w4850 , w4851 , w4852 , w4853 , w4854 , w4855 , w4856 , w4857 , w4858 , w4859 , w4860 , w4861 , w4862 , w4863 , w4864 , w4865 , w4866 , w4867 , w4868 , w4869 , w4870 , w4871 , w4872 , w4873 , w4874 , w4875 , w4876 , w4877 , w4878 , w4879 , w4880 , w4881 , w4882 , w4883 , w4884 , w4885 , w4886 , w4887 , w4888 , w4889 , w4890 , w4891 , w4892 , w4893 , w4894 , w4895 , w4896 , w4897 , w4898 , w4899 , w4900 , w4901 , w4902 , w4903 , w4904 , w4905 , w4906 , w4907 , w4908 , w4909 , w4910 , w4911 , w4912 , w4913 , w4914 , w4915 , w4916 , w4917 , w4918 , w4919 , w4920 , w4921 , w4922 , w4923 , w4924 , w4925 , w4926 , w4927 , w4928 , w4929 , w4930 , w4931 , w4932 , w4933 , w4934 , w4935 , w4936 , w4937 , w4938 , w4939 , w4940 , w4941 , w4942 , w4943 , w4944 , w4945 , w4946 , w4947 , w4948 , w4949 , w4950 , w4951 , w4952 , w4953 , w4954 , w4955 , w4956 , w4957 , w4958 , w4959 , w4960 , w4961 , w4962 , w4963 , w4964 , w4965 , w4966 , w4967 , w4968 , w4969 , w4970 , w4971 , w4972 , w4973 , w4974 , w4975 , w4976 , w4977 , w4978 , w4979 , w4980 , w4981 , w4982 , w4983 , w4984 , w4985 , w4986 , w4987 , w4988 , w4989 , w4990 , w4991 , w4992 , w4993 , w4994 , w4995 , w4996 , w4997 , w4998 , w4999 , w5000 , w5001 , w5002 , w5003 , w5004 , w5005 , w5006 , w5007 , w5008 , w5009 , w5010 , w5011 , w5012 , w5013 , w5014 , w5015 , w5016 , w5017 , w5018 , w5019 , w5020 , w5021 , w5022 , w5023 , w5024 , w5025 , w5026 , w5027 , w5028 , w5029 , w5030 , w5031 , w5032 , w5033 , w5034 , w5035 , w5036 , w5037 , w5038 , w5039 , w5040 , w5041 , w5042 , w5043 , w5044 , w5045 , w5046 , w5047 , w5048 , w5049 , w5050 , w5051 , w5052 , w5053 , w5054 , w5055 , w5056 , w5057 , w5058 , w5059 , w5060 , w5061 , w5062 , w5063 , w5064 , w5065 , w5066 , w5067 , w5068 , w5069 , w5070 , w5071 , w5072 , w5073 , w5074 , w5075 , w5076 , w5077 , w5078 , w5079 , w5080 , w5081 , w5082 , w5083 , w5084 , w5085 , w5086 , w5087 , w5088 , w5089 , w5090 , w5091 , w5092 , w5093 , w5094 , w5095 , w5096 , w5097 , w5098 , w5099 , w5100 , w5101 , w5102 , w5103 , w5104 , w5105 , w5106 , w5107 , w5108 , w5109 , w5110 , w5111 , w5112 , w5113 , w5114 , w5115 , w5116 , w5117 , w5118 , w5119 , w5120 , w5121 , w5122 , w5123 , w5124 , w5125 , w5126 , w5127 , w5128 , w5129 , w5130 , w5131 , w5132 , w5133 , w5134 , w5135 , w5136 , w5137 , w5138 , w5139 , w5140 , w5141 , w5142 , w5143 , w5144 , w5145 , w5146 , w5147 , w5148 , w5149 , w5150 , w5151 , w5152 , w5153 , w5154 , w5155 , w5156 , w5157 , w5158 , w5159 , w5160 , w5161 , w5162 , w5163 , w5164 , w5165 , w5166 , w5167 , w5168 , w5169 , w5170 , w5171 , w5172 , w5173 , w5174 , w5175 , w5176 , w5177 , w5178 , w5179 , w5180 , w5181 , w5182 , w5183 , w5184 , w5185 , w5186 , w5187 , w5188 , w5189 , w5190 , w5191 , w5192 , w5193 , w5194 , w5195 , w5196 , w5197 , w5198 , w5199 , w5200 , w5201 , w5202 , w5203 , w5204 , w5205 , w5206 , w5207 , w5208 , w5209 , w5210 , w5211 , w5212 , w5213 , w5214 , w5215 , w5216 , w5217 , w5218 , w5219 , w5220 , w5221 , w5222 , w5223 , w5224 , w5225 , w5226 , w5227 , w5228 , w5229 , w5230 , w5231 , w5232 , w5233 , w5234 , w5235 , w5236 , w5237 , w5238 , w5239 , w5240 , w5241 , w5242 , w5243 , w5244 , w5245 , w5246 , w5247 , w5248 , w5249 , w5250 , w5251 , w5252 , w5253 , w5254 , w5255 , w5256 , w5257 , w5258 , w5259 , w5260 , w5261 , w5262 , w5263 , w5264 , w5265 , w5266 , w5267 , w5268 , w5269 , w5270 , w5271 , w5272 , w5273 , w5274 , w5275 , w5276 , w5277 , w5278 , w5279 , w5280 , w5281 , w5282 , w5283 , w5284 , w5285 , w5286 , w5287 , w5288 , w5289 , w5290 , w5291 , w5292 , w5293 , w5294 , w5295 , w5296 , w5297 , w5298 , w5299 , w5300 , w5301 , w5302 , w5303 , w5304 , w5305 , w5306 , w5307 , w5308 , w5309 , w5310 , w5311 , w5312 , w5313 , w5314 , w5315 , w5316 , w5317 , w5318 , w5319 , w5320 , w5321 , w5322 , w5323 , w5324 , w5325 , w5326 , w5327 , w5328 , w5329 , w5330 , w5331 , w5332 , w5333 , w5334 , w5335 , w5336 , w5337 , w5338 , w5339 , w5340 , w5341 , w5342 , w5343 , w5344 , w5345 , w5346 , w5347 , w5348 , w5349 , w5350 , w5351 , w5352 , w5353 , w5354 , w5355 , w5356 , w5357 , w5358 , w5359 , w5360 , w5361 , w5362 , w5363 , w5364 , w5365 , w5366 , w5367 , w5368 , w5369 , w5370 , w5371 , w5372 , w5373 , w5374 , w5375 , w5376 , w5377 , w5378 , w5379 , w5380 , w5381 , w5382 , w5383 , w5384 , w5385 , w5386 , w5387 , w5388 , w5389 , w5390 , w5391 , w5392 , w5393 , w5394 , w5395 , w5396 , w5397 , w5398 , w5399 , w5400 , w5401 , w5402 , w5403 , w5404 , w5405 , w5406 , w5407 , w5408 , w5409 , w5410 , w5411 , w5412 , w5413 , w5414 , w5415 , w5416 , w5417 , w5418 , w5419 , w5420 , w5421 , w5422 , w5423 , w5424 , w5425 , w5426 , w5427 , w5428 , w5429 , w5430 , w5431 , w5432 , w5433 , w5434 , w5435 , w5436 , w5437 , w5438 , w5439 , w5440 , w5441 , w5442 , w5443 , w5444 , w5445 , w5446 , w5447 , w5448 , w5449 , w5450 , w5451 , w5452 , w5453 , w5454 , w5455 , w5456 , w5457 , w5458 , w5459 , w5460 , w5461 , w5462 , w5463 , w5464 , w5465 , w5466 , w5467 , w5468 , w5469 , w5470 , w5471 , w5472 , w5473 , w5474 , w5475 , w5476 , w5477 , w5478 , w5479 , w5480 , w5481 , w5482 , w5483 , w5484 , w5485 , w5486 , w5487 , w5488 , w5489 , w5490 , w5491 , w5492 , w5493 , w5494 , w5495 , w5496 , w5497 , w5498 , w5499 , w5500 , w5501 , w5502 , w5503 , w5504 , w5505 , w5506 , w5507 , w5508 , w5509 , w5510 , w5511 , w5512 , w5513 , w5514 , w5515 , w5516 , w5517 , w5518 , w5519 , w5520 , w5521 , w5522 , w5523 , w5524 , w5525 , w5526 , w5527 , w5528 , w5529 , w5530 , w5531 , w5532 , w5533 , w5534 , w5535 , w5536 , w5537 , w5538 , w5539 , w5540 , w5541 , w5542 , w5543 , w5544 , w5545 , w5546 , w5547 , w5548 , w5549 , w5550 , w5551 , w5552 , w5553 , w5554 , w5555 , w5556 , w5557 , w5558 , w5559 , w5560 , w5561 , w5562 , w5563 , w5564 , w5565 , w5566 , w5567 , w5568 , w5569 , w5570 , w5571 , w5572 , w5573 , w5574 , w5575 , w5576 , w5577 , w5578 , w5579 , w5580 , w5581 , w5582 , w5583 , w5584 , w5585 , w5586 , w5587 , w5588 , w5589 , w5590 , w5591 , w5592 , w5593 , w5594 , w5595 , w5596 , w5597 , w5598 , w5599 , w5600 , w5601 , w5602 , w5603 , w5604 , w5605 , w5606 , w5607 , w5608 , w5609 , w5610 , w5611 , w5612 , w5613 , w5614 , w5615 , w5616 , w5617 , w5618 , w5619 , w5620 , w5621 , w5622 , w5623 , w5624 , w5625 , w5626 , w5627 , w5628 , w5629 , w5630 , w5631 , w5632 , w5633 , w5634 , w5635 , w5636 , w5637 , w5638 , w5639 , w5640 , w5641 , w5642 , w5643 , w5644 , w5645 , w5646 , w5647 , w5648 , w5649 , w5650 , w5651 , w5652 , w5653 , w5654 , w5655 , w5656 , w5657 , w5658 , w5659 , w5660 , w5661 , w5662 , w5663 , w5664 , w5665 , w5666 , w5667 , w5668 , w5669 , w5670 , w5671 , w5672 , w5673 , w5674 , w5675 , w5676 , w5677 , w5678 , w5679 , w5680 , w5681 , w5682 , w5683 , w5684 , w5685 , w5686 , w5687 , w5688 , w5689 , w5690 , w5691 , w5692 , w5693 , w5694 , w5695 , w5696 , w5697 , w5698 , w5699 , w5700 , w5701 , w5702 , w5703 , w5704 , w5705 , w5706 , w5707 , w5708 , w5709 , w5710 , w5711 , w5712 , w5713 , w5714 , w5715 , w5716 , w5717 , w5718 , w5719 , w5720 , w5721 , w5722 , w5723 , w5724 , w5725 , w5726 , w5727 , w5728 , w5729 , w5730 , w5731 , w5732 , w5733 , w5734 , w5735 , w5736 , w5737 , w5738 , w5739 , w5740 , w5741 , w5742 , w5743 , w5744 , w5745 , w5746 , w5747 , w5748 , w5749 , w5750 , w5751 , w5752 , w5753 , w5754 , w5755 , w5756 , w5757 , w5758 , w5759 , w5760 , w5761 , w5762 , w5763 , w5764 , w5765 , w5766 , w5767 , w5768 , w5769 , w5770 , w5771 , w5772 , w5773 , w5774 , w5775 , w5776 , w5777 , w5778 , w5779 , w5780 , w5781 , w5782 , w5783 , w5784 , w5785 , w5786 , w5787 , w5788 , w5789 , w5790 , w5791 , w5792 , w5793 , w5794 , w5795 , w5796 , w5797 , w5798 , w5799 , w5800 , w5801 , w5802 , w5803 , w5804 , w5805 , w5806 , w5807 , w5808 , w5809 , w5810 , w5811 , w5812 , w5813 , w5814 , w5815 , w5816 , w5817 , w5818 , w5819 , w5820 , w5821 , w5822 , w5823 , w5824 , w5825 , w5826 , w5827 , w5828 , w5829 , w5830 , w5831 , w5832 , w5833 , w5834 , w5835 , w5836 , w5837 , w5838 , w5839 , w5840 , w5841 , w5842 , w5843 , w5844 , w5845 , w5846 , w5847 , w5848 , w5849 , w5850 , w5851 , w5852 , w5853 , w5854 , w5855 , w5856 , w5857 , w5858 , w5859 , w5860 , w5861 , w5862 , w5863 , w5864 , w5865 , w5866 , w5867 , w5868 , w5869 , w5870 , w5871 , w5872 , w5873 , w5874 , w5875 , w5876 , w5877 , w5878 , w5879 , w5880 , w5881 , w5882 , w5883 , w5884 , w5885 , w5886 , w5887 , w5888 , w5889 , w5890 , w5891 , w5892 , w5893 , w5894 , w5895 , w5896 , w5897 , w5898 , w5899 , w5900 , w5901 , w5902 , w5903 , w5904 , w5905 , w5906 , w5907 , w5908 , w5909 , w5910 , w5911 , w5912 , w5913 , w5914 , w5915 , w5916 , w5917 , w5918 , w5919 , w5920 , w5921 , w5922 , w5923 , w5924 , w5925 , w5926 , w5927 , w5928 , w5929 , w5930 , w5931 , w5932 , w5933 , w5934 , w5935 , w5936 , w5937 , w5938 , w5939 , w5940 , w5941 , w5942 , w5943 , w5944 , w5945 , w5946 , w5947 , w5948 , w5949 , w5950 , w5951 , w5952 , w5953 , w5954 , w5955 , w5956 , w5957 , w5958 , w5959 , w5960 , w5961 , w5962 , w5963 , w5964 , w5965 , w5966 , w5967 , w5968 , w5969 , w5970 , w5971 , w5972 , w5973 , w5974 , w5975 , w5976 , w5977 , w5978 , w5979 , w5980 , w5981 , w5982 , w5983 , w5984 , w5985 , w5986 , w5987 , w5988 , w5989 , w5990 , w5991 , w5992 , w5993 , w5994 , w5995 , w5996 , w5997 , w5998 , w5999 , w6000 , w6001 , w6002 , w6003 , w6004 , w6005 , w6006 , w6007 , w6008 , w6009 , w6010 , w6011 , w6012 , w6013 , w6014 , w6015 , w6016 , w6017 , w6018 , w6019 , w6020 , w6021 , w6022 , w6023 , w6024 , w6025 , w6026 , w6027 , w6028 , w6029 , w6030 , w6031 , w6032 , w6033 , w6034 , w6035 , w6036 , w6037 , w6038 , w6039 , w6040 , w6041 , w6042 , w6043 , w6044 , w6045 , w6046 , w6047 , w6048 , w6049 , w6050 , w6051 , w6052 , w6053 , w6054 , w6055 , w6056 , w6057 , w6058 , w6059 , w6060 , w6061 , w6062 , w6063 , w6064 , w6065 , w6066 , w6067 , w6068 , w6069 , w6070 , w6071 , w6072 , w6073 , w6074 , w6075 , w6076 , w6077 , w6078 , w6079 , w6080 , w6081 , w6082 , w6083 , w6084 , w6085 , w6086 , w6087 , w6088 , w6089 , w6090 , w6091 , w6092 , w6093 , w6094 , w6095 , w6096 , w6097 , w6098 , w6099 , w6100 , w6101 , w6102 , w6103 , w6104 , w6105 , w6106 , w6107 , w6108 , w6109 , w6110 , w6111 , w6112 , w6113 , w6114 , w6115 , w6116 , w6117 , w6118 , w6119 , w6120 , w6121 , w6122 , w6123 , w6124 , w6125 , w6126 , w6127 , w6128 , w6129 , w6130 , w6131 , w6132 , w6133 , w6134 , w6135 , w6136 , w6137 , w6138 , w6139 , w6140 , w6141 , w6142 , w6143 , w6144 , w6145 , w6146 , w6147 , w6148 , w6149 , w6150 , w6151 , w6152 , w6153 , w6154 , w6155 , w6156 , w6157 , w6158 , w6159 , w6160 , w6161 , w6162 , w6163 , w6164 , w6165 , w6166 , w6167 , w6168 , w6169 , w6170 , w6171 , w6172 , w6173 , w6174 , w6175 , w6176 , w6177 , w6178 , w6179 , w6180 , w6181 , w6182 , w6183 , w6184 , w6185 , w6186 , w6187 , w6188 , w6189 , w6190 , w6191 , w6192 , w6193 , w6194 , w6195 , w6196 , w6197 , w6198 , w6199 , w6200 , w6201 , w6202 , w6203 , w6204 , w6205 , w6206 , w6207 , w6208 , w6209 , w6210 , w6211 , w6212 , w6213 , w6214 , w6215 , w6216 , w6217 , w6218 , w6219 , w6220 , w6221 , w6222 , w6223 , w6224 , w6225 , w6226 , w6227 , w6228 , w6229 , w6230 , w6231 , w6232 , w6233 , w6234 , w6235 , w6236 , w6237 , w6238 , w6239 , w6240 , w6241 , w6242 , w6243 , w6244 , w6245 , w6246 , w6247 , w6248 , w6249 , w6250 , w6251 , w6252 , w6253 , w6254 , w6255 , w6256 , w6257 , w6258 , w6259 , w6260 , w6261 , w6262 , w6263 , w6264 , w6265 , w6266 , w6267 , w6268 , w6269 , w6270 , w6271 , w6272 , w6273 , w6274 , w6275 , w6276 , w6277 , w6278 , w6279 , w6280 , w6281 , w6282 , w6283 , w6284 , w6285 , w6286 , w6287 , w6288 , w6289 , w6290 , w6291 , w6292 , w6293 , w6294 , w6295 , w6296 , w6297 , w6298 , w6299 , w6300 , w6301 , w6302 , w6303 , w6304 , w6305 , w6306 , w6307 , w6308 , w6309 , w6310 , w6311 , w6312 , w6313 , w6314 , w6315 , w6316 , w6317 , w6318 , w6319 , w6320 , w6321 , w6322 , w6323 , w6324 , w6325 , w6326 , w6327 , w6328 , w6329 , w6330 , w6331 , w6332 , w6333 , w6334 , w6335 , w6336 , w6337 , w6338 , w6339 , w6340 , w6341 , w6342 , w6343 , w6344 , w6345 , w6346 , w6347 , w6348 , w6349 , w6350 , w6351 , w6352 , w6353 , w6354 , w6355 , w6356 , w6357 , w6358 , w6359 , w6360 , w6361 , w6362 , w6363 , w6364 , w6365 , w6366 , w6367 , w6368 , w6369 , w6370 , w6371 , w6372 , w6373 , w6374 , w6375 , w6376 , w6377 , w6378 , w6379 , w6380 , w6381 , w6382 , w6383 , w6384 , w6385 , w6386 , w6387 , w6388 , w6389 , w6390 , w6391 , w6392 , w6393 , w6394 , w6395 , w6396 , w6397 , w6398 , w6399 , w6400 , w6401 , w6402 , w6403 , w6404 , w6405 , w6406 , w6407 , w6408 , w6409 , w6410 , w6411 , w6412 , w6413 , w6414 , w6415 , w6416 , w6417 , w6418 , w6419 , w6420 , w6421 , w6422 , w6423 , w6424 , w6425 , w6426 , w6427 , w6428 , w6429 , w6430 , w6431 , w6432 , w6433 , w6434 , w6435 , w6436 , w6437 , w6438 , w6439 , w6440 , w6441 , w6442 , w6443 , w6444 , w6445 , w6446 , w6447 , w6448 , w6449 , w6450 , w6451 , w6452 , w6453 , w6454 , w6455 , w6456 , w6457 , w6458 , w6459 , w6460 , w6461 , w6462 , w6463 , w6464 , w6465 , w6466 , w6467 , w6468 , w6469 , w6470 , w6471 , w6472 , w6473 , w6474 , w6475 , w6476 , w6477 , w6478 , w6479 , w6480 , w6481 , w6482 , w6483 , w6484 , w6485 , w6486 , w6487 , w6488 , w6489 , w6490 , w6491 , w6492 , w6493 , w6494 , w6495 , w6496 , w6497 , w6498 , w6499 , w6500 , w6501 , w6502 , w6503 , w6504 , w6505 , w6506 , w6507 , w6508 , w6509 , w6510 , w6511 , w6512 , w6513 , w6514 , w6515 , w6516 , w6517 , w6518 , w6519 , w6520 , w6521 , w6522 , w6523 , w6524 , w6525 , w6526 , w6527 , w6528 , w6529 , w6530 , w6531 , w6532 , w6533 , w6534 , w6535 , w6536 , w6537 , w6538 , w6539 , w6540 , w6541 , w6542 , w6543 , w6544 , w6545 , w6546 , w6547 , w6548 , w6549 , w6550 , w6551 , w6552 , w6553 , w6554 , w6555 , w6556 , w6557 , w6558 , w6559 , w6560 , w6561 , w6562 , w6563 , w6564 , w6565 , w6566 , w6567 , w6568 , w6569 , w6570 , w6571 , w6572 , w6573 , w6574 , w6575 , w6576 , w6577 , w6578 , w6579 , w6580 , w6581 , w6582 , w6583 , w6584 , w6585 , w6586 , w6587 , w6588 , w6589 , w6590 , w6591 , w6592 , w6593 , w6594 , w6595 , w6596 , w6597 , w6598 , w6599 , w6600 , w6601 , w6602 , w6603 , w6604 , w6605 , w6606 , w6607 , w6608 , w6609 , w6610 , w6611 , w6612 , w6613 , w6614 , w6615 , w6616 , w6617 , w6618 , w6619 , w6620 , w6621 , w6622 , w6623 , w6624 , w6625 , w6626 , w6627 , w6628 , w6629 , w6630 , w6631 , w6632 , w6633 , w6634 , w6635 , w6636 , w6637 , w6638 , w6639 , w6640 , w6641 , w6642 , w6643 , w6644 , w6645 , w6646 , w6647 , w6648 , w6649 , w6650 , w6651 , w6652 , w6653 , w6654 , w6655 , w6656 , w6657 , w6658 , w6659 , w6660 , w6661 , w6662 , w6663 , w6664 , w6665 , w6666 , w6667 , w6668 , w6669 , w6670 , w6671 , w6672 , w6673 , w6674 , w6675 , w6676 , w6677 , w6678 , w6679 , w6680 , w6681 , w6682 , w6683 , w6684 , w6685 , w6686 , w6687 , w6688 , w6689 , w6690 , w6691 , w6692 , w6693 , w6694 , w6695 , w6696 , w6697 , w6698 , w6699 , w6700 , w6701 , w6702 , w6703 , w6704 , w6705 , w6706 , w6707 , w6708 , w6709 , w6710 , w6711 , w6712 , w6713 , w6714 , w6715 , w6716 , w6717 , w6718 , w6719 , w6720 , w6721 , w6722 , w6723 , w6724 , w6725 , w6726 , w6727 , w6728 , w6729 , w6730 , w6731 , w6732 , w6733 , w6734 , w6735 , w6736 , w6737 , w6738 , w6739 , w6740 , w6741 , w6742 , w6743 , w6744 , w6745 , w6746 , w6747 , w6748 , w6749 , w6750 , w6751 , w6752 , w6753 , w6754 , w6755 , w6756 , w6757 , w6758 , w6759 , w6760 , w6761 , w6762 , w6763 , w6764 , w6765 , w6766 , w6767 , w6768 , w6769 , w6770 , w6771 , w6772 , w6773 , w6774 , w6775 , w6776 , w6777 , w6778 , w6779 , w6780 , w6781 , w6782 , w6783 , w6784 , w6785 , w6786 , w6787 , w6788 , w6789 , w6790 , w6791 , w6792 , w6793 , w6794 , w6795 , w6796 , w6797 , w6798 , w6799 , w6800 , w6801 , w6802 , w6803 , w6804 , w6805 , w6806 , w6807 , w6808 , w6809 , w6810 , w6811 , w6812 , w6813 , w6814 , w6815 , w6816 , w6817 , w6818 , w6819 , w6820 , w6821 , w6822 , w6823 , w6824 , w6825 , w6826 , w6827 , w6828 , w6829 , w6830 , w6831 , w6832 , w6833 , w6834 , w6835 , w6836 , w6837 , w6838 , w6839 , w6840 , w6841 , w6842 , w6843 , w6844 , w6845 , w6846 , w6847 , w6848 , w6849 , w6850 , w6851 , w6852 , w6853 , w6854 , w6855 , w6856 , w6857 , w6858 , w6859 , w6860 , w6861 , w6862 , w6863 , w6864 , w6865 , w6866 , w6867 , w6868 , w6869 , w6870 , w6871 , w6872 , w6873 , w6874 , w6875 , w6876 , w6877 , w6878 , w6879 , w6880 , w6881 , w6882 , w6883 , w6884 , w6885 , w6886 , w6887 , w6888 , w6889 , w6890 , w6891 , w6892 , w6893 , w6894 , w6895 , w6896 , w6897 , w6898 , w6899 , w6900 , w6901 , w6902 , w6903 , w6904 , w6905 , w6906 , w6907 , w6908 , w6909 , w6910 , w6911 , w6912 , w6913 , w6914 , w6915 , w6916 , w6917 , w6918 , w6919 , w6920 , w6921 , w6922 , w6923 , w6924 , w6925 , w6926 , w6927 , w6928 , w6929 , w6930 , w6931 , w6932 , w6933 , w6934 , w6935 , w6936 , w6937 , w6938 , w6939 , w6940 , w6941 , w6942 , w6943 , w6944 , w6945 , w6946 , w6947 , w6948 , w6949 , w6950 , w6951 , w6952 , w6953 , w6954 , w6955 , w6956 , w6957 , w6958 , w6959 , w6960 , w6961 , w6962 , w6963 , w6964 , w6965 , w6966 , w6967 , w6968 , w6969 , w6970 , w6971 , w6972 , w6973 , w6974 , w6975 , w6976 , w6977 , w6978 , w6979 , w6980 , w6981 , w6982 , w6983 , w6984 , w6985 , w6986 , w6987 , w6988 , w6989 , w6990 , w6991 , w6992 , w6993 , w6994 , w6995 , w6996 , w6997 , w6998 , w6999 , w7000 , w7001 , w7002 , w7003 , w7004 , w7005 , w7006 , w7007 , w7008 , w7009 , w7010 , w7011 , w7012 , w7013 , w7014 , w7015 , w7016 , w7017 , w7018 , w7019 , w7020 , w7021 , w7022 , w7023 , w7024 , w7025 , w7026 , w7027 , w7028 , w7029 , w7030 , w7031 , w7032 , w7033 , w7034 , w7035 , w7036 , w7037 , w7038 , w7039 , w7040 , w7041 , w7042 , w7043 , w7044 , w7045 , w7046 , w7047 , w7048 , w7049 , w7050 , w7051 , w7052 , w7053 , w7054 , w7055 , w7056 , w7057 , w7058 , w7059 , w7060 , w7061 , w7062 , w7063 , w7064 , w7065 , w7066 , w7067 , w7068 , w7069 , w7070 , w7071 , w7072 , w7073 , w7074 , w7075 , w7076 , w7077 , w7078 , w7079 , w7080 , w7081 , w7082 , w7083 , w7084 , w7085 , w7086 , w7087 , w7088 , w7089 , w7090 , w7091 , w7092 , w7093 , w7094 , w7095 , w7096 , w7097 , w7098 , w7099 , w7100 , w7101 , w7102 , w7103 , w7104 , w7105 , w7106 , w7107 , w7108 , w7109 , w7110 , w7111 , w7112 , w7113 , w7114 , w7115 , w7116 , w7117 , w7118 , w7119 , w7120 , w7121 , w7122 , w7123 , w7124 , w7125 , w7126 , w7127 , w7128 , w7129 , w7130 , w7131 , w7132 , w7133 , w7134 , w7135 , w7136 , w7137 , w7138 , w7139 , w7140 , w7141 , w7142 , w7143 , w7144 , w7145 , w7146 , w7147 , w7148 , w7149 , w7150 , w7151 , w7152 , w7153 , w7154 , w7155 , w7156 , w7157 , w7158 , w7159 , w7160 , w7161 , w7162 , w7163 , w7164 , w7165 , w7166 , w7167 , w7168 , w7169 , w7170 , w7171 , w7172 , w7173 , w7174 , w7175 , w7176 , w7177 , w7178 , w7179 , w7180 , w7181 , w7182 , w7183 , w7184 , w7185 , w7186 , w7187 , w7188 , w7189 , w7190 , w7191 , w7192 , w7193 , w7194 , w7195 , w7196 , w7197 , w7198 , w7199 , w7200 , w7201 , w7202 , w7203 , w7204 , w7205 , w7206 , w7207 , w7208 , w7209 , w7210 , w7211 , w7212 , w7213 , w7214 , w7215 , w7216 , w7217 , w7218 , w7219 , w7220 , w7221 , w7222 , w7223 , w7224 , w7225 , w7226 , w7227 , w7228 , w7229 , w7230 , w7231 , w7232 , w7233 , w7234 , w7235 , w7236 , w7237 , w7238 , w7239 , w7240 , w7241 , w7242 , w7243 , w7244 , w7245 , w7246 , w7247 , w7248 , w7249 , w7250 , w7251 , w7252 , w7253 , w7254 , w7255 , w7256 , w7257 , w7258 , w7259 , w7260 , w7261 , w7262 , w7263 , w7264 , w7265 , w7266 , w7267 , w7268 , w7269 , w7270 , w7271 , w7272 , w7273 , w7274 , w7275 , w7276 , w7277 , w7278 , w7279 , w7280 , w7281 , w7282 , w7283 , w7284 , w7285 , w7286 , w7287 , w7288 , w7289 , w7290 , w7291 , w7292 , w7293 , w7294 , w7295 , w7296 , w7297 , w7298 , w7299 , w7300 , w7301 , w7302 , w7303 , w7304 , w7305 , w7306 , w7307 , w7308 , w7309 , w7310 , w7311 , w7312 , w7313 , w7314 , w7315 , w7316 , w7317 , w7318 , w7319 , w7320 , w7321 , w7322 , w7323 , w7324 , w7325 , w7326 , w7327 , w7328 , w7329 , w7330 , w7331 , w7332 , w7333 , w7334 , w7335 , w7336 , w7337 , w7338 , w7339 , w7340 , w7341 , w7342 , w7343 , w7344 , w7345 , w7346 , w7347 , w7348 , w7349 , w7350 , w7351 , w7352 , w7353 , w7354 , w7355 , w7356 , w7357 , w7358 , w7359 , w7360 , w7361 , w7362 , w7363 , w7364 , w7365 , w7366 , w7367 , w7368 , w7369 , w7370 , w7371 , w7372 , w7373 , w7374 , w7375 , w7376 , w7377 , w7378 , w7379 , w7380 , w7381 , w7382 , w7383 , w7384 , w7385 , w7386 , w7387 , w7388 , w7389 , w7390 , w7391 , w7392 , w7393 , w7394 , w7395 , w7396 , w7397 , w7398 , w7399 , w7400 , w7401 , w7402 , w7403 , w7404 , w7405 , w7406 , w7407 , w7408 , w7409 , w7410 , w7411 , w7412 , w7413 , w7414 , w7415 , w7416 , w7417 , w7418 , w7419 , w7420 , w7421 , w7422 , w7423 , w7424 , w7425 , w7426 , w7427 , w7428 , w7429 , w7430 , w7431 , w7432 , w7433 , w7434 , w7435 , w7436 , w7437 , w7438 , w7439 , w7440 , w7441 , w7442 , w7443 , w7444 , w7445 , w7446 , w7447 , w7448 , w7449 , w7450 , w7451 , w7452 , w7453 , w7454 , w7455 , w7456 , w7457 , w7458 , w7459 , w7460 , w7461 , w7462 , w7463 , w7464 , w7465 , w7466 , w7467 , w7468 , w7469 , w7470 , w7471 , w7472 , w7473 , w7474 , w7475 , w7476 , w7477 , w7478 , w7479 , w7480 , w7481 , w7482 , w7483 , w7484 , w7485 , w7486 , w7487 , w7488 , w7489 , w7490 , w7491 , w7492 , w7493 , w7494 , w7495 , w7496 , w7497 , w7498 , w7499 , w7500 , w7501 , w7502 , w7503 , w7504 , w7505 , w7506 , w7507 , w7508 , w7509 , w7510 , w7511 , w7512 , w7513 , w7514 , w7515 , w7516 , w7517 , w7518 , w7519 , w7520 , w7521 , w7522 , w7523 , w7524 , w7525 , w7526 , w7527 , w7528 , w7529 , w7530 , w7531 , w7532 , w7533 , w7534 , w7535 , w7536 , w7537 , w7538 , w7539 , w7540 , w7541 , w7542 , w7543 , w7544 , w7545 , w7546 , w7547 , w7548 , w7549 , w7550 , w7551 , w7552 , w7553 , w7554 , w7555 , w7556 , w7557 , w7558 , w7559 , w7560 , w7561 , w7562 , w7563 , w7564 , w7565 , w7566 , w7567 , w7568 , w7569 , w7570 , w7571 , w7572 , w7573 , w7574 , w7575 , w7576 , w7577 , w7578 , w7579 , w7580 , w7581 , w7582 , w7583 , w7584 , w7585 , w7586 , w7587 , w7588 , w7589 , w7590 , w7591 , w7592 , w7593 , w7594 , w7595 , w7596 , w7597 , w7598 , w7599 , w7600 , w7601 , w7602 , w7603 , w7604 , w7605 , w7606 , w7607 , w7608 , w7609 , w7610 , w7611 , w7612 , w7613 , w7614 , w7615 , w7616 , w7617 , w7618 , w7619 , w7620 , w7621 , w7622 , w7623 , w7624 , w7625 , w7626 , w7627 , w7628 , w7629 , w7630 , w7631 , w7632 , w7633 , w7634 , w7635 , w7636 , w7637 , w7638 , w7639 , w7640 , w7641 , w7642 , w7643 , w7644 , w7645 , w7646 , w7647 , w7648 , w7649 , w7650 , w7651 , w7652 , w7653 , w7654 , w7655 , w7656 , w7657 , w7658 , w7659 , w7660 , w7661 , w7662 , w7663 , w7664 , w7665 , w7666 , w7667 , w7668 , w7669 , w7670 , w7671 , w7672 , w7673 , w7674 , w7675 , w7676 , w7677 , w7678 , w7679 , w7680 , w7681 , w7682 , w7683 , w7684 , w7685 , w7686 , w7687 , w7688 , w7689 , w7690 , w7691 , w7692 , w7693 , w7694 , w7695 , w7696 , w7697 , w7698 , w7699 , w7700 , w7701 , w7702 , w7703 , w7704 , w7705 , w7706 , w7707 , w7708 , w7709 , w7710 , w7711 , w7712 , w7713 , w7714 , w7715 , w7716 , w7717 , w7718 , w7719 , w7720 , w7721 , w7722 , w7723 , w7724 , w7725 , w7726 , w7727 , w7728 , w7729 , w7730 , w7731 , w7732 , w7733 , w7734 , w7735 , w7736 , w7737 , w7738 , w7739 , w7740 , w7741 , w7742 , w7743 , w7744 , w7745 , w7746 , w7747 , w7748 , w7749 , w7750 , w7751 , w7752 , w7753 , w7754 , w7755 , w7756 , w7757 , w7758 , w7759 , w7760 , w7761 , w7762 , w7763 , w7764 , w7765 , w7766 , w7767 , w7768 , w7769 , w7770 , w7771 , w7772 , w7773 , w7774 , w7775 , w7776 , w7777 , w7778 , w7779 , w7780 , w7781 , w7782 , w7783 , w7784 , w7785 , w7786 , w7787 , w7788 , w7789 , w7790 , w7791 , w7792 , w7793 , w7794 , w7795 , w7796 , w7797 , w7798 , w7799 , w7800 , w7801 , w7802 , w7803 , w7804 , w7805 , w7806 , w7807 , w7808 , w7809 , w7810 , w7811 , w7812 , w7813 , w7814 , w7815 , w7816 , w7817 , w7818 , w7819 , w7820 , w7821 , w7822 , w7823 , w7824 , w7825 , w7826 , w7827 , w7828 , w7829 , w7830 , w7831 , w7832 , w7833 , w7834 , w7835 , w7836 , w7837 , w7838 , w7839 , w7840 , w7841 , w7842 , w7843 , w7844 , w7845 , w7846 , w7847 , w7848 , w7849 , w7850 , w7851 , w7852 , w7853 , w7854 , w7855 , w7856 , w7857 , w7858 , w7859 , w7860 , w7861 , w7862 , w7863 , w7864 , w7865 , w7866 , w7867 , w7868 , w7869 , w7870 , w7871 , w7872 , w7873 , w7874 , w7875 , w7876 , w7877 , w7878 , w7879 , w7880 , w7881 , w7882 , w7883 , w7884 , w7885 , w7886 , w7887 , w7888 , w7889 , w7890 , w7891 , w7892 , w7893 , w7894 , w7895 , w7896 , w7897 , w7898 , w7899 , w7900 , w7901 , w7902 , w7903 , w7904 , w7905 , w7906 , w7907 , w7908 , w7909 , w7910 , w7911 , w7912 , w7913 , w7914 , w7915 , w7916 , w7917 , w7918 , w7919 , w7920 , w7921 , w7922 , w7923 , w7924 , w7925 , w7926 , w7927 , w7928 , w7929 , w7930 , w7931 , w7932 , w7933 , w7934 , w7935 , w7936 , w7937 , w7938 , w7939 , w7940 , w7941 , w7942 , w7943 , w7944 , w7945 , w7946 , w7947 , w7948 , w7949 , w7950 , w7951 , w7952 , w7953 , w7954 , w7955 , w7956 , w7957 , w7958 , w7959 , w7960 , w7961 , w7962 , w7963 , w7964 , w7965 , w7966 , w7967 , w7968 , w7969 , w7970 , w7971 , w7972 , w7973 , w7974 , w7975 , w7976 , w7977 , w7978 , w7979 , w7980 , w7981 , w7982 , w7983 , w7984 , w7985 , w7986 , w7987 , w7988 , w7989 , w7990 , w7991 , w7992 , w7993 , w7994 , w7995 , w7996 , w7997 , w7998 , w7999 , w8000 , w8001 , w8002 , w8003 , w8004 , w8005 , w8006 , w8007 , w8008 , w8009 , w8010 , w8011 , w8012 , w8013 , w8014 , w8015 , w8016 , w8017 , w8018 , w8019 , w8020 , w8021 , w8022 , w8023 , w8024 , w8025 , w8026 , w8027 , w8028 , w8029 , w8030 , w8031 , w8032 , w8033 , w8034 , w8035 , w8036 , w8037 , w8038 , w8039 , w8040 , w8041 , w8042 , w8043 , w8044 , w8045 , w8046 , w8047 , w8048 , w8049 , w8050 , w8051 , w8052 , w8053 , w8054 , w8055 , w8056 , w8057 , w8058 , w8059 , w8060 , w8061 , w8062 , w8063 , w8064 , w8065 , w8066 , w8067 , w8068 , w8069 , w8070 , w8071 , w8072 , w8073 , w8074 , w8075 , w8076 , w8077 , w8078 , w8079 , w8080 , w8081 , w8082 , w8083 , w8084 , w8085 , w8086 , w8087 , w8088 , w8089 , w8090 , w8091 , w8092 , w8093 , w8094 , w8095 , w8096 , w8097 , w8098 , w8099 , w8100 , w8101 , w8102 , w8103 , w8104 , w8105 , w8106 , w8107 , w8108 , w8109 , w8110 , w8111 , w8112 , w8113 , w8114 , w8115 , w8116 , w8117 , w8118 , w8119 , w8120 , w8121 , w8122 , w8123 , w8124 , w8125 , w8126 , w8127 , w8128 , w8129 , w8130 , w8131 , w8132 , w8133 , w8134 , w8135 , w8136 , w8137 , w8138 , w8139 , w8140 , w8141 , w8142 , w8143 , w8144 , w8145 , w8146 , w8147 , w8148 , w8149 , w8150 , w8151 , w8152 , w8153 , w8154 , w8155 , w8156 , w8157 , w8158 , w8159 , w8160 , w8161 , w8162 , w8163 , w8164 , w8165 , w8166 , w8167 , w8168 , w8169 , w8170 , w8171 , w8172 , w8173 , w8174 , w8175 , w8176 , w8177 , w8178 , w8179 , w8180 , w8181 , w8182 , w8183 , w8184 , w8185 , w8186 , w8187 , w8188 , w8189 , w8190 , w8191 , w8192 , w8193 , w8194 , w8195 , w8196 , w8197 , w8198 , w8199 , w8200 , w8201 , w8202 , w8203 , w8204 , w8205 , w8206 , w8207 , w8208 , w8209 , w8210 , w8211 , w8212 , w8213 , w8214 , w8215 , w8216 , w8217 , w8218 , w8219 , w8220 , w8221 , w8222 , w8223 , w8224 , w8225 , w8226 , w8227 , w8228 , w8229 , w8230 , w8231 , w8232 , w8233 , w8234 , w8235 , w8236 , w8237 , w8238 , w8239 , w8240 , w8241 , w8242 , w8243 , w8244 , w8245 , w8246 , w8247 , w8248 , w8249 , w8250 , w8251 , w8252 , w8253 , w8254 , w8255 , w8256 , w8257 , w8258 , w8259 , w8260 , w8261 , w8262 , w8263 , w8264 , w8265 , w8266 , w8267 , w8268 , w8269 , w8270 , w8271 , w8272 , w8273 , w8274 , w8275 , w8276 , w8277 , w8278 , w8279 , w8280 , w8281 , w8282 , w8283 , w8284 , w8285 , w8286 , w8287 , w8288 , w8289 , w8290 , w8291 , w8292 , w8293 , w8294 , w8295 , w8296 , w8297 , w8298 , w8299 , w8300 , w8301 , w8302 , w8303 , w8304 , w8305 , w8306 , w8307 , w8308 , w8309 , w8310 , w8311 , w8312 , w8313 , w8314 , w8315 , w8316 , w8317 , w8318 , w8319 , w8320 , w8321 , w8322 , w8323 , w8324 , w8325 , w8326 , w8327 , w8328 , w8329 , w8330 , w8331 , w8332 , w8333 , w8334 , w8335 , w8336 , w8337 , w8338 , w8339 , w8340 , w8341 , w8342 , w8343 , w8344 , w8345 , w8346 , w8347 , w8348 , w8349 , w8350 , w8351 , w8352 , w8353 , w8354 , w8355 , w8356 , w8357 , w8358 , w8359 , w8360 , w8361 , w8362 , w8363 , w8364 , w8365 , w8366 , w8367 , w8368 , w8369 , w8370 , w8371 , w8372 , w8373 , w8374 , w8375 , w8376 , w8377 , w8378 , w8379 , w8380 , w8381 , w8382 , w8383 , w8384 , w8385 , w8386 , w8387 , w8388 , w8389 , w8390 , w8391 , w8392 , w8393 , w8394 , w8395 , w8396 , w8397 , w8398 , w8399 , w8400 , w8401 , w8402 , w8403 , w8404 , w8405 , w8406 , w8407 , w8408 , w8409 , w8410 , w8411 , w8412 , w8413 , w8414 , w8415 , w8416 , w8417 , w8418 , w8419 , w8420 , w8421 , w8422 , w8423 , w8424 , w8425 , w8426 , w8427 , w8428 , w8429 , w8430 , w8431 , w8432 , w8433 , w8434 , w8435 , w8436 , w8437 , w8438 , w8439 , w8440 , w8441 , w8442 , w8443 , w8444 , w8445 , w8446 , w8447 , w8448 , w8449 , w8450 , w8451 , w8452 , w8453 , w8454 , w8455 , w8456 , w8457 , w8458 , w8459 , w8460 , w8461 , w8462 , w8463 , w8464 , w8465 , w8466 , w8467 , w8468 , w8469 , w8470 , w8471 , w8472 , w8473 , w8474 , w8475 , w8476 , w8477 , w8478 , w8479 , w8480 , w8481 , w8482 , w8483 , w8484 , w8485 , w8486 , w8487 , w8488 , w8489 , w8490 , w8491 , w8492 , w8493 , w8494 , w8495 , w8496 , w8497 , w8498 , w8499 , w8500 , w8501 , w8502 , w8503 , w8504 , w8505 , w8506 , w8507 , w8508 , w8509 , w8510 , w8511 , w8512 , w8513 , w8514 , w8515 , w8516 , w8517 , w8518 , w8519 , w8520 , w8521 , w8522 , w8523 , w8524 , w8525 , w8526 , w8527 , w8528 , w8529 , w8530 , w8531 , w8532 , w8533 , w8534 , w8535 , w8536 , w8537 , w8538 , w8539 , w8540 , w8541 , w8542 , w8543 , w8544 , w8545 , w8546 , w8547 , w8548 , w8549 , w8550 , w8551 , w8552 , w8553 , w8554 , w8555 , w8556 , w8557 , w8558 , w8559 , w8560 , w8561 , w8562 , w8563 , w8564 , w8565 , w8566 , w8567 , w8568 , w8569 , w8570 , w8571 , w8572 , w8573 , w8574 , w8575 , w8576 , w8577 , w8578 , w8579 , w8580 , w8581 , w8582 , w8583 , w8584 , w8585 , w8586 , w8587 , w8588 , w8589 , w8590 , w8591 , w8592 , w8593 , w8594 , w8595 , w8596 , w8597 , w8598 , w8599 , w8600 , w8601 , w8602 , w8603 , w8604 , w8605 , w8606 , w8607 , w8608 , w8609 , w8610 , w8611 , w8612 , w8613 , w8614 , w8615 , w8616 , w8617 , w8618 , w8619 , w8620 , w8621 , w8622 , w8623 , w8624 , w8625 , w8626 , w8627 , w8628 , w8629 , w8630 , w8631 , w8632 , w8633 , w8634 , w8635 , w8636 , w8637 , w8638 , w8639 , w8640 , w8641 , w8642 , w8643 , w8644 , w8645 , w8646 , w8647 , w8648 , w8649 , w8650 , w8651 , w8652 , w8653 , w8654 , w8655 , w8656 , w8657 , w8658 , w8659 , w8660 , w8661 , w8662 , w8663 , w8664 , w8665 , w8666 , w8667 , w8668 , w8669 , w8670 , w8671 , w8672 , w8673 , w8674 , w8675 , w8676 , w8677 , w8678 , w8679 , w8680 , w8681 , w8682 , w8683 , w8684 , w8685 , w8686 , w8687 , w8688 , w8689 , w8690 , w8691 , w8692 , w8693 , w8694 , w8695 , w8696 , w8697 , w8698 , w8699 , w8700 , w8701 , w8702 , w8703 , w8704 , w8705 , w8706 , w8707 , w8708 , w8709 , w8710 , w8711 , w8712 , w8713 , w8714 , w8715 , w8716 , w8717 , w8718 , w8719 , w8720 , w8721 , w8722 , w8723 , w8724 , w8725 , w8726 , w8727 , w8728 , w8729 , w8730 , w8731 , w8732 , w8733 , w8734 , w8735 , w8736 , w8737 , w8738 , w8739 , w8740 , w8741 , w8742 , w8743 , w8744 , w8745 , w8746 , w8747 , w8748 , w8749 , w8750 , w8751 , w8752 , w8753 , w8754 , w8755 , w8756 , w8757 , w8758 , w8759 , w8760 , w8761 , w8762 , w8763 , w8764 , w8765 , w8766 , w8767 , w8768 , w8769 , w8770 , w8771 , w8772 , w8773 , w8774 , w8775 , w8776 , w8777 , w8778 , w8779 , w8780 , w8781 , w8782 , w8783 , w8784 , w8785 , w8786 , w8787 , w8788 , w8789 , w8790 , w8791 , w8792 , w8793 , w8794 , w8795 , w8796 , w8797 , w8798 , w8799 , w8800 , w8801 , w8802 , w8803 , w8804 , w8805 , w8806 , w8807 , w8808 , w8809 , w8810 , w8811 , w8812 , w8813 , w8814 , w8815 , w8816 , w8817 , w8818 , w8819 , w8820 , w8821 , w8822 , w8823 , w8824 , w8825 , w8826 , w8827 , w8828 , w8829 , w8830 , w8831 , w8832 , w8833 , w8834 , w8835 , w8836 , w8837 , w8838 , w8839 , w8840 , w8841 , w8842 , w8843 , w8844 , w8845 , w8846 , w8847 , w8848 , w8849 , w8850 , w8851 , w8852 , w8853 , w8854 , w8855 , w8856 , w8857 , w8858 , w8859 , w8860 , w8861 , w8862 , w8863 , w8864 , w8865 , w8866 , w8867 , w8868 , w8869 , w8870 , w8871 , w8872 , w8873 , w8874 , w8875 , w8876 , w8877 , w8878 , w8879 , w8880 , w8881 , w8882 , w8883 , w8884 , w8885 , w8886 , w8887 , w8888 , w8889 , w8890 , w8891 , w8892 , w8893 , w8894 , w8895 , w8896 , w8897 , w8898 , w8899 , w8900 , w8901 , w8902 , w8903 , w8904 , w8905 , w8906 , w8907 , w8908 , w8909 , w8910 , w8911 , w8912 , w8913 , w8914 , w8915 , w8916 , w8917 , w8918 , w8919 , w8920 , w8921 , w8922 , w8923 , w8924 , w8925 , w8926 , w8927 , w8928 , w8929 , w8930 , w8931 , w8932 , w8933 , w8934 , w8935 , w8936 , w8937 , w8938 , w8939 , w8940 , w8941 , w8942 , w8943 , w8944 , w8945 , w8946 , w8947 , w8948 , w8949 , w8950 , w8951 , w8952 , w8953 , w8954 , w8955 , w8956 , w8957 , w8958 , w8959 , w8960 , w8961 , w8962 , w8963 , w8964 , w8965 , w8966 , w8967 , w8968 , w8969 , w8970 , w8971 , w8972 , w8973 , w8974 , w8975 , w8976 , w8977 , w8978 , w8979 , w8980 , w8981 , w8982 , w8983 , w8984 , w8985 , w8986 , w8987 , w8988 , w8989 , w8990 , w8991 , w8992 , w8993 , w8994 , w8995 , w8996 , w8997 , w8998 , w8999 , w9000 , w9001 , w9002 , w9003 , w9004 , w9005 , w9006 , w9007 , w9008 , w9009 , w9010 , w9011 , w9012 , w9013 , w9014 , w9015 , w9016 , w9017 , w9018 , w9019 , w9020 , w9021 , w9022 , w9023 , w9024 , w9025 , w9026 , w9027 , w9028 , w9029 , w9030 , w9031 , w9032 , w9033 , w9034 , w9035 , w9036 , w9037 , w9038 , w9039 , w9040 , w9041 , w9042 , w9043 , w9044 , w9045 , w9046 , w9047 , w9048 , w9049 , w9050 , w9051 , w9052 , w9053 , w9054 , w9055 , w9056 , w9057 , w9058 , w9059 , w9060 , w9061 , w9062 , w9063 , w9064 , w9065 , w9066 , w9067 , w9068 , w9069 , w9070 , w9071 , w9072 , w9073 , w9074 , w9075 , w9076 , w9077 , w9078 , w9079 , w9080 , w9081 , w9082 , w9083 , w9084 , w9085 , w9086 , w9087 , w9088 , w9089 , w9090 , w9091 , w9092 , w9093 , w9094 , w9095 , w9096 , w9097 , w9098 , w9099 , w9100 , w9101 , w9102 , w9103 , w9104 , w9105 , w9106 , w9107 , w9108 , w9109 , w9110 , w9111 , w9112 , w9113 , w9114 , w9115 , w9116 , w9117 , w9118 , w9119 , w9120 , w9121 , w9122 , w9123 , w9124 , w9125 , w9126 , w9127 , w9128 , w9129 , w9130 , w9131 , w9132 , w9133 , w9134 , w9135 , w9136 , w9137 , w9138 , w9139 , w9140 , w9141 , w9142 , w9143 , w9144 , w9145 , w9146 , w9147 , w9148 , w9149 , w9150 , w9151 , w9152 , w9153 , w9154 , w9155 , w9156 , w9157 , w9158 , w9159 , w9160 , w9161 , w9162 , w9163 , w9164 , w9165 , w9166 , w9167 , w9168 , w9169 , w9170 , w9171 , w9172 , w9173 , w9174 , w9175 , w9176 , w9177 , w9178 , w9179 , w9180 , w9181 , w9182 , w9183 , w9184 , w9185 , w9186 , w9187 , w9188 , w9189 , w9190 , w9191 , w9192 , w9193 , w9194 , w9195 , w9196 , w9197 , w9198 , w9199 , w9200 , w9201 , w9202 , w9203 , w9204 , w9205 , w9206 , w9207 , w9208 , w9209 , w9210 , w9211 , w9212 , w9213 , w9214 , w9215 , w9216 , w9217 , w9218 , w9219 , w9220 , w9221 , w9222 , w9223 , w9224 , w9225 , w9226 , w9227 , w9228 , w9229 , w9230 , w9231 , w9232 , w9233 , w9234 , w9235 , w9236 , w9237 , w9238 , w9239 , w9240 , w9241 , w9242 , w9243 , w9244 , w9245 , w9246 , w9247 , w9248 , w9249 , w9250 , w9251 , w9252 , w9253 , w9254 , w9255 , w9256 , w9257 , w9258 , w9259 , w9260 , w9261 , w9262 , w9263 , w9264 , w9265 , w9266 , w9267 , w9268 , w9269 , w9270 , w9271 , w9272 , w9273 , w9274 , w9275 , w9276 , w9277 , w9278 , w9279 , w9280 , w9281 , w9282 , w9283 , w9284 , w9285 , w9286 , w9287 , w9288 , w9289 , w9290 , w9291 , w9292 , w9293 , w9294 , w9295 , w9296 , w9297 , w9298 , w9299 , w9300 , w9301 , w9302 , w9303 , w9304 , w9305 , w9306 , w9307 , w9308 , w9309 , w9310 , w9311 , w9312 , w9313 , w9314 , w9315 , w9316 , w9317 , w9318 , w9319 , w9320 , w9321 , w9322 , w9323 , w9324 , w9325 , w9326 , w9327 , w9328 , w9329 , w9330 , w9331 , w9332 , w9333 , w9334 , w9335 , w9336 , w9337 , w9338 , w9339 , w9340 , w9341 , w9342 , w9343 , w9344 , w9345 , w9346 , w9347 , w9348 , w9349 , w9350 , w9351 , w9352 , w9353 , w9354 , w9355 , w9356 , w9357 , w9358 , w9359 , w9360 , w9361 , w9362 , w9363 , w9364 , w9365 , w9366 , w9367 , w9368 , w9369 , w9370 , w9371 , w9372 , w9373 , w9374 , w9375 , w9376 , w9377 , w9378 , w9379 , w9380 , w9381 , w9382 , w9383 , w9384 , w9385 , w9386 , w9387 , w9388 , w9389 , w9390 , w9391 , w9392 , w9393 , w9394 , w9395 , w9396 , w9397 , w9398 , w9399 , w9400 , w9401 , w9402 , w9403 , w9404 , w9405 , w9406 , w9407 , w9408 , w9409 , w9410 , w9411 , w9412 , w9413 , w9414 , w9415 , w9416 , w9417 , w9418 , w9419 , w9420 , w9421 , w9422 , w9423 , w9424 , w9425 , w9426 , w9427 , w9428 , w9429 , w9430 , w9431 , w9432 , w9433 , w9434 , w9435 , w9436 , w9437 , w9438 , w9439 , w9440 , w9441 , w9442 , w9443 , w9444 , w9445 , w9446 , w9447 , w9448 , w9449 , w9450 , w9451 , w9452 , w9453 , w9454 , w9455 , w9456 , w9457 , w9458 , w9459 , w9460 , w9461 , w9462 , w9463 , w9464 , w9465 , w9466 , w9467 , w9468 , w9469 , w9470 , w9471 , w9472 , w9473 , w9474 , w9475 , w9476 , w9477 , w9478 , w9479 , w9480 , w9481 , w9482 , w9483 , w9484 , w9485 , w9486 , w9487 , w9488 , w9489 , w9490 , w9491 , w9492 , w9493 , w9494 , w9495 , w9496 , w9497 , w9498 , w9499 , w9500 , w9501 , w9502 , w9503 , w9504 , w9505 , w9506 , w9507 , w9508 , w9509 , w9510 , w9511 , w9512 , w9513 , w9514 , w9515 , w9516 , w9517 , w9518 , w9519 , w9520 , w9521 , w9522 , w9523 , w9524 , w9525 , w9526 , w9527 , w9528 , w9529 , w9530 , w9531 , w9532 , w9533 , w9534 , w9535 , w9536 , w9537 , w9538 , w9539 , w9540 , w9541 , w9542 , w9543 , w9544 , w9545 , w9546 , w9547 , w9548 , w9549 , w9550 , w9551 , w9552 , w9553 , w9554 , w9555 , w9556 , w9557 , w9558 , w9559 , w9560 , w9561 , w9562 , w9563 , w9564 , w9565 , w9566 , w9567 , w9568 , w9569 , w9570 , w9571 , w9572 , w9573 , w9574 , w9575 , w9576 , w9577 , w9578 , w9579 , w9580 , w9581 , w9582 , w9583 , w9584 , w9585 , w9586 , w9587 , w9588 , w9589 , w9590 , w9591 , w9592 , w9593 , w9594 , w9595 , w9596 , w9597 , w9598 , w9599 , w9600 , w9601 , w9602 , w9603 , w9604 , w9605 , w9606 , w9607 , w9608 , w9609 , w9610 , w9611 , w9612 , w9613 , w9614 , w9615 , w9616 , w9617 , w9618 , w9619 , w9620 , w9621 , w9622 , w9623 , w9624 , w9625 , w9626 , w9627 , w9628 , w9629 , w9630 , w9631 , w9632 , w9633 , w9634 , w9635 , w9636 , w9637 , w9638 , w9639 , w9640 , w9641 , w9642 , w9643 , w9644 , w9645 , w9646 , w9647 , w9648 , w9649 , w9650 , w9651 , w9652 , w9653 , w9654 , w9655 , w9656 , w9657 , w9658 , w9659 , w9660 , w9661 , w9662 , w9663 , w9664 , w9665 , w9666 , w9667 , w9668 , w9669 , w9670 , w9671 , w9672 , w9673 , w9674 , w9675 , w9676 , w9677 , w9678 , w9679 , w9680 , w9681 , w9682 , w9683 , w9684 , w9685 , w9686 , w9687 , w9688 , w9689 , w9690 , w9691 , w9692 , w9693 , w9694 , w9695 , w9696 , w9697 , w9698 , w9699 , w9700 , w9701 , w9702 , w9703 , w9704 , w9705 , w9706 , w9707 , w9708 , w9709 , w9710 , w9711 , w9712 , w9713 , w9714 , w9715 , w9716 , w9717 , w9718 , w9719 , w9720 , w9721 , w9722 , w9723 , w9724 , w9725 , w9726 , w9727 , w9728 , w9729 , w9730 , w9731 , w9732 , w9733 , w9734 , w9735 , w9736 , w9737 , w9738 , w9739 , w9740 , w9741 , w9742 , w9743 , w9744 , w9745 , w9746 , w9747 , w9748 , w9749 , w9750 , w9751 , w9752 , w9753 , w9754 , w9755 , w9756 , w9757 , w9758 , w9759 , w9760 , w9761 , w9762 , w9763 , w9764 , w9765 , w9766 , w9767 , w9768 , w9769 , w9770 , w9771 , w9772 , w9773 , w9774 , w9775 , w9776 , w9777 , w9778 , w9779 , w9780 , w9781 , w9782 , w9783 , w9784 , w9785 , w9786 , w9787 , w9788 , w9789 , w9790 , w9791 , w9792 , w9793 , w9794 , w9795 , w9796 , w9797 , w9798 , w9799 , w9800 , w9801 , w9802 , w9803 , w9804 , w9805 , w9806 , w9807 , w9808 , w9809 , w9810 , w9811 , w9812 , w9813 , w9814 , w9815 , w9816 , w9817 , w9818 , w9819 , w9820 , w9821 , w9822 , w9823 , w9824 , w9825 , w9826 , w9827 , w9828 , w9829 , w9830 , w9831 , w9832 , w9833 , w9834 , w9835 , w9836 , w9837 , w9838 , w9839 , w9840 , w9841 , w9842 , w9843 , w9844 , w9845 , w9846 , w9847 , w9848 , w9849 , w9850 , w9851 , w9852 , w9853 , w9854 , w9855 , w9856 , w9857 , w9858 , w9859 , w9860 , w9861 , w9862 , w9863 , w9864 , w9865 , w9866 , w9867 , w9868 , w9869 , w9870 , w9871 , w9872 , w9873 , w9874 , w9875 , w9876 , w9877 , w9878 , w9879 , w9880 , w9881 , w9882 , w9883 , w9884 , w9885 , w9886 , w9887 , w9888 , w9889 , w9890 , w9891 , w9892 , w9893 , w9894 , w9895 , w9896 , w9897 , w9898 , w9899 , w9900 , w9901 , w9902 , w9903 , w9904 , w9905 , w9906 , w9907 , w9908 , w9909 , w9910 , w9911 , w9912 , w9913 , w9914 , w9915 , w9916 , w9917 , w9918 , w9919 , w9920 , w9921 , w9922 , w9923 , w9924 , w9925 , w9926 , w9927 , w9928 , w9929 , w9930 , w9931 , w9932 , w9933 , w9934 , w9935 , w9936 , w9937 , w9938 , w9939 , w9940 , w9941 , w9942 , w9943 , w9944 , w9945 , w9946 , w9947 , w9948 , w9949 , w9950 , w9951 , w9952 , w9953 , w9954 , w9955 , w9956 , w9957 , w9958 , w9959 , w9960 , w9961 , w9962 , w9963 , w9964 , w9965 , w9966 , w9967 , w9968 , w9969 , w9970 , w9971 , w9972 , w9973 , w9974 , w9975 , w9976 , w9977 , w9978 , w9979 , w9980 , w9981 , w9982 , w9983 , w9984 , w9985 , w9986 , w9987 , w9988 , w9989 , w9990 , w9991 , w9992 , w9993 , w9994 , w9995 , w9996 , w9997 , w9998 , w9999 , w10000 , w10001 , w10002 , w10003 , w10004 , w10005 , w10006 , w10007 , w10008 , w10009 , w10010 , w10011 , w10012 , w10013 , w10014 , w10015 , w10016 , w10017 , w10018 , w10019 , w10020 , w10021 , w10022 , w10023 , w10024 , w10025 , w10026 , w10027 , w10028 , w10029 , w10030 , w10031 , w10032 , w10033 , w10034 , w10035 , w10036 , w10037 , w10038 , w10039 , w10040 , w10041 , w10042 , w10043 , w10044 , w10045 , w10046 , w10047 , w10048 , w10049 , w10050 , w10051 , w10052 , w10053 , w10054 , w10055 , w10056 , w10057 , w10058 , w10059 , w10060 , w10061 , w10062 , w10063 , w10064 , w10065 , w10066 , w10067 , w10068 , w10069 , w10070 , w10071 , w10072 , w10073 , w10074 , w10075 , w10076 , w10077 , w10078 , w10079 , w10080 , w10081 , w10082 , w10083 , w10084 , w10085 , w10086 , w10087 , w10088 , w10089 , w10090 , w10091 , w10092 , w10093 , w10094 , w10095 , w10096 , w10097 , w10098 , w10099 , w10100 , w10101 , w10102 , w10103 , w10104 , w10105 , w10106 , w10107 , w10108 , w10109 , w10110 , w10111 , w10112 , w10113 , w10114 , w10115 , w10116 , w10117 , w10118 , w10119 , w10120 , w10121 , w10122 , w10123 , w10124 , w10125 , w10126 , w10127 , w10128 , w10129 , w10130 , w10131 , w10132 , w10133 , w10134 , w10135 , w10136 , w10137 , w10138 , w10139 , w10140 , w10141 , w10142 , w10143 , w10144 , w10145 , w10146 , w10147 , w10148 , w10149 , w10150 , w10151 , w10152 , w10153 , w10154 , w10155 , w10156 , w10157 , w10158 , w10159 , w10160 , w10161 , w10162 , w10163 , w10164 , w10165 , w10166 , w10167 , w10168 , w10169 , w10170 , w10171 , w10172 , w10173 , w10174 , w10175 , w10176 , w10177 , w10178 , w10179 , w10180 , w10181 , w10182 , w10183 , w10184 , w10185 , w10186 , w10187 , w10188 , w10189 , w10190 , w10191 , w10192 , w10193 , w10194 , w10195 , w10196 , w10197 , w10198 , w10199 , w10200 , w10201 , w10202 , w10203 , w10204 , w10205 , w10206 , w10207 , w10208 , w10209 , w10210 , w10211 , w10212 , w10213 , w10214 , w10215 , w10216 , w10217 , w10218 , w10219 , w10220 , w10221 , w10222 , w10223 , w10224 , w10225 , w10226 , w10227 , w10228 , w10229 , w10230 , w10231 , w10232 , w10233 , w10234 , w10235 , w10236 , w10237 , w10238 , w10239 , w10240 , w10241 , w10242 , w10243 , w10244 , w10245 , w10246 , w10247 , w10248 , w10249 , w10250 , w10251 , w10252 , w10253 , w10254 , w10255 , w10256 , w10257 , w10258 , w10259 , w10260 , w10261 , w10262 , w10263 , w10264 , w10265 , w10266 , w10267 , w10268 , w10269 , w10270 , w10271 , w10272 , w10273 , w10274 , w10275 , w10276 , w10277 , w10278 , w10279 , w10280 , w10281 , w10282 , w10283 , w10284 , w10285 , w10286 , w10287 , w10288 , w10289 , w10290 , w10291 , w10292 , w10293 , w10294 , w10295 , w10296 , w10297 , w10298 , w10299 , w10300 , w10301 , w10302 , w10303 , w10304 , w10305 , w10306 , w10307 , w10308 , w10309 , w10310 , w10311 , w10312 , w10313 , w10314 , w10315 , w10316 , w10317 , w10318 , w10319 , w10320 , w10321 , w10322 , w10323 , w10324 , w10325 , w10326 , w10327 , w10328 , w10329 , w10330 , w10331 , w10332 , w10333 , w10334 , w10335 , w10336 , w10337 , w10338 , w10339 , w10340 , w10341 , w10342 , w10343 , w10344 , w10345 , w10346 , w10347 , w10348 , w10349 , w10350 , w10351 , w10352 , w10353 , w10354 , w10355 , w10356 , w10357 , w10358 , w10359 , w10360 , w10361 , w10362 , w10363 , w10364 , w10365 , w10366 , w10367 , w10368 , w10369 , w10370 , w10371 , w10372 , w10373 , w10374 , w10375 , w10376 , w10377 , w10378 , w10379 , w10380 , w10381 , w10382 , w10383 , w10384 , w10385 , w10386 , w10387 , w10388 , w10389 , w10390 , w10391 , w10392 , w10393 , w10394 , w10395 , w10396 , w10397 , w10398 , w10399 , w10400 , w10401 , w10402 , w10403 , w10404 , w10405 , w10406 , w10407 , w10408 , w10409 , w10410 , w10411 , w10412 , w10413 , w10414 , w10415 , w10416 , w10417 , w10418 , w10419 , w10420 , w10421 , w10422 , w10423 , w10424 , w10425 , w10426 , w10427 , w10428 , w10429 , w10430 , w10431 , w10432 , w10433 , w10434 , w10435 , w10436 , w10437 , w10438 , w10439 , w10440 , w10441 , w10442 , w10443 , w10444 , w10445 , w10446 , w10447 , w10448 , w10449 , w10450 , w10451 , w10452 , w10453 , w10454 , w10455 , w10456 , w10457 , w10458 , w10459 , w10460 , w10461 , w10462 , w10463 , w10464 , w10465 , w10466 , w10467 , w10468 , w10469 , w10470 , w10471 , w10472 , w10473 , w10474 , w10475 , w10476 , w10477 , w10478 , w10479 , w10480 , w10481 , w10482 , w10483 , w10484 , w10485 , w10486 , w10487 , w10488 , w10489 , w10490 , w10491 , w10492 , w10493 , w10494 , w10495 , w10496 , w10497 , w10498 , w10499 , w10500 , w10501 , w10502 , w10503 , w10504 , w10505 , w10506 , w10507 , w10508 , w10509 , w10510 , w10511 , w10512 , w10513 , w10514 , w10515 , w10516 , w10517 , w10518 , w10519 , w10520 , w10521 , w10522 , w10523 , w10524 , w10525 , w10526 , w10527 , w10528 , w10529 , w10530 , w10531 , w10532 , w10533 , w10534 , w10535 , w10536 , w10537 , w10538 , w10539 , w10540 , w10541 , w10542 , w10543 , w10544 , w10545 , w10546 , w10547 , w10548 , w10549 , w10550 , w10551 , w10552 , w10553 , w10554 , w10555 , w10556 , w10557 , w10558 , w10559 , w10560 , w10561 , w10562 , w10563 , w10564 , w10565 , w10566 , w10567 , w10568 , w10569 , w10570 , w10571 , w10572 , w10573 , w10574 , w10575 , w10576 , w10577 , w10578 , w10579 , w10580 , w10581 , w10582 , w10583 , w10584 , w10585 , w10586 , w10587 , w10588 , w10589 , w10590 , w10591 , w10592 , w10593 , w10594 , w10595 , w10596 , w10597 , w10598 , w10599 , w10600 , w10601 , w10602 , w10603 , w10604 , w10605 , w10606 , w10607 , w10608 , w10609 , w10610 , w10611 , w10612 , w10613 , w10614 , w10615 , w10616 , w10617 , w10618 , w10619 , w10620 , w10621 , w10622 , w10623 , w10624 , w10625 , w10626 , w10627 , w10628 , w10629 , w10630 , w10631 , w10632 , w10633 , w10634 , w10635 , w10636 , w10637 , w10638 , w10639 , w10640 , w10641 , w10642 , w10643 , w10644 , w10645 , w10646 , w10647 , w10648 , w10649 , w10650 , w10651 , w10652 , w10653 , w10654 , w10655 , w10656 , w10657 , w10658 , w10659 , w10660 , w10661 , w10662 , w10663 , w10664 , w10665 , w10666 , w10667 , w10668 , w10669 , w10670 , w10671 , w10672 , w10673 , w10674 , w10675 , w10676 , w10677 , w10678 , w10679 , w10680 , w10681 , w10682 , w10683 , w10684 , w10685 , w10686 , w10687 , w10688 , w10689 , w10690 , w10691 , w10692 , w10693 , w10694 , w10695 , w10696 , w10697 , w10698 , w10699 , w10700 , w10701 , w10702 , w10703 , w10704 , w10705 , w10706 , w10707 , w10708 , w10709 , w10710 , w10711 , w10712 , w10713 , w10714 , w10715 , w10716 , w10717 , w10718 , w10719 , w10720 , w10721 , w10722 , w10723 , w10724 , w10725 , w10726 , w10727 , w10728 , w10729 , w10730 , w10731 , w10732 , w10733 , w10734 , w10735 , w10736 , w10737 , w10738 , w10739 , w10740 , w10741 , w10742 , w10743 , w10744 , w10745 , w10746 , w10747 , w10748 , w10749 , w10750 , w10751 , w10752 , w10753 , w10754 , w10755 , w10756 , w10757 , w10758 , w10759 , w10760 , w10761 , w10762 , w10763 , w10764 , w10765 , w10766 , w10767 , w10768 , w10769 , w10770 , w10771 , w10772 , w10773 , w10774 , w10775 , w10776 , w10777 , w10778 , w10779 , w10780 , w10781 , w10782 , w10783 , w10784 , w10785 , w10786 , w10787 , w10788 , w10789 , w10790 , w10791 , w10792 , w10793 , w10794 , w10795 , w10796 , w10797 , w10798 , w10799 , w10800 , w10801 , w10802 , w10803 , w10804 , w10805 , w10806 , w10807 , w10808 , w10809 , w10810 , w10811 , w10812 , w10813 , w10814 , w10815 , w10816 , w10817 , w10818 , w10819 , w10820 , w10821 , w10822 , w10823 , w10824 , w10825 , w10826 , w10827 , w10828 , w10829 , w10830 , w10831 , w10832 , w10833 , w10834 , w10835 , w10836 , w10837 , w10838 , w10839 , w10840 , w10841 , w10842 , w10843 , w10844 , w10845 , w10846 , w10847 , w10848 , w10849 , w10850 , w10851 , w10852 , w10853 , w10854 , w10855 , w10856 , w10857 , w10858 , w10859 , w10860 , w10861 , w10862 , w10863 , w10864 , w10865 , w10866 , w10867 , w10868 , w10869 , w10870 , w10871 , w10872 , w10873 , w10874 , w10875 , w10876 , w10877 , w10878 , w10879 , w10880 , w10881 , w10882 , w10883 , w10884 , w10885 , w10886 , w10887 , w10888 , w10889 , w10890 , w10891 , w10892 , w10893 , w10894 , w10895 , w10896 , w10897 , w10898 , w10899 , w10900 , w10901 , w10902 , w10903 , w10904 , w10905 , w10906 , w10907 , w10908 , w10909 , w10910 , w10911 , w10912 , w10913 , w10914 , w10915 , w10916 , w10917 , w10918 , w10919 , w10920 , w10921 , w10922 , w10923 , w10924 , w10925 , w10926 , w10927 , w10928 , w10929 , w10930 , w10931 , w10932 , w10933 , w10934 , w10935 , w10936 , w10937 , w10938 , w10939 , w10940 , w10941 , w10942 , w10943 , w10944 , w10945 , w10946 , w10947 , w10948 , w10949 , w10950 , w10951 , w10952 , w10953 , w10954 , w10955 , w10956 , w10957 , w10958 , w10959 , w10960 , w10961 , w10962 , w10963 , w10964 , w10965 , w10966 , w10967 , w10968 , w10969 , w10970 , w10971 , w10972 , w10973 , w10974 , w10975 , w10976 , w10977 , w10978 , w10979 , w10980 , w10981 , w10982 , w10983 , w10984 , w10985 , w10986 , w10987 , w10988 , w10989 , w10990 , w10991 , w10992 , w10993 , w10994 , w10995 , w10996 , w10997 , w10998 , w10999 , w11000 , w11001 , w11002 , w11003 , w11004 , w11005 , w11006 , w11007 , w11008 , w11009 , w11010 , w11011 , w11012 , w11013 , w11014 , w11015 , w11016 , w11017 , w11018 , w11019 , w11020 , w11021 , w11022 , w11023 , w11024 , w11025 , w11026 , w11027 , w11028 , w11029 , w11030 , w11031 , w11032 , w11033 , w11034 , w11035 , w11036 , w11037 , w11038 , w11039 , w11040 , w11041 , w11042 , w11043 , w11044 , w11045 , w11046 , w11047 , w11048 , w11049 , w11050 , w11051 , w11052 , w11053 , w11054 , w11055 , w11056 , w11057 , w11058 , w11059 , w11060 , w11061 , w11062 , w11063 , w11064 , w11065 , w11066 , w11067 , w11068 , w11069 , w11070 , w11071 , w11072 , w11073 , w11074 , w11075 , w11076 , w11077 , w11078 , w11079 , w11080 , w11081 , w11082 , w11083 , w11084 , w11085 , w11086 , w11087 , w11088 , w11089 , w11090 , w11091 , w11092 , w11093 , w11094 , w11095 , w11096 , w11097 , w11098 , w11099 , w11100 , w11101 , w11102 , w11103 , w11104 , w11105 , w11106 , w11107 , w11108 , w11109 , w11110 , w11111 , w11112 , w11113 , w11114 , w11115 , w11116 , w11117 , w11118 , w11119 , w11120 , w11121 , w11122 , w11123 , w11124 , w11125 , w11126 , w11127 , w11128 , w11129 , w11130 , w11131 , w11132 , w11133 , w11134 , w11135 , w11136 , w11137 , w11138 , w11139 , w11140 , w11141 , w11142 , w11143 , w11144 , w11145 , w11146 , w11147 , w11148 , w11149 , w11150 , w11151 , w11152 , w11153 , w11154 , w11155 , w11156 , w11157 , w11158 , w11159 , w11160 , w11161 , w11162 , w11163 , w11164 , w11165 , w11166 , w11167 , w11168 , w11169 , w11170 , w11171 , w11172 , w11173 , w11174 , w11175 , w11176 , w11177 , w11178 , w11179 , w11180 , w11181 , w11182 , w11183 , w11184 , w11185 , w11186 , w11187 , w11188 , w11189 , w11190 , w11191 , w11192 , w11193 , w11194 , w11195 , w11196 , w11197 , w11198 , w11199 , w11200 , w11201 , w11202 , w11203 , w11204 , w11205 , w11206 , w11207 , w11208 , w11209 , w11210 , w11211 , w11212 , w11213 , w11214 , w11215 , w11216 , w11217 , w11218 , w11219 , w11220 , w11221 , w11222 , w11223 , w11224 , w11225 , w11226 , w11227 , w11228 , w11229 , w11230 , w11231 , w11232 , w11233 , w11234 , w11235 , w11236 , w11237 , w11238 , w11239 , w11240 , w11241 , w11242 , w11243 , w11244 , w11245 , w11246 , w11247 , w11248 , w11249 , w11250 , w11251 , w11252 , w11253 , w11254 , w11255 , w11256 , w11257 , w11258 , w11259 , w11260 , w11261 , w11262 , w11263 , w11264 , w11265 , w11266 , w11267 , w11268 , w11269 , w11270 , w11271 , w11272 , w11273 , w11274 , w11275 , w11276 , w11277 , w11278 , w11279 , w11280 , w11281 , w11282 , w11283 , w11284 , w11285 , w11286 , w11287 , w11288 , w11289 , w11290 , w11291 , w11292 , w11293 , w11294 , w11295 , w11296 , w11297 , w11298 , w11299 , w11300 , w11301 , w11302 , w11303 , w11304 , w11305 , w11306 , w11307 , w11308 , w11309 , w11310 , w11311 , w11312 , w11313 , w11314 , w11315 , w11316 , w11317 , w11318 , w11319 , w11320 , w11321 , w11322 , w11323 , w11324 , w11325 , w11326 , w11327 , w11328 , w11329 , w11330 , w11331 , w11332 , w11333 , w11334 , w11335 , w11336 , w11337 , w11338 , w11339 , w11340 , w11341 , w11342 , w11343 , w11344 , w11345 , w11346 , w11347 , w11348 , w11349 , w11350 , w11351 , w11352 , w11353 , w11354 , w11355 , w11356 , w11357 , w11358 , w11359 , w11360 , w11361 , w11362 , w11363 , w11364 , w11365 , w11366 , w11367 , w11368 , w11369 , w11370 , w11371 , w11372 , w11373 , w11374 , w11375 , w11376 , w11377 , w11378 , w11379 , w11380 , w11381 , w11382 , w11383 , w11384 , w11385 , w11386 , w11387 , w11388 , w11389 , w11390 , w11391 , w11392 , w11393 , w11394 , w11395 , w11396 , w11397 , w11398 , w11399 , w11400 , w11401 , w11402 , w11403 , w11404 , w11405 , w11406 , w11407 , w11408 , w11409 , w11410 , w11411 , w11412 , w11413 , w11414 , w11415 , w11416 , w11417 , w11418 , w11419 , w11420 , w11421 , w11422 , w11423 , w11424 , w11425 , w11426 , w11427 , w11428 , w11429 , w11430 , w11431 , w11432 , w11433 , w11434 , w11435 , w11436 , w11437 , w11438 , w11439 , w11440 , w11441 , w11442 , w11443 , w11444 , w11445 , w11446 , w11447 , w11448 , w11449 , w11450 , w11451 , w11452 , w11453 , w11454 , w11455 , w11456 , w11457 , w11458 , w11459 , w11460 , w11461 , w11462 , w11463 , w11464 , w11465 , w11466 , w11467 , w11468 , w11469 , w11470 , w11471 , w11472 , w11473 , w11474 , w11475 , w11476 , w11477 , w11478 , w11479 , w11480 , w11481 , w11482 , w11483 , w11484 , w11485 , w11486 , w11487 , w11488 , w11489 , w11490 , w11491 , w11492 , w11493 , w11494 , w11495 , w11496 , w11497 , w11498 , w11499 , w11500 , w11501 , w11502 , w11503 , w11504 , w11505 , w11506 , w11507 , w11508 , w11509 , w11510 , w11511 , w11512 , w11513 , w11514 , w11515 , w11516 , w11517 , w11518 , w11519 , w11520 , w11521 , w11522 , w11523 , w11524 , w11525 , w11526 , w11527 , w11528 , w11529 , w11530 , w11531 , w11532 , w11533 , w11534 , w11535 , w11536 , w11537 , w11538 , w11539 , w11540 , w11541 , w11542 , w11543 , w11544 , w11545 , w11546 , w11547 , w11548 , w11549 , w11550 , w11551 , w11552 , w11553 , w11554 , w11555 , w11556 , w11557 , w11558 , w11559 , w11560 , w11561 , w11562 , w11563 , w11564 , w11565 , w11566 , w11567 , w11568 , w11569 , w11570 , w11571 , w11572 , w11573 , w11574 , w11575 , w11576 , w11577 , w11578 , w11579 , w11580 , w11581 , w11582 , w11583 , w11584 , w11585 , w11586 , w11587 , w11588 , w11589 , w11590 , w11591 , w11592 , w11593 , w11594 , w11595 , w11596 , w11597 , w11598 , w11599 , w11600 , w11601 , w11602 , w11603 , w11604 , w11605 , w11606 , w11607 , w11608 , w11609 , w11610 , w11611 , w11612 , w11613 , w11614 , w11615 , w11616 , w11617 , w11618 , w11619 , w11620 , w11621 , w11622 , w11623 , w11624 , w11625 , w11626 , w11627 , w11628 , w11629 , w11630 , w11631 , w11632 , w11633 , w11634 , w11635 , w11636 , w11637 , w11638 , w11639 , w11640 , w11641 , w11642 , w11643 , w11644 , w11645 , w11646 , w11647 , w11648 , w11649 , w11650 , w11651 , w11652 , w11653 , w11654 , w11655 , w11656 , w11657 , w11658 , w11659 , w11660 , w11661 , w11662 , w11663 , w11664 , w11665 , w11666 , w11667 , w11668 , w11669 , w11670 , w11671 , w11672 , w11673 , w11674 , w11675 , w11676 , w11677 , w11678 , w11679 , w11680 , w11681 , w11682 , w11683 , w11684 , w11685 , w11686 , w11687 , w11688 , w11689 , w11690 , w11691 , w11692 , w11693 , w11694 , w11695 , w11696 , w11697 , w11698 , w11699 , w11700 , w11701 , w11702 , w11703 , w11704 , w11705 , w11706 , w11707 , w11708 , w11709 , w11710 , w11711 , w11712 , w11713 , w11714 , w11715 , w11716 , w11717 , w11718 , w11719 , w11720 , w11721 , w11722 , w11723 , w11724 , w11725 , w11726 , w11727 , w11728 , w11729 , w11730 , w11731 , w11732 , w11733 , w11734 , w11735 , w11736 , w11737 , w11738 , w11739 , w11740 , w11741 , w11742 , w11743 , w11744 , w11745 , w11746 , w11747 , w11748 , w11749 , w11750 , w11751 , w11752 , w11753 , w11754 , w11755 , w11756 , w11757 , w11758 , w11759 , w11760 , w11761 , w11762 , w11763 , w11764 , w11765 , w11766 , w11767 , w11768 , w11769 , w11770 , w11771 , w11772 , w11773 , w11774 , w11775 , w11776 , w11777 , w11778 , w11779 , w11780 , w11781 , w11782 , w11783 , w11784 , w11785 , w11786 , w11787 , w11788 , w11789 , w11790 , w11791 , w11792 , w11793 , w11794 , w11795 , w11796 , w11797 , w11798 , w11799 , w11800 , w11801 , w11802 , w11803 , w11804 , w11805 , w11806 , w11807 , w11808 , w11809 , w11810 , w11811 , w11812 , w11813 , w11814 , w11815 , w11816 , w11817 , w11818 , w11819 , w11820 , w11821 , w11822 , w11823 , w11824 , w11825 , w11826 , w11827 , w11828 , w11829 , w11830 , w11831 , w11832 , w11833 , w11834 , w11835 , w11836 , w11837 , w11838 , w11839 , w11840 , w11841 , w11842 , w11843 , w11844 , w11845 , w11846 , w11847 , w11848 , w11849 , w11850 , w11851 , w11852 , w11853 , w11854 , w11855 , w11856 , w11857 , w11858 , w11859 , w11860 , w11861 , w11862 , w11863 , w11864 , w11865 , w11866 , w11867 , w11868 , w11869 , w11870 , w11871 , w11872 , w11873 , w11874 , w11875 , w11876 , w11877 , w11878 , w11879 , w11880 , w11881 , w11882 , w11883 , w11884 , w11885 , w11886 , w11887 , w11888 , w11889 , w11890 , w11891 , w11892 , w11893 , w11894 , w11895 , w11896 , w11897 , w11898 , w11899 , w11900 , w11901 , w11902 , w11903 , w11904 , w11905 , w11906 , w11907 , w11908 , w11909 , w11910 , w11911 , w11912 , w11913 , w11914 , w11915 , w11916 , w11917 , w11918 , w11919 , w11920 , w11921 , w11922 , w11923 , w11924 , w11925 , w11926 , w11927 , w11928 , w11929 , w11930 , w11931 , w11932 , w11933 , w11934 , w11935 , w11936 , w11937 , w11938 , w11939 , w11940 , w11941 , w11942 , w11943 , w11944 , w11945 , w11946 , w11947 , w11948 , w11949 , w11950 , w11951 , w11952 , w11953 , w11954 , w11955 , w11956 , w11957 , w11958 , w11959 , w11960 , w11961 , w11962 , w11963 , w11964 , w11965 , w11966 , w11967 , w11968 , w11969 , w11970 , w11971 , w11972 , w11973 , w11974 , w11975 , w11976 , w11977 , w11978 , w11979 , w11980 , w11981 , w11982 , w11983 , w11984 , w11985 , w11986 , w11987 , w11988 , w11989 , w11990 , w11991 , w11992 , w11993 , w11994 , w11995 , w11996 , w11997 , w11998 , w11999 , w12000 , w12001 , w12002 , w12003 , w12004 , w12005 , w12006 , w12007 , w12008 , w12009 , w12010 , w12011 , w12012 , w12013 , w12014 , w12015 , w12016 , w12017 , w12018 , w12019 , w12020 , w12021 , w12022 , w12023 , w12024 , w12025 , w12026 , w12027 , w12028 , w12029 , w12030 , w12031 , w12032 , w12033 , w12034 , w12035 , w12036 , w12037 , w12038 , w12039 , w12040 , w12041 , w12042 , w12043 , w12044 , w12045 , w12046 , w12047 , w12048 , w12049 , w12050 , w12051 , w12052 , w12053 , w12054 , w12055 , w12056 , w12057 , w12058 , w12059 , w12060 , w12061 , w12062 , w12063 , w12064 , w12065 , w12066 , w12067 , w12068 , w12069 , w12070 , w12071 , w12072 , w12073 , w12074 , w12075 , w12076 , w12077 , w12078 , w12079 , w12080 , w12081 , w12082 , w12083 , w12084 , w12085 , w12086 , w12087 , w12088 , w12089 , w12090 , w12091 , w12092 , w12093 , w12094 , w12095 , w12096 , w12097 , w12098 , w12099 , w12100 , w12101 , w12102 , w12103 , w12104 , w12105 , w12106 , w12107 , w12108 , w12109 , w12110 , w12111 , w12112 , w12113 , w12114 , w12115 , w12116 , w12117 , w12118 , w12119 , w12120 , w12121 , w12122 , w12123 , w12124 , w12125 , w12126 , w12127 , w12128 , w12129 , w12130 , w12131 , w12132 , w12133 , w12134 , w12135 , w12136 , w12137 , w12138 , w12139 , w12140 , w12141 , w12142 , w12143 , w12144 , w12145 , w12146 , w12147 , w12148 , w12149 , w12150 , w12151 , w12152 , w12153 , w12154 , w12155 , w12156 , w12157 , w12158 , w12159 , w12160 , w12161 , w12162 , w12163 , w12164 , w12165 , w12166 , w12167 , w12168 , w12169 , w12170 , w12171 , w12172 , w12173 , w12174 , w12175 , w12176 , w12177 , w12178 , w12179 , w12180 , w12181 , w12182 , w12183 , w12184 , w12185 , w12186 , w12187 , w12188 , w12189 , w12190 , w12191 , w12192 , w12193 , w12194 , w12195 , w12196 , w12197 , w12198 , w12199 , w12200 , w12201 , w12202 , w12203 , w12204 , w12205 , w12206 , w12207 , w12208 , w12209 , w12210 , w12211 , w12212 , w12213 , w12214 , w12215 , w12216 , w12217 , w12218 , w12219 , w12220 , w12221 , w12222 , w12223 , w12224 , w12225 , w12226 , w12227 , w12228 , w12229 , w12230 , w12231 , w12232 , w12233 , w12234 , w12235 , w12236 , w12237 , w12238 , w12239 , w12240 , w12241 , w12242 , w12243 , w12244 , w12245 , w12246 , w12247 , w12248 , w12249 , w12250 , w12251 , w12252 , w12253 , w12254 , w12255 , w12256 , w12257 , w12258 , w12259 , w12260 , w12261 , w12262 , w12263 , w12264 , w12265 , w12266 , w12267 , w12268 , w12269 , w12270 , w12271 , w12272 , w12273 , w12274 , w12275 , w12276 , w12277 , w12278 , w12279 , w12280 , w12281 , w12282 , w12283 , w12284 , w12285 , w12286 , w12287 , w12288 , w12289 , w12290 , w12291 , w12292 , w12293 , w12294 , w12295 , w12296 , w12297 , w12298 , w12299 , w12300 , w12301 , w12302 , w12303 , w12304 , w12305 , w12306 , w12307 , w12308 , w12309 , w12310 , w12311 , w12312 , w12313 , w12314 , w12315 , w12316 , w12317 , w12318 , w12319 , w12320 , w12321 , w12322 , w12323 , w12324 , w12325 , w12326 , w12327 , w12328 , w12329 , w12330 , w12331 , w12332 , w12333 , w12334 , w12335 , w12336 , w12337 , w12338 , w12339 , w12340 , w12341 , w12342 , w12343 , w12344 , w12345 , w12346 , w12347 , w12348 , w12349 , w12350 , w12351 , w12352 , w12353 , w12354 , w12355 , w12356 , w12357 , w12358 , w12359 , w12360 , w12361 , w12362 , w12363 , w12364 , w12365 , w12366 , w12367 , w12368 , w12369 , w12370 , w12371 , w12372 , w12373 , w12374 , w12375 , w12376 , w12377 , w12378 , w12379 , w12380 , w12381 , w12382 , w12383 , w12384 , w12385 , w12386 , w12387 , w12388 , w12389 , w12390 , w12391 , w12392 , w12393 , w12394 , w12395 , w12396 , w12397 , w12398 , w12399 , w12400 , w12401 , w12402 , w12403 , w12404 , w12405 , w12406 , w12407 , w12408 , w12409 , w12410 , w12411 , w12412 , w12413 , w12414 , w12415 , w12416 , w12417 , w12418 , w12419 , w12420 , w12421 , w12422 , w12423 , w12424 , w12425 , w12426 , w12427 , w12428 , w12429 , w12430 , w12431 , w12432 , w12433 , w12434 , w12435 , w12436 , w12437 , w12438 , w12439 , w12440 , w12441 , w12442 , w12443 , w12444 , w12445 , w12446 , w12447 , w12448 , w12449 , w12450 , w12451 , w12452 , w12453 , w12454 , w12455 , w12456 , w12457 , w12458 , w12459 , w12460 , w12461 , w12462 , w12463 , w12464 , w12465 , w12466 , w12467 , w12468 , w12469 , w12470 , w12471 , w12472 , w12473 , w12474 , w12475 , w12476 , w12477 , w12478 , w12479 , w12480 , w12481 , w12482 , w12483 , w12484 , w12485 , w12486 , w12487 , w12488 , w12489 , w12490 , w12491 , w12492 , w12493 , w12494 , w12495 , w12496 , w12497 , w12498 , w12499 , w12500 , w12501 , w12502 , w12503 , w12504 , w12505 , w12506 , w12507 , w12508 , w12509 , w12510 , w12511 , w12512 , w12513 , w12514 , w12515 , w12516 , w12517 , w12518 , w12519 , w12520 , w12521 , w12522 , w12523 , w12524 , w12525 , w12526 , w12527 , w12528 , w12529 , w12530 , w12531 , w12532 , w12533 , w12534 , w12535 , w12536 , w12537 , w12538 , w12539 , w12540 , w12541 , w12542 , w12543 , w12544 , w12545 , w12546 , w12547 , w12548 , w12549 , w12550 , w12551 , w12552 , w12553 , w12554 , w12555 , w12556 , w12557 , w12558 , w12559 , w12560 , w12561 , w12562 , w12563 , w12564 , w12565 , w12566 , w12567 , w12568 , w12569 , w12570 , w12571 , w12572 , w12573 , w12574 , w12575 , w12576 , w12577 , w12578 , w12579 , w12580 , w12581 , w12582 , w12583 , w12584 , w12585 , w12586 , w12587 , w12588 , w12589 , w12590 , w12591 , w12592 , w12593 , w12594 , w12595 , w12596 , w12597 , w12598 , w12599 , w12600 , w12601 , w12602 , w12603 , w12604 , w12605 , w12606 , w12607 , w12608 , w12609 , w12610 , w12611 , w12612 , w12613 , w12614 , w12615 , w12616 , w12617 , w12618 , w12619 , w12620 , w12621 , w12622 , w12623 , w12624 , w12625 , w12626 , w12627 , w12628 , w12629 , w12630 , w12631 , w12632 , w12633 , w12634 , w12635 , w12636 , w12637 , w12638 , w12639 , w12640 , w12641 , w12642 , w12643 , w12644 , w12645 , w12646 , w12647 , w12648 , w12649 , w12650 , w12651 , w12652 , w12653 , w12654 , w12655 , w12656 , w12657 , w12658 , w12659 , w12660 , w12661 , w12662 , w12663 , w12664 , w12665 , w12666 , w12667 , w12668 , w12669 , w12670 , w12671 , w12672 , w12673 , w12674 , w12675 , w12676 , w12677 , w12678 , w12679 , w12680 , w12681 , w12682 , w12683 , w12684 , w12685 , w12686 , w12687 , w12688 , w12689 , w12690 , w12691 , w12692 , w12693 , w12694 , w12695 , w12696 , w12697 , w12698 , w12699 , w12700 , w12701 , w12702 , w12703 , w12704 , w12705 , w12706 , w12707 , w12708 , w12709 , w12710 , w12711 , w12712 , w12713 , w12714 , w12715 , w12716 , w12717 , w12718 , w12719 , w12720 , w12721 , w12722 , w12723 , w12724 , w12725 , w12726 , w12727 , w12728 , w12729 , w12730 , w12731 , w12732 , w12733 , w12734 , w12735 , w12736 , w12737 , w12738 , w12739 , w12740 , w12741 , w12742 , w12743 , w12744 , w12745 , w12746 , w12747 , w12748 , w12749 , w12750 , w12751 , w12752 , w12753 , w12754 , w12755 , w12756 , w12757 , w12758 , w12759 , w12760 , w12761 , w12762 , w12763 , w12764 , w12765 , w12766 , w12767 , w12768 , w12769 , w12770 , w12771 , w12772 , w12773 , w12774 , w12775 , w12776 , w12777 , w12778 , w12779 , w12780 , w12781 , w12782 , w12783 , w12784 , w12785 , w12786 , w12787 , w12788 , w12789 , w12790 , w12791 , w12792 , w12793 , w12794 , w12795 , w12796 , w12797 , w12798 , w12799 , w12800 , w12801 , w12802 , w12803 , w12804 , w12805 , w12806 , w12807 , w12808 , w12809 , w12810 , w12811 , w12812 , w12813 , w12814 , w12815 , w12816 , w12817 , w12818 , w12819 , w12820 , w12821 , w12822 , w12823 , w12824 , w12825 , w12826 , w12827 , w12828 , w12829 , w12830 , w12831 , w12832 , w12833 , w12834 , w12835 , w12836 , w12837 , w12838 , w12839 , w12840 , w12841 , w12842 , w12843 , w12844 , w12845 , w12846 , w12847 , w12848 , w12849 , w12850 , w12851 , w12852 , w12853 , w12854 , w12855 , w12856 , w12857 , w12858 , w12859 , w12860 , w12861 , w12862 , w12863 , w12864 , w12865 , w12866 , w12867 , w12868 , w12869 , w12870 , w12871 , w12872 , w12873 , w12874 , w12875 , w12876 , w12877 , w12878 , w12879 , w12880 , w12881 , w12882 , w12883 , w12884 , w12885 , w12886 , w12887 , w12888 , w12889 , w12890 , w12891 , w12892 , w12893 , w12894 , w12895 , w12896 , w12897 , w12898 , w12899 , w12900 , w12901 , w12902 , w12903 , w12904 , w12905 , w12906 , w12907 , w12908 , w12909 , w12910 , w12911 , w12912 , w12913 , w12914 , w12915 , w12916 , w12917 , w12918 , w12919 , w12920 , w12921 , w12922 , w12923 , w12924 , w12925 , w12926 , w12927 , w12928 , w12929 , w12930 , w12931 , w12932 , w12933 , w12934 , w12935 , w12936 , w12937 , w12938 , w12939 , w12940 , w12941 , w12942 , w12943 , w12944 , w12945 , w12946 , w12947 , w12948 , w12949 , w12950 , w12951 , w12952 , w12953 , w12954 , w12955 , w12956 , w12957 , w12958 , w12959 , w12960 , w12961 , w12962 , w12963 , w12964 , w12965 , w12966 , w12967 , w12968 , w12969 , w12970 , w12971 , w12972 , w12973 , w12974 , w12975 , w12976 , w12977 , w12978 , w12979 , w12980 , w12981 , w12982 , w12983 , w12984 , w12985 , w12986 , w12987 , w12988 , w12989 , w12990 , w12991 , w12992 , w12993 , w12994 , w12995 , w12996 , w12997 , w12998 , w12999 , w13000 , w13001 , w13002 , w13003 , w13004 , w13005 , w13006 , w13007 , w13008 , w13009 , w13010 , w13011 , w13012 , w13013 , w13014 , w13015 , w13016 , w13017 , w13018 , w13019 , w13020 , w13021 , w13022 , w13023 , w13024 , w13025 , w13026 , w13027 , w13028 , w13029 , w13030 , w13031 , w13032 , w13033 , w13034 , w13035 , w13036 , w13037 , w13038 , w13039 , w13040 , w13041 , w13042 , w13043 , w13044 , w13045 , w13046 , w13047 , w13048 , w13049 , w13050 , w13051 , w13052 , w13053 , w13054 , w13055 , w13056 , w13057 , w13058 , w13059 , w13060 , w13061 , w13062 , w13063 , w13064 , w13065 , w13066 , w13067 , w13068 , w13069 , w13070 , w13071 , w13072 , w13073 , w13074 , w13075 , w13076 , w13077 , w13078 , w13079 , w13080 , w13081 , w13082 , w13083 , w13084 , w13085 , w13086 , w13087 , w13088 , w13089 , w13090 , w13091 , w13092 , w13093 , w13094 , w13095 , w13096 , w13097 , w13098 , w13099 , w13100 , w13101 , w13102 , w13103 , w13104 , w13105 , w13106 , w13107 , w13108 , w13109 , w13110 , w13111 , w13112 , w13113 , w13114 , w13115 , w13116 , w13117 , w13118 , w13119 , w13120 , w13121 , w13122 , w13123 , w13124 , w13125 , w13126 , w13127 , w13128 , w13129 , w13130 , w13131 , w13132 , w13133 , w13134 , w13135 , w13136 , w13137 , w13138 , w13139 , w13140 , w13141 , w13142 , w13143 , w13144 , w13145 , w13146 , w13147 , w13148 , w13149 , w13150 , w13151 , w13152 , w13153 , w13154 , w13155 , w13156 , w13157 , w13158 , w13159 , w13160 , w13161 , w13162 , w13163 , w13164 , w13165 , w13166 , w13167 , w13168 , w13169 , w13170 , w13171 , w13172 , w13173 , w13174 , w13175 , w13176 , w13177 , w13178 , w13179 , w13180 , w13181 , w13182 , w13183 , w13184 , w13185 , w13186 , w13187 , w13188 , w13189 , w13190 , w13191 , w13192 , w13193 , w13194 , w13195 , w13196 , w13197 , w13198 , w13199 , w13200 , w13201 , w13202 , w13203 , w13204 , w13205 , w13206 , w13207 , w13208 , w13209 , w13210 , w13211 , w13212 , w13213 , w13214 , w13215 , w13216 , w13217 , w13218 , w13219 , w13220 , w13221 , w13222 , w13223 , w13224 , w13225 , w13226 , w13227 , w13228 , w13229 , w13230 , w13231 , w13232 , w13233 , w13234 , w13235 , w13236 , w13237 , w13238 , w13239 , w13240 , w13241 , w13242 , w13243 , w13244 , w13245 , w13246 , w13247 , w13248 , w13249 , w13250 , w13251 , w13252 , w13253 , w13254 , w13255 , w13256 , w13257 , w13258 , w13259 , w13260 , w13261 , w13262 , w13263 , w13264 , w13265 , w13266 , w13267 , w13268 , w13269 , w13270 , w13271 , w13272 , w13273 , w13274 , w13275 , w13276 , w13277 , w13278 , w13279 , w13280 , w13281 , w13282 , w13283 , w13284 , w13285 , w13286 , w13287 , w13288 , w13289 , w13290 , w13291 , w13292 , w13293 , w13294 , w13295 , w13296 , w13297 , w13298 , w13299 , w13300 , w13301 , w13302 , w13303 , w13304 , w13305 , w13306 , w13307 , w13308 , w13309 , w13310 , w13311 , w13312 , w13313 , w13314 , w13315 , w13316 , w13317 , w13318 , w13319 , w13320 , w13321 , w13322 , w13323 , w13324 , w13325 , w13326 , w13327 , w13328 , w13329 , w13330 , w13331 , w13332 , w13333 , w13334 , w13335 , w13336 , w13337 , w13338 , w13339 , w13340 , w13341 , w13342 , w13343 , w13344 , w13345 , w13346 , w13347 , w13348 , w13349 , w13350 , w13351 , w13352 , w13353 , w13354 , w13355 , w13356 , w13357 , w13358 , w13359 , w13360 , w13361 , w13362 , w13363 , w13364 , w13365 , w13366 , w13367 , w13368 , w13369 , w13370 , w13371 , w13372 , w13373 , w13374 , w13375 , w13376 , w13377 , w13378 , w13379 , w13380 , w13381 , w13382 , w13383 , w13384 , w13385 , w13386 , w13387 , w13388 , w13389 , w13390 , w13391 , w13392 , w13393 , w13394 , w13395 , w13396 , w13397 , w13398 , w13399 , w13400 , w13401 , w13402 , w13403 , w13404 , w13405 , w13406 , w13407 , w13408 , w13409 , w13410 , w13411 , w13412 , w13413 , w13414 , w13415 , w13416 , w13417 , w13418 , w13419 , w13420 , w13421 , w13422 , w13423 , w13424 , w13425 , w13426 , w13427 , w13428 , w13429 , w13430 , w13431 , w13432 , w13433 , w13434 , w13435 , w13436 , w13437 , w13438 , w13439 , w13440 , w13441 , w13442 , w13443 , w13444 , w13445 , w13446 , w13447 , w13448 , w13449 , w13450 , w13451 , w13452 , w13453 , w13454 , w13455 , w13456 , w13457 , w13458 , w13459 , w13460 , w13461 , w13462 , w13463 , w13464 , w13465 , w13466 , w13467 , w13468 , w13469 , w13470 , w13471 , w13472 , w13473 , w13474 , w13475 , w13476 , w13477 , w13478 , w13479 , w13480 , w13481 , w13482 , w13483 , w13484 , w13485 , w13486 , w13487 , w13488 , w13489 , w13490 , w13491 , w13492 , w13493 , w13494 , w13495 , w13496 , w13497 , w13498 , w13499 , w13500 , w13501 , w13502 , w13503 , w13504 , w13505 , w13506 , w13507 , w13508 , w13509 , w13510 , w13511 , w13512 , w13513 , w13514 , w13515 , w13516 , w13517 , w13518 , w13519 , w13520 , w13521 , w13522 , w13523 , w13524 , w13525 , w13526 , w13527 , w13528 , w13529 , w13530 , w13531 , w13532 , w13533 , w13534 , w13535 , w13536 , w13537 , w13538 , w13539 , w13540 , w13541 , w13542 , w13543 , w13544 , w13545 , w13546 , w13547 , w13548 , w13549 , w13550 , w13551 , w13552 , w13553 , w13554 , w13555 , w13556 , w13557 , w13558 , w13559 , w13560 , w13561 , w13562 , w13563 , w13564 , w13565 , w13566 , w13567 , w13568 , w13569 , w13570 , w13571 , w13572 , w13573 , w13574 , w13575 , w13576 , w13577 , w13578 , w13579 , w13580 , w13581 , w13582 , w13583 , w13584 , w13585 , w13586 , w13587 , w13588 , w13589 , w13590 , w13591 , w13592 , w13593 , w13594 , w13595 , w13596 , w13597 , w13598 , w13599 , w13600 , w13601 , w13602 , w13603 , w13604 , w13605 , w13606 , w13607 , w13608 , w13609 , w13610 , w13611 , w13612 , w13613 , w13614 , w13615 , w13616 , w13617 , w13618 , w13619 , w13620 , w13621 , w13622 , w13623 , w13624 , w13625 , w13626 , w13627 , w13628 , w13629 , w13630 , w13631 , w13632 , w13633 , w13634 , w13635 , w13636 , w13637 , w13638 , w13639 , w13640 , w13641 , w13642 , w13643 , w13644 , w13645 , w13646 , w13647 , w13648 , w13649 , w13650 , w13651 , w13652 , w13653 , w13654 , w13655 , w13656 , w13657 , w13658 , w13659 , w13660 , w13661 , w13662 , w13663 , w13664 , w13665 , w13666 , w13667 , w13668 , w13669 , w13670 , w13671 , w13672 , w13673 , w13674 , w13675 , w13676 , w13677 , w13678 , w13679 , w13680 , w13681 , w13682 , w13683 , w13684 , w13685 , w13686 , w13687 , w13688 , w13689 , w13690 , w13691 , w13692 , w13693 , w13694 , w13695 , w13696 , w13697 , w13698 , w13699 , w13700 , w13701 , w13702 , w13703 , w13704 , w13705 , w13706 , w13707 , w13708 , w13709 , w13710 , w13711 , w13712 , w13713 , w13714 , w13715 , w13716 , w13717 , w13718 , w13719 , w13720 , w13721 , w13722 , w13723 , w13724 , w13725 , w13726 , w13727 , w13728 , w13729 , w13730 , w13731 , w13732 , w13733 , w13734 , w13735 , w13736 , w13737 , w13738 , w13739 , w13740 , w13741 , w13742 , w13743 , w13744 , w13745 , w13746 , w13747 , w13748 , w13749 , w13750 , w13751 , w13752 , w13753 , w13754 , w13755 , w13756 , w13757 , w13758 , w13759 , w13760 , w13761 , w13762 , w13763 , w13764 , w13765 , w13766 , w13767 , w13768 , w13769 , w13770 , w13771 , w13772 , w13773 , w13774 , w13775 , w13776 , w13777 , w13778 , w13779 , w13780 , w13781 , w13782 , w13783 , w13784 , w13785 , w13786 , w13787 , w13788 , w13789 , w13790 , w13791 , w13792 , w13793 , w13794 , w13795 , w13796 , w13797 , w13798 , w13799 , w13800 , w13801 , w13802 , w13803 , w13804 , w13805 , w13806 , w13807 , w13808 , w13809 , w13810 , w13811 , w13812 , w13813 , w13814 , w13815 , w13816 , w13817 , w13818 , w13819 , w13820 , w13821 , w13822 , w13823 , w13824 , w13825 , w13826 , w13827 , w13828 , w13829 , w13830 , w13831 , w13832 , w13833 , w13834 , w13835 , w13836 , w13837 , w13838 , w13839 , w13840 , w13841 , w13842 , w13843 , w13844 , w13845 , w13846 , w13847 , w13848 , w13849 , w13850 , w13851 , w13852 , w13853 , w13854 , w13855 , w13856 , w13857 , w13858 , w13859 , w13860 , w13861 , w13862 , w13863 , w13864 , w13865 , w13866 , w13867 , w13868 , w13869 , w13870 , w13871 , w13872 , w13873 , w13874 , w13875 , w13876 , w13877 , w13878 , w13879 , w13880 , w13881 , w13882 , w13883 , w13884 , w13885 , w13886 , w13887 , w13888 , w13889 , w13890 , w13891 , w13892 , w13893 , w13894 , w13895 , w13896 , w13897 , w13898 , w13899 , w13900 , w13901 , w13902 , w13903 , w13904 , w13905 , w13906 , w13907 , w13908 , w13909 , w13910 , w13911 , w13912 , w13913 , w13914 , w13915 , w13916 , w13917 , w13918 , w13919 , w13920 , w13921 , w13922 , w13923 , w13924 , w13925 , w13926 , w13927 , w13928 , w13929 , w13930 , w13931 , w13932 , w13933 , w13934 , w13935 , w13936 , w13937 , w13938 , w13939 , w13940 , w13941 , w13942 , w13943 , w13944 , w13945 , w13946 , w13947 , w13948 , w13949 , w13950 , w13951 , w13952 , w13953 , w13954 , w13955 , w13956 , w13957 , w13958 , w13959 , w13960 , w13961 , w13962 , w13963 , w13964 , w13965 , w13966 , w13967 , w13968 , w13969 , w13970 , w13971 , w13972 , w13973 , w13974 , w13975 , w13976 , w13977 , w13978 , w13979 , w13980 , w13981 , w13982 , w13983 , w13984 , w13985 , w13986 , w13987 , w13988 , w13989 , w13990 , w13991 , w13992 , w13993 , w13994 , w13995 , w13996 , w13997 , w13998 , w13999 , w14000 , w14001 , w14002 , w14003 , w14004 , w14005 , w14006 , w14007 , w14008 , w14009 , w14010 , w14011 , w14012 , w14013 , w14014 , w14015 , w14016 , w14017 , w14018 , w14019 , w14020 , w14021 , w14022 , w14023 , w14024 , w14025 , w14026 , w14027 , w14028 , w14029 , w14030 , w14031 , w14032 , w14033 , w14034 , w14035 , w14036 , w14037 , w14038 , w14039 , w14040 , w14041 , w14042 , w14043 , w14044 , w14045 , w14046 , w14047 , w14048 , w14049 , w14050 , w14051 , w14052 , w14053 , w14054 , w14055 , w14056 , w14057 , w14058 , w14059 , w14060 , w14061 , w14062 , w14063 , w14064 , w14065 , w14066 , w14067 , w14068 , w14069 , w14070 , w14071 , w14072 , w14073 , w14074 , w14075 , w14076 , w14077 , w14078 , w14079 , w14080 , w14081 , w14082 , w14083 , w14084 , w14085 , w14086 , w14087 , w14088 , w14089 , w14090 , w14091 , w14092 , w14093 , w14094 , w14095 , w14096 , w14097 , w14098 , w14099 , w14100 , w14101 , w14102 , w14103 , w14104 , w14105 , w14106 , w14107 , w14108 , w14109 , w14110 , w14111 , w14112 , w14113 , w14114 , w14115 , w14116 , w14117 , w14118 , w14119 , w14120 , w14121 , w14122 , w14123 , w14124 , w14125 , w14126 , w14127 , w14128 , w14129 , w14130 , w14131 , w14132 , w14133 , w14134 , w14135 , w14136 , w14137 , w14138 , w14139 , w14140 , w14141 , w14142 , w14143 , w14144 , w14145 , w14146 , w14147 , w14148 , w14149 , w14150 , w14151 , w14152 , w14153 , w14154 , w14155 , w14156 , w14157 , w14158 , w14159 , w14160 , w14161 , w14162 , w14163 , w14164 , w14165 , w14166 , w14167 , w14168 , w14169 , w14170 , w14171 , w14172 , w14173 , w14174 , w14175 , w14176 , w14177 , w14178 , w14179 , w14180 , w14181 , w14182 , w14183 , w14184 , w14185 , w14186 , w14187 , w14188 , w14189 , w14190 , w14191 , w14192 , w14193 , w14194 , w14195 , w14196 , w14197 , w14198 , w14199 , w14200 , w14201 , w14202 , w14203 , w14204 , w14205 , w14206 , w14207 , w14208 , w14209 , w14210 , w14211 , w14212 , w14213 , w14214 , w14215 , w14216 , w14217 , w14218 , w14219 , w14220 , w14221 , w14222 , w14223 , w14224 , w14225 , w14226 , w14227 , w14228 , w14229 , w14230 , w14231 , w14232 , w14233 , w14234 , w14235 , w14236 , w14237 , w14238 , w14239 , w14240 , w14241 , w14242 , w14243 , w14244 , w14245 , w14246 , w14247 , w14248 , w14249 , w14250 , w14251 , w14252 , w14253 , w14254 , w14255 , w14256 , w14257 , w14258 , w14259 , w14260 , w14261 , w14262 , w14263 , w14264 , w14265 , w14266 , w14267 , w14268 , w14269 , w14270 , w14271 , w14272 , w14273 , w14274 , w14275 , w14276 , w14277 , w14278 , w14279 , w14280 , w14281 , w14282 , w14283 , w14284 , w14285 , w14286 , w14287 , w14288 , w14289 , w14290 , w14291 , w14292 , w14293 , w14294 , w14295 , w14296 , w14297 , w14298 , w14299 , w14300 , w14301 , w14302 , w14303 , w14304 , w14305 , w14306 , w14307 , w14308 , w14309 , w14310 , w14311 , w14312 , w14313 , w14314 , w14315 , w14316 , w14317 , w14318 , w14319 , w14320 , w14321 , w14322 , w14323 , w14324 , w14325 , w14326 , w14327 , w14328 , w14329 , w14330 , w14331 , w14332 , w14333 , w14334 , w14335 , w14336 , w14337 , w14338 , w14339 , w14340 , w14341 , w14342 , w14343 , w14344 , w14345 , w14346 , w14347 , w14348 , w14349 , w14350 , w14351 , w14352 , w14353 , w14354 , w14355 , w14356 , w14357 , w14358 , w14359 , w14360 , w14361 , w14362 , w14363 , w14364 , w14365 , w14366 , w14367 , w14368 , w14369 , w14370 , w14371 , w14372 , w14373 , w14374 , w14375 , w14376 , w14377 , w14378 , w14379 , w14380 , w14381 , w14382 , w14383 , w14384 , w14385 , w14386 , w14387 , w14388 , w14389 , w14390 , w14391 , w14392 , w14393 , w14394 , w14395 , w14396 , w14397 , w14398 , w14399 , w14400 , w14401 , w14402 , w14403 , w14404 , w14405 , w14406 , w14407 , w14408 , w14409 , w14410 , w14411 , w14412 , w14413 , w14414 , w14415 , w14416 , w14417 , w14418 , w14419 , w14420 , w14421 , w14422 , w14423 , w14424 , w14425 , w14426 , w14427 , w14428 , w14429 , w14430 , w14431 , w14432 , w14433 , w14434 , w14435 , w14436 , w14437 , w14438 , w14439 , w14440 , w14441 , w14442 , w14443 , w14444 , w14445 , w14446 , w14447 , w14448 , w14449 , w14450 , w14451 , w14452 , w14453 , w14454 , w14455 , w14456 , w14457 , w14458 , w14459 , w14460 , w14461 , w14462 , w14463 , w14464 , w14465 , w14466 , w14467 , w14468 , w14469 , w14470 , w14471 , w14472 , w14473 , w14474 , w14475 , w14476 , w14477 , w14478 , w14479 , w14480 , w14481 , w14482 , w14483 , w14484 , w14485 , w14486 , w14487 , w14488 , w14489 , w14490 , w14491 , w14492 , w14493 , w14494 , w14495 , w14496 , w14497 , w14498 , w14499 , w14500 , w14501 , w14502 , w14503 , w14504 , w14505 , w14506 , w14507 , w14508 , w14509 , w14510 , w14511 , w14512 , w14513 , w14514 , w14515 , w14516 , w14517 , w14518 , w14519 , w14520 , w14521 , w14522 , w14523 , w14524 , w14525 , w14526 , w14527 , w14528 , w14529 , w14530 , w14531 , w14532 , w14533 , w14534 , w14535 , w14536 , w14537 , w14538 , w14539 , w14540 , w14541 , w14542 , w14543 , w14544 , w14545 , w14546 , w14547 , w14548 , w14549 , w14550 , w14551 , w14552 , w14553 , w14554 , w14555 , w14556 , w14557 , w14558 , w14559 , w14560 , w14561 , w14562 , w14563 , w14564 , w14565 , w14566 , w14567 , w14568 , w14569 , w14570 , w14571 , w14572 , w14573 , w14574 , w14575 , w14576 , w14577 , w14578 , w14579 , w14580 , w14581 , w14582 , w14583 , w14584 , w14585 , w14586 , w14587 , w14588 , w14589 , w14590 , w14591 , w14592 , w14593 , w14594 , w14595 , w14596 , w14597 , w14598 , w14599 , w14600 , w14601 , w14602 , w14603 , w14604 , w14605 , w14606 , w14607 , w14608 , w14609 , w14610 , w14611 , w14612 , w14613 , w14614 , w14615 , w14616 , w14617 , w14618 , w14619 , w14620 , w14621 , w14622 , w14623 , w14624 , w14625 , w14626 , w14627 , w14628 , w14629 , w14630 , w14631 , w14632 , w14633 , w14634 , w14635 , w14636 , w14637 , w14638 , w14639 , w14640 , w14641 , w14642 , w14643 , w14644 , w14645 , w14646 , w14647 , w14648 , w14649 , w14650 , w14651 , w14652 , w14653 , w14654 , w14655 , w14656 , w14657 , w14658 , w14659 , w14660 , w14661 , w14662 , w14663 , w14664 , w14665 , w14666 , w14667 , w14668 , w14669 , w14670 , w14671 , w14672 , w14673 , w14674 , w14675 , w14676 , w14677 , w14678 , w14679 , w14680 , w14681 , w14682 , w14683 , w14684 , w14685 , w14686 , w14687 , w14688 , w14689 , w14690 , w14691 , w14692 , w14693 , w14694 , w14695 , w14696 , w14697 , w14698 , w14699 , w14700 , w14701 , w14702 , w14703 , w14704 , w14705 , w14706 , w14707 , w14708 , w14709 , w14710 , w14711 , w14712 , w14713 , w14714 , w14715 , w14716 , w14717 , w14718 , w14719 , w14720 , w14721 , w14722 , w14723 , w14724 , w14725 , w14726 , w14727 , w14728 , w14729 , w14730 , w14731 , w14732 , w14733 , w14734 , w14735 , w14736 , w14737 , w14738 , w14739 , w14740 , w14741 , w14742 , w14743 , w14744 , w14745 , w14746 , w14747 , w14748 , w14749 , w14750 , w14751 , w14752 , w14753 , w14754 , w14755 , w14756 , w14757 , w14758 , w14759 , w14760 , w14761 , w14762 , w14763 , w14764 , w14765 , w14766 , w14767 , w14768 , w14769 , w14770 , w14771 , w14772 , w14773 , w14774 , w14775 , w14776 , w14777 , w14778 , w14779 , w14780 , w14781 , w14782 , w14783 , w14784 , w14785 , w14786 , w14787 , w14788 , w14789 , w14790 , w14791 , w14792 , w14793 , w14794 , w14795 , w14796 , w14797 , w14798 , w14799 , w14800 , w14801 , w14802 , w14803 , w14804 , w14805 , w14806 , w14807 , w14808 , w14809 , w14810 , w14811 , w14812 , w14813 , w14814 , w14815 , w14816 , w14817 , w14818 , w14819 , w14820 , w14821 , w14822 , w14823 , w14824 , w14825 , w14826 , w14827 , w14828 , w14829 , w14830 , w14831 , w14832 , w14833 , w14834 , w14835 , w14836 , w14837 , w14838 , w14839 , w14840 , w14841 , w14842 , w14843 , w14844 , w14845 , w14846 , w14847 , w14848 , w14849 , w14850 , w14851 , w14852 , w14853 , w14854 , w14855 , w14856 , w14857 , w14858 , w14859 , w14860 , w14861 , w14862 , w14863 , w14864 , w14865 , w14866 , w14867 , w14868 , w14869 , w14870 , w14871 , w14872 , w14873 , w14874 , w14875 , w14876 , w14877 , w14878 , w14879 , w14880 , w14881 , w14882 , w14883 , w14884 , w14885 , w14886 , w14887 , w14888 , w14889 , w14890 , w14891 , w14892 , w14893 , w14894 , w14895 , w14896 , w14897 , w14898 , w14899 , w14900 , w14901 , w14902 , w14903 , w14904 , w14905 , w14906 , w14907 , w14908 , w14909 , w14910 , w14911 , w14912 , w14913 , w14914 , w14915 , w14916 , w14917 , w14918 , w14919 , w14920 , w14921 , w14922 , w14923 , w14924 , w14925 , w14926 , w14927 , w14928 , w14929 , w14930 , w14931 , w14932 , w14933 , w14934 , w14935 , w14936 , w14937 , w14938 , w14939 , w14940 , w14941 , w14942 , w14943 , w14944 , w14945 , w14946 , w14947 , w14948 , w14949 , w14950 , w14951 , w14952 , w14953 , w14954 , w14955 , w14956 , w14957 , w14958 , w14959 , w14960 , w14961 , w14962 , w14963 , w14964 , w14965 , w14966 , w14967 , w14968 , w14969 , w14970 , w14971 , w14972 , w14973 , w14974 , w14975 , w14976 , w14977 , w14978 , w14979 , w14980 , w14981 , w14982 , w14983 , w14984 , w14985 , w14986 , w14987 , w14988 , w14989 , w14990 , w14991 , w14992 , w14993 , w14994 , w14995 , w14996 , w14997 , w14998 , w14999 , w15000 , w15001 , w15002 , w15003 , w15004 , w15005 , w15006 , w15007 , w15008 , w15009 , w15010 , w15011 , w15012 , w15013 , w15014 , w15015 , w15016 , w15017 , w15018 , w15019 , w15020 , w15021 , w15022 , w15023 , w15024 , w15025 , w15026 , w15027 , w15028 , w15029 , w15030 , w15031 , w15032 , w15033 , w15034 , w15035 , w15036 , w15037 , w15038 , w15039 , w15040 , w15041 , w15042 , w15043 , w15044 , w15045 , w15046 , w15047 , w15048 , w15049 , w15050 , w15051 , w15052 , w15053 , w15054 , w15055 , w15056 , w15057 , w15058 , w15059 , w15060 , w15061 , w15062 , w15063 , w15064 , w15065 , w15066 , w15067 , w15068 , w15069 , w15070 , w15071 , w15072 , w15073 , w15074 , w15075 , w15076 , w15077 , w15078 , w15079 , w15080 , w15081 , w15082 , w15083 , w15084 , w15085 , w15086 , w15087 , w15088 , w15089 , w15090 , w15091 , w15092 , w15093 , w15094 , w15095 , w15096 , w15097 , w15098 , w15099 , w15100 , w15101 , w15102 , w15103 , w15104 , w15105 , w15106 , w15107 , w15108 , w15109 , w15110 , w15111 , w15112 , w15113 , w15114 , w15115 , w15116 , w15117 , w15118 , w15119 , w15120 , w15121 , w15122 , w15123 , w15124 , w15125 , w15126 , w15127 , w15128 , w15129 , w15130 , w15131 , w15132 , w15133 , w15134 , w15135 , w15136 , w15137 , w15138 , w15139 , w15140 , w15141 , w15142 , w15143 , w15144 , w15145 , w15146 , w15147 , w15148 , w15149 , w15150 , w15151 , w15152 , w15153 , w15154 , w15155 , w15156 , w15157 , w15158 , w15159 , w15160 , w15161 , w15162 , w15163 , w15164 , w15165 , w15166 , w15167 , w15168 , w15169 , w15170 , w15171 , w15172 , w15173 , w15174 , w15175 , w15176 , w15177 , w15178 , w15179 , w15180 , w15181 , w15182 , w15183 , w15184 , w15185 , w15186 , w15187 , w15188 , w15189 , w15190 , w15191 , w15192 , w15193 , w15194 , w15195 , w15196 , w15197 , w15198 , w15199 , w15200 , w15201 , w15202 , w15203 , w15204 , w15205 , w15206 , w15207 , w15208 , w15209 , w15210 , w15211 , w15212 , w15213 , w15214 , w15215 , w15216 , w15217 , w15218 , w15219 , w15220 , w15221 , w15222 , w15223 , w15224 , w15225 , w15226 , w15227 , w15228 , w15229 , w15230 , w15231 , w15232 , w15233 , w15234 , w15235 , w15236 , w15237 , w15238 , w15239 , w15240 , w15241 , w15242 , w15243 , w15244 , w15245 , w15246 , w15247 , w15248 , w15249 , w15250 , w15251 , w15252 , w15253 , w15254 , w15255 , w15256 , w15257 , w15258 , w15259 , w15260 , w15261 , w15262 , w15263 , w15264 , w15265 , w15266 , w15267 , w15268 , w15269 , w15270 , w15271 , w15272 , w15273 , w15274 , w15275 , w15276 , w15277 , w15278 , w15279 , w15280 , w15281 , w15282 , w15283 , w15284 , w15285 , w15286 , w15287 , w15288 , w15289 , w15290 , w15291 , w15292 , w15293 , w15294 , w15295 , w15296 , w15297 , w15298 , w15299 , w15300 , w15301 , w15302 , w15303 , w15304 , w15305 , w15306 , w15307 , w15308 , w15309 , w15310 , w15311 , w15312 , w15313 , w15314 , w15315 , w15316 , w15317 , w15318 , w15319 , w15320 , w15321 , w15322 , w15323 , w15324 , w15325 , w15326 , w15327 , w15328 , w15329 , w15330 , w15331 , w15332 , w15333 , w15334 , w15335 , w15336 , w15337 , w15338 , w15339 , w15340 , w15341 , w15342 , w15343 , w15344 , w15345 , w15346 , w15347 , w15348 , w15349 , w15350 , w15351 , w15352 , w15353 , w15354 , w15355 , w15356 , w15357 , w15358 , w15359 , w15360 , w15361 , w15362 , w15363 , w15364 , w15365 , w15366 , w15367 , w15368 , w15369 , w15370 , w15371 , w15372 , w15373 , w15374 , w15375 , w15376 , w15377 , w15378 , w15379 , w15380 , w15381 , w15382 , w15383 , w15384 , w15385 , w15386 , w15387 , w15388 , w15389 , w15390 , w15391 , w15392 , w15393 , w15394 , w15395 , w15396 , w15397 , w15398 , w15399 , w15400 , w15401 , w15402 , w15403 , w15404 , w15405 , w15406 , w15407 , w15408 , w15409 , w15410 , w15411 , w15412 , w15413 , w15414 , w15415 , w15416 , w15417 , w15418 , w15419 , w15420 , w15421 , w15422 , w15423 , w15424 , w15425 , w15426 , w15427 , w15428 , w15429 , w15430 , w15431 , w15432 , w15433 , w15434 , w15435 , w15436 , w15437 , w15438 , w15439 , w15440 , w15441 , w15442 , w15443 , w15444 , w15445 , w15446 , w15447 , w15448 , w15449 , w15450 , w15451 , w15452 , w15453 , w15454 , w15455 , w15456 , w15457 , w15458 , w15459 , w15460 , w15461 , w15462 , w15463 , w15464 , w15465 , w15466 , w15467 , w15468 , w15469 , w15470 , w15471 , w15472 , w15473 , w15474 , w15475 , w15476 , w15477 , w15478 , w15479 , w15480 , w15481 , w15482 , w15483 , w15484 , w15485 , w15486 , w15487 , w15488 , w15489 , w15490 , w15491 , w15492 , w15493 , w15494 , w15495 , w15496 , w15497 , w15498 , w15499 , w15500 , w15501 , w15502 , w15503 , w15504 , w15505 , w15506 , w15507 , w15508 , w15509 , w15510 , w15511 , w15512 , w15513 , w15514 , w15515 , w15516 , w15517 , w15518 , w15519 , w15520 , w15521 , w15522 , w15523 , w15524 , w15525 , w15526 , w15527 , w15528 , w15529 , w15530 , w15531 , w15532 , w15533 , w15534 , w15535 , w15536 , w15537 , w15538 , w15539 , w15540 , w15541 , w15542 , w15543 , w15544 , w15545 , w15546 , w15547 , w15548 , w15549 , w15550 , w15551 , w15552 , w15553 , w15554 , w15555 , w15556 , w15557 , w15558 , w15559 , w15560 , w15561 , w15562 , w15563 , w15564 , w15565 , w15566 , w15567 , w15568 , w15569 , w15570 , w15571 , w15572 , w15573 , w15574 , w15575 , w15576 , w15577 , w15578 , w15579 , w15580 , w15581 , w15582 , w15583 , w15584 , w15585 , w15586 , w15587 , w15588 , w15589 , w15590 , w15591 , w15592 , w15593 , w15594 , w15595 , w15596 , w15597 , w15598 , w15599 , w15600 , w15601 , w15602 , w15603 , w15604 , w15605 , w15606 , w15607 , w15608 , w15609 , w15610 , w15611 , w15612 , w15613 , w15614 , w15615 , w15616 , w15617 , w15618 , w15619 , w15620 , w15621 , w15622 , w15623 , w15624 , w15625 , w15626 , w15627 , w15628 , w15629 , w15630 , w15631 , w15632 , w15633 , w15634 , w15635 , w15636 , w15637 , w15638 , w15639 , w15640 , w15641 , w15642 , w15643 , w15644 , w15645 , w15646 , w15647 , w15648 , w15649 , w15650 , w15651 , w15652 , w15653 , w15654 , w15655 , w15656 , w15657 , w15658 , w15659 , w15660 , w15661 , w15662 , w15663 , w15664 , w15665 , w15666 , w15667 , w15668 , w15669 , w15670 , w15671 , w15672 , w15673 , w15674 , w15675 , w15676 , w15677 , w15678 , w15679 , w15680 , w15681 , w15682 , w15683 , w15684 , w15685 , w15686 , w15687 , w15688 , w15689 , w15690 , w15691 , w15692 , w15693 , w15694 , w15695 , w15696 , w15697 , w15698 , w15699 , w15700 , w15701 , w15702 , w15703 , w15704 , w15705 , w15706 , w15707 , w15708 , w15709 , w15710 , w15711 , w15712 , w15713 , w15714 , w15715 , w15716 , w15717 , w15718 , w15719 , w15720 , w15721 , w15722 , w15723 , w15724 , w15725 , w15726 , w15727 , w15728 , w15729 , w15730 , w15731 , w15732 , w15733 , w15734 , w15735 , w15736 , w15737 , w15738 , w15739 , w15740 , w15741 , w15742 , w15743 , w15744 , w15745 , w15746 , w15747 , w15748 , w15749 , w15750 , w15751 , w15752 , w15753 , w15754 , w15755 , w15756 , w15757 , w15758 , w15759 , w15760 , w15761 , w15762 , w15763 , w15764 , w15765 , w15766 , w15767 , w15768 , w15769 , w15770 , w15771 , w15772 , w15773 , w15774 , w15775 , w15776 , w15777 , w15778 , w15779 , w15780 , w15781 , w15782 , w15783 , w15784 , w15785 , w15786 , w15787 , w15788 , w15789 , w15790 , w15791 , w15792 , w15793 , w15794 , w15795 , w15796 , w15797 , w15798 , w15799 , w15800 , w15801 , w15802 , w15803 , w15804 , w15805 , w15806 , w15807 , w15808 , w15809 , w15810 , w15811 , w15812 , w15813 , w15814 , w15815 , w15816 , w15817 , w15818 , w15819 , w15820 , w15821 , w15822 , w15823 , w15824 , w15825 , w15826 , w15827 , w15828 , w15829 , w15830 , w15831 , w15832 , w15833 , w15834 , w15835 , w15836 , w15837 , w15838 , w15839 , w15840 , w15841 , w15842 , w15843 , w15844 , w15845 , w15846 , w15847 , w15848 , w15849 , w15850 , w15851 , w15852 , w15853 , w15854 , w15855 , w15856 , w15857 , w15858 , w15859 , w15860 , w15861 , w15862 , w15863 , w15864 , w15865 , w15866 , w15867 , w15868 , w15869 , w15870 , w15871 , w15872 , w15873 , w15874 , w15875 , w15876 , w15877 , w15878 , w15879 , w15880 , w15881 , w15882 , w15883 , w15884 , w15885 , w15886 , w15887 , w15888 , w15889 , w15890 , w15891 , w15892 , w15893 , w15894 , w15895 , w15896 , w15897 , w15898 , w15899 , w15900 , w15901 , w15902 , w15903 , w15904 , w15905 , w15906 , w15907 , w15908 , w15909 , w15910 , w15911 , w15912 , w15913 , w15914 , w15915 , w15916 , w15917 , w15918 , w15919 , w15920 , w15921 , w15922 , w15923 , w15924 , w15925 , w15926 , w15927 , w15928 , w15929 , w15930 , w15931 , w15932 , w15933 , w15934 , w15935 , w15936 , w15937 , w15938 , w15939 , w15940 , w15941 , w15942 , w15943 , w15944 , w15945 , w15946 , w15947 , w15948 , w15949 , w15950 , w15951 , w15952 , w15953 , w15954 , w15955 , w15956 , w15957 , w15958 , w15959 , w15960 , w15961 , w15962 , w15963 , w15964 , w15965 , w15966 , w15967 , w15968 , w15969 , w15970 , w15971 , w15972 , w15973 , w15974 , w15975 , w15976 , w15977 , w15978 , w15979 , w15980 , w15981 , w15982 , w15983 , w15984 , w15985 , w15986 , w15987 , w15988 , w15989 , w15990 , w15991 , w15992 , w15993 , w15994 , w15995 , w15996 , w15997 , w15998 , w15999 , w16000 , w16001 , w16002 , w16003 , w16004 , w16005 , w16006 , w16007 , w16008 , w16009 , w16010 , w16011 , w16012 , w16013 , w16014 , w16015 , w16016 , w16017 , w16018 , w16019 , w16020 , w16021 , w16022 , w16023 , w16024 , w16025 , w16026 , w16027 , w16028 , w16029 , w16030 , w16031 , w16032 , w16033 , w16034 , w16035 , w16036 , w16037 , w16038 , w16039 , w16040 , w16041 , w16042 , w16043 , w16044 , w16045 , w16046 , w16047 , w16048 , w16049 , w16050 , w16051 , w16052 , w16053 , w16054 , w16055 , w16056 , w16057 , w16058 , w16059 , w16060 , w16061 , w16062 , w16063 , w16064 , w16065 , w16066 , w16067 , w16068 , w16069 , w16070 , w16071 , w16072 , w16073 , w16074 , w16075 , w16076 , w16077 , w16078 , w16079 , w16080 , w16081 , w16082 , w16083 , w16084 , w16085 , w16086 , w16087 , w16088 , w16089 , w16090 , w16091 , w16092 , w16093 , w16094 , w16095 , w16096 , w16097 , w16098 , w16099 , w16100 , w16101 , w16102 , w16103 , w16104 , w16105 , w16106 , w16107 , w16108 , w16109 , w16110 , w16111 , w16112 , w16113 , w16114 , w16115 , w16116 , w16117 , w16118 , w16119 , w16120 , w16121 , w16122 , w16123 , w16124 , w16125 , w16126 , w16127 , w16128 , w16129 , w16130 , w16131 , w16132 , w16133 , w16134 , w16135 , w16136 , w16137 , w16138 , w16139 , w16140 , w16141 , w16142 , w16143 , w16144 , w16145 , w16146 , w16147 , w16148 , w16149 , w16150 , w16151 , w16152 , w16153 , w16154 , w16155 , w16156 , w16157 , w16158 , w16159 , w16160 , w16161 , w16162 , w16163 , w16164 , w16165 , w16166 , w16167 , w16168 , w16169 , w16170 , w16171 , w16172 , w16173 , w16174 , w16175 , w16176 , w16177 , w16178 , w16179 , w16180 , w16181 , w16182 , w16183 , w16184 , w16185 , w16186 , w16187 , w16188 , w16189 , w16190 , w16191 , w16192 , w16193 , w16194 , w16195 , w16196 , w16197 , w16198 , w16199 , w16200 , w16201 , w16202 , w16203 , w16204 , w16205 , w16206 , w16207 , w16208 , w16209 , w16210 , w16211 , w16212 , w16213 , w16214 , w16215 , w16216 , w16217 , w16218 , w16219 , w16220 , w16221 , w16222 , w16223 , w16224 , w16225 , w16226 , w16227 , w16228 , w16229 , w16230 , w16231 , w16232 , w16233 , w16234 , w16235 , w16236 , w16237 , w16238 , w16239 , w16240 , w16241 , w16242 , w16243 , w16244 , w16245 , w16246 , w16247 , w16248 , w16249 , w16250 , w16251 , w16252 , w16253 , w16254 , w16255 , w16256 , w16257 , w16258 , w16259 , w16260 , w16261 , w16262 , w16263 , w16264 , w16265 , w16266 , w16267 , w16268 , w16269 , w16270 , w16271 , w16272 , w16273 , w16274 , w16275 , w16276 , w16277 , w16278 , w16279 , w16280 , w16281 , w16282 , w16283 , w16284 , w16285 , w16286 , w16287 , w16288 , w16289 , w16290 , w16291 , w16292 , w16293 , w16294 , w16295 , w16296 , w16297 , w16298 , w16299 , w16300 , w16301 , w16302 , w16303 , w16304 , w16305 , w16306 , w16307 , w16308 , w16309 , w16310 , w16311 , w16312 , w16313 , w16314 , w16315 , w16316 , w16317 , w16318 , w16319 , w16320 , w16321 , w16322 , w16323 , w16324 , w16325 , w16326 , w16327 , w16328 , w16329 , w16330 , w16331 , w16332 , w16333 , w16334 , w16335 , w16336 , w16337 , w16338 , w16339 , w16340 , w16341 , w16342 , w16343 , w16344 , w16345 , w16346 , w16347 , w16348 , w16349 , w16350 , w16351 , w16352 , w16353 , w16354 , w16355 , w16356 , w16357 , w16358 , w16359 , w16360 , w16361 , w16362 , w16363 , w16364 , w16365 , w16366 , w16367 , w16368 , w16369 , w16370 , w16371 , w16372 , w16373 , w16374 , w16375 , w16376 , w16377 , w16378 , w16379 , w16380 , w16381 , w16382 , w16383 , w16384 , w16385 , w16386 , w16387 , w16388 , w16389 , w16390 , w16391 , w16392 , w16393 , w16394 , w16395 , w16396 , w16397 , w16398 , w16399 , w16400 , w16401 , w16402 , w16403 , w16404 , w16405 , w16406 , w16407 , w16408 , w16409 , w16410 , w16411 , w16412 , w16413 , w16414 , w16415 , w16416 , w16417 , w16418 , w16419 , w16420 , w16421 , w16422 , w16423 , w16424 , w16425 , w16426 , w16427 , w16428 , w16429 , w16430 , w16431 , w16432 , w16433 , w16434 , w16435 , w16436 , w16437 , w16438 , w16439 , w16440 , w16441 , w16442 , w16443 , w16444 , w16445 , w16446 , w16447 , w16448 , w16449 , w16450 , w16451 , w16452 , w16453 , w16454 , w16455 , w16456 , w16457 , w16458 , w16459 , w16460 , w16461 , w16462 , w16463 , w16464 , w16465 , w16466 , w16467 , w16468 , w16469 , w16470 , w16471 , w16472 , w16473 , w16474 , w16475 , w16476 , w16477 , w16478 , w16479 , w16480 , w16481 , w16482 , w16483 , w16484 , w16485 , w16486 , w16487 , w16488 , w16489 , w16490 , w16491 , w16492 , w16493 , w16494 , w16495 , w16496 , w16497 , w16498 , w16499 , w16500 , w16501 , w16502 , w16503 , w16504 , w16505 , w16506 , w16507 , w16508 , w16509 , w16510 , w16511 , w16512 , w16513 , w16514 , w16515 , w16516 , w16517 , w16518 , w16519 , w16520 , w16521 , w16522 , w16523 , w16524 , w16525 , w16526 , w16527 , w16528 , w16529 , w16530 , w16531 , w16532 , w16533 , w16534 , w16535 , w16536 , w16537 , w16538 , w16539 , w16540 , w16541 , w16542 , w16543 , w16544 , w16545 , w16546 , w16547 , w16548 , w16549 , w16550 , w16551 , w16552 , w16553 , w16554 , w16555 , w16556 , w16557 , w16558 , w16559 , w16560 , w16561 , w16562 , w16563 , w16564 , w16565 , w16566 , w16567 , w16568 , w16569 , w16570 , w16571 , w16572 , w16573 , w16574 , w16575 , w16576 , w16577 , w16578 , w16579 , w16580 , w16581 , w16582 , w16583 , w16584 , w16585 , w16586 , w16587 , w16588 , w16589 , w16590 , w16591 , w16592 , w16593 , w16594 , w16595 , w16596 , w16597 , w16598 , w16599 , w16600 , w16601 , w16602 , w16603 , w16604 , w16605 , w16606 , w16607 , w16608 , w16609 , w16610 , w16611 , w16612 , w16613 , w16614 , w16615 , w16616 , w16617 , w16618 , w16619 , w16620 , w16621 , w16622 , w16623 , w16624 , w16625 , w16626 , w16627 , w16628 , w16629 , w16630 , w16631 , w16632 , w16633 , w16634 , w16635 , w16636 , w16637 , w16638 , w16639 , w16640 , w16641 , w16642 , w16643 , w16644 , w16645 , w16646 , w16647 , w16648 , w16649 , w16650 , w16651 , w16652 , w16653 , w16654 , w16655 , w16656 , w16657 , w16658 , w16659 , w16660 , w16661 , w16662 , w16663 , w16664 , w16665 , w16666 , w16667 , w16668 , w16669 , w16670 , w16671 , w16672 , w16673 , w16674 , w16675 , w16676 , w16677 , w16678 , w16679 , w16680 , w16681 , w16682 , w16683 , w16684 , w16685 , w16686 , w16687 , w16688 , w16689 , w16690 , w16691 , w16692 , w16693 , w16694 , w16695 , w16696 , w16697 , w16698 , w16699 , w16700 , w16701 , w16702 , w16703 , w16704 , w16705 , w16706 , w16707 , w16708 , w16709 , w16710 , w16711 , w16712 , w16713 , w16714 , w16715 , w16716 , w16717 , w16718 , w16719 , w16720 , w16721 , w16722 , w16723 , w16724 , w16725 , w16726 , w16727 , w16728 , w16729 , w16730 , w16731 , w16732 , w16733 , w16734 , w16735 , w16736 , w16737 , w16738 , w16739 , w16740 , w16741 , w16742 , w16743 , w16744 , w16745 , w16746 , w16747 , w16748 , w16749 , w16750 , w16751 , w16752 , w16753 , w16754 , w16755 , w16756 , w16757 , w16758 , w16759 , w16760 , w16761 , w16762 , w16763 , w16764 , w16765 , w16766 , w16767 , w16768 , w16769 , w16770 , w16771 , w16772 , w16773 , w16774 , w16775 , w16776 , w16777 , w16778 , w16779 , w16780 , w16781 , w16782 , w16783 , w16784 , w16785 , w16786 , w16787 , w16788 , w16789 , w16790 , w16791 , w16792 , w16793 , w16794 , w16795 , w16796 , w16797 , w16798 , w16799 , w16800 , w16801 , w16802 , w16803 , w16804 , w16805 , w16806 , w16807 , w16808 , w16809 , w16810 , w16811 , w16812 , w16813 , w16814 , w16815 , w16816 , w16817 , w16818 , w16819 , w16820 , w16821 , w16822 , w16823 , w16824 , w16825 , w16826 , w16827 , w16828 , w16829 , w16830 , w16831 , w16832 , w16833 , w16834 , w16835 , w16836 , w16837 , w16838 , w16839 , w16840 , w16841 , w16842 , w16843 , w16844 , w16845 , w16846 , w16847 , w16848 , w16849 , w16850 , w16851 , w16852 , w16853 , w16854 , w16855 , w16856 , w16857 , w16858 , w16859 , w16860 , w16861 , w16862 , w16863 , w16864 , w16865 , w16866 , w16867 , w16868 , w16869 , w16870 , w16871 , w16872 , w16873 , w16874 , w16875 , w16876 , w16877 , w16878 , w16879 , w16880 , w16881 , w16882 , w16883 , w16884 , w16885 , w16886 , w16887 , w16888 , w16889 , w16890 , w16891 , w16892 , w16893 , w16894 , w16895 , w16896 , w16897 , w16898 , w16899 , w16900 , w16901 , w16902 , w16903 , w16904 , w16905 , w16906 , w16907 , w16908 , w16909 , w16910 , w16911 , w16912 , w16913 , w16914 , w16915 , w16916 , w16917 , w16918 , w16919 , w16920 , w16921 , w16922 , w16923 , w16924 , w16925 , w16926 , w16927 , w16928 , w16929 , w16930 , w16931 , w16932 , w16933 , w16934 , w16935 , w16936 , w16937 , w16938 , w16939 , w16940 , w16941 , w16942 , w16943 , w16944 , w16945 , w16946 , w16947 , w16948 , w16949 , w16950 , w16951 , w16952 , w16953 , w16954 , w16955 , w16956 , w16957 , w16958 , w16959 , w16960 , w16961 , w16962 , w16963 , w16964 , w16965 , w16966 , w16967 , w16968 , w16969 , w16970 , w16971 , w16972 , w16973 , w16974 , w16975 , w16976 , w16977 , w16978 , w16979 , w16980 , w16981 , w16982 , w16983 , w16984 , w16985 , w16986 , w16987 , w16988 , w16989 , w16990 , w16991 , w16992 , w16993 , w16994 , w16995 , w16996 , w16997 , w16998 , w16999 , w17000 , w17001 , w17002 , w17003 , w17004 , w17005 , w17006 , w17007 , w17008 , w17009 , w17010 , w17011 , w17012 , w17013 , w17014 , w17015 , w17016 , w17017 , w17018 , w17019 , w17020 , w17021 , w17022 , w17023 , w17024 , w17025 , w17026 , w17027 , w17028 , w17029 , w17030 , w17031 , w17032 , w17033 , w17034 , w17035 , w17036 , w17037 , w17038 , w17039 , w17040 , w17041 , w17042 , w17043 , w17044 , w17045 , w17046 , w17047 , w17048 , w17049 , w17050 , w17051 , w17052 , w17053 , w17054 , w17055 , w17056 , w17057 , w17058 , w17059 , w17060 , w17061 , w17062 , w17063 , w17064 , w17065 , w17066 , w17067 , w17068 , w17069 , w17070 , w17071 , w17072 , w17073 , w17074 , w17075 , w17076 , w17077 , w17078 , w17079 , w17080 , w17081 , w17082 , w17083 , w17084 , w17085 , w17086 , w17087 , w17088 , w17089 , w17090 , w17091 , w17092 , w17093 , w17094 , w17095 , w17096 , w17097 , w17098 , w17099 , w17100 , w17101 , w17102 , w17103 , w17104 , w17105 , w17106 , w17107 , w17108 , w17109 , w17110 , w17111 , w17112 , w17113 , w17114 , w17115 , w17116 , w17117 , w17118 , w17119 , w17120 , w17121 , w17122 , w17123 , w17124 , w17125 , w17126 , w17127 , w17128 , w17129 , w17130 , w17131 , w17132 , w17133 , w17134 , w17135 , w17136 , w17137 , w17138 , w17139 , w17140 , w17141 , w17142 , w17143 , w17144 , w17145 , w17146 , w17147 , w17148 , w17149 , w17150 , w17151 , w17152 , w17153 , w17154 , w17155 , w17156 , w17157 , w17158 , w17159 , w17160 , w17161 , w17162 , w17163 , w17164 , w17165 , w17166 , w17167 , w17168 , w17169 , w17170 , w17171 , w17172 , w17173 , w17174 , w17175 , w17176 , w17177 , w17178 , w17179 , w17180 , w17181 , w17182 , w17183 , w17184 , w17185 , w17186 , w17187 , w17188 , w17189 , w17190 , w17191 , w17192 , w17193 , w17194 , w17195 , w17196 , w17197 , w17198 , w17199 , w17200 , w17201 , w17202 , w17203 , w17204 , w17205 , w17206 , w17207 , w17208 , w17209 , w17210 , w17211 , w17212 , w17213 , w17214 , w17215 , w17216 , w17217 , w17218 , w17219 , w17220 , w17221 , w17222 , w17223 , w17224 , w17225 , w17226 , w17227 , w17228 , w17229 , w17230 , w17231 , w17232 , w17233 , w17234 , w17235 , w17236 , w17237 , w17238 , w17239 , w17240 , w17241 , w17242 , w17243 , w17244 , w17245 , w17246 , w17247 , w17248 , w17249 , w17250 , w17251 , w17252 , w17253 , w17254 , w17255 , w17256 , w17257 , w17258 , w17259 , w17260 , w17261 , w17262 , w17263 , w17264 , w17265 , w17266 , w17267 , w17268 , w17269 , w17270 , w17271 , w17272 , w17273 , w17274 , w17275 , w17276 , w17277 , w17278 , w17279 , w17280 , w17281 , w17282 , w17283 , w17284 , w17285 , w17286 , w17287 , w17288 , w17289 , w17290 , w17291 , w17292 , w17293 , w17294 , w17295 , w17296 , w17297 , w17298 , w17299 , w17300 , w17301 , w17302 , w17303 , w17304 , w17305 , w17306 , w17307 , w17308 , w17309 , w17310 , w17311 , w17312 , w17313 , w17314 , w17315 , w17316 , w17317 , w17318 , w17319 , w17320 , w17321 , w17322 , w17323 , w17324 , w17325 , w17326 , w17327 , w17328 , w17329 , w17330 , w17331 , w17332 , w17333 , w17334 , w17335 , w17336 , w17337 , w17338 , w17339 , w17340 , w17341 , w17342 , w17343 , w17344 , w17345 , w17346 , w17347 , w17348 , w17349 , w17350 , w17351 , w17352 , w17353 , w17354 , w17355 , w17356 , w17357 , w17358 , w17359 , w17360 , w17361 , w17362 , w17363 , w17364 , w17365 , w17366 , w17367 , w17368 , w17369 , w17370 , w17371 , w17372 , w17373 , w17374 , w17375 , w17376 , w17377 , w17378 , w17379 , w17380 , w17381 , w17382 , w17383 , w17384 , w17385 , w17386 , w17387 , w17388 , w17389 , w17390 , w17391 , w17392 , w17393 , w17394 , w17395 , w17396 , w17397 , w17398 , w17399 , w17400 , w17401 , w17402 , w17403 , w17404 , w17405 , w17406 , w17407 , w17408 , w17409 , w17410 , w17411 , w17412 , w17413 , w17414 , w17415 , w17416 , w17417 , w17418 , w17419 , w17420 , w17421 , w17422 , w17423 , w17424 , w17425 , w17426 , w17427 , w17428 , w17429 , w17430 , w17431 , w17432 , w17433 , w17434 , w17435 , w17436 , w17437 , w17438 , w17439 , w17440 , w17441 , w17442 , w17443 , w17444 , w17445 , w17446 , w17447 , w17448 , w17449 , w17450 , w17451 , w17452 , w17453 , w17454 , w17455 , w17456 , w17457 , w17458 , w17459 , w17460 , w17461 , w17462 , w17463 , w17464 , w17465 , w17466 , w17467 , w17468 , w17469 , w17470 , w17471 , w17472 , w17473 , w17474 , w17475 , w17476 , w17477 , w17478 , w17479 , w17480 , w17481 , w17482 , w17483 , w17484 , w17485 , w17486 , w17487 , w17488 , w17489 , w17490 , w17491 , w17492 , w17493 , w17494 , w17495 , w17496 , w17497 ;
  assign zero = 0;
  assign w129 = \pi126 | \pi127 ;
  assign w130 = \pi124 | \pi125 ;
  assign w131 = \pi126 ^ \pi127 ;
  assign w132 = ( \pi127 & w130 ) | ( \pi127 & ~w131 ) | ( w130 & ~w131 ) ;
  assign w133 = \pi122 | \pi123 ;
  assign w134 = ( \pi124 & ~\pi125 ) | ( \pi124 & \pi127 ) | ( ~\pi125 & \pi127 ) ;
  assign w135 = ( \pi124 & ~\pi127 ) | ( \pi124 & w133 ) | ( ~\pi127 & w133 ) ;
  assign w136 = ~\pi126 & w135 ;
  assign w137 = ~w134 & w136 ;
  assign w138 = \pi125 ^ w132 ;
  assign w139 = ~\pi124 & w133 ;
  assign w140 = \pi124 & ~w132 ;
  assign w141 = ( w138 & w139 ) | ( w138 & w140 ) | ( w139 & w140 ) ;
  assign w142 = \pi126 ^ w130 ;
  assign w143 = \pi127 & ~w142 ;
  assign w144 = ( ~w137 & w141 ) | ( ~w137 & w143 ) | ( w141 & w143 ) ;
  assign w145 = w137 | w144 ;
  assign w146 = \pi120 | \pi121 ;
  assign w147 = \pi126 | w130 ;
  assign w148 = \pi122 | w146 ;
  assign w149 = \pi126 & ~\pi127 ;
  assign w150 = ( ~w147 & w148 ) | ( ~w147 & w149 ) | ( w148 & w149 ) ;
  assign w151 = \pi122 & \pi123 ;
  assign w152 = ~w132 & w151 ;
  assign w153 = ( \pi122 & w150 ) | ( \pi122 & w151 ) | ( w150 & w151 ) ;
  assign w154 = ( ~w145 & w152 ) | ( ~w145 & w153 ) | ( w152 & w153 ) ;
  assign w155 = w132 & ~w146 ;
  assign w156 = \pi123 ^ w145 ;
  assign w157 = ( \pi123 & ~w145 ) | ( \pi123 & w150 ) | ( ~w145 & w150 ) ;
  assign w158 = ( ~\pi122 & w156 ) | ( ~\pi122 & w157 ) | ( w156 & w157 ) ;
  assign w159 = w155 | w158 ;
  assign w160 = ( w154 & ~w155 ) | ( w154 & w159 ) | ( ~w155 & w159 ) ;
  assign w161 = \pi124 & ~w133 ;
  assign w162 = ( \pi125 & ~\pi126 ) | ( \pi125 & w161 ) | ( ~\pi126 & w161 ) ;
  assign w163 = ( \pi124 & \pi126 ) | ( \pi124 & w162 ) | ( \pi126 & w162 ) ;
  assign w164 = ( \pi127 & ~w133 ) | ( \pi127 & w162 ) | ( ~w133 & w162 ) ;
  assign w165 = w163 ^ w164 ;
  assign w166 = ( \pi125 & \pi126 ) | ( \pi125 & ~w160 ) | ( \pi126 & ~w160 ) ;
  assign w167 = \pi124 ^ w133 ;
  assign w168 = ( \pi126 & w166 ) | ( \pi126 & ~w167 ) | ( w166 & ~w167 ) ;
  assign w169 = ( ~\pi127 & w160 ) | ( ~\pi127 & w168 ) | ( w160 & w168 ) ;
  assign w170 = ~\pi126 & w169 ;
  assign w171 = ( \pi125 & ~\pi126 ) | ( \pi125 & \pi127 ) | ( ~\pi126 & \pi127 ) ;
  assign w172 = ( \pi124 & \pi126 ) | ( \pi124 & \pi127 ) | ( \pi126 & \pi127 ) ;
  assign w173 = \pi125 ^ w172 ;
  assign w174 = \pi124 | w133 ;
  assign w175 = ( w171 & w173 ) | ( w171 & ~w174 ) | ( w173 & ~w174 ) ;
  assign w176 = w171 ^ w175 ;
  assign w177 = ( \pi125 & \pi126 ) | ( \pi125 & \pi127 ) | ( \pi126 & \pi127 ) ;
  assign w178 = ( \pi125 & \pi127 ) | ( \pi125 & w133 ) | ( \pi127 & w133 ) ;
  assign w179 = ( \pi124 & \pi126 ) | ( \pi124 & w178 ) | ( \pi126 & w178 ) ;
  assign w180 = \pi126 ^ w179 ;
  assign w181 = w177 & w180 ;
  assign w182 = w170 | w176 ;
  assign w183 = ( w160 & w165 ) | ( w160 & w182 ) | ( w165 & w182 ) ;
  assign w184 = ( w181 & ~w182 ) | ( w181 & w183 ) | ( ~w182 & w183 ) ;
  assign w185 = w182 | w184 ;
  assign w186 = \pi118 | \pi119 ;
  assign w187 = ( \pi120 & w145 ) | ( \pi120 & ~w186 ) | ( w145 & ~w186 ) ;
  assign w188 = ( ~\pi120 & w145 ) | ( ~\pi120 & w185 ) | ( w145 & w185 ) ;
  assign w189 = w187 & w188 ;
  assign w190 = \pi120 & ~w185 ;
  assign w191 = ( ~\pi120 & w141 ) | ( ~\pi120 & w186 ) | ( w141 & w186 ) ;
  assign w192 = ( w137 & ~w141 ) | ( w137 & w143 ) | ( ~w141 & w143 ) ;
  assign w193 = ( w190 & w191 ) | ( w190 & ~w192 ) | ( w191 & ~w192 ) ;
  assign w194 = ~w141 & w193 ;
  assign w195 = ~\pi120 & w185 ;
  assign w196 = \pi121 ^ w195 ;
  assign w197 = w194 | w196 ;
  assign w198 = ( \pi124 & \pi125 ) | ( \pi124 & \pi127 ) | ( \pi125 & \pi127 ) ;
  assign w199 = ( \pi127 & w133 ) | ( \pi127 & w198 ) | ( w133 & w198 ) ;
  assign w200 = \pi126 | w160 ;
  assign w201 = ( ~\pi124 & \pi127 ) | ( ~\pi124 & w133 ) | ( \pi127 & w133 ) ;
  assign w202 = ( w198 & ~w200 ) | ( w198 & w201 ) | ( ~w200 & w201 ) ;
  assign w203 = ~w199 & w202 ;
  assign w204 = \pi125 ^ \pi127 ;
  assign w205 = ( ~\pi124 & w133 ) | ( ~\pi124 & w204 ) | ( w133 & w204 ) ;
  assign w206 = ( ~\pi124 & w160 ) | ( ~\pi124 & w205 ) | ( w160 & w205 ) ;
  assign w207 = ~\pi124 & w178 ;
  assign w208 = ( w204 & ~w206 ) | ( w204 & w207 ) | ( ~w206 & w207 ) ;
  assign w209 = ( \pi126 & w203 ) | ( \pi126 & w208 ) | ( w203 & w208 ) ;
  assign w210 = w203 | w209 ;
  assign w211 = w146 & w185 ;
  assign w212 = ( w185 & w210 ) | ( w185 & ~w211 ) | ( w210 & ~w211 ) ;
  assign w213 = \pi122 ^ w212 ;
  assign w214 = ~w189 & w197 ;
  assign w215 = ( ~w132 & w213 ) | ( ~w132 & w214 ) | ( w213 & w214 ) ;
  assign w216 = w145 | w150 ;
  assign w217 = ( \pi122 & w145 ) | ( \pi122 & ~w150 ) | ( w145 & ~w150 ) ;
  assign w218 = ( \pi122 & w132 ) | ( \pi122 & ~w148 ) | ( w132 & ~w148 ) ;
  assign w219 = ( w216 & ~w217 ) | ( w216 & w218 ) | ( ~w217 & w218 ) ;
  assign w220 = w185 & ~w219 ;
  assign w221 = ~\pi122 & w145 ;
  assign w222 = \pi123 ^ w221 ;
  assign w223 = w220 ^ w222 ;
  assign w224 = ( w160 & w165 ) | ( w160 & w215 ) | ( w165 & w215 ) ;
  assign w225 = ~w129 & w224 ;
  assign w226 = w160 ^ w165 ;
  assign w227 = ( w185 & w215 ) | ( w185 & ~w226 ) | ( w215 & ~w226 ) ;
  assign w228 = ( ~w129 & w223 ) | ( ~w129 & w227 ) | ( w223 & w227 ) ;
  assign w229 = ( ~w129 & w225 ) | ( ~w129 & w228 ) | ( w225 & w228 ) ;
  assign w230 = ( w189 & ~w197 ) | ( w189 & w223 ) | ( ~w197 & w223 ) ;
  assign w231 = ( w132 & ~w213 ) | ( w132 & w230 ) | ( ~w213 & w230 ) ;
  assign w232 = w223 & ~w231 ;
  assign w233 = ( w129 & w160 ) | ( w129 & w165 ) | ( w160 & w165 ) ;
  assign w234 = ( w165 & ~w185 ) | ( w165 & w233 ) | ( ~w185 & w233 ) ;
  assign w235 = w160 & w234 ;
  assign w236 = w233 ^ w235 ;
  assign w237 = ( \pi124 & ~\pi126 ) | ( \pi124 & \pi127 ) | ( ~\pi126 & \pi127 ) ;
  assign w238 = ( \pi125 & ~w133 ) | ( \pi125 & w237 ) | ( ~w133 & w237 ) ;
  assign w239 = \pi126 & ~w238 ;
  assign w240 = ( \pi124 & ~w160 ) | ( \pi124 & w238 ) | ( ~w160 & w238 ) ;
  assign w241 = ~\pi124 & \pi127 ;
  assign w242 = w240 & w241 ;
  assign w243 = ( w239 & w240 ) | ( w239 & w242 ) | ( w240 & w242 ) ;
  assign w244 = w232 | w243 ;
  assign w245 = ( w229 & ~w232 ) | ( w229 & w236 ) | ( ~w232 & w236 ) ;
  assign w246 = w244 | w245 ;
  assign w247 = ( \pi116 & ~\pi117 ) | ( \pi116 & \pi118 ) | ( ~\pi117 & \pi118 ) ;
  assign w248 = \pi117 | w247 ;
  assign w249 = \pi118 & w246 ;
  assign w250 = w248 | w249 ;
  assign w251 = ( w185 & w249 ) | ( w185 & ~w250 ) | ( w249 & ~w250 ) ;
  assign w252 = ( w160 & w165 ) | ( w160 & w170 ) | ( w165 & w170 ) ;
  assign w253 = ( ~w170 & w248 ) | ( ~w170 & w252 ) | ( w248 & w252 ) ;
  assign w254 = ( w176 & w181 ) | ( w176 & ~w252 ) | ( w181 & ~w252 ) ;
  assign w255 = ( w252 & w253 ) | ( w252 & w254 ) | ( w253 & w254 ) ;
  assign w256 = w253 & ~w255 ;
  assign w257 = ( \pi119 & ~w246 ) | ( \pi119 & w256 ) | ( ~w246 & w256 ) ;
  assign w258 = \pi118 ^ \pi119 ;
  assign w259 = w246 & ~w258 ;
  assign w260 = w257 | w259 ;
  assign w261 = ( w145 & w251 ) | ( w145 & ~w260 ) | ( w251 & ~w260 ) ;
  assign w262 = w145 & w261 ;
  assign w263 = ( w145 & w251 ) | ( w145 & w260 ) | ( w251 & w260 ) ;
  assign w264 = w260 & ~w263 ;
  assign w265 = w185 & ~w243 ;
  assign w266 = ~w232 & w265 ;
  assign w267 = ~w245 & w266 ;
  assign w268 = w186 & w246 ;
  assign w269 = ( w246 & w267 ) | ( w246 & ~w268 ) | ( w267 & ~w268 ) ;
  assign w270 = \pi120 ^ w269 ;
  assign w271 = w264 | w270 ;
  assign w272 = ( w132 & w262 ) | ( w132 & ~w271 ) | ( w262 & ~w271 ) ;
  assign w273 = w132 & w272 ;
  assign w274 = ( ~w132 & w262 ) | ( ~w132 & w271 ) | ( w262 & w271 ) ;
  assign w275 = ~w262 & w274 ;
  assign w276 = ( w189 & ~w194 ) | ( w189 & w246 ) | ( ~w194 & w246 ) ;
  assign w277 = ~w189 & w276 ;
  assign w278 = \pi121 ^ w277 ;
  assign w279 = w195 ^ w278 ;
  assign w280 = w275 | w279 ;
  assign w281 = ~w273 & w280 ;
  assign w282 = ( w189 & ~w197 ) | ( w189 & w246 ) | ( ~w197 & w246 ) ;
  assign w283 = w132 ^ w282 ;
  assign w284 = w246 & w283 ;
  assign w285 = w213 ^ w284 ;
  assign w286 = w215 & ~w223 ;
  assign w287 = w232 | w285 ;
  assign w288 = ( ~w223 & w246 ) | ( ~w223 & w286 ) | ( w246 & w286 ) ;
  assign w289 = ( ~w286 & w287 ) | ( ~w286 & w288 ) | ( w287 & w288 ) ;
  assign w290 = ( ~w129 & w281 ) | ( ~w129 & w289 ) | ( w281 & w289 ) ;
  assign w291 = ~w129 & w290 ;
  assign w292 = ( w273 & w280 ) | ( w273 & w285 ) | ( w280 & w285 ) ;
  assign w293 = ~w273 & w292 ;
  assign w294 = w129 & ~w232 ;
  assign w295 = ( w215 & w223 ) | ( w215 & w246 ) | ( w223 & w246 ) ;
  assign w296 = ( w223 & w294 ) | ( w223 & w295 ) | ( w294 & w295 ) ;
  assign w297 = w294 & w296 ;
  assign w298 = ( w185 & ~w219 ) | ( w185 & w243 ) | ( ~w219 & w243 ) ;
  assign w299 = ( ~\pi122 & w145 ) | ( ~\pi122 & w243 ) | ( w145 & w243 ) ;
  assign w300 = w298 ^ w299 ;
  assign w301 = \pi123 ^ w300 ;
  assign w302 = ~w243 & w301 ;
  assign w303 = ~w232 & w302 ;
  assign w304 = ~w245 & w303 ;
  assign w305 = w293 | w304 ;
  assign w306 = ( w291 & ~w293 ) | ( w291 & w297 ) | ( ~w293 & w297 ) ;
  assign w307 = w305 | w306 ;
  assign w308 = ( ~\pi115 & \pi116 ) | ( ~\pi115 & w246 ) | ( \pi116 & w246 ) ;
  assign w309 = ( ~\pi114 & \pi116 ) | ( ~\pi114 & w308 ) | ( \pi116 & w308 ) ;
  assign w310 = ( ~\pi116 & w246 ) | ( ~\pi116 & w307 ) | ( w246 & w307 ) ;
  assign w311 = w309 & w310 ;
  assign w312 = ( w232 & w236 ) | ( w232 & ~w243 ) | ( w236 & ~w243 ) ;
  assign w313 = \pi115 & ~w312 ;
  assign w314 = \pi114 | \pi116 ;
  assign w315 = ( ~w312 & w313 ) | ( ~w312 & w314 ) | ( w313 & w314 ) ;
  assign w316 = ~w243 & w315 ;
  assign w317 = ~w229 & w316 ;
  assign w318 = ( \pi116 & w307 ) | ( \pi116 & ~w316 ) | ( w307 & ~w316 ) ;
  assign w319 = w317 & ~w318 ;
  assign w320 = ~\pi116 & w307 ;
  assign w321 = \pi117 ^ w320 ;
  assign w322 = w319 | w321 ;
  assign w323 = ( w185 & w311 ) | ( w185 & ~w322 ) | ( w311 & ~w322 ) ;
  assign w324 = w185 & w323 ;
  assign w325 = ( ~w185 & w311 ) | ( ~w185 & w322 ) | ( w311 & w322 ) ;
  assign w326 = ~w311 & w325 ;
  assign w327 = w246 & ~w304 ;
  assign w328 = ~w293 & w327 ;
  assign w329 = ~w306 & w328 ;
  assign w330 = \pi117 & w307 ;
  assign w331 = ( \pi116 & w307 ) | ( \pi116 & ~w330 ) | ( w307 & ~w330 ) ;
  assign w332 = ( ~\pi116 & w329 ) | ( ~\pi116 & w331 ) | ( w329 & w331 ) ;
  assign w333 = \pi118 ^ w332 ;
  assign w334 = w326 | w333 ;
  assign w335 = ( w145 & w324 ) | ( w145 & ~w334 ) | ( w324 & ~w334 ) ;
  assign w336 = w145 & w335 ;
  assign w337 = ~\pi118 & w246 ;
  assign w338 = \pi119 ^ w337 ;
  assign w339 = ( ~w246 & w256 ) | ( ~w246 & w337 ) | ( w256 & w337 ) ;
  assign w340 = ~w251 & w307 ;
  assign w341 = ~w339 & w340 ;
  assign w342 = w338 ^ w341 ;
  assign w343 = ( ~w145 & w324 ) | ( ~w145 & w334 ) | ( w324 & w334 ) ;
  assign w344 = ~w324 & w343 ;
  assign w345 = w342 | w344 ;
  assign w346 = ( w132 & w336 ) | ( w132 & ~w345 ) | ( w336 & ~w345 ) ;
  assign w347 = w132 & w346 ;
  assign w348 = w262 | w264 ;
  assign w349 = w307 & ~w348 ;
  assign w350 = w270 ^ w349 ;
  assign w351 = ( ~w132 & w336 ) | ( ~w132 & w345 ) | ( w336 & w345 ) ;
  assign w352 = ~w336 & w351 ;
  assign w353 = w350 | w352 ;
  assign w354 = ~w347 & w353 ;
  assign w355 = w273 | w275 ;
  assign w356 = w307 & ~w355 ;
  assign w357 = w279 ^ w356 ;
  assign w358 = ( ~w293 & w354 ) | ( ~w293 & w357 ) | ( w354 & w357 ) ;
  assign w359 = w281 & ~w358 ;
  assign w360 = ~w285 & w307 ;
  assign w361 = ( w358 & ~w359 ) | ( w358 & w360 ) | ( ~w359 & w360 ) ;
  assign w362 = w293 | w361 ;
  assign w363 = ~w129 & w362 ;
  assign w364 = ( w347 & w353 ) | ( w347 & w357 ) | ( w353 & w357 ) ;
  assign w365 = ~w347 & w364 ;
  assign w366 = ( w129 & w281 ) | ( w129 & w285 ) | ( w281 & w285 ) ;
  assign w367 = ( w285 & ~w307 ) | ( w285 & w366 ) | ( ~w307 & w366 ) ;
  assign w368 = w281 & w367 ;
  assign w369 = w366 ^ w368 ;
  assign w370 = ( w246 & w283 ) | ( w246 & w304 ) | ( w283 & w304 ) ;
  assign w371 = w213 ^ w370 ;
  assign w372 = ~w304 & w371 ;
  assign w373 = ~w293 & w372 ;
  assign w374 = ~w306 & w373 ;
  assign w375 = w365 | w374 ;
  assign w376 = ( w363 & ~w365 ) | ( w363 & w369 ) | ( ~w365 & w369 ) ;
  assign w377 = w375 | w376 ;
  assign w378 = ( ~\pi113 & \pi114 ) | ( ~\pi113 & w307 ) | ( \pi114 & w307 ) ;
  assign w379 = ( ~\pi112 & \pi114 ) | ( ~\pi112 & w378 ) | ( \pi114 & w378 ) ;
  assign w380 = ( ~\pi114 & w307 ) | ( ~\pi114 & w377 ) | ( w307 & w377 ) ;
  assign w381 = w379 & w380 ;
  assign w382 = ( w293 & w297 ) | ( w293 & ~w304 ) | ( w297 & ~w304 ) ;
  assign w383 = \pi113 & ~w382 ;
  assign w384 = \pi112 | \pi114 ;
  assign w385 = ( ~w382 & w383 ) | ( ~w382 & w384 ) | ( w383 & w384 ) ;
  assign w386 = ~w304 & w385 ;
  assign w387 = ~w291 & w386 ;
  assign w388 = ( \pi114 & w377 ) | ( \pi114 & ~w386 ) | ( w377 & ~w386 ) ;
  assign w389 = w387 & ~w388 ;
  assign w390 = ~\pi114 & w377 ;
  assign w391 = \pi115 ^ w390 ;
  assign w392 = w389 | w391 ;
  assign w393 = ( w246 & w381 ) | ( w246 & ~w392 ) | ( w381 & ~w392 ) ;
  assign w394 = w246 & w393 ;
  assign w395 = ( ~w246 & w381 ) | ( ~w246 & w392 ) | ( w381 & w392 ) ;
  assign w396 = ~w381 & w395 ;
  assign w397 = w307 & ~w374 ;
  assign w398 = ~w365 & w397 ;
  assign w399 = ~w376 & w398 ;
  assign w400 = \pi115 & w377 ;
  assign w401 = ( \pi114 & w377 ) | ( \pi114 & ~w400 ) | ( w377 & ~w400 ) ;
  assign w402 = ( ~\pi114 & w399 ) | ( ~\pi114 & w401 ) | ( w399 & w401 ) ;
  assign w403 = \pi116 ^ w402 ;
  assign w404 = w396 | w403 ;
  assign w405 = ( w185 & w394 ) | ( w185 & ~w404 ) | ( w394 & ~w404 ) ;
  assign w406 = w185 & w405 ;
  assign w407 = ( w311 & ~w319 ) | ( w311 & w377 ) | ( ~w319 & w377 ) ;
  assign w408 = ~w311 & w407 ;
  assign w409 = \pi117 ^ w408 ;
  assign w410 = w320 ^ w409 ;
  assign w411 = ( ~w185 & w394 ) | ( ~w185 & w404 ) | ( w394 & w404 ) ;
  assign w412 = ~w394 & w411 ;
  assign w413 = w410 | w412 ;
  assign w414 = ( w145 & w406 ) | ( w145 & ~w413 ) | ( w406 & ~w413 ) ;
  assign w415 = w145 & w414 ;
  assign w416 = w324 | w326 ;
  assign w417 = w377 & ~w416 ;
  assign w418 = w333 ^ w417 ;
  assign w419 = ( ~w145 & w406 ) | ( ~w145 & w413 ) | ( w406 & w413 ) ;
  assign w420 = ~w406 & w419 ;
  assign w421 = w418 | w420 ;
  assign w422 = ( w132 & w415 ) | ( w132 & ~w421 ) | ( w415 & ~w421 ) ;
  assign w423 = w132 & w422 ;
  assign w424 = w336 | w344 ;
  assign w425 = w377 & ~w424 ;
  assign w426 = w342 ^ w425 ;
  assign w427 = ( ~w132 & w415 ) | ( ~w132 & w421 ) | ( w415 & w421 ) ;
  assign w428 = ~w415 & w427 ;
  assign w429 = w426 | w428 ;
  assign w430 = ~w423 & w429 ;
  assign w431 = w347 | w352 ;
  assign w432 = w377 & ~w431 ;
  assign w433 = w350 ^ w432 ;
  assign w434 = ( ~w365 & w430 ) | ( ~w365 & w433 ) | ( w430 & w433 ) ;
  assign w435 = w354 & ~w434 ;
  assign w436 = ~w357 & w377 ;
  assign w437 = ( w434 & ~w435 ) | ( w434 & w436 ) | ( ~w435 & w436 ) ;
  assign w438 = w365 | w437 ;
  assign w439 = ~w129 & w438 ;
  assign w440 = ( w423 & w429 ) | ( w423 & w433 ) | ( w429 & w433 ) ;
  assign w441 = ~w423 & w440 ;
  assign w442 = ( w129 & w354 ) | ( w129 & w357 ) | ( w354 & w357 ) ;
  assign w443 = ( w357 & ~w377 ) | ( w357 & w442 ) | ( ~w377 & w442 ) ;
  assign w444 = w354 & w443 ;
  assign w445 = w442 ^ w444 ;
  assign w446 = ( w273 & w275 ) | ( w273 & w307 ) | ( w275 & w307 ) ;
  assign w447 = w307 & ~w446 ;
  assign w448 = w279 ^ w447 ;
  assign w449 = ( ~w369 & w374 ) | ( ~w369 & w448 ) | ( w374 & w448 ) ;
  assign w450 = ~w374 & w449 ;
  assign w451 = ( ~w363 & w365 ) | ( ~w363 & w450 ) | ( w365 & w450 ) ;
  assign w452 = ~w365 & w451 ;
  assign w453 = w441 | w452 ;
  assign w454 = ( w439 & ~w441 ) | ( w439 & w445 ) | ( ~w441 & w445 ) ;
  assign w455 = w453 | w454 ;
  assign w456 = ( ~\pi111 & \pi112 ) | ( ~\pi111 & w377 ) | ( \pi112 & w377 ) ;
  assign w457 = ( ~\pi110 & \pi112 ) | ( ~\pi110 & w456 ) | ( \pi112 & w456 ) ;
  assign w458 = ( ~\pi112 & w377 ) | ( ~\pi112 & w455 ) | ( w377 & w455 ) ;
  assign w459 = w457 & w458 ;
  assign w460 = ( w365 & w369 ) | ( w365 & ~w374 ) | ( w369 & ~w374 ) ;
  assign w461 = \pi111 & ~w460 ;
  assign w462 = \pi110 | \pi112 ;
  assign w463 = ( ~w460 & w461 ) | ( ~w460 & w462 ) | ( w461 & w462 ) ;
  assign w464 = ~w374 & w463 ;
  assign w465 = ~w363 & w464 ;
  assign w466 = ( \pi112 & w455 ) | ( \pi112 & ~w464 ) | ( w455 & ~w464 ) ;
  assign w467 = w465 & ~w466 ;
  assign w468 = ~\pi112 & w455 ;
  assign w469 = \pi113 ^ w468 ;
  assign w470 = w467 | w469 ;
  assign w471 = ( w307 & w459 ) | ( w307 & ~w470 ) | ( w459 & ~w470 ) ;
  assign w472 = w307 & w471 ;
  assign w473 = ( ~w307 & w459 ) | ( ~w307 & w470 ) | ( w459 & w470 ) ;
  assign w474 = ~w459 & w473 ;
  assign w475 = w377 & ~w452 ;
  assign w476 = ~w441 & w475 ;
  assign w477 = ~w454 & w476 ;
  assign w478 = \pi113 & w455 ;
  assign w479 = ( \pi112 & w455 ) | ( \pi112 & ~w478 ) | ( w455 & ~w478 ) ;
  assign w480 = ( ~\pi112 & w477 ) | ( ~\pi112 & w479 ) | ( w477 & w479 ) ;
  assign w481 = \pi114 ^ w480 ;
  assign w482 = w474 | w481 ;
  assign w483 = ( w246 & w472 ) | ( w246 & ~w482 ) | ( w472 & ~w482 ) ;
  assign w484 = w246 & w483 ;
  assign w485 = ( w381 & ~w389 ) | ( w381 & w455 ) | ( ~w389 & w455 ) ;
  assign w486 = ~w381 & w485 ;
  assign w487 = \pi115 ^ w486 ;
  assign w488 = w390 ^ w487 ;
  assign w489 = ( ~w246 & w472 ) | ( ~w246 & w482 ) | ( w472 & w482 ) ;
  assign w490 = ~w472 & w489 ;
  assign w491 = w488 | w490 ;
  assign w492 = ( w185 & w484 ) | ( w185 & ~w491 ) | ( w484 & ~w491 ) ;
  assign w493 = w185 & w492 ;
  assign w494 = w394 | w396 ;
  assign w495 = w455 & ~w494 ;
  assign w496 = w403 ^ w495 ;
  assign w497 = ( ~w185 & w484 ) | ( ~w185 & w491 ) | ( w484 & w491 ) ;
  assign w498 = ~w484 & w497 ;
  assign w499 = w496 | w498 ;
  assign w500 = ( w145 & w493 ) | ( w145 & ~w499 ) | ( w493 & ~w499 ) ;
  assign w501 = w145 & w500 ;
  assign w502 = w406 | w412 ;
  assign w503 = w455 & ~w502 ;
  assign w504 = w410 ^ w503 ;
  assign w505 = ( ~w145 & w493 ) | ( ~w145 & w499 ) | ( w493 & w499 ) ;
  assign w506 = ~w493 & w505 ;
  assign w507 = w504 | w506 ;
  assign w508 = ( w132 & w501 ) | ( w132 & ~w507 ) | ( w501 & ~w507 ) ;
  assign w509 = w132 & w508 ;
  assign w510 = w415 | w420 ;
  assign w511 = w455 & ~w510 ;
  assign w512 = w418 ^ w511 ;
  assign w513 = ( ~w132 & w501 ) | ( ~w132 & w507 ) | ( w501 & w507 ) ;
  assign w514 = ~w501 & w513 ;
  assign w515 = w512 | w514 ;
  assign w516 = ~w509 & w515 ;
  assign w517 = w423 | w428 ;
  assign w518 = w455 & ~w517 ;
  assign w519 = w426 ^ w518 ;
  assign w520 = ( ~w441 & w516 ) | ( ~w441 & w519 ) | ( w516 & w519 ) ;
  assign w521 = w430 & ~w520 ;
  assign w522 = ~w433 & w455 ;
  assign w523 = ( w520 & ~w521 ) | ( w520 & w522 ) | ( ~w521 & w522 ) ;
  assign w524 = w441 | w523 ;
  assign w525 = ~w129 & w524 ;
  assign w526 = ( w509 & w515 ) | ( w509 & w519 ) | ( w515 & w519 ) ;
  assign w527 = ~w509 & w526 ;
  assign w528 = ( w129 & w430 ) | ( w129 & w433 ) | ( w430 & w433 ) ;
  assign w529 = ( w433 & ~w455 ) | ( w433 & w528 ) | ( ~w455 & w528 ) ;
  assign w530 = w430 & w529 ;
  assign w531 = w528 ^ w530 ;
  assign w532 = ( w347 & w352 ) | ( w347 & w377 ) | ( w352 & w377 ) ;
  assign w533 = w377 & ~w532 ;
  assign w534 = w350 ^ w533 ;
  assign w535 = ( ~w445 & w452 ) | ( ~w445 & w534 ) | ( w452 & w534 ) ;
  assign w536 = ~w452 & w535 ;
  assign w537 = ( ~w439 & w441 ) | ( ~w439 & w536 ) | ( w441 & w536 ) ;
  assign w538 = ~w441 & w537 ;
  assign w539 = w527 | w538 ;
  assign w540 = ( w525 & ~w527 ) | ( w525 & w531 ) | ( ~w527 & w531 ) ;
  assign w541 = w539 | w540 ;
  assign w542 = ( ~\pi109 & \pi110 ) | ( ~\pi109 & w455 ) | ( \pi110 & w455 ) ;
  assign w543 = ( ~\pi108 & \pi110 ) | ( ~\pi108 & w542 ) | ( \pi110 & w542 ) ;
  assign w544 = ( ~\pi110 & w455 ) | ( ~\pi110 & w541 ) | ( w455 & w541 ) ;
  assign w545 = w543 & w544 ;
  assign w546 = ( w441 & w445 ) | ( w441 & ~w452 ) | ( w445 & ~w452 ) ;
  assign w547 = \pi109 & ~w546 ;
  assign w548 = \pi108 | \pi110 ;
  assign w549 = ( ~w546 & w547 ) | ( ~w546 & w548 ) | ( w547 & w548 ) ;
  assign w550 = ~w452 & w549 ;
  assign w551 = ~w439 & w550 ;
  assign w552 = ( \pi110 & w541 ) | ( \pi110 & ~w550 ) | ( w541 & ~w550 ) ;
  assign w553 = w551 & ~w552 ;
  assign w554 = ~\pi110 & w541 ;
  assign w555 = \pi111 ^ w554 ;
  assign w556 = w553 | w555 ;
  assign w557 = ( w377 & w545 ) | ( w377 & ~w556 ) | ( w545 & ~w556 ) ;
  assign w558 = w377 & w557 ;
  assign w559 = ( ~w377 & w545 ) | ( ~w377 & w556 ) | ( w545 & w556 ) ;
  assign w560 = ~w545 & w559 ;
  assign w561 = w455 & ~w538 ;
  assign w562 = ~w527 & w561 ;
  assign w563 = ~w540 & w562 ;
  assign w564 = \pi111 & w541 ;
  assign w565 = ( \pi110 & w541 ) | ( \pi110 & ~w564 ) | ( w541 & ~w564 ) ;
  assign w566 = ( ~\pi110 & w563 ) | ( ~\pi110 & w565 ) | ( w563 & w565 ) ;
  assign w567 = \pi112 ^ w566 ;
  assign w568 = w560 | w567 ;
  assign w569 = ( w307 & w558 ) | ( w307 & ~w568 ) | ( w558 & ~w568 ) ;
  assign w570 = w307 & w569 ;
  assign w571 = ( ~w307 & w558 ) | ( ~w307 & w568 ) | ( w558 & w568 ) ;
  assign w572 = ~w558 & w571 ;
  assign w573 = ( w459 & ~w467 ) | ( w459 & w541 ) | ( ~w467 & w541 ) ;
  assign w574 = ~w459 & w573 ;
  assign w575 = \pi113 ^ w574 ;
  assign w576 = w468 ^ w575 ;
  assign w577 = w572 | w576 ;
  assign w578 = ( w246 & w570 ) | ( w246 & ~w577 ) | ( w570 & ~w577 ) ;
  assign w579 = w246 & w578 ;
  assign w580 = w472 | w474 ;
  assign w581 = w541 & ~w580 ;
  assign w582 = w481 ^ w581 ;
  assign w583 = ( ~w246 & w570 ) | ( ~w246 & w577 ) | ( w570 & w577 ) ;
  assign w584 = ~w570 & w583 ;
  assign w585 = w582 | w584 ;
  assign w586 = ( w185 & w579 ) | ( w185 & ~w585 ) | ( w579 & ~w585 ) ;
  assign w587 = w185 & w586 ;
  assign w588 = w484 | w490 ;
  assign w589 = w541 & ~w588 ;
  assign w590 = w488 ^ w589 ;
  assign w591 = ( ~w185 & w579 ) | ( ~w185 & w585 ) | ( w579 & w585 ) ;
  assign w592 = ~w579 & w591 ;
  assign w593 = w590 | w592 ;
  assign w594 = ( w145 & w587 ) | ( w145 & ~w593 ) | ( w587 & ~w593 ) ;
  assign w595 = w145 & w594 ;
  assign w596 = w493 | w498 ;
  assign w597 = w541 & ~w596 ;
  assign w598 = w496 ^ w597 ;
  assign w599 = ( ~w145 & w587 ) | ( ~w145 & w593 ) | ( w587 & w593 ) ;
  assign w600 = ~w587 & w599 ;
  assign w601 = w598 | w600 ;
  assign w602 = ( w132 & w595 ) | ( w132 & ~w601 ) | ( w595 & ~w601 ) ;
  assign w603 = w132 & w602 ;
  assign w604 = w501 | w506 ;
  assign w605 = w541 & ~w604 ;
  assign w606 = w504 ^ w605 ;
  assign w607 = ( ~w132 & w595 ) | ( ~w132 & w601 ) | ( w595 & w601 ) ;
  assign w608 = ~w595 & w607 ;
  assign w609 = w606 | w608 ;
  assign w610 = ~w603 & w609 ;
  assign w611 = w509 | w514 ;
  assign w612 = w541 & ~w611 ;
  assign w613 = w512 ^ w612 ;
  assign w614 = ( ~w527 & w610 ) | ( ~w527 & w613 ) | ( w610 & w613 ) ;
  assign w615 = w516 & ~w614 ;
  assign w616 = ~w519 & w541 ;
  assign w617 = ( w614 & ~w615 ) | ( w614 & w616 ) | ( ~w615 & w616 ) ;
  assign w618 = w527 | w617 ;
  assign w619 = ~w129 & w618 ;
  assign w620 = ( w603 & w609 ) | ( w603 & w613 ) | ( w609 & w613 ) ;
  assign w621 = ~w603 & w620 ;
  assign w622 = ( w129 & w516 ) | ( w129 & w519 ) | ( w516 & w519 ) ;
  assign w623 = ( w519 & ~w541 ) | ( w519 & w622 ) | ( ~w541 & w622 ) ;
  assign w624 = w516 & w623 ;
  assign w625 = w622 ^ w624 ;
  assign w626 = ( w423 & w428 ) | ( w423 & w455 ) | ( w428 & w455 ) ;
  assign w627 = w455 & ~w626 ;
  assign w628 = w426 ^ w627 ;
  assign w629 = ( ~w531 & w538 ) | ( ~w531 & w628 ) | ( w538 & w628 ) ;
  assign w630 = ~w538 & w629 ;
  assign w631 = ( ~w525 & w527 ) | ( ~w525 & w630 ) | ( w527 & w630 ) ;
  assign w632 = ~w527 & w631 ;
  assign w633 = w621 | w632 ;
  assign w634 = ( w619 & ~w621 ) | ( w619 & w625 ) | ( ~w621 & w625 ) ;
  assign w635 = w633 | w634 ;
  assign w636 = ( ~\pi107 & \pi108 ) | ( ~\pi107 & w541 ) | ( \pi108 & w541 ) ;
  assign w637 = ( ~\pi106 & \pi108 ) | ( ~\pi106 & w636 ) | ( \pi108 & w636 ) ;
  assign w638 = ( ~\pi108 & w541 ) | ( ~\pi108 & w635 ) | ( w541 & w635 ) ;
  assign w639 = w637 & w638 ;
  assign w640 = ( w527 & w531 ) | ( w527 & ~w538 ) | ( w531 & ~w538 ) ;
  assign w641 = \pi107 & ~w640 ;
  assign w642 = \pi106 | \pi108 ;
  assign w643 = ( ~w640 & w641 ) | ( ~w640 & w642 ) | ( w641 & w642 ) ;
  assign w644 = ~w538 & w643 ;
  assign w645 = ~w525 & w644 ;
  assign w646 = ( \pi108 & w635 ) | ( \pi108 & ~w644 ) | ( w635 & ~w644 ) ;
  assign w647 = w645 & ~w646 ;
  assign w648 = ~\pi108 & w635 ;
  assign w649 = \pi109 ^ w648 ;
  assign w650 = w647 | w649 ;
  assign w651 = ( w455 & w639 ) | ( w455 & ~w650 ) | ( w639 & ~w650 ) ;
  assign w652 = w455 & w651 ;
  assign w653 = ( ~w455 & w639 ) | ( ~w455 & w650 ) | ( w639 & w650 ) ;
  assign w654 = ~w639 & w653 ;
  assign w655 = w541 & ~w632 ;
  assign w656 = ~w621 & w655 ;
  assign w657 = ~w634 & w656 ;
  assign w658 = \pi109 & w635 ;
  assign w659 = ( \pi108 & w635 ) | ( \pi108 & ~w658 ) | ( w635 & ~w658 ) ;
  assign w660 = ( ~\pi108 & w657 ) | ( ~\pi108 & w659 ) | ( w657 & w659 ) ;
  assign w661 = \pi110 ^ w660 ;
  assign w662 = w654 | w661 ;
  assign w663 = ( w377 & w652 ) | ( w377 & ~w662 ) | ( w652 & ~w662 ) ;
  assign w664 = w377 & w663 ;
  assign w665 = ( w545 & ~w553 ) | ( w545 & w635 ) | ( ~w553 & w635 ) ;
  assign w666 = ~w545 & w665 ;
  assign w667 = \pi111 ^ w666 ;
  assign w668 = w554 ^ w667 ;
  assign w669 = ( ~w377 & w652 ) | ( ~w377 & w662 ) | ( w652 & w662 ) ;
  assign w670 = ~w652 & w669 ;
  assign w671 = w668 | w670 ;
  assign w672 = ( w307 & w664 ) | ( w307 & ~w671 ) | ( w664 & ~w671 ) ;
  assign w673 = w307 & w672 ;
  assign w674 = w558 | w560 ;
  assign w675 = w635 & ~w674 ;
  assign w676 = w567 ^ w675 ;
  assign w677 = ( ~w307 & w664 ) | ( ~w307 & w671 ) | ( w664 & w671 ) ;
  assign w678 = ~w664 & w677 ;
  assign w679 = w676 | w678 ;
  assign w680 = ( w246 & w673 ) | ( w246 & ~w679 ) | ( w673 & ~w679 ) ;
  assign w681 = w246 & w680 ;
  assign w682 = ( ~w246 & w673 ) | ( ~w246 & w679 ) | ( w673 & w679 ) ;
  assign w683 = ~w673 & w682 ;
  assign w684 = w570 | w572 ;
  assign w685 = w635 & ~w684 ;
  assign w686 = w576 ^ w685 ;
  assign w687 = w683 | w686 ;
  assign w688 = ( w185 & w681 ) | ( w185 & ~w687 ) | ( w681 & ~w687 ) ;
  assign w689 = w185 & w688 ;
  assign w690 = w579 | w584 ;
  assign w691 = w635 & ~w690 ;
  assign w692 = w582 ^ w691 ;
  assign w693 = ( ~w185 & w681 ) | ( ~w185 & w687 ) | ( w681 & w687 ) ;
  assign w694 = ~w681 & w693 ;
  assign w695 = w692 | w694 ;
  assign w696 = ( w145 & w689 ) | ( w145 & ~w695 ) | ( w689 & ~w695 ) ;
  assign w697 = w145 & w696 ;
  assign w698 = w587 | w592 ;
  assign w699 = w635 & ~w698 ;
  assign w700 = w590 ^ w699 ;
  assign w701 = ( ~w145 & w689 ) | ( ~w145 & w695 ) | ( w689 & w695 ) ;
  assign w702 = ~w689 & w701 ;
  assign w703 = w700 | w702 ;
  assign w704 = ( w132 & w697 ) | ( w132 & ~w703 ) | ( w697 & ~w703 ) ;
  assign w705 = w132 & w704 ;
  assign w706 = w595 | w600 ;
  assign w707 = w635 & ~w706 ;
  assign w708 = w598 ^ w707 ;
  assign w709 = ( ~w132 & w697 ) | ( ~w132 & w703 ) | ( w697 & w703 ) ;
  assign w710 = ~w697 & w709 ;
  assign w711 = w708 | w710 ;
  assign w712 = ~w705 & w711 ;
  assign w713 = w603 | w608 ;
  assign w714 = w635 & ~w713 ;
  assign w715 = w606 ^ w714 ;
  assign w716 = ( ~w621 & w712 ) | ( ~w621 & w715 ) | ( w712 & w715 ) ;
  assign w717 = w610 & ~w716 ;
  assign w718 = ~w613 & w635 ;
  assign w719 = ( w716 & ~w717 ) | ( w716 & w718 ) | ( ~w717 & w718 ) ;
  assign w720 = w621 | w719 ;
  assign w721 = ~w129 & w720 ;
  assign w722 = ( w705 & w711 ) | ( w705 & w715 ) | ( w711 & w715 ) ;
  assign w723 = ~w705 & w722 ;
  assign w724 = ( w129 & w610 ) | ( w129 & w613 ) | ( w610 & w613 ) ;
  assign w725 = ( w613 & ~w635 ) | ( w613 & w724 ) | ( ~w635 & w724 ) ;
  assign w726 = w610 & w725 ;
  assign w727 = w724 ^ w726 ;
  assign w728 = ( w509 & w514 ) | ( w509 & w541 ) | ( w514 & w541 ) ;
  assign w729 = w541 & ~w728 ;
  assign w730 = w512 ^ w729 ;
  assign w731 = ( ~w625 & w632 ) | ( ~w625 & w730 ) | ( w632 & w730 ) ;
  assign w732 = ~w632 & w731 ;
  assign w733 = ( ~w619 & w621 ) | ( ~w619 & w732 ) | ( w621 & w732 ) ;
  assign w734 = ~w621 & w733 ;
  assign w735 = w723 | w734 ;
  assign w736 = ( w721 & ~w723 ) | ( w721 & w727 ) | ( ~w723 & w727 ) ;
  assign w737 = w735 | w736 ;
  assign w738 = ( ~\pi105 & \pi106 ) | ( ~\pi105 & w635 ) | ( \pi106 & w635 ) ;
  assign w739 = ( ~\pi104 & \pi106 ) | ( ~\pi104 & w738 ) | ( \pi106 & w738 ) ;
  assign w740 = ( ~\pi106 & w635 ) | ( ~\pi106 & w737 ) | ( w635 & w737 ) ;
  assign w741 = w739 & w740 ;
  assign w742 = ( w621 & w625 ) | ( w621 & ~w632 ) | ( w625 & ~w632 ) ;
  assign w743 = \pi105 & ~w742 ;
  assign w744 = \pi104 | \pi106 ;
  assign w745 = ( ~w742 & w743 ) | ( ~w742 & w744 ) | ( w743 & w744 ) ;
  assign w746 = ~w632 & w745 ;
  assign w747 = ~w619 & w746 ;
  assign w748 = ( \pi106 & w737 ) | ( \pi106 & ~w746 ) | ( w737 & ~w746 ) ;
  assign w749 = w747 & ~w748 ;
  assign w750 = ~\pi106 & w737 ;
  assign w751 = \pi107 ^ w750 ;
  assign w752 = w749 | w751 ;
  assign w753 = ( w541 & w741 ) | ( w541 & ~w752 ) | ( w741 & ~w752 ) ;
  assign w754 = w541 & w753 ;
  assign w755 = ( ~w541 & w741 ) | ( ~w541 & w752 ) | ( w741 & w752 ) ;
  assign w756 = ~w741 & w755 ;
  assign w757 = w635 & ~w734 ;
  assign w758 = ~w723 & w757 ;
  assign w759 = ~w736 & w758 ;
  assign w760 = \pi107 & w737 ;
  assign w761 = ( \pi106 & w737 ) | ( \pi106 & ~w760 ) | ( w737 & ~w760 ) ;
  assign w762 = ( ~\pi106 & w759 ) | ( ~\pi106 & w761 ) | ( w759 & w761 ) ;
  assign w763 = \pi108 ^ w762 ;
  assign w764 = w756 | w763 ;
  assign w765 = ( w455 & w754 ) | ( w455 & ~w764 ) | ( w754 & ~w764 ) ;
  assign w766 = w455 & w765 ;
  assign w767 = ( w639 & ~w647 ) | ( w639 & w737 ) | ( ~w647 & w737 ) ;
  assign w768 = ~w639 & w767 ;
  assign w769 = \pi109 ^ w768 ;
  assign w770 = w648 ^ w769 ;
  assign w771 = ( ~w455 & w754 ) | ( ~w455 & w764 ) | ( w754 & w764 ) ;
  assign w772 = ~w754 & w771 ;
  assign w773 = w770 | w772 ;
  assign w774 = ( w377 & w766 ) | ( w377 & ~w773 ) | ( w766 & ~w773 ) ;
  assign w775 = w377 & w774 ;
  assign w776 = w652 | w654 ;
  assign w777 = w737 & ~w776 ;
  assign w778 = w661 ^ w777 ;
  assign w779 = ( ~w377 & w766 ) | ( ~w377 & w773 ) | ( w766 & w773 ) ;
  assign w780 = ~w766 & w779 ;
  assign w781 = w778 | w780 ;
  assign w782 = ( w307 & w775 ) | ( w307 & ~w781 ) | ( w775 & ~w781 ) ;
  assign w783 = w307 & w782 ;
  assign w784 = w664 | w670 ;
  assign w785 = w737 & ~w784 ;
  assign w786 = w668 ^ w785 ;
  assign w787 = ( ~w307 & w775 ) | ( ~w307 & w781 ) | ( w775 & w781 ) ;
  assign w788 = ~w775 & w787 ;
  assign w789 = w786 | w788 ;
  assign w790 = ( w246 & w783 ) | ( w246 & ~w789 ) | ( w783 & ~w789 ) ;
  assign w791 = w246 & w790 ;
  assign w792 = w673 | w678 ;
  assign w793 = w737 & ~w792 ;
  assign w794 = w676 ^ w793 ;
  assign w795 = ( ~w246 & w783 ) | ( ~w246 & w789 ) | ( w783 & w789 ) ;
  assign w796 = ~w783 & w795 ;
  assign w797 = w794 | w796 ;
  assign w798 = ( w185 & w791 ) | ( w185 & ~w797 ) | ( w791 & ~w797 ) ;
  assign w799 = w185 & w798 ;
  assign w800 = ( ~w185 & w791 ) | ( ~w185 & w797 ) | ( w791 & w797 ) ;
  assign w801 = ~w791 & w800 ;
  assign w802 = w681 | w683 ;
  assign w803 = w737 & ~w802 ;
  assign w804 = w686 ^ w803 ;
  assign w805 = w801 | w804 ;
  assign w806 = ( w145 & w799 ) | ( w145 & ~w805 ) | ( w799 & ~w805 ) ;
  assign w807 = w145 & w806 ;
  assign w808 = w689 | w694 ;
  assign w809 = w737 & ~w808 ;
  assign w810 = w692 ^ w809 ;
  assign w811 = ( ~w145 & w799 ) | ( ~w145 & w805 ) | ( w799 & w805 ) ;
  assign w812 = ~w799 & w811 ;
  assign w813 = w810 | w812 ;
  assign w814 = ( w132 & w807 ) | ( w132 & ~w813 ) | ( w807 & ~w813 ) ;
  assign w815 = w132 & w814 ;
  assign w816 = w697 | w702 ;
  assign w817 = w737 & ~w816 ;
  assign w818 = w700 ^ w817 ;
  assign w819 = ( ~w132 & w807 ) | ( ~w132 & w813 ) | ( w807 & w813 ) ;
  assign w820 = ~w807 & w819 ;
  assign w821 = w818 | w820 ;
  assign w822 = ~w815 & w821 ;
  assign w823 = w705 | w710 ;
  assign w824 = w737 & ~w823 ;
  assign w825 = w708 ^ w824 ;
  assign w826 = ( ~w723 & w822 ) | ( ~w723 & w825 ) | ( w822 & w825 ) ;
  assign w827 = w712 & ~w826 ;
  assign w828 = ~w715 & w737 ;
  assign w829 = ( w826 & ~w827 ) | ( w826 & w828 ) | ( ~w827 & w828 ) ;
  assign w830 = w723 | w829 ;
  assign w831 = ~w129 & w830 ;
  assign w832 = ( w815 & w821 ) | ( w815 & w825 ) | ( w821 & w825 ) ;
  assign w833 = ~w815 & w832 ;
  assign w834 = ( w129 & w712 ) | ( w129 & w715 ) | ( w712 & w715 ) ;
  assign w835 = ( w715 & ~w737 ) | ( w715 & w834 ) | ( ~w737 & w834 ) ;
  assign w836 = w712 & w835 ;
  assign w837 = w834 ^ w836 ;
  assign w838 = ( w603 & w608 ) | ( w603 & w635 ) | ( w608 & w635 ) ;
  assign w839 = w635 & ~w838 ;
  assign w840 = w606 ^ w839 ;
  assign w841 = ( ~w727 & w734 ) | ( ~w727 & w840 ) | ( w734 & w840 ) ;
  assign w842 = ~w734 & w841 ;
  assign w843 = ( ~w721 & w723 ) | ( ~w721 & w842 ) | ( w723 & w842 ) ;
  assign w844 = ~w723 & w843 ;
  assign w845 = w833 | w844 ;
  assign w846 = ( w831 & ~w833 ) | ( w831 & w837 ) | ( ~w833 & w837 ) ;
  assign w847 = w845 | w846 ;
  assign w848 = ( ~\pi103 & \pi104 ) | ( ~\pi103 & w737 ) | ( \pi104 & w737 ) ;
  assign w849 = ( ~\pi102 & \pi104 ) | ( ~\pi102 & w848 ) | ( \pi104 & w848 ) ;
  assign w850 = ( ~\pi104 & w737 ) | ( ~\pi104 & w847 ) | ( w737 & w847 ) ;
  assign w851 = w849 & w850 ;
  assign w852 = ( w723 & w727 ) | ( w723 & ~w734 ) | ( w727 & ~w734 ) ;
  assign w853 = \pi103 & ~w852 ;
  assign w854 = \pi102 | \pi104 ;
  assign w855 = ( ~w852 & w853 ) | ( ~w852 & w854 ) | ( w853 & w854 ) ;
  assign w856 = ~w734 & w855 ;
  assign w857 = ~w721 & w856 ;
  assign w858 = ( \pi104 & w847 ) | ( \pi104 & ~w856 ) | ( w847 & ~w856 ) ;
  assign w859 = w857 & ~w858 ;
  assign w860 = ~\pi104 & w847 ;
  assign w861 = \pi105 ^ w860 ;
  assign w862 = w859 | w861 ;
  assign w863 = ( w635 & w851 ) | ( w635 & ~w862 ) | ( w851 & ~w862 ) ;
  assign w864 = w635 & w863 ;
  assign w865 = ( ~w635 & w851 ) | ( ~w635 & w862 ) | ( w851 & w862 ) ;
  assign w866 = ~w851 & w865 ;
  assign w867 = w737 & ~w844 ;
  assign w868 = ~w833 & w867 ;
  assign w869 = ~w846 & w868 ;
  assign w870 = \pi105 & w847 ;
  assign w871 = ( \pi104 & w847 ) | ( \pi104 & ~w870 ) | ( w847 & ~w870 ) ;
  assign w872 = ( ~\pi104 & w869 ) | ( ~\pi104 & w871 ) | ( w869 & w871 ) ;
  assign w873 = \pi106 ^ w872 ;
  assign w874 = w866 | w873 ;
  assign w875 = ( w541 & w864 ) | ( w541 & ~w874 ) | ( w864 & ~w874 ) ;
  assign w876 = w541 & w875 ;
  assign w877 = ( w741 & ~w749 ) | ( w741 & w847 ) | ( ~w749 & w847 ) ;
  assign w878 = ~w741 & w877 ;
  assign w879 = \pi107 ^ w878 ;
  assign w880 = w750 ^ w879 ;
  assign w881 = ( ~w541 & w864 ) | ( ~w541 & w874 ) | ( w864 & w874 ) ;
  assign w882 = ~w864 & w881 ;
  assign w883 = w880 | w882 ;
  assign w884 = ( w455 & w876 ) | ( w455 & ~w883 ) | ( w876 & ~w883 ) ;
  assign w885 = w455 & w884 ;
  assign w886 = w754 | w756 ;
  assign w887 = w847 & ~w886 ;
  assign w888 = w763 ^ w887 ;
  assign w889 = ( ~w455 & w876 ) | ( ~w455 & w883 ) | ( w876 & w883 ) ;
  assign w890 = ~w876 & w889 ;
  assign w891 = w888 | w890 ;
  assign w892 = ( w377 & w885 ) | ( w377 & ~w891 ) | ( w885 & ~w891 ) ;
  assign w893 = w377 & w892 ;
  assign w894 = w766 | w772 ;
  assign w895 = w847 & ~w894 ;
  assign w896 = w770 ^ w895 ;
  assign w897 = ( ~w377 & w885 ) | ( ~w377 & w891 ) | ( w885 & w891 ) ;
  assign w898 = ~w885 & w897 ;
  assign w899 = w896 | w898 ;
  assign w900 = ( w307 & w893 ) | ( w307 & ~w899 ) | ( w893 & ~w899 ) ;
  assign w901 = w307 & w900 ;
  assign w902 = w775 | w780 ;
  assign w903 = w847 & ~w902 ;
  assign w904 = w778 ^ w903 ;
  assign w905 = ( ~w307 & w893 ) | ( ~w307 & w899 ) | ( w893 & w899 ) ;
  assign w906 = ~w893 & w905 ;
  assign w907 = w904 | w906 ;
  assign w908 = ( w246 & w901 ) | ( w246 & ~w907 ) | ( w901 & ~w907 ) ;
  assign w909 = w246 & w908 ;
  assign w910 = w783 | w788 ;
  assign w911 = w847 & ~w910 ;
  assign w912 = w786 ^ w911 ;
  assign w913 = ( ~w246 & w901 ) | ( ~w246 & w907 ) | ( w901 & w907 ) ;
  assign w914 = ~w901 & w913 ;
  assign w915 = w912 | w914 ;
  assign w916 = ( w185 & w909 ) | ( w185 & ~w915 ) | ( w909 & ~w915 ) ;
  assign w917 = w185 & w916 ;
  assign w918 = w791 | w796 ;
  assign w919 = w847 & ~w918 ;
  assign w920 = w794 ^ w919 ;
  assign w921 = ( ~w185 & w909 ) | ( ~w185 & w915 ) | ( w909 & w915 ) ;
  assign w922 = ~w909 & w921 ;
  assign w923 = w920 | w922 ;
  assign w924 = ( w145 & w917 ) | ( w145 & ~w923 ) | ( w917 & ~w923 ) ;
  assign w925 = w145 & w924 ;
  assign w926 = ( ~w145 & w917 ) | ( ~w145 & w923 ) | ( w917 & w923 ) ;
  assign w927 = ~w917 & w926 ;
  assign w928 = w799 | w801 ;
  assign w929 = w847 & ~w928 ;
  assign w930 = w804 ^ w929 ;
  assign w931 = w927 | w930 ;
  assign w932 = ( w132 & w925 ) | ( w132 & ~w931 ) | ( w925 & ~w931 ) ;
  assign w933 = w132 & w932 ;
  assign w934 = w807 | w812 ;
  assign w935 = w847 & ~w934 ;
  assign w936 = w810 ^ w935 ;
  assign w937 = ( ~w132 & w925 ) | ( ~w132 & w931 ) | ( w925 & w931 ) ;
  assign w938 = ~w925 & w937 ;
  assign w939 = w936 | w938 ;
  assign w940 = ~w933 & w939 ;
  assign w941 = w815 | w820 ;
  assign w942 = w847 & ~w941 ;
  assign w943 = w818 ^ w942 ;
  assign w944 = ( ~w833 & w940 ) | ( ~w833 & w943 ) | ( w940 & w943 ) ;
  assign w945 = w822 & ~w944 ;
  assign w946 = ~w825 & w847 ;
  assign w947 = ( w944 & ~w945 ) | ( w944 & w946 ) | ( ~w945 & w946 ) ;
  assign w948 = w833 | w947 ;
  assign w949 = ~w129 & w948 ;
  assign w950 = ( w933 & w939 ) | ( w933 & w943 ) | ( w939 & w943 ) ;
  assign w951 = ~w933 & w950 ;
  assign w952 = ( w129 & w822 ) | ( w129 & w825 ) | ( w822 & w825 ) ;
  assign w953 = ( w825 & ~w847 ) | ( w825 & w952 ) | ( ~w847 & w952 ) ;
  assign w954 = w822 & w953 ;
  assign w955 = w952 ^ w954 ;
  assign w956 = ( w705 & w710 ) | ( w705 & w737 ) | ( w710 & w737 ) ;
  assign w957 = w737 & ~w956 ;
  assign w958 = w708 ^ w957 ;
  assign w959 = ( ~w837 & w844 ) | ( ~w837 & w958 ) | ( w844 & w958 ) ;
  assign w960 = ~w844 & w959 ;
  assign w961 = ( ~w831 & w833 ) | ( ~w831 & w960 ) | ( w833 & w960 ) ;
  assign w962 = ~w833 & w961 ;
  assign w963 = w951 | w962 ;
  assign w964 = ( w949 & ~w951 ) | ( w949 & w955 ) | ( ~w951 & w955 ) ;
  assign w965 = w963 | w964 ;
  assign w966 = ( ~\pi101 & \pi102 ) | ( ~\pi101 & w847 ) | ( \pi102 & w847 ) ;
  assign w967 = ( ~\pi100 & \pi102 ) | ( ~\pi100 & w966 ) | ( \pi102 & w966 ) ;
  assign w968 = ( ~\pi102 & w847 ) | ( ~\pi102 & w965 ) | ( w847 & w965 ) ;
  assign w969 = w967 & w968 ;
  assign w970 = ( w833 & w837 ) | ( w833 & ~w844 ) | ( w837 & ~w844 ) ;
  assign w971 = \pi101 & ~w970 ;
  assign w972 = \pi100 | \pi102 ;
  assign w973 = ( ~w970 & w971 ) | ( ~w970 & w972 ) | ( w971 & w972 ) ;
  assign w974 = ~w844 & w973 ;
  assign w975 = ~w831 & w974 ;
  assign w976 = ( \pi102 & w965 ) | ( \pi102 & ~w974 ) | ( w965 & ~w974 ) ;
  assign w977 = w975 & ~w976 ;
  assign w978 = ~\pi102 & w965 ;
  assign w979 = \pi103 ^ w978 ;
  assign w980 = w977 | w979 ;
  assign w981 = ( w737 & w969 ) | ( w737 & ~w980 ) | ( w969 & ~w980 ) ;
  assign w982 = w737 & w981 ;
  assign w983 = ( ~w737 & w969 ) | ( ~w737 & w980 ) | ( w969 & w980 ) ;
  assign w984 = ~w969 & w983 ;
  assign w985 = w847 & ~w962 ;
  assign w986 = ~w951 & w985 ;
  assign w987 = ~w964 & w986 ;
  assign w988 = \pi103 & w965 ;
  assign w989 = ( \pi102 & w965 ) | ( \pi102 & ~w988 ) | ( w965 & ~w988 ) ;
  assign w990 = ( ~\pi102 & w987 ) | ( ~\pi102 & w989 ) | ( w987 & w989 ) ;
  assign w991 = \pi104 ^ w990 ;
  assign w992 = w984 | w991 ;
  assign w993 = ( w635 & w982 ) | ( w635 & ~w992 ) | ( w982 & ~w992 ) ;
  assign w994 = w635 & w993 ;
  assign w995 = ( w851 & ~w859 ) | ( w851 & w965 ) | ( ~w859 & w965 ) ;
  assign w996 = ~w851 & w995 ;
  assign w997 = \pi105 ^ w996 ;
  assign w998 = w860 ^ w997 ;
  assign w999 = ( ~w635 & w982 ) | ( ~w635 & w992 ) | ( w982 & w992 ) ;
  assign w1000 = ~w982 & w999 ;
  assign w1001 = w998 | w1000 ;
  assign w1002 = ( w541 & w994 ) | ( w541 & ~w1001 ) | ( w994 & ~w1001 ) ;
  assign w1003 = w541 & w1002 ;
  assign w1004 = w864 | w866 ;
  assign w1005 = w965 & ~w1004 ;
  assign w1006 = w873 ^ w1005 ;
  assign w1007 = ( ~w541 & w994 ) | ( ~w541 & w1001 ) | ( w994 & w1001 ) ;
  assign w1008 = ~w994 & w1007 ;
  assign w1009 = w1006 | w1008 ;
  assign w1010 = ( w455 & w1003 ) | ( w455 & ~w1009 ) | ( w1003 & ~w1009 ) ;
  assign w1011 = w455 & w1010 ;
  assign w1012 = w876 | w882 ;
  assign w1013 = w965 & ~w1012 ;
  assign w1014 = w880 ^ w1013 ;
  assign w1015 = ( ~w455 & w1003 ) | ( ~w455 & w1009 ) | ( w1003 & w1009 ) ;
  assign w1016 = ~w1003 & w1015 ;
  assign w1017 = w1014 | w1016 ;
  assign w1018 = ( w377 & w1011 ) | ( w377 & ~w1017 ) | ( w1011 & ~w1017 ) ;
  assign w1019 = w377 & w1018 ;
  assign w1020 = w885 | w890 ;
  assign w1021 = w965 & ~w1020 ;
  assign w1022 = w888 ^ w1021 ;
  assign w1023 = ( ~w377 & w1011 ) | ( ~w377 & w1017 ) | ( w1011 & w1017 ) ;
  assign w1024 = ~w1011 & w1023 ;
  assign w1025 = w1022 | w1024 ;
  assign w1026 = ( w307 & w1019 ) | ( w307 & ~w1025 ) | ( w1019 & ~w1025 ) ;
  assign w1027 = w307 & w1026 ;
  assign w1028 = w893 | w898 ;
  assign w1029 = w965 & ~w1028 ;
  assign w1030 = w896 ^ w1029 ;
  assign w1031 = ( ~w307 & w1019 ) | ( ~w307 & w1025 ) | ( w1019 & w1025 ) ;
  assign w1032 = ~w1019 & w1031 ;
  assign w1033 = w1030 | w1032 ;
  assign w1034 = ( w246 & w1027 ) | ( w246 & ~w1033 ) | ( w1027 & ~w1033 ) ;
  assign w1035 = w246 & w1034 ;
  assign w1036 = w901 | w906 ;
  assign w1037 = w965 & ~w1036 ;
  assign w1038 = w904 ^ w1037 ;
  assign w1039 = ( ~w246 & w1027 ) | ( ~w246 & w1033 ) | ( w1027 & w1033 ) ;
  assign w1040 = ~w1027 & w1039 ;
  assign w1041 = w1038 | w1040 ;
  assign w1042 = ( w185 & w1035 ) | ( w185 & ~w1041 ) | ( w1035 & ~w1041 ) ;
  assign w1043 = w185 & w1042 ;
  assign w1044 = w909 | w914 ;
  assign w1045 = w965 & ~w1044 ;
  assign w1046 = w912 ^ w1045 ;
  assign w1047 = ( ~w185 & w1035 ) | ( ~w185 & w1041 ) | ( w1035 & w1041 ) ;
  assign w1048 = ~w1035 & w1047 ;
  assign w1049 = w1046 | w1048 ;
  assign w1050 = ( w145 & w1043 ) | ( w145 & ~w1049 ) | ( w1043 & ~w1049 ) ;
  assign w1051 = w145 & w1050 ;
  assign w1052 = w917 | w922 ;
  assign w1053 = w965 & ~w1052 ;
  assign w1054 = w920 ^ w1053 ;
  assign w1055 = ( ~w145 & w1043 ) | ( ~w145 & w1049 ) | ( w1043 & w1049 ) ;
  assign w1056 = ~w1043 & w1055 ;
  assign w1057 = w1054 | w1056 ;
  assign w1058 = ( w132 & w1051 ) | ( w132 & ~w1057 ) | ( w1051 & ~w1057 ) ;
  assign w1059 = w132 & w1058 ;
  assign w1060 = ( ~w132 & w1051 ) | ( ~w132 & w1057 ) | ( w1051 & w1057 ) ;
  assign w1061 = ~w1051 & w1060 ;
  assign w1062 = w925 | w927 ;
  assign w1063 = w965 & ~w1062 ;
  assign w1064 = w930 ^ w1063 ;
  assign w1065 = w1061 | w1064 ;
  assign w1066 = ~w1059 & w1065 ;
  assign w1067 = w933 | w938 ;
  assign w1068 = w965 & ~w1067 ;
  assign w1069 = w936 ^ w1068 ;
  assign w1070 = ( ~w951 & w1066 ) | ( ~w951 & w1069 ) | ( w1066 & w1069 ) ;
  assign w1071 = w940 & ~w1070 ;
  assign w1072 = ~w943 & w965 ;
  assign w1073 = ( w1070 & ~w1071 ) | ( w1070 & w1072 ) | ( ~w1071 & w1072 ) ;
  assign w1074 = w951 | w1073 ;
  assign w1075 = ~w129 & w1074 ;
  assign w1076 = ( w1059 & w1065 ) | ( w1059 & w1069 ) | ( w1065 & w1069 ) ;
  assign w1077 = ~w1059 & w1076 ;
  assign w1078 = ( w129 & w940 ) | ( w129 & w943 ) | ( w940 & w943 ) ;
  assign w1079 = ( w943 & ~w965 ) | ( w943 & w1078 ) | ( ~w965 & w1078 ) ;
  assign w1080 = w940 & w1079 ;
  assign w1081 = w1078 ^ w1080 ;
  assign w1082 = ( w815 & w820 ) | ( w815 & w847 ) | ( w820 & w847 ) ;
  assign w1083 = w847 & ~w1082 ;
  assign w1084 = w818 ^ w1083 ;
  assign w1085 = ( ~w955 & w962 ) | ( ~w955 & w1084 ) | ( w962 & w1084 ) ;
  assign w1086 = ~w962 & w1085 ;
  assign w1087 = ( ~w949 & w951 ) | ( ~w949 & w1086 ) | ( w951 & w1086 ) ;
  assign w1088 = ~w951 & w1087 ;
  assign w1089 = w1077 | w1088 ;
  assign w1090 = ( w1075 & ~w1077 ) | ( w1075 & w1081 ) | ( ~w1077 & w1081 ) ;
  assign w1091 = w1089 | w1090 ;
  assign w1092 = ( ~\pi099 & \pi100 ) | ( ~\pi099 & w965 ) | ( \pi100 & w965 ) ;
  assign w1093 = ( ~\pi098 & \pi100 ) | ( ~\pi098 & w1092 ) | ( \pi100 & w1092 ) ;
  assign w1094 = ( ~\pi100 & w965 ) | ( ~\pi100 & w1091 ) | ( w965 & w1091 ) ;
  assign w1095 = w1093 & w1094 ;
  assign w1096 = ( w951 & w955 ) | ( w951 & ~w962 ) | ( w955 & ~w962 ) ;
  assign w1097 = \pi099 & ~w1096 ;
  assign w1098 = \pi098 | \pi100 ;
  assign w1099 = ( ~w1096 & w1097 ) | ( ~w1096 & w1098 ) | ( w1097 & w1098 ) ;
  assign w1100 = ~w962 & w1099 ;
  assign w1101 = ~w949 & w1100 ;
  assign w1102 = ( \pi100 & w1091 ) | ( \pi100 & ~w1100 ) | ( w1091 & ~w1100 ) ;
  assign w1103 = w1101 & ~w1102 ;
  assign w1104 = ~\pi100 & w1091 ;
  assign w1105 = \pi101 ^ w1104 ;
  assign w1106 = w1103 | w1105 ;
  assign w1107 = ( w847 & w1095 ) | ( w847 & ~w1106 ) | ( w1095 & ~w1106 ) ;
  assign w1108 = w847 & w1107 ;
  assign w1109 = ( ~w847 & w1095 ) | ( ~w847 & w1106 ) | ( w1095 & w1106 ) ;
  assign w1110 = ~w1095 & w1109 ;
  assign w1111 = w965 & ~w1088 ;
  assign w1112 = ~w1077 & w1111 ;
  assign w1113 = ~w1090 & w1112 ;
  assign w1114 = \pi101 & w1091 ;
  assign w1115 = ( \pi100 & w1091 ) | ( \pi100 & ~w1114 ) | ( w1091 & ~w1114 ) ;
  assign w1116 = ( ~\pi100 & w1113 ) | ( ~\pi100 & w1115 ) | ( w1113 & w1115 ) ;
  assign w1117 = \pi102 ^ w1116 ;
  assign w1118 = w1110 | w1117 ;
  assign w1119 = ( w737 & w1108 ) | ( w737 & ~w1118 ) | ( w1108 & ~w1118 ) ;
  assign w1120 = w737 & w1119 ;
  assign w1121 = ( w969 & ~w977 ) | ( w969 & w1091 ) | ( ~w977 & w1091 ) ;
  assign w1122 = ~w969 & w1121 ;
  assign w1123 = \pi103 ^ w1122 ;
  assign w1124 = w978 ^ w1123 ;
  assign w1125 = ( ~w737 & w1108 ) | ( ~w737 & w1118 ) | ( w1108 & w1118 ) ;
  assign w1126 = ~w1108 & w1125 ;
  assign w1127 = w1124 | w1126 ;
  assign w1128 = ( w635 & w1120 ) | ( w635 & ~w1127 ) | ( w1120 & ~w1127 ) ;
  assign w1129 = w635 & w1128 ;
  assign w1130 = w982 | w984 ;
  assign w1131 = w1091 & ~w1130 ;
  assign w1132 = w991 ^ w1131 ;
  assign w1133 = ( ~w635 & w1120 ) | ( ~w635 & w1127 ) | ( w1120 & w1127 ) ;
  assign w1134 = ~w1120 & w1133 ;
  assign w1135 = w1132 | w1134 ;
  assign w1136 = ( w541 & w1129 ) | ( w541 & ~w1135 ) | ( w1129 & ~w1135 ) ;
  assign w1137 = w541 & w1136 ;
  assign w1138 = w994 | w1000 ;
  assign w1139 = w1091 & ~w1138 ;
  assign w1140 = w998 ^ w1139 ;
  assign w1141 = ( ~w541 & w1129 ) | ( ~w541 & w1135 ) | ( w1129 & w1135 ) ;
  assign w1142 = ~w1129 & w1141 ;
  assign w1143 = w1140 | w1142 ;
  assign w1144 = ( w455 & w1137 ) | ( w455 & ~w1143 ) | ( w1137 & ~w1143 ) ;
  assign w1145 = w455 & w1144 ;
  assign w1146 = w1003 | w1008 ;
  assign w1147 = w1091 & ~w1146 ;
  assign w1148 = w1006 ^ w1147 ;
  assign w1149 = ( ~w455 & w1137 ) | ( ~w455 & w1143 ) | ( w1137 & w1143 ) ;
  assign w1150 = ~w1137 & w1149 ;
  assign w1151 = w1148 | w1150 ;
  assign w1152 = ( w377 & w1145 ) | ( w377 & ~w1151 ) | ( w1145 & ~w1151 ) ;
  assign w1153 = w377 & w1152 ;
  assign w1154 = w1011 | w1016 ;
  assign w1155 = w1091 & ~w1154 ;
  assign w1156 = w1014 ^ w1155 ;
  assign w1157 = ( ~w377 & w1145 ) | ( ~w377 & w1151 ) | ( w1145 & w1151 ) ;
  assign w1158 = ~w1145 & w1157 ;
  assign w1159 = w1156 | w1158 ;
  assign w1160 = ( w307 & w1153 ) | ( w307 & ~w1159 ) | ( w1153 & ~w1159 ) ;
  assign w1161 = w307 & w1160 ;
  assign w1162 = w1019 | w1024 ;
  assign w1163 = w1091 & ~w1162 ;
  assign w1164 = w1022 ^ w1163 ;
  assign w1165 = ( ~w307 & w1153 ) | ( ~w307 & w1159 ) | ( w1153 & w1159 ) ;
  assign w1166 = ~w1153 & w1165 ;
  assign w1167 = w1164 | w1166 ;
  assign w1168 = ( w246 & w1161 ) | ( w246 & ~w1167 ) | ( w1161 & ~w1167 ) ;
  assign w1169 = w246 & w1168 ;
  assign w1170 = w1027 | w1032 ;
  assign w1171 = w1091 & ~w1170 ;
  assign w1172 = w1030 ^ w1171 ;
  assign w1173 = ( ~w246 & w1161 ) | ( ~w246 & w1167 ) | ( w1161 & w1167 ) ;
  assign w1174 = ~w1161 & w1173 ;
  assign w1175 = w1172 | w1174 ;
  assign w1176 = ( w185 & w1169 ) | ( w185 & ~w1175 ) | ( w1169 & ~w1175 ) ;
  assign w1177 = w185 & w1176 ;
  assign w1178 = w1035 | w1040 ;
  assign w1179 = w1091 & ~w1178 ;
  assign w1180 = w1038 ^ w1179 ;
  assign w1181 = ( ~w185 & w1169 ) | ( ~w185 & w1175 ) | ( w1169 & w1175 ) ;
  assign w1182 = ~w1169 & w1181 ;
  assign w1183 = w1180 | w1182 ;
  assign w1184 = ( w145 & w1177 ) | ( w145 & ~w1183 ) | ( w1177 & ~w1183 ) ;
  assign w1185 = w145 & w1184 ;
  assign w1186 = w1043 | w1048 ;
  assign w1187 = w1091 & ~w1186 ;
  assign w1188 = w1046 ^ w1187 ;
  assign w1189 = ( ~w145 & w1177 ) | ( ~w145 & w1183 ) | ( w1177 & w1183 ) ;
  assign w1190 = ~w1177 & w1189 ;
  assign w1191 = w1188 | w1190 ;
  assign w1192 = ( w132 & w1185 ) | ( w132 & ~w1191 ) | ( w1185 & ~w1191 ) ;
  assign w1193 = w132 & w1192 ;
  assign w1194 = w1051 | w1056 ;
  assign w1195 = w1091 & ~w1194 ;
  assign w1196 = w1054 ^ w1195 ;
  assign w1197 = ( ~w132 & w1185 ) | ( ~w132 & w1191 ) | ( w1185 & w1191 ) ;
  assign w1198 = ~w1185 & w1197 ;
  assign w1199 = w1196 | w1198 ;
  assign w1200 = ~w1193 & w1199 ;
  assign w1201 = w1059 | w1061 ;
  assign w1202 = w1091 & ~w1201 ;
  assign w1203 = w1064 ^ w1202 ;
  assign w1204 = ( ~w1077 & w1200 ) | ( ~w1077 & w1203 ) | ( w1200 & w1203 ) ;
  assign w1205 = w1066 & ~w1204 ;
  assign w1206 = ~w1069 & w1091 ;
  assign w1207 = ( w1204 & ~w1205 ) | ( w1204 & w1206 ) | ( ~w1205 & w1206 ) ;
  assign w1208 = w1077 | w1207 ;
  assign w1209 = ~w129 & w1208 ;
  assign w1210 = ( w1193 & w1199 ) | ( w1193 & w1203 ) | ( w1199 & w1203 ) ;
  assign w1211 = ~w1193 & w1210 ;
  assign w1212 = ( w129 & w1066 ) | ( w129 & w1069 ) | ( w1066 & w1069 ) ;
  assign w1213 = ( w1069 & ~w1091 ) | ( w1069 & w1212 ) | ( ~w1091 & w1212 ) ;
  assign w1214 = w1066 & w1213 ;
  assign w1215 = w1212 ^ w1214 ;
  assign w1216 = ( w933 & w938 ) | ( w933 & w965 ) | ( w938 & w965 ) ;
  assign w1217 = w965 & ~w1216 ;
  assign w1218 = w936 ^ w1217 ;
  assign w1219 = ( ~w1081 & w1088 ) | ( ~w1081 & w1218 ) | ( w1088 & w1218 ) ;
  assign w1220 = ~w1088 & w1219 ;
  assign w1221 = ( ~w1075 & w1077 ) | ( ~w1075 & w1220 ) | ( w1077 & w1220 ) ;
  assign w1222 = ~w1077 & w1221 ;
  assign w1223 = w1211 | w1222 ;
  assign w1224 = ( w1209 & ~w1211 ) | ( w1209 & w1215 ) | ( ~w1211 & w1215 ) ;
  assign w1225 = w1223 | w1224 ;
  assign w1226 = ( ~\pi097 & \pi098 ) | ( ~\pi097 & w1091 ) | ( \pi098 & w1091 ) ;
  assign w1227 = ( ~\pi096 & \pi098 ) | ( ~\pi096 & w1226 ) | ( \pi098 & w1226 ) ;
  assign w1228 = ( ~\pi098 & w1091 ) | ( ~\pi098 & w1225 ) | ( w1091 & w1225 ) ;
  assign w1229 = w1227 & w1228 ;
  assign w1230 = ( w1077 & w1081 ) | ( w1077 & ~w1088 ) | ( w1081 & ~w1088 ) ;
  assign w1231 = \pi097 & ~w1230 ;
  assign w1232 = \pi096 | \pi098 ;
  assign w1233 = ( ~w1230 & w1231 ) | ( ~w1230 & w1232 ) | ( w1231 & w1232 ) ;
  assign w1234 = ~w1088 & w1233 ;
  assign w1235 = ~w1075 & w1234 ;
  assign w1236 = ( \pi098 & w1225 ) | ( \pi098 & ~w1234 ) | ( w1225 & ~w1234 ) ;
  assign w1237 = w1235 & ~w1236 ;
  assign w1238 = ~\pi098 & w1225 ;
  assign w1239 = \pi099 ^ w1238 ;
  assign w1240 = w1237 | w1239 ;
  assign w1241 = ( w965 & w1229 ) | ( w965 & ~w1240 ) | ( w1229 & ~w1240 ) ;
  assign w1242 = w965 & w1241 ;
  assign w1243 = ( ~w965 & w1229 ) | ( ~w965 & w1240 ) | ( w1229 & w1240 ) ;
  assign w1244 = ~w1229 & w1243 ;
  assign w1245 = w1091 & ~w1222 ;
  assign w1246 = ~w1211 & w1245 ;
  assign w1247 = ~w1224 & w1246 ;
  assign w1248 = \pi099 & w1225 ;
  assign w1249 = ( \pi098 & w1225 ) | ( \pi098 & ~w1248 ) | ( w1225 & ~w1248 ) ;
  assign w1250 = ( ~\pi098 & w1247 ) | ( ~\pi098 & w1249 ) | ( w1247 & w1249 ) ;
  assign w1251 = \pi100 ^ w1250 ;
  assign w1252 = w1244 | w1251 ;
  assign w1253 = ( w847 & w1242 ) | ( w847 & ~w1252 ) | ( w1242 & ~w1252 ) ;
  assign w1254 = w847 & w1253 ;
  assign w1255 = ( w1095 & ~w1103 ) | ( w1095 & w1225 ) | ( ~w1103 & w1225 ) ;
  assign w1256 = ~w1095 & w1255 ;
  assign w1257 = \pi101 ^ w1256 ;
  assign w1258 = w1104 ^ w1257 ;
  assign w1259 = ( ~w847 & w1242 ) | ( ~w847 & w1252 ) | ( w1242 & w1252 ) ;
  assign w1260 = ~w1242 & w1259 ;
  assign w1261 = w1258 | w1260 ;
  assign w1262 = ( w737 & w1254 ) | ( w737 & ~w1261 ) | ( w1254 & ~w1261 ) ;
  assign w1263 = w737 & w1262 ;
  assign w1264 = w1108 | w1110 ;
  assign w1265 = w1225 & ~w1264 ;
  assign w1266 = w1117 ^ w1265 ;
  assign w1267 = ( ~w737 & w1254 ) | ( ~w737 & w1261 ) | ( w1254 & w1261 ) ;
  assign w1268 = ~w1254 & w1267 ;
  assign w1269 = w1266 | w1268 ;
  assign w1270 = ( w635 & w1263 ) | ( w635 & ~w1269 ) | ( w1263 & ~w1269 ) ;
  assign w1271 = w635 & w1270 ;
  assign w1272 = w1120 | w1126 ;
  assign w1273 = w1225 & ~w1272 ;
  assign w1274 = w1124 ^ w1273 ;
  assign w1275 = ( ~w635 & w1263 ) | ( ~w635 & w1269 ) | ( w1263 & w1269 ) ;
  assign w1276 = ~w1263 & w1275 ;
  assign w1277 = w1274 | w1276 ;
  assign w1278 = ( w541 & w1271 ) | ( w541 & ~w1277 ) | ( w1271 & ~w1277 ) ;
  assign w1279 = w541 & w1278 ;
  assign w1280 = w1129 | w1134 ;
  assign w1281 = w1225 & ~w1280 ;
  assign w1282 = w1132 ^ w1281 ;
  assign w1283 = ( ~w541 & w1271 ) | ( ~w541 & w1277 ) | ( w1271 & w1277 ) ;
  assign w1284 = ~w1271 & w1283 ;
  assign w1285 = w1282 | w1284 ;
  assign w1286 = ( w455 & w1279 ) | ( w455 & ~w1285 ) | ( w1279 & ~w1285 ) ;
  assign w1287 = w455 & w1286 ;
  assign w1288 = w1137 | w1142 ;
  assign w1289 = w1225 & ~w1288 ;
  assign w1290 = w1140 ^ w1289 ;
  assign w1291 = ( ~w455 & w1279 ) | ( ~w455 & w1285 ) | ( w1279 & w1285 ) ;
  assign w1292 = ~w1279 & w1291 ;
  assign w1293 = w1290 | w1292 ;
  assign w1294 = ( w377 & w1287 ) | ( w377 & ~w1293 ) | ( w1287 & ~w1293 ) ;
  assign w1295 = w377 & w1294 ;
  assign w1296 = w1145 | w1150 ;
  assign w1297 = w1225 & ~w1296 ;
  assign w1298 = w1148 ^ w1297 ;
  assign w1299 = ( ~w377 & w1287 ) | ( ~w377 & w1293 ) | ( w1287 & w1293 ) ;
  assign w1300 = ~w1287 & w1299 ;
  assign w1301 = w1298 | w1300 ;
  assign w1302 = ( w307 & w1295 ) | ( w307 & ~w1301 ) | ( w1295 & ~w1301 ) ;
  assign w1303 = w307 & w1302 ;
  assign w1304 = w1153 | w1158 ;
  assign w1305 = w1225 & ~w1304 ;
  assign w1306 = w1156 ^ w1305 ;
  assign w1307 = ( ~w307 & w1295 ) | ( ~w307 & w1301 ) | ( w1295 & w1301 ) ;
  assign w1308 = ~w1295 & w1307 ;
  assign w1309 = w1306 | w1308 ;
  assign w1310 = ( w246 & w1303 ) | ( w246 & ~w1309 ) | ( w1303 & ~w1309 ) ;
  assign w1311 = w246 & w1310 ;
  assign w1312 = w1161 | w1166 ;
  assign w1313 = w1225 & ~w1312 ;
  assign w1314 = w1164 ^ w1313 ;
  assign w1315 = ( ~w246 & w1303 ) | ( ~w246 & w1309 ) | ( w1303 & w1309 ) ;
  assign w1316 = ~w1303 & w1315 ;
  assign w1317 = w1314 | w1316 ;
  assign w1318 = ( w185 & w1311 ) | ( w185 & ~w1317 ) | ( w1311 & ~w1317 ) ;
  assign w1319 = w185 & w1318 ;
  assign w1320 = w1169 | w1174 ;
  assign w1321 = w1225 & ~w1320 ;
  assign w1322 = w1172 ^ w1321 ;
  assign w1323 = ( ~w185 & w1311 ) | ( ~w185 & w1317 ) | ( w1311 & w1317 ) ;
  assign w1324 = ~w1311 & w1323 ;
  assign w1325 = w1322 | w1324 ;
  assign w1326 = ( w145 & w1319 ) | ( w145 & ~w1325 ) | ( w1319 & ~w1325 ) ;
  assign w1327 = w145 & w1326 ;
  assign w1328 = w1177 | w1182 ;
  assign w1329 = w1225 & ~w1328 ;
  assign w1330 = w1180 ^ w1329 ;
  assign w1331 = ( ~w145 & w1319 ) | ( ~w145 & w1325 ) | ( w1319 & w1325 ) ;
  assign w1332 = ~w1319 & w1331 ;
  assign w1333 = w1330 | w1332 ;
  assign w1334 = ( w132 & w1327 ) | ( w132 & ~w1333 ) | ( w1327 & ~w1333 ) ;
  assign w1335 = w132 & w1334 ;
  assign w1336 = w1185 | w1190 ;
  assign w1337 = w1225 & ~w1336 ;
  assign w1338 = w1188 ^ w1337 ;
  assign w1339 = ( ~w132 & w1327 ) | ( ~w132 & w1333 ) | ( w1327 & w1333 ) ;
  assign w1340 = ~w1327 & w1339 ;
  assign w1341 = w1338 | w1340 ;
  assign w1342 = ~w1335 & w1341 ;
  assign w1343 = w1193 | w1198 ;
  assign w1344 = w1225 & ~w1343 ;
  assign w1345 = w1196 ^ w1344 ;
  assign w1346 = ( ~w1211 & w1342 ) | ( ~w1211 & w1345 ) | ( w1342 & w1345 ) ;
  assign w1347 = w1200 & ~w1346 ;
  assign w1348 = ~w1203 & w1225 ;
  assign w1349 = ( w1346 & ~w1347 ) | ( w1346 & w1348 ) | ( ~w1347 & w1348 ) ;
  assign w1350 = w1211 | w1349 ;
  assign w1351 = ~w129 & w1350 ;
  assign w1352 = ( w1335 & w1341 ) | ( w1335 & w1345 ) | ( w1341 & w1345 ) ;
  assign w1353 = ~w1335 & w1352 ;
  assign w1354 = ( w129 & w1200 ) | ( w129 & w1203 ) | ( w1200 & w1203 ) ;
  assign w1355 = ( w1203 & ~w1225 ) | ( w1203 & w1354 ) | ( ~w1225 & w1354 ) ;
  assign w1356 = w1200 & w1355 ;
  assign w1357 = w1354 ^ w1356 ;
  assign w1358 = ( w1059 & w1061 ) | ( w1059 & w1091 ) | ( w1061 & w1091 ) ;
  assign w1359 = w1091 & ~w1358 ;
  assign w1360 = w1064 ^ w1359 ;
  assign w1361 = ( ~w1215 & w1222 ) | ( ~w1215 & w1360 ) | ( w1222 & w1360 ) ;
  assign w1362 = ~w1222 & w1361 ;
  assign w1363 = ( ~w1209 & w1211 ) | ( ~w1209 & w1362 ) | ( w1211 & w1362 ) ;
  assign w1364 = ~w1211 & w1363 ;
  assign w1365 = w1353 | w1364 ;
  assign w1366 = ( w1351 & ~w1353 ) | ( w1351 & w1357 ) | ( ~w1353 & w1357 ) ;
  assign w1367 = w1365 | w1366 ;
  assign w1368 = ( ~\pi095 & \pi096 ) | ( ~\pi095 & w1225 ) | ( \pi096 & w1225 ) ;
  assign w1369 = ( ~\pi094 & \pi096 ) | ( ~\pi094 & w1368 ) | ( \pi096 & w1368 ) ;
  assign w1370 = ( ~\pi096 & w1225 ) | ( ~\pi096 & w1367 ) | ( w1225 & w1367 ) ;
  assign w1371 = w1369 & w1370 ;
  assign w1372 = ( w1211 & w1215 ) | ( w1211 & ~w1222 ) | ( w1215 & ~w1222 ) ;
  assign w1373 = \pi095 & ~w1372 ;
  assign w1374 = \pi094 | \pi096 ;
  assign w1375 = ( ~w1372 & w1373 ) | ( ~w1372 & w1374 ) | ( w1373 & w1374 ) ;
  assign w1376 = ~w1222 & w1375 ;
  assign w1377 = ~w1209 & w1376 ;
  assign w1378 = ( \pi096 & w1367 ) | ( \pi096 & ~w1376 ) | ( w1367 & ~w1376 ) ;
  assign w1379 = w1377 & ~w1378 ;
  assign w1380 = ~\pi096 & w1367 ;
  assign w1381 = \pi097 ^ w1380 ;
  assign w1382 = w1379 | w1381 ;
  assign w1383 = ( w1091 & w1371 ) | ( w1091 & ~w1382 ) | ( w1371 & ~w1382 ) ;
  assign w1384 = w1091 & w1383 ;
  assign w1385 = ( ~w1091 & w1371 ) | ( ~w1091 & w1382 ) | ( w1371 & w1382 ) ;
  assign w1386 = ~w1371 & w1385 ;
  assign w1387 = w1225 & ~w1364 ;
  assign w1388 = ~w1353 & w1387 ;
  assign w1389 = ~w1366 & w1388 ;
  assign w1390 = \pi097 & w1367 ;
  assign w1391 = ( \pi096 & w1367 ) | ( \pi096 & ~w1390 ) | ( w1367 & ~w1390 ) ;
  assign w1392 = ( ~\pi096 & w1389 ) | ( ~\pi096 & w1391 ) | ( w1389 & w1391 ) ;
  assign w1393 = \pi098 ^ w1392 ;
  assign w1394 = w1386 | w1393 ;
  assign w1395 = ( w965 & w1384 ) | ( w965 & ~w1394 ) | ( w1384 & ~w1394 ) ;
  assign w1396 = w965 & w1395 ;
  assign w1397 = ( w1229 & ~w1237 ) | ( w1229 & w1367 ) | ( ~w1237 & w1367 ) ;
  assign w1398 = ~w1229 & w1397 ;
  assign w1399 = \pi099 ^ w1398 ;
  assign w1400 = w1238 ^ w1399 ;
  assign w1401 = ( ~w965 & w1384 ) | ( ~w965 & w1394 ) | ( w1384 & w1394 ) ;
  assign w1402 = ~w1384 & w1401 ;
  assign w1403 = w1400 | w1402 ;
  assign w1404 = ( w847 & w1396 ) | ( w847 & ~w1403 ) | ( w1396 & ~w1403 ) ;
  assign w1405 = w847 & w1404 ;
  assign w1406 = w1242 | w1244 ;
  assign w1407 = w1367 & ~w1406 ;
  assign w1408 = w1251 ^ w1407 ;
  assign w1409 = ( ~w847 & w1396 ) | ( ~w847 & w1403 ) | ( w1396 & w1403 ) ;
  assign w1410 = ~w1396 & w1409 ;
  assign w1411 = w1408 | w1410 ;
  assign w1412 = ( w737 & w1405 ) | ( w737 & ~w1411 ) | ( w1405 & ~w1411 ) ;
  assign w1413 = w737 & w1412 ;
  assign w1414 = w1254 | w1260 ;
  assign w1415 = w1367 & ~w1414 ;
  assign w1416 = w1258 ^ w1415 ;
  assign w1417 = ( ~w737 & w1405 ) | ( ~w737 & w1411 ) | ( w1405 & w1411 ) ;
  assign w1418 = ~w1405 & w1417 ;
  assign w1419 = w1416 | w1418 ;
  assign w1420 = ( w635 & w1413 ) | ( w635 & ~w1419 ) | ( w1413 & ~w1419 ) ;
  assign w1421 = w635 & w1420 ;
  assign w1422 = w1263 | w1268 ;
  assign w1423 = w1367 & ~w1422 ;
  assign w1424 = w1266 ^ w1423 ;
  assign w1425 = ( ~w635 & w1413 ) | ( ~w635 & w1419 ) | ( w1413 & w1419 ) ;
  assign w1426 = ~w1413 & w1425 ;
  assign w1427 = w1424 | w1426 ;
  assign w1428 = ( w541 & w1421 ) | ( w541 & ~w1427 ) | ( w1421 & ~w1427 ) ;
  assign w1429 = w541 & w1428 ;
  assign w1430 = w1271 | w1276 ;
  assign w1431 = w1367 & ~w1430 ;
  assign w1432 = w1274 ^ w1431 ;
  assign w1433 = ( ~w541 & w1421 ) | ( ~w541 & w1427 ) | ( w1421 & w1427 ) ;
  assign w1434 = ~w1421 & w1433 ;
  assign w1435 = w1432 | w1434 ;
  assign w1436 = ( w455 & w1429 ) | ( w455 & ~w1435 ) | ( w1429 & ~w1435 ) ;
  assign w1437 = w455 & w1436 ;
  assign w1438 = w1279 | w1284 ;
  assign w1439 = w1367 & ~w1438 ;
  assign w1440 = w1282 ^ w1439 ;
  assign w1441 = ( ~w455 & w1429 ) | ( ~w455 & w1435 ) | ( w1429 & w1435 ) ;
  assign w1442 = ~w1429 & w1441 ;
  assign w1443 = w1440 | w1442 ;
  assign w1444 = ( w377 & w1437 ) | ( w377 & ~w1443 ) | ( w1437 & ~w1443 ) ;
  assign w1445 = w377 & w1444 ;
  assign w1446 = w1287 | w1292 ;
  assign w1447 = w1367 & ~w1446 ;
  assign w1448 = w1290 ^ w1447 ;
  assign w1449 = ( ~w377 & w1437 ) | ( ~w377 & w1443 ) | ( w1437 & w1443 ) ;
  assign w1450 = ~w1437 & w1449 ;
  assign w1451 = w1448 | w1450 ;
  assign w1452 = ( w307 & w1445 ) | ( w307 & ~w1451 ) | ( w1445 & ~w1451 ) ;
  assign w1453 = w307 & w1452 ;
  assign w1454 = w1295 | w1300 ;
  assign w1455 = w1367 & ~w1454 ;
  assign w1456 = w1298 ^ w1455 ;
  assign w1457 = ( ~w307 & w1445 ) | ( ~w307 & w1451 ) | ( w1445 & w1451 ) ;
  assign w1458 = ~w1445 & w1457 ;
  assign w1459 = w1456 | w1458 ;
  assign w1460 = ( w246 & w1453 ) | ( w246 & ~w1459 ) | ( w1453 & ~w1459 ) ;
  assign w1461 = w246 & w1460 ;
  assign w1462 = w1303 | w1308 ;
  assign w1463 = w1367 & ~w1462 ;
  assign w1464 = w1306 ^ w1463 ;
  assign w1465 = ( ~w246 & w1453 ) | ( ~w246 & w1459 ) | ( w1453 & w1459 ) ;
  assign w1466 = ~w1453 & w1465 ;
  assign w1467 = w1464 | w1466 ;
  assign w1468 = ( w185 & w1461 ) | ( w185 & ~w1467 ) | ( w1461 & ~w1467 ) ;
  assign w1469 = w185 & w1468 ;
  assign w1470 = w1311 | w1316 ;
  assign w1471 = w1367 & ~w1470 ;
  assign w1472 = w1314 ^ w1471 ;
  assign w1473 = ( ~w185 & w1461 ) | ( ~w185 & w1467 ) | ( w1461 & w1467 ) ;
  assign w1474 = ~w1461 & w1473 ;
  assign w1475 = w1472 | w1474 ;
  assign w1476 = ( w145 & w1469 ) | ( w145 & ~w1475 ) | ( w1469 & ~w1475 ) ;
  assign w1477 = w145 & w1476 ;
  assign w1478 = w1319 | w1324 ;
  assign w1479 = w1367 & ~w1478 ;
  assign w1480 = w1322 ^ w1479 ;
  assign w1481 = ( ~w145 & w1469 ) | ( ~w145 & w1475 ) | ( w1469 & w1475 ) ;
  assign w1482 = ~w1469 & w1481 ;
  assign w1483 = w1480 | w1482 ;
  assign w1484 = ( w132 & w1477 ) | ( w132 & ~w1483 ) | ( w1477 & ~w1483 ) ;
  assign w1485 = w132 & w1484 ;
  assign w1486 = w1327 | w1332 ;
  assign w1487 = w1367 & ~w1486 ;
  assign w1488 = w1330 ^ w1487 ;
  assign w1489 = ( ~w132 & w1477 ) | ( ~w132 & w1483 ) | ( w1477 & w1483 ) ;
  assign w1490 = ~w1477 & w1489 ;
  assign w1491 = w1488 | w1490 ;
  assign w1492 = ~w1485 & w1491 ;
  assign w1493 = w1335 | w1340 ;
  assign w1494 = w1367 & ~w1493 ;
  assign w1495 = w1338 ^ w1494 ;
  assign w1496 = ( ~w1353 & w1492 ) | ( ~w1353 & w1495 ) | ( w1492 & w1495 ) ;
  assign w1497 = w1342 & ~w1496 ;
  assign w1498 = ~w1345 & w1367 ;
  assign w1499 = ( w1496 & ~w1497 ) | ( w1496 & w1498 ) | ( ~w1497 & w1498 ) ;
  assign w1500 = w1353 | w1499 ;
  assign w1501 = ~w129 & w1500 ;
  assign w1502 = ( w1485 & w1491 ) | ( w1485 & w1495 ) | ( w1491 & w1495 ) ;
  assign w1503 = ~w1485 & w1502 ;
  assign w1504 = ( w129 & w1342 ) | ( w129 & w1345 ) | ( w1342 & w1345 ) ;
  assign w1505 = ( w1345 & ~w1367 ) | ( w1345 & w1504 ) | ( ~w1367 & w1504 ) ;
  assign w1506 = w1342 & w1505 ;
  assign w1507 = w1504 ^ w1506 ;
  assign w1508 = ( w1193 & w1198 ) | ( w1193 & w1225 ) | ( w1198 & w1225 ) ;
  assign w1509 = w1225 & ~w1508 ;
  assign w1510 = w1196 ^ w1509 ;
  assign w1511 = ( ~w1357 & w1364 ) | ( ~w1357 & w1510 ) | ( w1364 & w1510 ) ;
  assign w1512 = ~w1364 & w1511 ;
  assign w1513 = ( ~w1351 & w1353 ) | ( ~w1351 & w1512 ) | ( w1353 & w1512 ) ;
  assign w1514 = ~w1353 & w1513 ;
  assign w1515 = w1503 | w1514 ;
  assign w1516 = ( w1501 & ~w1503 ) | ( w1501 & w1507 ) | ( ~w1503 & w1507 ) ;
  assign w1517 = w1515 | w1516 ;
  assign w1518 = ( ~\pi093 & \pi094 ) | ( ~\pi093 & w1367 ) | ( \pi094 & w1367 ) ;
  assign w1519 = ( ~\pi092 & \pi094 ) | ( ~\pi092 & w1518 ) | ( \pi094 & w1518 ) ;
  assign w1520 = ( ~\pi094 & w1367 ) | ( ~\pi094 & w1517 ) | ( w1367 & w1517 ) ;
  assign w1521 = w1519 & w1520 ;
  assign w1522 = ( w1353 & w1357 ) | ( w1353 & ~w1364 ) | ( w1357 & ~w1364 ) ;
  assign w1523 = \pi093 & ~w1522 ;
  assign w1524 = \pi092 | \pi094 ;
  assign w1525 = ( ~w1522 & w1523 ) | ( ~w1522 & w1524 ) | ( w1523 & w1524 ) ;
  assign w1526 = ~w1364 & w1525 ;
  assign w1527 = ~w1351 & w1526 ;
  assign w1528 = ( \pi094 & w1517 ) | ( \pi094 & ~w1526 ) | ( w1517 & ~w1526 ) ;
  assign w1529 = w1527 & ~w1528 ;
  assign w1530 = ~\pi094 & w1517 ;
  assign w1531 = \pi095 ^ w1530 ;
  assign w1532 = w1529 | w1531 ;
  assign w1533 = ( w1225 & w1521 ) | ( w1225 & ~w1532 ) | ( w1521 & ~w1532 ) ;
  assign w1534 = w1225 & w1533 ;
  assign w1535 = ( ~w1225 & w1521 ) | ( ~w1225 & w1532 ) | ( w1521 & w1532 ) ;
  assign w1536 = ~w1521 & w1535 ;
  assign w1537 = w1367 & ~w1514 ;
  assign w1538 = ~w1503 & w1537 ;
  assign w1539 = ~w1516 & w1538 ;
  assign w1540 = \pi095 & w1517 ;
  assign w1541 = ( \pi094 & w1517 ) | ( \pi094 & ~w1540 ) | ( w1517 & ~w1540 ) ;
  assign w1542 = ( ~\pi094 & w1539 ) | ( ~\pi094 & w1541 ) | ( w1539 & w1541 ) ;
  assign w1543 = \pi096 ^ w1542 ;
  assign w1544 = w1536 | w1543 ;
  assign w1545 = ( w1091 & w1534 ) | ( w1091 & ~w1544 ) | ( w1534 & ~w1544 ) ;
  assign w1546 = w1091 & w1545 ;
  assign w1547 = ( ~w1091 & w1534 ) | ( ~w1091 & w1544 ) | ( w1534 & w1544 ) ;
  assign w1548 = ~w1534 & w1547 ;
  assign w1549 = ( w1371 & ~w1379 ) | ( w1371 & w1517 ) | ( ~w1379 & w1517 ) ;
  assign w1550 = ~w1371 & w1549 ;
  assign w1551 = \pi097 ^ w1550 ;
  assign w1552 = w1380 ^ w1551 ;
  assign w1553 = w1548 | w1552 ;
  assign w1554 = ( w965 & w1546 ) | ( w965 & ~w1553 ) | ( w1546 & ~w1553 ) ;
  assign w1555 = w965 & w1554 ;
  assign w1556 = w1384 | w1386 ;
  assign w1557 = w1517 & ~w1556 ;
  assign w1558 = w1393 ^ w1557 ;
  assign w1559 = ( ~w965 & w1546 ) | ( ~w965 & w1553 ) | ( w1546 & w1553 ) ;
  assign w1560 = ~w1546 & w1559 ;
  assign w1561 = w1558 | w1560 ;
  assign w1562 = ( w847 & w1555 ) | ( w847 & ~w1561 ) | ( w1555 & ~w1561 ) ;
  assign w1563 = w847 & w1562 ;
  assign w1564 = w1396 | w1402 ;
  assign w1565 = w1517 & ~w1564 ;
  assign w1566 = w1400 ^ w1565 ;
  assign w1567 = ( ~w847 & w1555 ) | ( ~w847 & w1561 ) | ( w1555 & w1561 ) ;
  assign w1568 = ~w1555 & w1567 ;
  assign w1569 = w1566 | w1568 ;
  assign w1570 = ( w737 & w1563 ) | ( w737 & ~w1569 ) | ( w1563 & ~w1569 ) ;
  assign w1571 = w737 & w1570 ;
  assign w1572 = w1405 | w1410 ;
  assign w1573 = w1517 & ~w1572 ;
  assign w1574 = w1408 ^ w1573 ;
  assign w1575 = ( ~w737 & w1563 ) | ( ~w737 & w1569 ) | ( w1563 & w1569 ) ;
  assign w1576 = ~w1563 & w1575 ;
  assign w1577 = w1574 | w1576 ;
  assign w1578 = ( w635 & w1571 ) | ( w635 & ~w1577 ) | ( w1571 & ~w1577 ) ;
  assign w1579 = w635 & w1578 ;
  assign w1580 = w1413 | w1418 ;
  assign w1581 = w1517 & ~w1580 ;
  assign w1582 = w1416 ^ w1581 ;
  assign w1583 = ( ~w635 & w1571 ) | ( ~w635 & w1577 ) | ( w1571 & w1577 ) ;
  assign w1584 = ~w1571 & w1583 ;
  assign w1585 = w1582 | w1584 ;
  assign w1586 = ( w541 & w1579 ) | ( w541 & ~w1585 ) | ( w1579 & ~w1585 ) ;
  assign w1587 = w541 & w1586 ;
  assign w1588 = w1421 | w1426 ;
  assign w1589 = w1517 & ~w1588 ;
  assign w1590 = w1424 ^ w1589 ;
  assign w1591 = ( ~w541 & w1579 ) | ( ~w541 & w1585 ) | ( w1579 & w1585 ) ;
  assign w1592 = ~w1579 & w1591 ;
  assign w1593 = w1590 | w1592 ;
  assign w1594 = ( w455 & w1587 ) | ( w455 & ~w1593 ) | ( w1587 & ~w1593 ) ;
  assign w1595 = w455 & w1594 ;
  assign w1596 = w1429 | w1434 ;
  assign w1597 = w1517 & ~w1596 ;
  assign w1598 = w1432 ^ w1597 ;
  assign w1599 = ( ~w455 & w1587 ) | ( ~w455 & w1593 ) | ( w1587 & w1593 ) ;
  assign w1600 = ~w1587 & w1599 ;
  assign w1601 = w1598 | w1600 ;
  assign w1602 = ( w377 & w1595 ) | ( w377 & ~w1601 ) | ( w1595 & ~w1601 ) ;
  assign w1603 = w377 & w1602 ;
  assign w1604 = w1437 | w1442 ;
  assign w1605 = w1517 & ~w1604 ;
  assign w1606 = w1440 ^ w1605 ;
  assign w1607 = ( ~w377 & w1595 ) | ( ~w377 & w1601 ) | ( w1595 & w1601 ) ;
  assign w1608 = ~w1595 & w1607 ;
  assign w1609 = w1606 | w1608 ;
  assign w1610 = ( w307 & w1603 ) | ( w307 & ~w1609 ) | ( w1603 & ~w1609 ) ;
  assign w1611 = w307 & w1610 ;
  assign w1612 = w1445 | w1450 ;
  assign w1613 = w1517 & ~w1612 ;
  assign w1614 = w1448 ^ w1613 ;
  assign w1615 = ( ~w307 & w1603 ) | ( ~w307 & w1609 ) | ( w1603 & w1609 ) ;
  assign w1616 = ~w1603 & w1615 ;
  assign w1617 = w1614 | w1616 ;
  assign w1618 = ( w246 & w1611 ) | ( w246 & ~w1617 ) | ( w1611 & ~w1617 ) ;
  assign w1619 = w246 & w1618 ;
  assign w1620 = w1453 | w1458 ;
  assign w1621 = w1517 & ~w1620 ;
  assign w1622 = w1456 ^ w1621 ;
  assign w1623 = ( ~w246 & w1611 ) | ( ~w246 & w1617 ) | ( w1611 & w1617 ) ;
  assign w1624 = ~w1611 & w1623 ;
  assign w1625 = w1622 | w1624 ;
  assign w1626 = ( w185 & w1619 ) | ( w185 & ~w1625 ) | ( w1619 & ~w1625 ) ;
  assign w1627 = w185 & w1626 ;
  assign w1628 = w1461 | w1466 ;
  assign w1629 = w1517 & ~w1628 ;
  assign w1630 = w1464 ^ w1629 ;
  assign w1631 = ( ~w185 & w1619 ) | ( ~w185 & w1625 ) | ( w1619 & w1625 ) ;
  assign w1632 = ~w1619 & w1631 ;
  assign w1633 = w1630 | w1632 ;
  assign w1634 = ( w145 & w1627 ) | ( w145 & ~w1633 ) | ( w1627 & ~w1633 ) ;
  assign w1635 = w145 & w1634 ;
  assign w1636 = w1469 | w1474 ;
  assign w1637 = w1517 & ~w1636 ;
  assign w1638 = w1472 ^ w1637 ;
  assign w1639 = ( ~w145 & w1627 ) | ( ~w145 & w1633 ) | ( w1627 & w1633 ) ;
  assign w1640 = ~w1627 & w1639 ;
  assign w1641 = w1638 | w1640 ;
  assign w1642 = ( w132 & w1635 ) | ( w132 & ~w1641 ) | ( w1635 & ~w1641 ) ;
  assign w1643 = w132 & w1642 ;
  assign w1644 = w1477 | w1482 ;
  assign w1645 = w1517 & ~w1644 ;
  assign w1646 = w1480 ^ w1645 ;
  assign w1647 = ( ~w132 & w1635 ) | ( ~w132 & w1641 ) | ( w1635 & w1641 ) ;
  assign w1648 = ~w1635 & w1647 ;
  assign w1649 = w1646 | w1648 ;
  assign w1650 = ~w1643 & w1649 ;
  assign w1651 = w1485 | w1490 ;
  assign w1652 = w1517 & ~w1651 ;
  assign w1653 = w1488 ^ w1652 ;
  assign w1654 = ( ~w1503 & w1650 ) | ( ~w1503 & w1653 ) | ( w1650 & w1653 ) ;
  assign w1655 = w1492 & ~w1654 ;
  assign w1656 = ~w1495 & w1517 ;
  assign w1657 = ( w1654 & ~w1655 ) | ( w1654 & w1656 ) | ( ~w1655 & w1656 ) ;
  assign w1658 = w1503 | w1657 ;
  assign w1659 = ~w129 & w1658 ;
  assign w1660 = ( w1643 & w1649 ) | ( w1643 & w1653 ) | ( w1649 & w1653 ) ;
  assign w1661 = ~w1643 & w1660 ;
  assign w1662 = ( w129 & w1492 ) | ( w129 & w1495 ) | ( w1492 & w1495 ) ;
  assign w1663 = ( w1495 & ~w1517 ) | ( w1495 & w1662 ) | ( ~w1517 & w1662 ) ;
  assign w1664 = w1492 & w1663 ;
  assign w1665 = w1662 ^ w1664 ;
  assign w1666 = ( w1335 & w1340 ) | ( w1335 & w1367 ) | ( w1340 & w1367 ) ;
  assign w1667 = w1367 & ~w1666 ;
  assign w1668 = w1338 ^ w1667 ;
  assign w1669 = ( ~w1507 & w1514 ) | ( ~w1507 & w1668 ) | ( w1514 & w1668 ) ;
  assign w1670 = ~w1514 & w1669 ;
  assign w1671 = ( ~w1501 & w1503 ) | ( ~w1501 & w1670 ) | ( w1503 & w1670 ) ;
  assign w1672 = ~w1503 & w1671 ;
  assign w1673 = w1661 | w1672 ;
  assign w1674 = ( w1659 & ~w1661 ) | ( w1659 & w1665 ) | ( ~w1661 & w1665 ) ;
  assign w1675 = w1673 | w1674 ;
  assign w1676 = ( ~\pi091 & \pi092 ) | ( ~\pi091 & w1517 ) | ( \pi092 & w1517 ) ;
  assign w1677 = ( ~\pi090 & \pi092 ) | ( ~\pi090 & w1676 ) | ( \pi092 & w1676 ) ;
  assign w1678 = ( ~\pi092 & w1517 ) | ( ~\pi092 & w1675 ) | ( w1517 & w1675 ) ;
  assign w1679 = w1677 & w1678 ;
  assign w1680 = ( w1503 & w1507 ) | ( w1503 & ~w1514 ) | ( w1507 & ~w1514 ) ;
  assign w1681 = \pi091 & ~w1680 ;
  assign w1682 = \pi090 | \pi092 ;
  assign w1683 = ( ~w1680 & w1681 ) | ( ~w1680 & w1682 ) | ( w1681 & w1682 ) ;
  assign w1684 = ~w1514 & w1683 ;
  assign w1685 = ~w1501 & w1684 ;
  assign w1686 = ( \pi092 & w1675 ) | ( \pi092 & ~w1684 ) | ( w1675 & ~w1684 ) ;
  assign w1687 = w1685 & ~w1686 ;
  assign w1688 = ~\pi092 & w1675 ;
  assign w1689 = \pi093 ^ w1688 ;
  assign w1690 = w1687 | w1689 ;
  assign w1691 = ( w1367 & w1679 ) | ( w1367 & ~w1690 ) | ( w1679 & ~w1690 ) ;
  assign w1692 = w1367 & w1691 ;
  assign w1693 = ( ~w1367 & w1679 ) | ( ~w1367 & w1690 ) | ( w1679 & w1690 ) ;
  assign w1694 = ~w1679 & w1693 ;
  assign w1695 = w1517 & ~w1672 ;
  assign w1696 = ~w1661 & w1695 ;
  assign w1697 = ~w1674 & w1696 ;
  assign w1698 = \pi093 & w1675 ;
  assign w1699 = ( \pi092 & w1675 ) | ( \pi092 & ~w1698 ) | ( w1675 & ~w1698 ) ;
  assign w1700 = ( ~\pi092 & w1697 ) | ( ~\pi092 & w1699 ) | ( w1697 & w1699 ) ;
  assign w1701 = \pi094 ^ w1700 ;
  assign w1702 = w1694 | w1701 ;
  assign w1703 = ( w1225 & w1692 ) | ( w1225 & ~w1702 ) | ( w1692 & ~w1702 ) ;
  assign w1704 = w1225 & w1703 ;
  assign w1705 = ( w1521 & ~w1529 ) | ( w1521 & w1675 ) | ( ~w1529 & w1675 ) ;
  assign w1706 = ~w1521 & w1705 ;
  assign w1707 = \pi095 ^ w1706 ;
  assign w1708 = w1530 ^ w1707 ;
  assign w1709 = ( ~w1225 & w1692 ) | ( ~w1225 & w1702 ) | ( w1692 & w1702 ) ;
  assign w1710 = ~w1692 & w1709 ;
  assign w1711 = w1708 | w1710 ;
  assign w1712 = ( w1091 & w1704 ) | ( w1091 & ~w1711 ) | ( w1704 & ~w1711 ) ;
  assign w1713 = w1091 & w1712 ;
  assign w1714 = w1534 | w1536 ;
  assign w1715 = w1675 & ~w1714 ;
  assign w1716 = w1543 ^ w1715 ;
  assign w1717 = ( ~w1091 & w1704 ) | ( ~w1091 & w1711 ) | ( w1704 & w1711 ) ;
  assign w1718 = ~w1704 & w1717 ;
  assign w1719 = w1716 | w1718 ;
  assign w1720 = ( w965 & w1713 ) | ( w965 & ~w1719 ) | ( w1713 & ~w1719 ) ;
  assign w1721 = w965 & w1720 ;
  assign w1722 = ( ~w965 & w1713 ) | ( ~w965 & w1719 ) | ( w1713 & w1719 ) ;
  assign w1723 = ~w1713 & w1722 ;
  assign w1724 = w1546 | w1548 ;
  assign w1725 = w1675 & ~w1724 ;
  assign w1726 = w1552 ^ w1725 ;
  assign w1727 = w1723 | w1726 ;
  assign w1728 = ( w847 & w1721 ) | ( w847 & ~w1727 ) | ( w1721 & ~w1727 ) ;
  assign w1729 = w847 & w1728 ;
  assign w1730 = w1555 | w1560 ;
  assign w1731 = w1675 & ~w1730 ;
  assign w1732 = w1558 ^ w1731 ;
  assign w1733 = ( ~w847 & w1721 ) | ( ~w847 & w1727 ) | ( w1721 & w1727 ) ;
  assign w1734 = ~w1721 & w1733 ;
  assign w1735 = w1732 | w1734 ;
  assign w1736 = ( w737 & w1729 ) | ( w737 & ~w1735 ) | ( w1729 & ~w1735 ) ;
  assign w1737 = w737 & w1736 ;
  assign w1738 = w1563 | w1568 ;
  assign w1739 = w1675 & ~w1738 ;
  assign w1740 = w1566 ^ w1739 ;
  assign w1741 = ( ~w737 & w1729 ) | ( ~w737 & w1735 ) | ( w1729 & w1735 ) ;
  assign w1742 = ~w1729 & w1741 ;
  assign w1743 = w1740 | w1742 ;
  assign w1744 = ( w635 & w1737 ) | ( w635 & ~w1743 ) | ( w1737 & ~w1743 ) ;
  assign w1745 = w635 & w1744 ;
  assign w1746 = w1571 | w1576 ;
  assign w1747 = w1675 & ~w1746 ;
  assign w1748 = w1574 ^ w1747 ;
  assign w1749 = ( ~w635 & w1737 ) | ( ~w635 & w1743 ) | ( w1737 & w1743 ) ;
  assign w1750 = ~w1737 & w1749 ;
  assign w1751 = w1748 | w1750 ;
  assign w1752 = ( w541 & w1745 ) | ( w541 & ~w1751 ) | ( w1745 & ~w1751 ) ;
  assign w1753 = w541 & w1752 ;
  assign w1754 = w1579 | w1584 ;
  assign w1755 = w1675 & ~w1754 ;
  assign w1756 = w1582 ^ w1755 ;
  assign w1757 = ( ~w541 & w1745 ) | ( ~w541 & w1751 ) | ( w1745 & w1751 ) ;
  assign w1758 = ~w1745 & w1757 ;
  assign w1759 = w1756 | w1758 ;
  assign w1760 = ( w455 & w1753 ) | ( w455 & ~w1759 ) | ( w1753 & ~w1759 ) ;
  assign w1761 = w455 & w1760 ;
  assign w1762 = w1587 | w1592 ;
  assign w1763 = w1675 & ~w1762 ;
  assign w1764 = w1590 ^ w1763 ;
  assign w1765 = ( ~w455 & w1753 ) | ( ~w455 & w1759 ) | ( w1753 & w1759 ) ;
  assign w1766 = ~w1753 & w1765 ;
  assign w1767 = w1764 | w1766 ;
  assign w1768 = ( w377 & w1761 ) | ( w377 & ~w1767 ) | ( w1761 & ~w1767 ) ;
  assign w1769 = w377 & w1768 ;
  assign w1770 = w1595 | w1600 ;
  assign w1771 = w1675 & ~w1770 ;
  assign w1772 = w1598 ^ w1771 ;
  assign w1773 = ( ~w377 & w1761 ) | ( ~w377 & w1767 ) | ( w1761 & w1767 ) ;
  assign w1774 = ~w1761 & w1773 ;
  assign w1775 = w1772 | w1774 ;
  assign w1776 = ( w307 & w1769 ) | ( w307 & ~w1775 ) | ( w1769 & ~w1775 ) ;
  assign w1777 = w307 & w1776 ;
  assign w1778 = w1603 | w1608 ;
  assign w1779 = w1675 & ~w1778 ;
  assign w1780 = w1606 ^ w1779 ;
  assign w1781 = ( ~w307 & w1769 ) | ( ~w307 & w1775 ) | ( w1769 & w1775 ) ;
  assign w1782 = ~w1769 & w1781 ;
  assign w1783 = w1780 | w1782 ;
  assign w1784 = ( w246 & w1777 ) | ( w246 & ~w1783 ) | ( w1777 & ~w1783 ) ;
  assign w1785 = w246 & w1784 ;
  assign w1786 = w1611 | w1616 ;
  assign w1787 = w1675 & ~w1786 ;
  assign w1788 = w1614 ^ w1787 ;
  assign w1789 = ( ~w246 & w1777 ) | ( ~w246 & w1783 ) | ( w1777 & w1783 ) ;
  assign w1790 = ~w1777 & w1789 ;
  assign w1791 = w1788 | w1790 ;
  assign w1792 = ( w185 & w1785 ) | ( w185 & ~w1791 ) | ( w1785 & ~w1791 ) ;
  assign w1793 = w185 & w1792 ;
  assign w1794 = w1619 | w1624 ;
  assign w1795 = w1675 & ~w1794 ;
  assign w1796 = w1622 ^ w1795 ;
  assign w1797 = ( ~w185 & w1785 ) | ( ~w185 & w1791 ) | ( w1785 & w1791 ) ;
  assign w1798 = ~w1785 & w1797 ;
  assign w1799 = w1796 | w1798 ;
  assign w1800 = ( w145 & w1793 ) | ( w145 & ~w1799 ) | ( w1793 & ~w1799 ) ;
  assign w1801 = w145 & w1800 ;
  assign w1802 = w1627 | w1632 ;
  assign w1803 = w1675 & ~w1802 ;
  assign w1804 = w1630 ^ w1803 ;
  assign w1805 = ( ~w145 & w1793 ) | ( ~w145 & w1799 ) | ( w1793 & w1799 ) ;
  assign w1806 = ~w1793 & w1805 ;
  assign w1807 = w1804 | w1806 ;
  assign w1808 = ( w132 & w1801 ) | ( w132 & ~w1807 ) | ( w1801 & ~w1807 ) ;
  assign w1809 = w132 & w1808 ;
  assign w1810 = w1635 | w1640 ;
  assign w1811 = w1675 & ~w1810 ;
  assign w1812 = w1638 ^ w1811 ;
  assign w1813 = ( ~w132 & w1801 ) | ( ~w132 & w1807 ) | ( w1801 & w1807 ) ;
  assign w1814 = ~w1801 & w1813 ;
  assign w1815 = w1812 | w1814 ;
  assign w1816 = ~w1809 & w1815 ;
  assign w1817 = w1643 | w1648 ;
  assign w1818 = w1675 & ~w1817 ;
  assign w1819 = w1646 ^ w1818 ;
  assign w1820 = ( ~w1661 & w1816 ) | ( ~w1661 & w1819 ) | ( w1816 & w1819 ) ;
  assign w1821 = w1650 & ~w1820 ;
  assign w1822 = ~w1653 & w1675 ;
  assign w1823 = ( w1820 & ~w1821 ) | ( w1820 & w1822 ) | ( ~w1821 & w1822 ) ;
  assign w1824 = w1661 | w1823 ;
  assign w1825 = ~w129 & w1824 ;
  assign w1826 = ( w1809 & w1815 ) | ( w1809 & w1819 ) | ( w1815 & w1819 ) ;
  assign w1827 = ~w1809 & w1826 ;
  assign w1828 = ( w129 & w1650 ) | ( w129 & w1653 ) | ( w1650 & w1653 ) ;
  assign w1829 = ( w1653 & ~w1675 ) | ( w1653 & w1828 ) | ( ~w1675 & w1828 ) ;
  assign w1830 = w1650 & w1829 ;
  assign w1831 = w1828 ^ w1830 ;
  assign w1832 = ( w1485 & w1490 ) | ( w1485 & w1517 ) | ( w1490 & w1517 ) ;
  assign w1833 = w1517 & ~w1832 ;
  assign w1834 = w1488 ^ w1833 ;
  assign w1835 = ( ~w1665 & w1672 ) | ( ~w1665 & w1834 ) | ( w1672 & w1834 ) ;
  assign w1836 = ~w1672 & w1835 ;
  assign w1837 = ( ~w1659 & w1661 ) | ( ~w1659 & w1836 ) | ( w1661 & w1836 ) ;
  assign w1838 = ~w1661 & w1837 ;
  assign w1839 = w1827 | w1838 ;
  assign w1840 = ( w1825 & ~w1827 ) | ( w1825 & w1831 ) | ( ~w1827 & w1831 ) ;
  assign w1841 = w1839 | w1840 ;
  assign w1842 = ( ~\pi089 & \pi090 ) | ( ~\pi089 & w1675 ) | ( \pi090 & w1675 ) ;
  assign w1843 = ( ~\pi088 & \pi090 ) | ( ~\pi088 & w1842 ) | ( \pi090 & w1842 ) ;
  assign w1844 = ( ~\pi090 & w1675 ) | ( ~\pi090 & w1841 ) | ( w1675 & w1841 ) ;
  assign w1845 = w1843 & w1844 ;
  assign w1846 = ( w1661 & w1665 ) | ( w1661 & ~w1672 ) | ( w1665 & ~w1672 ) ;
  assign w1847 = \pi089 & ~w1846 ;
  assign w1848 = \pi088 | \pi090 ;
  assign w1849 = ( ~w1846 & w1847 ) | ( ~w1846 & w1848 ) | ( w1847 & w1848 ) ;
  assign w1850 = ~w1672 & w1849 ;
  assign w1851 = ~w1659 & w1850 ;
  assign w1852 = ( \pi090 & w1841 ) | ( \pi090 & ~w1850 ) | ( w1841 & ~w1850 ) ;
  assign w1853 = w1851 & ~w1852 ;
  assign w1854 = ~\pi090 & w1841 ;
  assign w1855 = \pi091 ^ w1854 ;
  assign w1856 = w1853 | w1855 ;
  assign w1857 = ( w1517 & w1845 ) | ( w1517 & ~w1856 ) | ( w1845 & ~w1856 ) ;
  assign w1858 = w1517 & w1857 ;
  assign w1859 = ( ~w1517 & w1845 ) | ( ~w1517 & w1856 ) | ( w1845 & w1856 ) ;
  assign w1860 = ~w1845 & w1859 ;
  assign w1861 = w1675 & ~w1838 ;
  assign w1862 = ~w1827 & w1861 ;
  assign w1863 = ~w1840 & w1862 ;
  assign w1864 = \pi091 & w1841 ;
  assign w1865 = ( \pi090 & w1841 ) | ( \pi090 & ~w1864 ) | ( w1841 & ~w1864 ) ;
  assign w1866 = ( ~\pi090 & w1863 ) | ( ~\pi090 & w1865 ) | ( w1863 & w1865 ) ;
  assign w1867 = \pi092 ^ w1866 ;
  assign w1868 = w1860 | w1867 ;
  assign w1869 = ( w1367 & w1858 ) | ( w1367 & ~w1868 ) | ( w1858 & ~w1868 ) ;
  assign w1870 = w1367 & w1869 ;
  assign w1871 = ( w1679 & ~w1687 ) | ( w1679 & w1841 ) | ( ~w1687 & w1841 ) ;
  assign w1872 = ~w1679 & w1871 ;
  assign w1873 = \pi093 ^ w1872 ;
  assign w1874 = w1688 ^ w1873 ;
  assign w1875 = ( ~w1367 & w1858 ) | ( ~w1367 & w1868 ) | ( w1858 & w1868 ) ;
  assign w1876 = ~w1858 & w1875 ;
  assign w1877 = w1874 | w1876 ;
  assign w1878 = ( w1225 & w1870 ) | ( w1225 & ~w1877 ) | ( w1870 & ~w1877 ) ;
  assign w1879 = w1225 & w1878 ;
  assign w1880 = w1692 | w1694 ;
  assign w1881 = w1841 & ~w1880 ;
  assign w1882 = w1701 ^ w1881 ;
  assign w1883 = ( ~w1225 & w1870 ) | ( ~w1225 & w1877 ) | ( w1870 & w1877 ) ;
  assign w1884 = ~w1870 & w1883 ;
  assign w1885 = w1882 | w1884 ;
  assign w1886 = ( w1091 & w1879 ) | ( w1091 & ~w1885 ) | ( w1879 & ~w1885 ) ;
  assign w1887 = w1091 & w1886 ;
  assign w1888 = w1704 | w1710 ;
  assign w1889 = w1841 & ~w1888 ;
  assign w1890 = w1708 ^ w1889 ;
  assign w1891 = ( ~w1091 & w1879 ) | ( ~w1091 & w1885 ) | ( w1879 & w1885 ) ;
  assign w1892 = ~w1879 & w1891 ;
  assign w1893 = w1890 | w1892 ;
  assign w1894 = ( w965 & w1887 ) | ( w965 & ~w1893 ) | ( w1887 & ~w1893 ) ;
  assign w1895 = w965 & w1894 ;
  assign w1896 = w1713 | w1718 ;
  assign w1897 = w1841 & ~w1896 ;
  assign w1898 = w1716 ^ w1897 ;
  assign w1899 = ( ~w965 & w1887 ) | ( ~w965 & w1893 ) | ( w1887 & w1893 ) ;
  assign w1900 = ~w1887 & w1899 ;
  assign w1901 = w1898 | w1900 ;
  assign w1902 = ( w847 & w1895 ) | ( w847 & ~w1901 ) | ( w1895 & ~w1901 ) ;
  assign w1903 = w847 & w1902 ;
  assign w1904 = ( ~w847 & w1895 ) | ( ~w847 & w1901 ) | ( w1895 & w1901 ) ;
  assign w1905 = ~w1895 & w1904 ;
  assign w1906 = w1721 | w1723 ;
  assign w1907 = w1841 & ~w1906 ;
  assign w1908 = w1726 ^ w1907 ;
  assign w1909 = w1905 | w1908 ;
  assign w1910 = ( w737 & w1903 ) | ( w737 & ~w1909 ) | ( w1903 & ~w1909 ) ;
  assign w1911 = w737 & w1910 ;
  assign w1912 = w1729 | w1734 ;
  assign w1913 = w1841 & ~w1912 ;
  assign w1914 = w1732 ^ w1913 ;
  assign w1915 = ( ~w737 & w1903 ) | ( ~w737 & w1909 ) | ( w1903 & w1909 ) ;
  assign w1916 = ~w1903 & w1915 ;
  assign w1917 = w1914 | w1916 ;
  assign w1918 = ( w635 & w1911 ) | ( w635 & ~w1917 ) | ( w1911 & ~w1917 ) ;
  assign w1919 = w635 & w1918 ;
  assign w1920 = w1737 | w1742 ;
  assign w1921 = w1841 & ~w1920 ;
  assign w1922 = w1740 ^ w1921 ;
  assign w1923 = ( ~w635 & w1911 ) | ( ~w635 & w1917 ) | ( w1911 & w1917 ) ;
  assign w1924 = ~w1911 & w1923 ;
  assign w1925 = w1922 | w1924 ;
  assign w1926 = ( w541 & w1919 ) | ( w541 & ~w1925 ) | ( w1919 & ~w1925 ) ;
  assign w1927 = w541 & w1926 ;
  assign w1928 = w1745 | w1750 ;
  assign w1929 = w1841 & ~w1928 ;
  assign w1930 = w1748 ^ w1929 ;
  assign w1931 = ( ~w541 & w1919 ) | ( ~w541 & w1925 ) | ( w1919 & w1925 ) ;
  assign w1932 = ~w1919 & w1931 ;
  assign w1933 = w1930 | w1932 ;
  assign w1934 = ( w455 & w1927 ) | ( w455 & ~w1933 ) | ( w1927 & ~w1933 ) ;
  assign w1935 = w455 & w1934 ;
  assign w1936 = w1753 | w1758 ;
  assign w1937 = w1841 & ~w1936 ;
  assign w1938 = w1756 ^ w1937 ;
  assign w1939 = ( ~w455 & w1927 ) | ( ~w455 & w1933 ) | ( w1927 & w1933 ) ;
  assign w1940 = ~w1927 & w1939 ;
  assign w1941 = w1938 | w1940 ;
  assign w1942 = ( w377 & w1935 ) | ( w377 & ~w1941 ) | ( w1935 & ~w1941 ) ;
  assign w1943 = w377 & w1942 ;
  assign w1944 = w1761 | w1766 ;
  assign w1945 = w1841 & ~w1944 ;
  assign w1946 = w1764 ^ w1945 ;
  assign w1947 = ( ~w377 & w1935 ) | ( ~w377 & w1941 ) | ( w1935 & w1941 ) ;
  assign w1948 = ~w1935 & w1947 ;
  assign w1949 = w1946 | w1948 ;
  assign w1950 = ( w307 & w1943 ) | ( w307 & ~w1949 ) | ( w1943 & ~w1949 ) ;
  assign w1951 = w307 & w1950 ;
  assign w1952 = w1769 | w1774 ;
  assign w1953 = w1841 & ~w1952 ;
  assign w1954 = w1772 ^ w1953 ;
  assign w1955 = ( ~w307 & w1943 ) | ( ~w307 & w1949 ) | ( w1943 & w1949 ) ;
  assign w1956 = ~w1943 & w1955 ;
  assign w1957 = w1954 | w1956 ;
  assign w1958 = ( w246 & w1951 ) | ( w246 & ~w1957 ) | ( w1951 & ~w1957 ) ;
  assign w1959 = w246 & w1958 ;
  assign w1960 = w1777 | w1782 ;
  assign w1961 = w1841 & ~w1960 ;
  assign w1962 = w1780 ^ w1961 ;
  assign w1963 = ( ~w246 & w1951 ) | ( ~w246 & w1957 ) | ( w1951 & w1957 ) ;
  assign w1964 = ~w1951 & w1963 ;
  assign w1965 = w1962 | w1964 ;
  assign w1966 = ( w185 & w1959 ) | ( w185 & ~w1965 ) | ( w1959 & ~w1965 ) ;
  assign w1967 = w185 & w1966 ;
  assign w1968 = w1785 | w1790 ;
  assign w1969 = w1841 & ~w1968 ;
  assign w1970 = w1788 ^ w1969 ;
  assign w1971 = ( ~w185 & w1959 ) | ( ~w185 & w1965 ) | ( w1959 & w1965 ) ;
  assign w1972 = ~w1959 & w1971 ;
  assign w1973 = w1970 | w1972 ;
  assign w1974 = ( w145 & w1967 ) | ( w145 & ~w1973 ) | ( w1967 & ~w1973 ) ;
  assign w1975 = w145 & w1974 ;
  assign w1976 = w1793 | w1798 ;
  assign w1977 = w1841 & ~w1976 ;
  assign w1978 = w1796 ^ w1977 ;
  assign w1979 = ( ~w145 & w1967 ) | ( ~w145 & w1973 ) | ( w1967 & w1973 ) ;
  assign w1980 = ~w1967 & w1979 ;
  assign w1981 = w1978 | w1980 ;
  assign w1982 = ( w132 & w1975 ) | ( w132 & ~w1981 ) | ( w1975 & ~w1981 ) ;
  assign w1983 = w132 & w1982 ;
  assign w1984 = w1801 | w1806 ;
  assign w1985 = w1841 & ~w1984 ;
  assign w1986 = w1804 ^ w1985 ;
  assign w1987 = ( ~w132 & w1975 ) | ( ~w132 & w1981 ) | ( w1975 & w1981 ) ;
  assign w1988 = ~w1975 & w1987 ;
  assign w1989 = w1986 | w1988 ;
  assign w1990 = ~w1983 & w1989 ;
  assign w1991 = w1809 | w1814 ;
  assign w1992 = w1841 & ~w1991 ;
  assign w1993 = w1812 ^ w1992 ;
  assign w1994 = ( ~w1827 & w1990 ) | ( ~w1827 & w1993 ) | ( w1990 & w1993 ) ;
  assign w1995 = w1816 & ~w1994 ;
  assign w1996 = ~w1819 & w1841 ;
  assign w1997 = ( w1994 & ~w1995 ) | ( w1994 & w1996 ) | ( ~w1995 & w1996 ) ;
  assign w1998 = w1827 | w1997 ;
  assign w1999 = ~w129 & w1998 ;
  assign w2000 = ( w1983 & w1989 ) | ( w1983 & w1993 ) | ( w1989 & w1993 ) ;
  assign w2001 = ~w1983 & w2000 ;
  assign w2002 = ( w129 & w1816 ) | ( w129 & w1819 ) | ( w1816 & w1819 ) ;
  assign w2003 = ( w1819 & ~w1841 ) | ( w1819 & w2002 ) | ( ~w1841 & w2002 ) ;
  assign w2004 = w1816 & w2003 ;
  assign w2005 = w2002 ^ w2004 ;
  assign w2006 = ( w1643 & w1648 ) | ( w1643 & w1675 ) | ( w1648 & w1675 ) ;
  assign w2007 = w1675 & ~w2006 ;
  assign w2008 = w1646 ^ w2007 ;
  assign w2009 = ( ~w1831 & w1838 ) | ( ~w1831 & w2008 ) | ( w1838 & w2008 ) ;
  assign w2010 = ~w1838 & w2009 ;
  assign w2011 = ( ~w1825 & w1827 ) | ( ~w1825 & w2010 ) | ( w1827 & w2010 ) ;
  assign w2012 = ~w1827 & w2011 ;
  assign w2013 = w2001 | w2012 ;
  assign w2014 = ( w1999 & ~w2001 ) | ( w1999 & w2005 ) | ( ~w2001 & w2005 ) ;
  assign w2015 = w2013 | w2014 ;
  assign w2016 = ( ~\pi087 & \pi088 ) | ( ~\pi087 & w1841 ) | ( \pi088 & w1841 ) ;
  assign w2017 = ( ~\pi086 & \pi088 ) | ( ~\pi086 & w2016 ) | ( \pi088 & w2016 ) ;
  assign w2018 = ( ~\pi088 & w1841 ) | ( ~\pi088 & w2015 ) | ( w1841 & w2015 ) ;
  assign w2019 = w2017 & w2018 ;
  assign w2020 = ( w1827 & w1831 ) | ( w1827 & ~w1838 ) | ( w1831 & ~w1838 ) ;
  assign w2021 = \pi087 & ~w2020 ;
  assign w2022 = \pi086 | \pi088 ;
  assign w2023 = ( ~w2020 & w2021 ) | ( ~w2020 & w2022 ) | ( w2021 & w2022 ) ;
  assign w2024 = ~w1838 & w2023 ;
  assign w2025 = ~w1825 & w2024 ;
  assign w2026 = ( \pi088 & w2015 ) | ( \pi088 & ~w2024 ) | ( w2015 & ~w2024 ) ;
  assign w2027 = w2025 & ~w2026 ;
  assign w2028 = ~\pi088 & w2015 ;
  assign w2029 = \pi089 ^ w2028 ;
  assign w2030 = w2027 | w2029 ;
  assign w2031 = ( w1675 & w2019 ) | ( w1675 & ~w2030 ) | ( w2019 & ~w2030 ) ;
  assign w2032 = w1675 & w2031 ;
  assign w2033 = ( ~w1675 & w2019 ) | ( ~w1675 & w2030 ) | ( w2019 & w2030 ) ;
  assign w2034 = ~w2019 & w2033 ;
  assign w2035 = w1841 & ~w2012 ;
  assign w2036 = ~w2001 & w2035 ;
  assign w2037 = ~w2014 & w2036 ;
  assign w2038 = \pi089 & w2015 ;
  assign w2039 = ( \pi088 & w2015 ) | ( \pi088 & ~w2038 ) | ( w2015 & ~w2038 ) ;
  assign w2040 = ( ~\pi088 & w2037 ) | ( ~\pi088 & w2039 ) | ( w2037 & w2039 ) ;
  assign w2041 = \pi090 ^ w2040 ;
  assign w2042 = w2034 | w2041 ;
  assign w2043 = ( w1517 & w2032 ) | ( w1517 & ~w2042 ) | ( w2032 & ~w2042 ) ;
  assign w2044 = w1517 & w2043 ;
  assign w2045 = ( w1845 & ~w1853 ) | ( w1845 & w2015 ) | ( ~w1853 & w2015 ) ;
  assign w2046 = ~w1845 & w2045 ;
  assign w2047 = \pi091 ^ w2046 ;
  assign w2048 = w1854 ^ w2047 ;
  assign w2049 = ( ~w1517 & w2032 ) | ( ~w1517 & w2042 ) | ( w2032 & w2042 ) ;
  assign w2050 = ~w2032 & w2049 ;
  assign w2051 = w2048 | w2050 ;
  assign w2052 = ( w1367 & w2044 ) | ( w1367 & ~w2051 ) | ( w2044 & ~w2051 ) ;
  assign w2053 = w1367 & w2052 ;
  assign w2054 = w1858 | w1860 ;
  assign w2055 = w2015 & ~w2054 ;
  assign w2056 = w1867 ^ w2055 ;
  assign w2057 = ( ~w1367 & w2044 ) | ( ~w1367 & w2051 ) | ( w2044 & w2051 ) ;
  assign w2058 = ~w2044 & w2057 ;
  assign w2059 = w2056 | w2058 ;
  assign w2060 = ( w1225 & w2053 ) | ( w1225 & ~w2059 ) | ( w2053 & ~w2059 ) ;
  assign w2061 = w1225 & w2060 ;
  assign w2062 = w1870 | w1876 ;
  assign w2063 = w2015 & ~w2062 ;
  assign w2064 = w1874 ^ w2063 ;
  assign w2065 = ( ~w1225 & w2053 ) | ( ~w1225 & w2059 ) | ( w2053 & w2059 ) ;
  assign w2066 = ~w2053 & w2065 ;
  assign w2067 = w2064 | w2066 ;
  assign w2068 = ( w1091 & w2061 ) | ( w1091 & ~w2067 ) | ( w2061 & ~w2067 ) ;
  assign w2069 = w1091 & w2068 ;
  assign w2070 = w1879 | w1884 ;
  assign w2071 = w2015 & ~w2070 ;
  assign w2072 = w1882 ^ w2071 ;
  assign w2073 = ( ~w1091 & w2061 ) | ( ~w1091 & w2067 ) | ( w2061 & w2067 ) ;
  assign w2074 = ~w2061 & w2073 ;
  assign w2075 = w2072 | w2074 ;
  assign w2076 = ( w965 & w2069 ) | ( w965 & ~w2075 ) | ( w2069 & ~w2075 ) ;
  assign w2077 = w965 & w2076 ;
  assign w2078 = w1887 | w1892 ;
  assign w2079 = w2015 & ~w2078 ;
  assign w2080 = w1890 ^ w2079 ;
  assign w2081 = ( ~w965 & w2069 ) | ( ~w965 & w2075 ) | ( w2069 & w2075 ) ;
  assign w2082 = ~w2069 & w2081 ;
  assign w2083 = w2080 | w2082 ;
  assign w2084 = ( w847 & w2077 ) | ( w847 & ~w2083 ) | ( w2077 & ~w2083 ) ;
  assign w2085 = w847 & w2084 ;
  assign w2086 = w1895 | w1900 ;
  assign w2087 = w2015 & ~w2086 ;
  assign w2088 = w1898 ^ w2087 ;
  assign w2089 = ( ~w847 & w2077 ) | ( ~w847 & w2083 ) | ( w2077 & w2083 ) ;
  assign w2090 = ~w2077 & w2089 ;
  assign w2091 = w2088 | w2090 ;
  assign w2092 = ( w737 & w2085 ) | ( w737 & ~w2091 ) | ( w2085 & ~w2091 ) ;
  assign w2093 = w737 & w2092 ;
  assign w2094 = ( ~w737 & w2085 ) | ( ~w737 & w2091 ) | ( w2085 & w2091 ) ;
  assign w2095 = ~w2085 & w2094 ;
  assign w2096 = w1903 | w1905 ;
  assign w2097 = w2015 & ~w2096 ;
  assign w2098 = w1908 ^ w2097 ;
  assign w2099 = w2095 | w2098 ;
  assign w2100 = ( w635 & w2093 ) | ( w635 & ~w2099 ) | ( w2093 & ~w2099 ) ;
  assign w2101 = w635 & w2100 ;
  assign w2102 = w1911 | w1916 ;
  assign w2103 = w2015 & ~w2102 ;
  assign w2104 = w1914 ^ w2103 ;
  assign w2105 = ( ~w635 & w2093 ) | ( ~w635 & w2099 ) | ( w2093 & w2099 ) ;
  assign w2106 = ~w2093 & w2105 ;
  assign w2107 = w2104 | w2106 ;
  assign w2108 = ( w541 & w2101 ) | ( w541 & ~w2107 ) | ( w2101 & ~w2107 ) ;
  assign w2109 = w541 & w2108 ;
  assign w2110 = w1919 | w1924 ;
  assign w2111 = w2015 & ~w2110 ;
  assign w2112 = w1922 ^ w2111 ;
  assign w2113 = ( ~w541 & w2101 ) | ( ~w541 & w2107 ) | ( w2101 & w2107 ) ;
  assign w2114 = ~w2101 & w2113 ;
  assign w2115 = w2112 | w2114 ;
  assign w2116 = ( w455 & w2109 ) | ( w455 & ~w2115 ) | ( w2109 & ~w2115 ) ;
  assign w2117 = w455 & w2116 ;
  assign w2118 = w1927 | w1932 ;
  assign w2119 = w2015 & ~w2118 ;
  assign w2120 = w1930 ^ w2119 ;
  assign w2121 = ( ~w455 & w2109 ) | ( ~w455 & w2115 ) | ( w2109 & w2115 ) ;
  assign w2122 = ~w2109 & w2121 ;
  assign w2123 = w2120 | w2122 ;
  assign w2124 = ( w377 & w2117 ) | ( w377 & ~w2123 ) | ( w2117 & ~w2123 ) ;
  assign w2125 = w377 & w2124 ;
  assign w2126 = w1935 | w1940 ;
  assign w2127 = w2015 & ~w2126 ;
  assign w2128 = w1938 ^ w2127 ;
  assign w2129 = ( ~w377 & w2117 ) | ( ~w377 & w2123 ) | ( w2117 & w2123 ) ;
  assign w2130 = ~w2117 & w2129 ;
  assign w2131 = w2128 | w2130 ;
  assign w2132 = ( w307 & w2125 ) | ( w307 & ~w2131 ) | ( w2125 & ~w2131 ) ;
  assign w2133 = w307 & w2132 ;
  assign w2134 = w1943 | w1948 ;
  assign w2135 = w2015 & ~w2134 ;
  assign w2136 = w1946 ^ w2135 ;
  assign w2137 = ( ~w307 & w2125 ) | ( ~w307 & w2131 ) | ( w2125 & w2131 ) ;
  assign w2138 = ~w2125 & w2137 ;
  assign w2139 = w2136 | w2138 ;
  assign w2140 = ( w246 & w2133 ) | ( w246 & ~w2139 ) | ( w2133 & ~w2139 ) ;
  assign w2141 = w246 & w2140 ;
  assign w2142 = w1951 | w1956 ;
  assign w2143 = w2015 & ~w2142 ;
  assign w2144 = w1954 ^ w2143 ;
  assign w2145 = ( ~w246 & w2133 ) | ( ~w246 & w2139 ) | ( w2133 & w2139 ) ;
  assign w2146 = ~w2133 & w2145 ;
  assign w2147 = w2144 | w2146 ;
  assign w2148 = ( w185 & w2141 ) | ( w185 & ~w2147 ) | ( w2141 & ~w2147 ) ;
  assign w2149 = w185 & w2148 ;
  assign w2150 = w1959 | w1964 ;
  assign w2151 = w2015 & ~w2150 ;
  assign w2152 = w1962 ^ w2151 ;
  assign w2153 = ( ~w185 & w2141 ) | ( ~w185 & w2147 ) | ( w2141 & w2147 ) ;
  assign w2154 = ~w2141 & w2153 ;
  assign w2155 = w2152 | w2154 ;
  assign w2156 = ( w145 & w2149 ) | ( w145 & ~w2155 ) | ( w2149 & ~w2155 ) ;
  assign w2157 = w145 & w2156 ;
  assign w2158 = w1967 | w1972 ;
  assign w2159 = w2015 & ~w2158 ;
  assign w2160 = w1970 ^ w2159 ;
  assign w2161 = ( ~w145 & w2149 ) | ( ~w145 & w2155 ) | ( w2149 & w2155 ) ;
  assign w2162 = ~w2149 & w2161 ;
  assign w2163 = w2160 | w2162 ;
  assign w2164 = ( w132 & w2157 ) | ( w132 & ~w2163 ) | ( w2157 & ~w2163 ) ;
  assign w2165 = w132 & w2164 ;
  assign w2166 = w1975 | w1980 ;
  assign w2167 = w2015 & ~w2166 ;
  assign w2168 = w1978 ^ w2167 ;
  assign w2169 = ( ~w132 & w2157 ) | ( ~w132 & w2163 ) | ( w2157 & w2163 ) ;
  assign w2170 = ~w2157 & w2169 ;
  assign w2171 = w2168 | w2170 ;
  assign w2172 = ~w2165 & w2171 ;
  assign w2173 = w1983 | w1988 ;
  assign w2174 = w2015 & ~w2173 ;
  assign w2175 = w1986 ^ w2174 ;
  assign w2176 = ( ~w2001 & w2172 ) | ( ~w2001 & w2175 ) | ( w2172 & w2175 ) ;
  assign w2177 = w1990 & ~w2176 ;
  assign w2178 = ~w1993 & w2015 ;
  assign w2179 = ( w2176 & ~w2177 ) | ( w2176 & w2178 ) | ( ~w2177 & w2178 ) ;
  assign w2180 = w2001 | w2179 ;
  assign w2181 = ~w129 & w2180 ;
  assign w2182 = ( w2165 & w2171 ) | ( w2165 & w2175 ) | ( w2171 & w2175 ) ;
  assign w2183 = ~w2165 & w2182 ;
  assign w2184 = ( w129 & w1990 ) | ( w129 & w1993 ) | ( w1990 & w1993 ) ;
  assign w2185 = ( w1993 & ~w2015 ) | ( w1993 & w2184 ) | ( ~w2015 & w2184 ) ;
  assign w2186 = w1990 & w2185 ;
  assign w2187 = w2184 ^ w2186 ;
  assign w2188 = ( w1809 & w1814 ) | ( w1809 & w1841 ) | ( w1814 & w1841 ) ;
  assign w2189 = w1841 & ~w2188 ;
  assign w2190 = w1812 ^ w2189 ;
  assign w2191 = ( ~w2005 & w2012 ) | ( ~w2005 & w2190 ) | ( w2012 & w2190 ) ;
  assign w2192 = ~w2012 & w2191 ;
  assign w2193 = ( ~w1999 & w2001 ) | ( ~w1999 & w2192 ) | ( w2001 & w2192 ) ;
  assign w2194 = ~w2001 & w2193 ;
  assign w2195 = w2183 | w2194 ;
  assign w2196 = ( w2181 & ~w2183 ) | ( w2181 & w2187 ) | ( ~w2183 & w2187 ) ;
  assign w2197 = w2195 | w2196 ;
  assign w2198 = ( ~\pi085 & \pi086 ) | ( ~\pi085 & w2015 ) | ( \pi086 & w2015 ) ;
  assign w2199 = ( ~\pi084 & \pi086 ) | ( ~\pi084 & w2198 ) | ( \pi086 & w2198 ) ;
  assign w2200 = ( ~\pi086 & w2015 ) | ( ~\pi086 & w2197 ) | ( w2015 & w2197 ) ;
  assign w2201 = w2199 & w2200 ;
  assign w2202 = ( w2001 & w2005 ) | ( w2001 & ~w2012 ) | ( w2005 & ~w2012 ) ;
  assign w2203 = \pi085 & ~w2202 ;
  assign w2204 = \pi084 | \pi086 ;
  assign w2205 = ( ~w2202 & w2203 ) | ( ~w2202 & w2204 ) | ( w2203 & w2204 ) ;
  assign w2206 = ~w2012 & w2205 ;
  assign w2207 = ~w1999 & w2206 ;
  assign w2208 = ( \pi086 & w2197 ) | ( \pi086 & ~w2206 ) | ( w2197 & ~w2206 ) ;
  assign w2209 = w2207 & ~w2208 ;
  assign w2210 = ~\pi086 & w2197 ;
  assign w2211 = \pi087 ^ w2210 ;
  assign w2212 = w2209 | w2211 ;
  assign w2213 = ( w1841 & w2201 ) | ( w1841 & ~w2212 ) | ( w2201 & ~w2212 ) ;
  assign w2214 = w1841 & w2213 ;
  assign w2215 = ( ~w1841 & w2201 ) | ( ~w1841 & w2212 ) | ( w2201 & w2212 ) ;
  assign w2216 = ~w2201 & w2215 ;
  assign w2217 = w2015 & ~w2194 ;
  assign w2218 = ~w2183 & w2217 ;
  assign w2219 = ~w2196 & w2218 ;
  assign w2220 = \pi087 & w2197 ;
  assign w2221 = ( \pi086 & w2197 ) | ( \pi086 & ~w2220 ) | ( w2197 & ~w2220 ) ;
  assign w2222 = ( ~\pi086 & w2219 ) | ( ~\pi086 & w2221 ) | ( w2219 & w2221 ) ;
  assign w2223 = \pi088 ^ w2222 ;
  assign w2224 = w2216 | w2223 ;
  assign w2225 = ( w1675 & w2214 ) | ( w1675 & ~w2224 ) | ( w2214 & ~w2224 ) ;
  assign w2226 = w1675 & w2225 ;
  assign w2227 = ( w2019 & ~w2027 ) | ( w2019 & w2197 ) | ( ~w2027 & w2197 ) ;
  assign w2228 = ~w2019 & w2227 ;
  assign w2229 = \pi089 ^ w2228 ;
  assign w2230 = w2028 ^ w2229 ;
  assign w2231 = ( ~w1675 & w2214 ) | ( ~w1675 & w2224 ) | ( w2214 & w2224 ) ;
  assign w2232 = ~w2214 & w2231 ;
  assign w2233 = w2230 | w2232 ;
  assign w2234 = ( w1517 & w2226 ) | ( w1517 & ~w2233 ) | ( w2226 & ~w2233 ) ;
  assign w2235 = w1517 & w2234 ;
  assign w2236 = w2032 | w2034 ;
  assign w2237 = w2197 & ~w2236 ;
  assign w2238 = w2041 ^ w2237 ;
  assign w2239 = ( ~w1517 & w2226 ) | ( ~w1517 & w2233 ) | ( w2226 & w2233 ) ;
  assign w2240 = ~w2226 & w2239 ;
  assign w2241 = w2238 | w2240 ;
  assign w2242 = ( w1367 & w2235 ) | ( w1367 & ~w2241 ) | ( w2235 & ~w2241 ) ;
  assign w2243 = w1367 & w2242 ;
  assign w2244 = w2044 | w2050 ;
  assign w2245 = w2197 & ~w2244 ;
  assign w2246 = w2048 ^ w2245 ;
  assign w2247 = ( ~w1367 & w2235 ) | ( ~w1367 & w2241 ) | ( w2235 & w2241 ) ;
  assign w2248 = ~w2235 & w2247 ;
  assign w2249 = w2246 | w2248 ;
  assign w2250 = ( w1225 & w2243 ) | ( w1225 & ~w2249 ) | ( w2243 & ~w2249 ) ;
  assign w2251 = w1225 & w2250 ;
  assign w2252 = w2053 | w2058 ;
  assign w2253 = w2197 & ~w2252 ;
  assign w2254 = w2056 ^ w2253 ;
  assign w2255 = ( ~w1225 & w2243 ) | ( ~w1225 & w2249 ) | ( w2243 & w2249 ) ;
  assign w2256 = ~w2243 & w2255 ;
  assign w2257 = w2254 | w2256 ;
  assign w2258 = ( w1091 & w2251 ) | ( w1091 & ~w2257 ) | ( w2251 & ~w2257 ) ;
  assign w2259 = w1091 & w2258 ;
  assign w2260 = w2061 | w2066 ;
  assign w2261 = w2197 & ~w2260 ;
  assign w2262 = w2064 ^ w2261 ;
  assign w2263 = ( ~w1091 & w2251 ) | ( ~w1091 & w2257 ) | ( w2251 & w2257 ) ;
  assign w2264 = ~w2251 & w2263 ;
  assign w2265 = w2262 | w2264 ;
  assign w2266 = ( w965 & w2259 ) | ( w965 & ~w2265 ) | ( w2259 & ~w2265 ) ;
  assign w2267 = w965 & w2266 ;
  assign w2268 = w2069 | w2074 ;
  assign w2269 = w2197 & ~w2268 ;
  assign w2270 = w2072 ^ w2269 ;
  assign w2271 = ( ~w965 & w2259 ) | ( ~w965 & w2265 ) | ( w2259 & w2265 ) ;
  assign w2272 = ~w2259 & w2271 ;
  assign w2273 = w2270 | w2272 ;
  assign w2274 = ( w847 & w2267 ) | ( w847 & ~w2273 ) | ( w2267 & ~w2273 ) ;
  assign w2275 = w847 & w2274 ;
  assign w2276 = w2077 | w2082 ;
  assign w2277 = w2197 & ~w2276 ;
  assign w2278 = w2080 ^ w2277 ;
  assign w2279 = ( ~w847 & w2267 ) | ( ~w847 & w2273 ) | ( w2267 & w2273 ) ;
  assign w2280 = ~w2267 & w2279 ;
  assign w2281 = w2278 | w2280 ;
  assign w2282 = ( w737 & w2275 ) | ( w737 & ~w2281 ) | ( w2275 & ~w2281 ) ;
  assign w2283 = w737 & w2282 ;
  assign w2284 = w2085 | w2090 ;
  assign w2285 = w2197 & ~w2284 ;
  assign w2286 = w2088 ^ w2285 ;
  assign w2287 = ( ~w737 & w2275 ) | ( ~w737 & w2281 ) | ( w2275 & w2281 ) ;
  assign w2288 = ~w2275 & w2287 ;
  assign w2289 = w2286 | w2288 ;
  assign w2290 = ( w635 & w2283 ) | ( w635 & ~w2289 ) | ( w2283 & ~w2289 ) ;
  assign w2291 = w635 & w2290 ;
  assign w2292 = ( ~w635 & w2283 ) | ( ~w635 & w2289 ) | ( w2283 & w2289 ) ;
  assign w2293 = ~w2283 & w2292 ;
  assign w2294 = w2093 | w2095 ;
  assign w2295 = w2197 & ~w2294 ;
  assign w2296 = w2098 ^ w2295 ;
  assign w2297 = w2293 | w2296 ;
  assign w2298 = ( w541 & w2291 ) | ( w541 & ~w2297 ) | ( w2291 & ~w2297 ) ;
  assign w2299 = w541 & w2298 ;
  assign w2300 = w2101 | w2106 ;
  assign w2301 = w2197 & ~w2300 ;
  assign w2302 = w2104 ^ w2301 ;
  assign w2303 = ( ~w541 & w2291 ) | ( ~w541 & w2297 ) | ( w2291 & w2297 ) ;
  assign w2304 = ~w2291 & w2303 ;
  assign w2305 = w2302 | w2304 ;
  assign w2306 = ( w455 & w2299 ) | ( w455 & ~w2305 ) | ( w2299 & ~w2305 ) ;
  assign w2307 = w455 & w2306 ;
  assign w2308 = w2109 | w2114 ;
  assign w2309 = w2197 & ~w2308 ;
  assign w2310 = w2112 ^ w2309 ;
  assign w2311 = ( ~w455 & w2299 ) | ( ~w455 & w2305 ) | ( w2299 & w2305 ) ;
  assign w2312 = ~w2299 & w2311 ;
  assign w2313 = w2310 | w2312 ;
  assign w2314 = ( w377 & w2307 ) | ( w377 & ~w2313 ) | ( w2307 & ~w2313 ) ;
  assign w2315 = w377 & w2314 ;
  assign w2316 = w2117 | w2122 ;
  assign w2317 = w2197 & ~w2316 ;
  assign w2318 = w2120 ^ w2317 ;
  assign w2319 = ( ~w377 & w2307 ) | ( ~w377 & w2313 ) | ( w2307 & w2313 ) ;
  assign w2320 = ~w2307 & w2319 ;
  assign w2321 = w2318 | w2320 ;
  assign w2322 = ( w307 & w2315 ) | ( w307 & ~w2321 ) | ( w2315 & ~w2321 ) ;
  assign w2323 = w307 & w2322 ;
  assign w2324 = w2125 | w2130 ;
  assign w2325 = w2197 & ~w2324 ;
  assign w2326 = w2128 ^ w2325 ;
  assign w2327 = ( ~w307 & w2315 ) | ( ~w307 & w2321 ) | ( w2315 & w2321 ) ;
  assign w2328 = ~w2315 & w2327 ;
  assign w2329 = w2326 | w2328 ;
  assign w2330 = ( w246 & w2323 ) | ( w246 & ~w2329 ) | ( w2323 & ~w2329 ) ;
  assign w2331 = w246 & w2330 ;
  assign w2332 = w2133 | w2138 ;
  assign w2333 = w2197 & ~w2332 ;
  assign w2334 = w2136 ^ w2333 ;
  assign w2335 = ( ~w246 & w2323 ) | ( ~w246 & w2329 ) | ( w2323 & w2329 ) ;
  assign w2336 = ~w2323 & w2335 ;
  assign w2337 = w2334 | w2336 ;
  assign w2338 = ( w185 & w2331 ) | ( w185 & ~w2337 ) | ( w2331 & ~w2337 ) ;
  assign w2339 = w185 & w2338 ;
  assign w2340 = w2141 | w2146 ;
  assign w2341 = w2197 & ~w2340 ;
  assign w2342 = w2144 ^ w2341 ;
  assign w2343 = ( ~w185 & w2331 ) | ( ~w185 & w2337 ) | ( w2331 & w2337 ) ;
  assign w2344 = ~w2331 & w2343 ;
  assign w2345 = w2342 | w2344 ;
  assign w2346 = ( w145 & w2339 ) | ( w145 & ~w2345 ) | ( w2339 & ~w2345 ) ;
  assign w2347 = w145 & w2346 ;
  assign w2348 = w2149 | w2154 ;
  assign w2349 = w2197 & ~w2348 ;
  assign w2350 = w2152 ^ w2349 ;
  assign w2351 = ( ~w145 & w2339 ) | ( ~w145 & w2345 ) | ( w2339 & w2345 ) ;
  assign w2352 = ~w2339 & w2351 ;
  assign w2353 = w2350 | w2352 ;
  assign w2354 = ( w132 & w2347 ) | ( w132 & ~w2353 ) | ( w2347 & ~w2353 ) ;
  assign w2355 = w132 & w2354 ;
  assign w2356 = w2157 | w2162 ;
  assign w2357 = w2197 & ~w2356 ;
  assign w2358 = w2160 ^ w2357 ;
  assign w2359 = ( ~w132 & w2347 ) | ( ~w132 & w2353 ) | ( w2347 & w2353 ) ;
  assign w2360 = ~w2347 & w2359 ;
  assign w2361 = w2358 | w2360 ;
  assign w2362 = ~w2355 & w2361 ;
  assign w2363 = w2165 | w2170 ;
  assign w2364 = w2197 & ~w2363 ;
  assign w2365 = w2168 ^ w2364 ;
  assign w2366 = ( ~w2183 & w2362 ) | ( ~w2183 & w2365 ) | ( w2362 & w2365 ) ;
  assign w2367 = w2172 & ~w2366 ;
  assign w2368 = ~w2175 & w2197 ;
  assign w2369 = ( w2366 & ~w2367 ) | ( w2366 & w2368 ) | ( ~w2367 & w2368 ) ;
  assign w2370 = w2183 | w2369 ;
  assign w2371 = ~w129 & w2370 ;
  assign w2372 = ( w2355 & w2361 ) | ( w2355 & w2365 ) | ( w2361 & w2365 ) ;
  assign w2373 = ~w2355 & w2372 ;
  assign w2374 = ( w129 & w2172 ) | ( w129 & w2175 ) | ( w2172 & w2175 ) ;
  assign w2375 = ( w2175 & ~w2197 ) | ( w2175 & w2374 ) | ( ~w2197 & w2374 ) ;
  assign w2376 = w2172 & w2375 ;
  assign w2377 = w2374 ^ w2376 ;
  assign w2378 = ( w1983 & w1988 ) | ( w1983 & w2015 ) | ( w1988 & w2015 ) ;
  assign w2379 = w2015 & ~w2378 ;
  assign w2380 = w1986 ^ w2379 ;
  assign w2381 = ( ~w2187 & w2194 ) | ( ~w2187 & w2380 ) | ( w2194 & w2380 ) ;
  assign w2382 = ~w2194 & w2381 ;
  assign w2383 = ( ~w2181 & w2183 ) | ( ~w2181 & w2382 ) | ( w2183 & w2382 ) ;
  assign w2384 = ~w2183 & w2383 ;
  assign w2385 = w2373 | w2384 ;
  assign w2386 = ( w2371 & ~w2373 ) | ( w2371 & w2377 ) | ( ~w2373 & w2377 ) ;
  assign w2387 = w2385 | w2386 ;
  assign w2388 = ( ~\pi083 & \pi084 ) | ( ~\pi083 & w2197 ) | ( \pi084 & w2197 ) ;
  assign w2389 = ( ~\pi082 & \pi084 ) | ( ~\pi082 & w2388 ) | ( \pi084 & w2388 ) ;
  assign w2390 = ( ~\pi084 & w2197 ) | ( ~\pi084 & w2387 ) | ( w2197 & w2387 ) ;
  assign w2391 = w2389 & w2390 ;
  assign w2392 = ( w2183 & w2187 ) | ( w2183 & ~w2194 ) | ( w2187 & ~w2194 ) ;
  assign w2393 = \pi083 & ~w2392 ;
  assign w2394 = \pi082 | \pi084 ;
  assign w2395 = ( ~w2392 & w2393 ) | ( ~w2392 & w2394 ) | ( w2393 & w2394 ) ;
  assign w2396 = ~w2194 & w2395 ;
  assign w2397 = ~w2181 & w2396 ;
  assign w2398 = ( \pi084 & w2387 ) | ( \pi084 & ~w2396 ) | ( w2387 & ~w2396 ) ;
  assign w2399 = w2397 & ~w2398 ;
  assign w2400 = ~\pi084 & w2387 ;
  assign w2401 = \pi085 ^ w2400 ;
  assign w2402 = w2399 | w2401 ;
  assign w2403 = ( w2015 & w2391 ) | ( w2015 & ~w2402 ) | ( w2391 & ~w2402 ) ;
  assign w2404 = w2015 & w2403 ;
  assign w2405 = ( ~w2015 & w2391 ) | ( ~w2015 & w2402 ) | ( w2391 & w2402 ) ;
  assign w2406 = ~w2391 & w2405 ;
  assign w2407 = w2197 & ~w2384 ;
  assign w2408 = ~w2373 & w2407 ;
  assign w2409 = ~w2386 & w2408 ;
  assign w2410 = \pi085 & w2387 ;
  assign w2411 = ( \pi084 & w2387 ) | ( \pi084 & ~w2410 ) | ( w2387 & ~w2410 ) ;
  assign w2412 = ( ~\pi084 & w2409 ) | ( ~\pi084 & w2411 ) | ( w2409 & w2411 ) ;
  assign w2413 = \pi086 ^ w2412 ;
  assign w2414 = w2406 | w2413 ;
  assign w2415 = ( w1841 & w2404 ) | ( w1841 & ~w2414 ) | ( w2404 & ~w2414 ) ;
  assign w2416 = w1841 & w2415 ;
  assign w2417 = ( w2201 & ~w2209 ) | ( w2201 & w2387 ) | ( ~w2209 & w2387 ) ;
  assign w2418 = ~w2201 & w2417 ;
  assign w2419 = \pi087 ^ w2418 ;
  assign w2420 = w2210 ^ w2419 ;
  assign w2421 = ( ~w1841 & w2404 ) | ( ~w1841 & w2414 ) | ( w2404 & w2414 ) ;
  assign w2422 = ~w2404 & w2421 ;
  assign w2423 = w2420 | w2422 ;
  assign w2424 = ( w1675 & w2416 ) | ( w1675 & ~w2423 ) | ( w2416 & ~w2423 ) ;
  assign w2425 = w1675 & w2424 ;
  assign w2426 = w2214 | w2216 ;
  assign w2427 = w2387 & ~w2426 ;
  assign w2428 = w2223 ^ w2427 ;
  assign w2429 = ( ~w1675 & w2416 ) | ( ~w1675 & w2423 ) | ( w2416 & w2423 ) ;
  assign w2430 = ~w2416 & w2429 ;
  assign w2431 = w2428 | w2430 ;
  assign w2432 = ( w1517 & w2425 ) | ( w1517 & ~w2431 ) | ( w2425 & ~w2431 ) ;
  assign w2433 = w1517 & w2432 ;
  assign w2434 = w2226 | w2232 ;
  assign w2435 = w2387 & ~w2434 ;
  assign w2436 = w2230 ^ w2435 ;
  assign w2437 = ( ~w1517 & w2425 ) | ( ~w1517 & w2431 ) | ( w2425 & w2431 ) ;
  assign w2438 = ~w2425 & w2437 ;
  assign w2439 = w2436 | w2438 ;
  assign w2440 = ( w1367 & w2433 ) | ( w1367 & ~w2439 ) | ( w2433 & ~w2439 ) ;
  assign w2441 = w1367 & w2440 ;
  assign w2442 = w2235 | w2240 ;
  assign w2443 = w2387 & ~w2442 ;
  assign w2444 = w2238 ^ w2443 ;
  assign w2445 = ( ~w1367 & w2433 ) | ( ~w1367 & w2439 ) | ( w2433 & w2439 ) ;
  assign w2446 = ~w2433 & w2445 ;
  assign w2447 = w2444 | w2446 ;
  assign w2448 = ( w1225 & w2441 ) | ( w1225 & ~w2447 ) | ( w2441 & ~w2447 ) ;
  assign w2449 = w1225 & w2448 ;
  assign w2450 = w2243 | w2248 ;
  assign w2451 = w2387 & ~w2450 ;
  assign w2452 = w2246 ^ w2451 ;
  assign w2453 = ( ~w1225 & w2441 ) | ( ~w1225 & w2447 ) | ( w2441 & w2447 ) ;
  assign w2454 = ~w2441 & w2453 ;
  assign w2455 = w2452 | w2454 ;
  assign w2456 = ( w1091 & w2449 ) | ( w1091 & ~w2455 ) | ( w2449 & ~w2455 ) ;
  assign w2457 = w1091 & w2456 ;
  assign w2458 = w2251 | w2256 ;
  assign w2459 = w2387 & ~w2458 ;
  assign w2460 = w2254 ^ w2459 ;
  assign w2461 = ( ~w1091 & w2449 ) | ( ~w1091 & w2455 ) | ( w2449 & w2455 ) ;
  assign w2462 = ~w2449 & w2461 ;
  assign w2463 = w2460 | w2462 ;
  assign w2464 = ( w965 & w2457 ) | ( w965 & ~w2463 ) | ( w2457 & ~w2463 ) ;
  assign w2465 = w965 & w2464 ;
  assign w2466 = w2259 | w2264 ;
  assign w2467 = w2387 & ~w2466 ;
  assign w2468 = w2262 ^ w2467 ;
  assign w2469 = ( ~w965 & w2457 ) | ( ~w965 & w2463 ) | ( w2457 & w2463 ) ;
  assign w2470 = ~w2457 & w2469 ;
  assign w2471 = w2468 | w2470 ;
  assign w2472 = ( w847 & w2465 ) | ( w847 & ~w2471 ) | ( w2465 & ~w2471 ) ;
  assign w2473 = w847 & w2472 ;
  assign w2474 = w2267 | w2272 ;
  assign w2475 = w2387 & ~w2474 ;
  assign w2476 = w2270 ^ w2475 ;
  assign w2477 = ( ~w847 & w2465 ) | ( ~w847 & w2471 ) | ( w2465 & w2471 ) ;
  assign w2478 = ~w2465 & w2477 ;
  assign w2479 = w2476 | w2478 ;
  assign w2480 = ( w737 & w2473 ) | ( w737 & ~w2479 ) | ( w2473 & ~w2479 ) ;
  assign w2481 = w737 & w2480 ;
  assign w2482 = w2275 | w2280 ;
  assign w2483 = w2387 & ~w2482 ;
  assign w2484 = w2278 ^ w2483 ;
  assign w2485 = ( ~w737 & w2473 ) | ( ~w737 & w2479 ) | ( w2473 & w2479 ) ;
  assign w2486 = ~w2473 & w2485 ;
  assign w2487 = w2484 | w2486 ;
  assign w2488 = ( w635 & w2481 ) | ( w635 & ~w2487 ) | ( w2481 & ~w2487 ) ;
  assign w2489 = w635 & w2488 ;
  assign w2490 = w2283 | w2288 ;
  assign w2491 = w2387 & ~w2490 ;
  assign w2492 = w2286 ^ w2491 ;
  assign w2493 = ( ~w635 & w2481 ) | ( ~w635 & w2487 ) | ( w2481 & w2487 ) ;
  assign w2494 = ~w2481 & w2493 ;
  assign w2495 = w2492 | w2494 ;
  assign w2496 = ( w541 & w2489 ) | ( w541 & ~w2495 ) | ( w2489 & ~w2495 ) ;
  assign w2497 = w541 & w2496 ;
  assign w2498 = ( ~w541 & w2489 ) | ( ~w541 & w2495 ) | ( w2489 & w2495 ) ;
  assign w2499 = ~w2489 & w2498 ;
  assign w2500 = w2291 | w2293 ;
  assign w2501 = w2387 & ~w2500 ;
  assign w2502 = w2296 ^ w2501 ;
  assign w2503 = w2499 | w2502 ;
  assign w2504 = ( w455 & w2497 ) | ( w455 & ~w2503 ) | ( w2497 & ~w2503 ) ;
  assign w2505 = w455 & w2504 ;
  assign w2506 = w2299 | w2304 ;
  assign w2507 = w2387 & ~w2506 ;
  assign w2508 = w2302 ^ w2507 ;
  assign w2509 = ( ~w455 & w2497 ) | ( ~w455 & w2503 ) | ( w2497 & w2503 ) ;
  assign w2510 = ~w2497 & w2509 ;
  assign w2511 = w2508 | w2510 ;
  assign w2512 = ( w377 & w2505 ) | ( w377 & ~w2511 ) | ( w2505 & ~w2511 ) ;
  assign w2513 = w377 & w2512 ;
  assign w2514 = w2307 | w2312 ;
  assign w2515 = w2387 & ~w2514 ;
  assign w2516 = w2310 ^ w2515 ;
  assign w2517 = ( ~w377 & w2505 ) | ( ~w377 & w2511 ) | ( w2505 & w2511 ) ;
  assign w2518 = ~w2505 & w2517 ;
  assign w2519 = w2516 | w2518 ;
  assign w2520 = ( w307 & w2513 ) | ( w307 & ~w2519 ) | ( w2513 & ~w2519 ) ;
  assign w2521 = w307 & w2520 ;
  assign w2522 = w2315 | w2320 ;
  assign w2523 = w2387 & ~w2522 ;
  assign w2524 = w2318 ^ w2523 ;
  assign w2525 = ( ~w307 & w2513 ) | ( ~w307 & w2519 ) | ( w2513 & w2519 ) ;
  assign w2526 = ~w2513 & w2525 ;
  assign w2527 = w2524 | w2526 ;
  assign w2528 = ( w246 & w2521 ) | ( w246 & ~w2527 ) | ( w2521 & ~w2527 ) ;
  assign w2529 = w246 & w2528 ;
  assign w2530 = w2323 | w2328 ;
  assign w2531 = w2387 & ~w2530 ;
  assign w2532 = w2326 ^ w2531 ;
  assign w2533 = ( ~w246 & w2521 ) | ( ~w246 & w2527 ) | ( w2521 & w2527 ) ;
  assign w2534 = ~w2521 & w2533 ;
  assign w2535 = w2532 | w2534 ;
  assign w2536 = ( w185 & w2529 ) | ( w185 & ~w2535 ) | ( w2529 & ~w2535 ) ;
  assign w2537 = w185 & w2536 ;
  assign w2538 = w2331 | w2336 ;
  assign w2539 = w2387 & ~w2538 ;
  assign w2540 = w2334 ^ w2539 ;
  assign w2541 = ( ~w185 & w2529 ) | ( ~w185 & w2535 ) | ( w2529 & w2535 ) ;
  assign w2542 = ~w2529 & w2541 ;
  assign w2543 = w2540 | w2542 ;
  assign w2544 = ( w145 & w2537 ) | ( w145 & ~w2543 ) | ( w2537 & ~w2543 ) ;
  assign w2545 = w145 & w2544 ;
  assign w2546 = w2339 | w2344 ;
  assign w2547 = w2387 & ~w2546 ;
  assign w2548 = w2342 ^ w2547 ;
  assign w2549 = ( ~w145 & w2537 ) | ( ~w145 & w2543 ) | ( w2537 & w2543 ) ;
  assign w2550 = ~w2537 & w2549 ;
  assign w2551 = w2548 | w2550 ;
  assign w2552 = ( w132 & w2545 ) | ( w132 & ~w2551 ) | ( w2545 & ~w2551 ) ;
  assign w2553 = w132 & w2552 ;
  assign w2554 = w2347 | w2352 ;
  assign w2555 = w2387 & ~w2554 ;
  assign w2556 = w2350 ^ w2555 ;
  assign w2557 = ( ~w132 & w2545 ) | ( ~w132 & w2551 ) | ( w2545 & w2551 ) ;
  assign w2558 = ~w2545 & w2557 ;
  assign w2559 = w2556 | w2558 ;
  assign w2560 = ~w2553 & w2559 ;
  assign w2561 = w2355 | w2360 ;
  assign w2562 = w2387 & ~w2561 ;
  assign w2563 = w2358 ^ w2562 ;
  assign w2564 = ( ~w2373 & w2560 ) | ( ~w2373 & w2563 ) | ( w2560 & w2563 ) ;
  assign w2565 = w2362 & ~w2564 ;
  assign w2566 = ~w2365 & w2387 ;
  assign w2567 = ( w2564 & ~w2565 ) | ( w2564 & w2566 ) | ( ~w2565 & w2566 ) ;
  assign w2568 = w2373 | w2567 ;
  assign w2569 = ~w129 & w2568 ;
  assign w2570 = ( w2553 & w2559 ) | ( w2553 & w2563 ) | ( w2559 & w2563 ) ;
  assign w2571 = ~w2553 & w2570 ;
  assign w2572 = ( w129 & w2362 ) | ( w129 & w2365 ) | ( w2362 & w2365 ) ;
  assign w2573 = ( w2365 & ~w2387 ) | ( w2365 & w2572 ) | ( ~w2387 & w2572 ) ;
  assign w2574 = w2362 & w2573 ;
  assign w2575 = w2572 ^ w2574 ;
  assign w2576 = ( w2165 & w2170 ) | ( w2165 & w2197 ) | ( w2170 & w2197 ) ;
  assign w2577 = w2197 & ~w2576 ;
  assign w2578 = w2168 ^ w2577 ;
  assign w2579 = ( ~w2377 & w2384 ) | ( ~w2377 & w2578 ) | ( w2384 & w2578 ) ;
  assign w2580 = ~w2384 & w2579 ;
  assign w2581 = ( ~w2371 & w2373 ) | ( ~w2371 & w2580 ) | ( w2373 & w2580 ) ;
  assign w2582 = ~w2373 & w2581 ;
  assign w2583 = w2571 | w2582 ;
  assign w2584 = ( w2569 & ~w2571 ) | ( w2569 & w2575 ) | ( ~w2571 & w2575 ) ;
  assign w2585 = w2583 | w2584 ;
  assign w2586 = ( ~\pi081 & \pi082 ) | ( ~\pi081 & w2387 ) | ( \pi082 & w2387 ) ;
  assign w2587 = ( ~\pi080 & \pi082 ) | ( ~\pi080 & w2586 ) | ( \pi082 & w2586 ) ;
  assign w2588 = ( ~\pi082 & w2387 ) | ( ~\pi082 & w2585 ) | ( w2387 & w2585 ) ;
  assign w2589 = w2587 & w2588 ;
  assign w2590 = ( w2373 & w2377 ) | ( w2373 & ~w2384 ) | ( w2377 & ~w2384 ) ;
  assign w2591 = \pi081 & ~w2590 ;
  assign w2592 = \pi080 | \pi082 ;
  assign w2593 = ( ~w2590 & w2591 ) | ( ~w2590 & w2592 ) | ( w2591 & w2592 ) ;
  assign w2594 = ~w2384 & w2593 ;
  assign w2595 = ~w2371 & w2594 ;
  assign w2596 = ( \pi082 & w2585 ) | ( \pi082 & ~w2594 ) | ( w2585 & ~w2594 ) ;
  assign w2597 = w2595 & ~w2596 ;
  assign w2598 = ~\pi082 & w2585 ;
  assign w2599 = \pi083 ^ w2598 ;
  assign w2600 = w2597 | w2599 ;
  assign w2601 = ( w2197 & w2589 ) | ( w2197 & ~w2600 ) | ( w2589 & ~w2600 ) ;
  assign w2602 = w2197 & w2601 ;
  assign w2603 = ( ~w2197 & w2589 ) | ( ~w2197 & w2600 ) | ( w2589 & w2600 ) ;
  assign w2604 = ~w2589 & w2603 ;
  assign w2605 = w2387 & ~w2582 ;
  assign w2606 = ~w2571 & w2605 ;
  assign w2607 = ~w2584 & w2606 ;
  assign w2608 = \pi083 & w2585 ;
  assign w2609 = ( \pi082 & w2585 ) | ( \pi082 & ~w2608 ) | ( w2585 & ~w2608 ) ;
  assign w2610 = ( ~\pi082 & w2607 ) | ( ~\pi082 & w2609 ) | ( w2607 & w2609 ) ;
  assign w2611 = \pi084 ^ w2610 ;
  assign w2612 = w2604 | w2611 ;
  assign w2613 = ( w2015 & w2602 ) | ( w2015 & ~w2612 ) | ( w2602 & ~w2612 ) ;
  assign w2614 = w2015 & w2613 ;
  assign w2615 = ( w2391 & ~w2399 ) | ( w2391 & w2585 ) | ( ~w2399 & w2585 ) ;
  assign w2616 = ~w2391 & w2615 ;
  assign w2617 = \pi085 ^ w2616 ;
  assign w2618 = w2400 ^ w2617 ;
  assign w2619 = ( ~w2015 & w2602 ) | ( ~w2015 & w2612 ) | ( w2602 & w2612 ) ;
  assign w2620 = ~w2602 & w2619 ;
  assign w2621 = w2618 | w2620 ;
  assign w2622 = ( w1841 & w2614 ) | ( w1841 & ~w2621 ) | ( w2614 & ~w2621 ) ;
  assign w2623 = w1841 & w2622 ;
  assign w2624 = w2404 | w2406 ;
  assign w2625 = w2585 & ~w2624 ;
  assign w2626 = w2413 ^ w2625 ;
  assign w2627 = ( ~w1841 & w2614 ) | ( ~w1841 & w2621 ) | ( w2614 & w2621 ) ;
  assign w2628 = ~w2614 & w2627 ;
  assign w2629 = w2626 | w2628 ;
  assign w2630 = ( w1675 & w2623 ) | ( w1675 & ~w2629 ) | ( w2623 & ~w2629 ) ;
  assign w2631 = w1675 & w2630 ;
  assign w2632 = w2416 | w2422 ;
  assign w2633 = w2585 & ~w2632 ;
  assign w2634 = w2420 ^ w2633 ;
  assign w2635 = ( ~w1675 & w2623 ) | ( ~w1675 & w2629 ) | ( w2623 & w2629 ) ;
  assign w2636 = ~w2623 & w2635 ;
  assign w2637 = w2634 | w2636 ;
  assign w2638 = ( w1517 & w2631 ) | ( w1517 & ~w2637 ) | ( w2631 & ~w2637 ) ;
  assign w2639 = w1517 & w2638 ;
  assign w2640 = w2425 | w2430 ;
  assign w2641 = w2585 & ~w2640 ;
  assign w2642 = w2428 ^ w2641 ;
  assign w2643 = ( ~w1517 & w2631 ) | ( ~w1517 & w2637 ) | ( w2631 & w2637 ) ;
  assign w2644 = ~w2631 & w2643 ;
  assign w2645 = w2642 | w2644 ;
  assign w2646 = ( w1367 & w2639 ) | ( w1367 & ~w2645 ) | ( w2639 & ~w2645 ) ;
  assign w2647 = w1367 & w2646 ;
  assign w2648 = w2433 | w2438 ;
  assign w2649 = w2585 & ~w2648 ;
  assign w2650 = w2436 ^ w2649 ;
  assign w2651 = ( ~w1367 & w2639 ) | ( ~w1367 & w2645 ) | ( w2639 & w2645 ) ;
  assign w2652 = ~w2639 & w2651 ;
  assign w2653 = w2650 | w2652 ;
  assign w2654 = ( w1225 & w2647 ) | ( w1225 & ~w2653 ) | ( w2647 & ~w2653 ) ;
  assign w2655 = w1225 & w2654 ;
  assign w2656 = w2441 | w2446 ;
  assign w2657 = w2585 & ~w2656 ;
  assign w2658 = w2444 ^ w2657 ;
  assign w2659 = ( ~w1225 & w2647 ) | ( ~w1225 & w2653 ) | ( w2647 & w2653 ) ;
  assign w2660 = ~w2647 & w2659 ;
  assign w2661 = w2658 | w2660 ;
  assign w2662 = ( w1091 & w2655 ) | ( w1091 & ~w2661 ) | ( w2655 & ~w2661 ) ;
  assign w2663 = w1091 & w2662 ;
  assign w2664 = w2449 | w2454 ;
  assign w2665 = w2585 & ~w2664 ;
  assign w2666 = w2452 ^ w2665 ;
  assign w2667 = ( ~w1091 & w2655 ) | ( ~w1091 & w2661 ) | ( w2655 & w2661 ) ;
  assign w2668 = ~w2655 & w2667 ;
  assign w2669 = w2666 | w2668 ;
  assign w2670 = ( w965 & w2663 ) | ( w965 & ~w2669 ) | ( w2663 & ~w2669 ) ;
  assign w2671 = w965 & w2670 ;
  assign w2672 = w2457 | w2462 ;
  assign w2673 = w2585 & ~w2672 ;
  assign w2674 = w2460 ^ w2673 ;
  assign w2675 = ( ~w965 & w2663 ) | ( ~w965 & w2669 ) | ( w2663 & w2669 ) ;
  assign w2676 = ~w2663 & w2675 ;
  assign w2677 = w2674 | w2676 ;
  assign w2678 = ( w847 & w2671 ) | ( w847 & ~w2677 ) | ( w2671 & ~w2677 ) ;
  assign w2679 = w847 & w2678 ;
  assign w2680 = w2465 | w2470 ;
  assign w2681 = w2585 & ~w2680 ;
  assign w2682 = w2468 ^ w2681 ;
  assign w2683 = ( ~w847 & w2671 ) | ( ~w847 & w2677 ) | ( w2671 & w2677 ) ;
  assign w2684 = ~w2671 & w2683 ;
  assign w2685 = w2682 | w2684 ;
  assign w2686 = ( w737 & w2679 ) | ( w737 & ~w2685 ) | ( w2679 & ~w2685 ) ;
  assign w2687 = w737 & w2686 ;
  assign w2688 = w2473 | w2478 ;
  assign w2689 = w2585 & ~w2688 ;
  assign w2690 = w2476 ^ w2689 ;
  assign w2691 = ( ~w737 & w2679 ) | ( ~w737 & w2685 ) | ( w2679 & w2685 ) ;
  assign w2692 = ~w2679 & w2691 ;
  assign w2693 = w2690 | w2692 ;
  assign w2694 = ( w635 & w2687 ) | ( w635 & ~w2693 ) | ( w2687 & ~w2693 ) ;
  assign w2695 = w635 & w2694 ;
  assign w2696 = w2481 | w2486 ;
  assign w2697 = w2585 & ~w2696 ;
  assign w2698 = w2484 ^ w2697 ;
  assign w2699 = ( ~w635 & w2687 ) | ( ~w635 & w2693 ) | ( w2687 & w2693 ) ;
  assign w2700 = ~w2687 & w2699 ;
  assign w2701 = w2698 | w2700 ;
  assign w2702 = ( w541 & w2695 ) | ( w541 & ~w2701 ) | ( w2695 & ~w2701 ) ;
  assign w2703 = w541 & w2702 ;
  assign w2704 = w2489 | w2494 ;
  assign w2705 = w2585 & ~w2704 ;
  assign w2706 = w2492 ^ w2705 ;
  assign w2707 = ( ~w541 & w2695 ) | ( ~w541 & w2701 ) | ( w2695 & w2701 ) ;
  assign w2708 = ~w2695 & w2707 ;
  assign w2709 = w2706 | w2708 ;
  assign w2710 = ( w455 & w2703 ) | ( w455 & ~w2709 ) | ( w2703 & ~w2709 ) ;
  assign w2711 = w455 & w2710 ;
  assign w2712 = ( ~w455 & w2703 ) | ( ~w455 & w2709 ) | ( w2703 & w2709 ) ;
  assign w2713 = ~w2703 & w2712 ;
  assign w2714 = w2497 | w2499 ;
  assign w2715 = w2585 & ~w2714 ;
  assign w2716 = w2502 ^ w2715 ;
  assign w2717 = w2713 | w2716 ;
  assign w2718 = ( w377 & w2711 ) | ( w377 & ~w2717 ) | ( w2711 & ~w2717 ) ;
  assign w2719 = w377 & w2718 ;
  assign w2720 = w2505 | w2510 ;
  assign w2721 = w2585 & ~w2720 ;
  assign w2722 = w2508 ^ w2721 ;
  assign w2723 = ( ~w377 & w2711 ) | ( ~w377 & w2717 ) | ( w2711 & w2717 ) ;
  assign w2724 = ~w2711 & w2723 ;
  assign w2725 = w2722 | w2724 ;
  assign w2726 = ( w307 & w2719 ) | ( w307 & ~w2725 ) | ( w2719 & ~w2725 ) ;
  assign w2727 = w307 & w2726 ;
  assign w2728 = w2513 | w2518 ;
  assign w2729 = w2585 & ~w2728 ;
  assign w2730 = w2516 ^ w2729 ;
  assign w2731 = ( ~w307 & w2719 ) | ( ~w307 & w2725 ) | ( w2719 & w2725 ) ;
  assign w2732 = ~w2719 & w2731 ;
  assign w2733 = w2730 | w2732 ;
  assign w2734 = ( w246 & w2727 ) | ( w246 & ~w2733 ) | ( w2727 & ~w2733 ) ;
  assign w2735 = w246 & w2734 ;
  assign w2736 = w2521 | w2526 ;
  assign w2737 = w2585 & ~w2736 ;
  assign w2738 = w2524 ^ w2737 ;
  assign w2739 = ( ~w246 & w2727 ) | ( ~w246 & w2733 ) | ( w2727 & w2733 ) ;
  assign w2740 = ~w2727 & w2739 ;
  assign w2741 = w2738 | w2740 ;
  assign w2742 = ( w185 & w2735 ) | ( w185 & ~w2741 ) | ( w2735 & ~w2741 ) ;
  assign w2743 = w185 & w2742 ;
  assign w2744 = w2529 | w2534 ;
  assign w2745 = w2585 & ~w2744 ;
  assign w2746 = w2532 ^ w2745 ;
  assign w2747 = ( ~w185 & w2735 ) | ( ~w185 & w2741 ) | ( w2735 & w2741 ) ;
  assign w2748 = ~w2735 & w2747 ;
  assign w2749 = w2746 | w2748 ;
  assign w2750 = ( w145 & w2743 ) | ( w145 & ~w2749 ) | ( w2743 & ~w2749 ) ;
  assign w2751 = w145 & w2750 ;
  assign w2752 = w2537 | w2542 ;
  assign w2753 = w2585 & ~w2752 ;
  assign w2754 = w2540 ^ w2753 ;
  assign w2755 = ( ~w145 & w2743 ) | ( ~w145 & w2749 ) | ( w2743 & w2749 ) ;
  assign w2756 = ~w2743 & w2755 ;
  assign w2757 = w2754 | w2756 ;
  assign w2758 = ( w132 & w2751 ) | ( w132 & ~w2757 ) | ( w2751 & ~w2757 ) ;
  assign w2759 = w132 & w2758 ;
  assign w2760 = w2545 | w2550 ;
  assign w2761 = w2585 & ~w2760 ;
  assign w2762 = w2548 ^ w2761 ;
  assign w2763 = ( ~w132 & w2751 ) | ( ~w132 & w2757 ) | ( w2751 & w2757 ) ;
  assign w2764 = ~w2751 & w2763 ;
  assign w2765 = w2762 | w2764 ;
  assign w2766 = ~w2759 & w2765 ;
  assign w2767 = w2553 | w2558 ;
  assign w2768 = w2585 & ~w2767 ;
  assign w2769 = w2556 ^ w2768 ;
  assign w2770 = ( ~w2571 & w2766 ) | ( ~w2571 & w2769 ) | ( w2766 & w2769 ) ;
  assign w2771 = w2560 & ~w2770 ;
  assign w2772 = ~w2563 & w2585 ;
  assign w2773 = ( w2770 & ~w2771 ) | ( w2770 & w2772 ) | ( ~w2771 & w2772 ) ;
  assign w2774 = w2571 | w2773 ;
  assign w2775 = ~w129 & w2774 ;
  assign w2776 = ( w2759 & w2765 ) | ( w2759 & w2769 ) | ( w2765 & w2769 ) ;
  assign w2777 = ~w2759 & w2776 ;
  assign w2778 = ( w129 & w2560 ) | ( w129 & w2563 ) | ( w2560 & w2563 ) ;
  assign w2779 = ( w2563 & ~w2585 ) | ( w2563 & w2778 ) | ( ~w2585 & w2778 ) ;
  assign w2780 = w2560 & w2779 ;
  assign w2781 = w2778 ^ w2780 ;
  assign w2782 = ( w2355 & w2360 ) | ( w2355 & w2387 ) | ( w2360 & w2387 ) ;
  assign w2783 = w2387 & ~w2782 ;
  assign w2784 = w2358 ^ w2783 ;
  assign w2785 = ( ~w2575 & w2582 ) | ( ~w2575 & w2784 ) | ( w2582 & w2784 ) ;
  assign w2786 = ~w2582 & w2785 ;
  assign w2787 = ( ~w2569 & w2571 ) | ( ~w2569 & w2786 ) | ( w2571 & w2786 ) ;
  assign w2788 = ~w2571 & w2787 ;
  assign w2789 = w2777 | w2788 ;
  assign w2790 = ( w2775 & ~w2777 ) | ( w2775 & w2781 ) | ( ~w2777 & w2781 ) ;
  assign w2791 = w2789 | w2790 ;
  assign w2792 = ( ~\pi079 & \pi080 ) | ( ~\pi079 & w2585 ) | ( \pi080 & w2585 ) ;
  assign w2793 = ( ~\pi078 & \pi080 ) | ( ~\pi078 & w2792 ) | ( \pi080 & w2792 ) ;
  assign w2794 = ( ~\pi080 & w2585 ) | ( ~\pi080 & w2791 ) | ( w2585 & w2791 ) ;
  assign w2795 = w2793 & w2794 ;
  assign w2796 = ( w2571 & w2575 ) | ( w2571 & ~w2582 ) | ( w2575 & ~w2582 ) ;
  assign w2797 = \pi079 & ~w2796 ;
  assign w2798 = \pi078 | \pi080 ;
  assign w2799 = ( ~w2796 & w2797 ) | ( ~w2796 & w2798 ) | ( w2797 & w2798 ) ;
  assign w2800 = ~w2582 & w2799 ;
  assign w2801 = ~w2569 & w2800 ;
  assign w2802 = ( \pi080 & w2791 ) | ( \pi080 & ~w2800 ) | ( w2791 & ~w2800 ) ;
  assign w2803 = w2801 & ~w2802 ;
  assign w2804 = ~\pi080 & w2791 ;
  assign w2805 = \pi081 ^ w2804 ;
  assign w2806 = w2803 | w2805 ;
  assign w2807 = ( w2387 & w2795 ) | ( w2387 & ~w2806 ) | ( w2795 & ~w2806 ) ;
  assign w2808 = w2387 & w2807 ;
  assign w2809 = ( ~w2387 & w2795 ) | ( ~w2387 & w2806 ) | ( w2795 & w2806 ) ;
  assign w2810 = ~w2795 & w2809 ;
  assign w2811 = w2585 & ~w2788 ;
  assign w2812 = ~w2777 & w2811 ;
  assign w2813 = ~w2790 & w2812 ;
  assign w2814 = \pi081 & w2791 ;
  assign w2815 = ( \pi080 & w2791 ) | ( \pi080 & ~w2814 ) | ( w2791 & ~w2814 ) ;
  assign w2816 = ( ~\pi080 & w2813 ) | ( ~\pi080 & w2815 ) | ( w2813 & w2815 ) ;
  assign w2817 = \pi082 ^ w2816 ;
  assign w2818 = w2810 | w2817 ;
  assign w2819 = ( w2197 & w2808 ) | ( w2197 & ~w2818 ) | ( w2808 & ~w2818 ) ;
  assign w2820 = w2197 & w2819 ;
  assign w2821 = ( w2589 & ~w2597 ) | ( w2589 & w2791 ) | ( ~w2597 & w2791 ) ;
  assign w2822 = ~w2589 & w2821 ;
  assign w2823 = \pi083 ^ w2822 ;
  assign w2824 = w2598 ^ w2823 ;
  assign w2825 = ( ~w2197 & w2808 ) | ( ~w2197 & w2818 ) | ( w2808 & w2818 ) ;
  assign w2826 = ~w2808 & w2825 ;
  assign w2827 = w2824 | w2826 ;
  assign w2828 = ( w2015 & w2820 ) | ( w2015 & ~w2827 ) | ( w2820 & ~w2827 ) ;
  assign w2829 = w2015 & w2828 ;
  assign w2830 = w2602 | w2604 ;
  assign w2831 = w2791 & ~w2830 ;
  assign w2832 = w2611 ^ w2831 ;
  assign w2833 = ( ~w2015 & w2820 ) | ( ~w2015 & w2827 ) | ( w2820 & w2827 ) ;
  assign w2834 = ~w2820 & w2833 ;
  assign w2835 = w2832 | w2834 ;
  assign w2836 = ( w1841 & w2829 ) | ( w1841 & ~w2835 ) | ( w2829 & ~w2835 ) ;
  assign w2837 = w1841 & w2836 ;
  assign w2838 = w2614 | w2620 ;
  assign w2839 = w2791 & ~w2838 ;
  assign w2840 = w2618 ^ w2839 ;
  assign w2841 = ( ~w1841 & w2829 ) | ( ~w1841 & w2835 ) | ( w2829 & w2835 ) ;
  assign w2842 = ~w2829 & w2841 ;
  assign w2843 = w2840 | w2842 ;
  assign w2844 = ( w1675 & w2837 ) | ( w1675 & ~w2843 ) | ( w2837 & ~w2843 ) ;
  assign w2845 = w1675 & w2844 ;
  assign w2846 = w2623 | w2628 ;
  assign w2847 = w2791 & ~w2846 ;
  assign w2848 = w2626 ^ w2847 ;
  assign w2849 = ( ~w1675 & w2837 ) | ( ~w1675 & w2843 ) | ( w2837 & w2843 ) ;
  assign w2850 = ~w2837 & w2849 ;
  assign w2851 = w2848 | w2850 ;
  assign w2852 = ( w1517 & w2845 ) | ( w1517 & ~w2851 ) | ( w2845 & ~w2851 ) ;
  assign w2853 = w1517 & w2852 ;
  assign w2854 = w2631 | w2636 ;
  assign w2855 = w2791 & ~w2854 ;
  assign w2856 = w2634 ^ w2855 ;
  assign w2857 = ( ~w1517 & w2845 ) | ( ~w1517 & w2851 ) | ( w2845 & w2851 ) ;
  assign w2858 = ~w2845 & w2857 ;
  assign w2859 = w2856 | w2858 ;
  assign w2860 = ( w1367 & w2853 ) | ( w1367 & ~w2859 ) | ( w2853 & ~w2859 ) ;
  assign w2861 = w1367 & w2860 ;
  assign w2862 = w2639 | w2644 ;
  assign w2863 = w2791 & ~w2862 ;
  assign w2864 = w2642 ^ w2863 ;
  assign w2865 = ( ~w1367 & w2853 ) | ( ~w1367 & w2859 ) | ( w2853 & w2859 ) ;
  assign w2866 = ~w2853 & w2865 ;
  assign w2867 = w2864 | w2866 ;
  assign w2868 = ( w1225 & w2861 ) | ( w1225 & ~w2867 ) | ( w2861 & ~w2867 ) ;
  assign w2869 = w1225 & w2868 ;
  assign w2870 = w2647 | w2652 ;
  assign w2871 = w2791 & ~w2870 ;
  assign w2872 = w2650 ^ w2871 ;
  assign w2873 = ( ~w1225 & w2861 ) | ( ~w1225 & w2867 ) | ( w2861 & w2867 ) ;
  assign w2874 = ~w2861 & w2873 ;
  assign w2875 = w2872 | w2874 ;
  assign w2876 = ( w1091 & w2869 ) | ( w1091 & ~w2875 ) | ( w2869 & ~w2875 ) ;
  assign w2877 = w1091 & w2876 ;
  assign w2878 = w2655 | w2660 ;
  assign w2879 = w2791 & ~w2878 ;
  assign w2880 = w2658 ^ w2879 ;
  assign w2881 = ( ~w1091 & w2869 ) | ( ~w1091 & w2875 ) | ( w2869 & w2875 ) ;
  assign w2882 = ~w2869 & w2881 ;
  assign w2883 = w2880 | w2882 ;
  assign w2884 = ( w965 & w2877 ) | ( w965 & ~w2883 ) | ( w2877 & ~w2883 ) ;
  assign w2885 = w965 & w2884 ;
  assign w2886 = w2663 | w2668 ;
  assign w2887 = w2791 & ~w2886 ;
  assign w2888 = w2666 ^ w2887 ;
  assign w2889 = ( ~w965 & w2877 ) | ( ~w965 & w2883 ) | ( w2877 & w2883 ) ;
  assign w2890 = ~w2877 & w2889 ;
  assign w2891 = w2888 | w2890 ;
  assign w2892 = ( w847 & w2885 ) | ( w847 & ~w2891 ) | ( w2885 & ~w2891 ) ;
  assign w2893 = w847 & w2892 ;
  assign w2894 = w2671 | w2676 ;
  assign w2895 = w2791 & ~w2894 ;
  assign w2896 = w2674 ^ w2895 ;
  assign w2897 = ( ~w847 & w2885 ) | ( ~w847 & w2891 ) | ( w2885 & w2891 ) ;
  assign w2898 = ~w2885 & w2897 ;
  assign w2899 = w2896 | w2898 ;
  assign w2900 = ( w737 & w2893 ) | ( w737 & ~w2899 ) | ( w2893 & ~w2899 ) ;
  assign w2901 = w737 & w2900 ;
  assign w2902 = w2679 | w2684 ;
  assign w2903 = w2791 & ~w2902 ;
  assign w2904 = w2682 ^ w2903 ;
  assign w2905 = ( ~w737 & w2893 ) | ( ~w737 & w2899 ) | ( w2893 & w2899 ) ;
  assign w2906 = ~w2893 & w2905 ;
  assign w2907 = w2904 | w2906 ;
  assign w2908 = ( w635 & w2901 ) | ( w635 & ~w2907 ) | ( w2901 & ~w2907 ) ;
  assign w2909 = w635 & w2908 ;
  assign w2910 = w2687 | w2692 ;
  assign w2911 = w2791 & ~w2910 ;
  assign w2912 = w2690 ^ w2911 ;
  assign w2913 = ( ~w635 & w2901 ) | ( ~w635 & w2907 ) | ( w2901 & w2907 ) ;
  assign w2914 = ~w2901 & w2913 ;
  assign w2915 = w2912 | w2914 ;
  assign w2916 = ( w541 & w2909 ) | ( w541 & ~w2915 ) | ( w2909 & ~w2915 ) ;
  assign w2917 = w541 & w2916 ;
  assign w2918 = w2695 | w2700 ;
  assign w2919 = w2791 & ~w2918 ;
  assign w2920 = w2698 ^ w2919 ;
  assign w2921 = ( ~w541 & w2909 ) | ( ~w541 & w2915 ) | ( w2909 & w2915 ) ;
  assign w2922 = ~w2909 & w2921 ;
  assign w2923 = w2920 | w2922 ;
  assign w2924 = ( w455 & w2917 ) | ( w455 & ~w2923 ) | ( w2917 & ~w2923 ) ;
  assign w2925 = w455 & w2924 ;
  assign w2926 = w2703 | w2708 ;
  assign w2927 = w2791 & ~w2926 ;
  assign w2928 = w2706 ^ w2927 ;
  assign w2929 = ( ~w455 & w2917 ) | ( ~w455 & w2923 ) | ( w2917 & w2923 ) ;
  assign w2930 = ~w2917 & w2929 ;
  assign w2931 = w2928 | w2930 ;
  assign w2932 = ( w377 & w2925 ) | ( w377 & ~w2931 ) | ( w2925 & ~w2931 ) ;
  assign w2933 = w377 & w2932 ;
  assign w2934 = ( ~w377 & w2925 ) | ( ~w377 & w2931 ) | ( w2925 & w2931 ) ;
  assign w2935 = ~w2925 & w2934 ;
  assign w2936 = w2711 | w2713 ;
  assign w2937 = w2791 & ~w2936 ;
  assign w2938 = w2716 ^ w2937 ;
  assign w2939 = w2935 | w2938 ;
  assign w2940 = ( w307 & w2933 ) | ( w307 & ~w2939 ) | ( w2933 & ~w2939 ) ;
  assign w2941 = w307 & w2940 ;
  assign w2942 = w2719 | w2724 ;
  assign w2943 = w2791 & ~w2942 ;
  assign w2944 = w2722 ^ w2943 ;
  assign w2945 = ( ~w307 & w2933 ) | ( ~w307 & w2939 ) | ( w2933 & w2939 ) ;
  assign w2946 = ~w2933 & w2945 ;
  assign w2947 = w2944 | w2946 ;
  assign w2948 = ( w246 & w2941 ) | ( w246 & ~w2947 ) | ( w2941 & ~w2947 ) ;
  assign w2949 = w246 & w2948 ;
  assign w2950 = w2727 | w2732 ;
  assign w2951 = w2791 & ~w2950 ;
  assign w2952 = w2730 ^ w2951 ;
  assign w2953 = ( ~w246 & w2941 ) | ( ~w246 & w2947 ) | ( w2941 & w2947 ) ;
  assign w2954 = ~w2941 & w2953 ;
  assign w2955 = w2952 | w2954 ;
  assign w2956 = ( w185 & w2949 ) | ( w185 & ~w2955 ) | ( w2949 & ~w2955 ) ;
  assign w2957 = w185 & w2956 ;
  assign w2958 = w2735 | w2740 ;
  assign w2959 = w2791 & ~w2958 ;
  assign w2960 = w2738 ^ w2959 ;
  assign w2961 = ( ~w185 & w2949 ) | ( ~w185 & w2955 ) | ( w2949 & w2955 ) ;
  assign w2962 = ~w2949 & w2961 ;
  assign w2963 = w2960 | w2962 ;
  assign w2964 = ( w145 & w2957 ) | ( w145 & ~w2963 ) | ( w2957 & ~w2963 ) ;
  assign w2965 = w145 & w2964 ;
  assign w2966 = w2743 | w2748 ;
  assign w2967 = w2791 & ~w2966 ;
  assign w2968 = w2746 ^ w2967 ;
  assign w2969 = ( ~w145 & w2957 ) | ( ~w145 & w2963 ) | ( w2957 & w2963 ) ;
  assign w2970 = ~w2957 & w2969 ;
  assign w2971 = w2968 | w2970 ;
  assign w2972 = ( w132 & w2965 ) | ( w132 & ~w2971 ) | ( w2965 & ~w2971 ) ;
  assign w2973 = w132 & w2972 ;
  assign w2974 = w2751 | w2756 ;
  assign w2975 = w2791 & ~w2974 ;
  assign w2976 = w2754 ^ w2975 ;
  assign w2977 = ( ~w132 & w2965 ) | ( ~w132 & w2971 ) | ( w2965 & w2971 ) ;
  assign w2978 = ~w2965 & w2977 ;
  assign w2979 = w2976 | w2978 ;
  assign w2980 = ~w2973 & w2979 ;
  assign w2981 = w2759 | w2764 ;
  assign w2982 = w2791 & ~w2981 ;
  assign w2983 = w2762 ^ w2982 ;
  assign w2984 = ( ~w2777 & w2980 ) | ( ~w2777 & w2983 ) | ( w2980 & w2983 ) ;
  assign w2985 = w2766 & ~w2984 ;
  assign w2986 = ~w2769 & w2791 ;
  assign w2987 = ( w2984 & ~w2985 ) | ( w2984 & w2986 ) | ( ~w2985 & w2986 ) ;
  assign w2988 = w2777 | w2987 ;
  assign w2989 = ~w129 & w2988 ;
  assign w2990 = ( w2973 & w2979 ) | ( w2973 & w2983 ) | ( w2979 & w2983 ) ;
  assign w2991 = ~w2973 & w2990 ;
  assign w2992 = ( w129 & w2766 ) | ( w129 & w2769 ) | ( w2766 & w2769 ) ;
  assign w2993 = ( w2769 & ~w2791 ) | ( w2769 & w2992 ) | ( ~w2791 & w2992 ) ;
  assign w2994 = w2766 & w2993 ;
  assign w2995 = w2992 ^ w2994 ;
  assign w2996 = ( w2553 & w2558 ) | ( w2553 & w2585 ) | ( w2558 & w2585 ) ;
  assign w2997 = w2585 & ~w2996 ;
  assign w2998 = w2556 ^ w2997 ;
  assign w2999 = ( ~w2781 & w2788 ) | ( ~w2781 & w2998 ) | ( w2788 & w2998 ) ;
  assign w3000 = ~w2788 & w2999 ;
  assign w3001 = ( ~w2775 & w2777 ) | ( ~w2775 & w3000 ) | ( w2777 & w3000 ) ;
  assign w3002 = ~w2777 & w3001 ;
  assign w3003 = w2991 | w3002 ;
  assign w3004 = ( w2989 & ~w2991 ) | ( w2989 & w2995 ) | ( ~w2991 & w2995 ) ;
  assign w3005 = w3003 | w3004 ;
  assign w3006 = ( ~\pi077 & \pi078 ) | ( ~\pi077 & w2791 ) | ( \pi078 & w2791 ) ;
  assign w3007 = ( ~\pi076 & \pi078 ) | ( ~\pi076 & w3006 ) | ( \pi078 & w3006 ) ;
  assign w3008 = ( ~\pi078 & w2791 ) | ( ~\pi078 & w3005 ) | ( w2791 & w3005 ) ;
  assign w3009 = w3007 & w3008 ;
  assign w3010 = ( w2777 & w2781 ) | ( w2777 & ~w2788 ) | ( w2781 & ~w2788 ) ;
  assign w3011 = \pi077 & ~w3010 ;
  assign w3012 = \pi076 | \pi078 ;
  assign w3013 = ( ~w3010 & w3011 ) | ( ~w3010 & w3012 ) | ( w3011 & w3012 ) ;
  assign w3014 = ~w2788 & w3013 ;
  assign w3015 = ~w2775 & w3014 ;
  assign w3016 = ( \pi078 & w3005 ) | ( \pi078 & ~w3014 ) | ( w3005 & ~w3014 ) ;
  assign w3017 = w3015 & ~w3016 ;
  assign w3018 = ~\pi078 & w3005 ;
  assign w3019 = \pi079 ^ w3018 ;
  assign w3020 = w3017 | w3019 ;
  assign w3021 = ( w2585 & w3009 ) | ( w2585 & ~w3020 ) | ( w3009 & ~w3020 ) ;
  assign w3022 = w2585 & w3021 ;
  assign w3023 = ( ~w2585 & w3009 ) | ( ~w2585 & w3020 ) | ( w3009 & w3020 ) ;
  assign w3024 = ~w3009 & w3023 ;
  assign w3025 = w2791 & ~w3002 ;
  assign w3026 = ~w2991 & w3025 ;
  assign w3027 = ~w3004 & w3026 ;
  assign w3028 = \pi079 & w3005 ;
  assign w3029 = ( \pi078 & w3005 ) | ( \pi078 & ~w3028 ) | ( w3005 & ~w3028 ) ;
  assign w3030 = ( ~\pi078 & w3027 ) | ( ~\pi078 & w3029 ) | ( w3027 & w3029 ) ;
  assign w3031 = \pi080 ^ w3030 ;
  assign w3032 = w3024 | w3031 ;
  assign w3033 = ( w2387 & w3022 ) | ( w2387 & ~w3032 ) | ( w3022 & ~w3032 ) ;
  assign w3034 = w2387 & w3033 ;
  assign w3035 = ( w2795 & ~w2803 ) | ( w2795 & w3005 ) | ( ~w2803 & w3005 ) ;
  assign w3036 = ~w2795 & w3035 ;
  assign w3037 = \pi081 ^ w3036 ;
  assign w3038 = w2804 ^ w3037 ;
  assign w3039 = ( ~w2387 & w3022 ) | ( ~w2387 & w3032 ) | ( w3022 & w3032 ) ;
  assign w3040 = ~w3022 & w3039 ;
  assign w3041 = w3038 | w3040 ;
  assign w3042 = ( w2197 & w3034 ) | ( w2197 & ~w3041 ) | ( w3034 & ~w3041 ) ;
  assign w3043 = w2197 & w3042 ;
  assign w3044 = w2808 | w2810 ;
  assign w3045 = w3005 & ~w3044 ;
  assign w3046 = w2817 ^ w3045 ;
  assign w3047 = ( ~w2197 & w3034 ) | ( ~w2197 & w3041 ) | ( w3034 & w3041 ) ;
  assign w3048 = ~w3034 & w3047 ;
  assign w3049 = w3046 | w3048 ;
  assign w3050 = ( w2015 & w3043 ) | ( w2015 & ~w3049 ) | ( w3043 & ~w3049 ) ;
  assign w3051 = w2015 & w3050 ;
  assign w3052 = w2820 | w2826 ;
  assign w3053 = w3005 & ~w3052 ;
  assign w3054 = w2824 ^ w3053 ;
  assign w3055 = ( ~w2015 & w3043 ) | ( ~w2015 & w3049 ) | ( w3043 & w3049 ) ;
  assign w3056 = ~w3043 & w3055 ;
  assign w3057 = w3054 | w3056 ;
  assign w3058 = ( w1841 & w3051 ) | ( w1841 & ~w3057 ) | ( w3051 & ~w3057 ) ;
  assign w3059 = w1841 & w3058 ;
  assign w3060 = w2829 | w2834 ;
  assign w3061 = w3005 & ~w3060 ;
  assign w3062 = w2832 ^ w3061 ;
  assign w3063 = ( ~w1841 & w3051 ) | ( ~w1841 & w3057 ) | ( w3051 & w3057 ) ;
  assign w3064 = ~w3051 & w3063 ;
  assign w3065 = w3062 | w3064 ;
  assign w3066 = ( w1675 & w3059 ) | ( w1675 & ~w3065 ) | ( w3059 & ~w3065 ) ;
  assign w3067 = w1675 & w3066 ;
  assign w3068 = w2837 | w2842 ;
  assign w3069 = w3005 & ~w3068 ;
  assign w3070 = w2840 ^ w3069 ;
  assign w3071 = ( ~w1675 & w3059 ) | ( ~w1675 & w3065 ) | ( w3059 & w3065 ) ;
  assign w3072 = ~w3059 & w3071 ;
  assign w3073 = w3070 | w3072 ;
  assign w3074 = ( w1517 & w3067 ) | ( w1517 & ~w3073 ) | ( w3067 & ~w3073 ) ;
  assign w3075 = w1517 & w3074 ;
  assign w3076 = w2845 | w2850 ;
  assign w3077 = w3005 & ~w3076 ;
  assign w3078 = w2848 ^ w3077 ;
  assign w3079 = ( ~w1517 & w3067 ) | ( ~w1517 & w3073 ) | ( w3067 & w3073 ) ;
  assign w3080 = ~w3067 & w3079 ;
  assign w3081 = w3078 | w3080 ;
  assign w3082 = ( w1367 & w3075 ) | ( w1367 & ~w3081 ) | ( w3075 & ~w3081 ) ;
  assign w3083 = w1367 & w3082 ;
  assign w3084 = w2853 | w2858 ;
  assign w3085 = w3005 & ~w3084 ;
  assign w3086 = w2856 ^ w3085 ;
  assign w3087 = ( ~w1367 & w3075 ) | ( ~w1367 & w3081 ) | ( w3075 & w3081 ) ;
  assign w3088 = ~w3075 & w3087 ;
  assign w3089 = w3086 | w3088 ;
  assign w3090 = ( w1225 & w3083 ) | ( w1225 & ~w3089 ) | ( w3083 & ~w3089 ) ;
  assign w3091 = w1225 & w3090 ;
  assign w3092 = w2861 | w2866 ;
  assign w3093 = w3005 & ~w3092 ;
  assign w3094 = w2864 ^ w3093 ;
  assign w3095 = ( ~w1225 & w3083 ) | ( ~w1225 & w3089 ) | ( w3083 & w3089 ) ;
  assign w3096 = ~w3083 & w3095 ;
  assign w3097 = w3094 | w3096 ;
  assign w3098 = ( w1091 & w3091 ) | ( w1091 & ~w3097 ) | ( w3091 & ~w3097 ) ;
  assign w3099 = w1091 & w3098 ;
  assign w3100 = w2869 | w2874 ;
  assign w3101 = w3005 & ~w3100 ;
  assign w3102 = w2872 ^ w3101 ;
  assign w3103 = ( ~w1091 & w3091 ) | ( ~w1091 & w3097 ) | ( w3091 & w3097 ) ;
  assign w3104 = ~w3091 & w3103 ;
  assign w3105 = w3102 | w3104 ;
  assign w3106 = ( w965 & w3099 ) | ( w965 & ~w3105 ) | ( w3099 & ~w3105 ) ;
  assign w3107 = w965 & w3106 ;
  assign w3108 = w2877 | w2882 ;
  assign w3109 = w3005 & ~w3108 ;
  assign w3110 = w2880 ^ w3109 ;
  assign w3111 = ( ~w965 & w3099 ) | ( ~w965 & w3105 ) | ( w3099 & w3105 ) ;
  assign w3112 = ~w3099 & w3111 ;
  assign w3113 = w3110 | w3112 ;
  assign w3114 = ( w847 & w3107 ) | ( w847 & ~w3113 ) | ( w3107 & ~w3113 ) ;
  assign w3115 = w847 & w3114 ;
  assign w3116 = w2885 | w2890 ;
  assign w3117 = w3005 & ~w3116 ;
  assign w3118 = w2888 ^ w3117 ;
  assign w3119 = ( ~w847 & w3107 ) | ( ~w847 & w3113 ) | ( w3107 & w3113 ) ;
  assign w3120 = ~w3107 & w3119 ;
  assign w3121 = w3118 | w3120 ;
  assign w3122 = ( w737 & w3115 ) | ( w737 & ~w3121 ) | ( w3115 & ~w3121 ) ;
  assign w3123 = w737 & w3122 ;
  assign w3124 = w2893 | w2898 ;
  assign w3125 = w3005 & ~w3124 ;
  assign w3126 = w2896 ^ w3125 ;
  assign w3127 = ( ~w737 & w3115 ) | ( ~w737 & w3121 ) | ( w3115 & w3121 ) ;
  assign w3128 = ~w3115 & w3127 ;
  assign w3129 = w3126 | w3128 ;
  assign w3130 = ( w635 & w3123 ) | ( w635 & ~w3129 ) | ( w3123 & ~w3129 ) ;
  assign w3131 = w635 & w3130 ;
  assign w3132 = w2901 | w2906 ;
  assign w3133 = w3005 & ~w3132 ;
  assign w3134 = w2904 ^ w3133 ;
  assign w3135 = ( ~w635 & w3123 ) | ( ~w635 & w3129 ) | ( w3123 & w3129 ) ;
  assign w3136 = ~w3123 & w3135 ;
  assign w3137 = w3134 | w3136 ;
  assign w3138 = ( w541 & w3131 ) | ( w541 & ~w3137 ) | ( w3131 & ~w3137 ) ;
  assign w3139 = w541 & w3138 ;
  assign w3140 = w2909 | w2914 ;
  assign w3141 = w3005 & ~w3140 ;
  assign w3142 = w2912 ^ w3141 ;
  assign w3143 = ( ~w541 & w3131 ) | ( ~w541 & w3137 ) | ( w3131 & w3137 ) ;
  assign w3144 = ~w3131 & w3143 ;
  assign w3145 = w3142 | w3144 ;
  assign w3146 = ( w455 & w3139 ) | ( w455 & ~w3145 ) | ( w3139 & ~w3145 ) ;
  assign w3147 = w455 & w3146 ;
  assign w3148 = w2917 | w2922 ;
  assign w3149 = w3005 & ~w3148 ;
  assign w3150 = w2920 ^ w3149 ;
  assign w3151 = ( ~w455 & w3139 ) | ( ~w455 & w3145 ) | ( w3139 & w3145 ) ;
  assign w3152 = ~w3139 & w3151 ;
  assign w3153 = w3150 | w3152 ;
  assign w3154 = ( w377 & w3147 ) | ( w377 & ~w3153 ) | ( w3147 & ~w3153 ) ;
  assign w3155 = w377 & w3154 ;
  assign w3156 = w2925 | w2930 ;
  assign w3157 = w3005 & ~w3156 ;
  assign w3158 = w2928 ^ w3157 ;
  assign w3159 = ( ~w377 & w3147 ) | ( ~w377 & w3153 ) | ( w3147 & w3153 ) ;
  assign w3160 = ~w3147 & w3159 ;
  assign w3161 = w3158 | w3160 ;
  assign w3162 = ( w307 & w3155 ) | ( w307 & ~w3161 ) | ( w3155 & ~w3161 ) ;
  assign w3163 = w307 & w3162 ;
  assign w3164 = ( ~w307 & w3155 ) | ( ~w307 & w3161 ) | ( w3155 & w3161 ) ;
  assign w3165 = ~w3155 & w3164 ;
  assign w3166 = w2933 | w2935 ;
  assign w3167 = w3005 & ~w3166 ;
  assign w3168 = w2938 ^ w3167 ;
  assign w3169 = w3165 | w3168 ;
  assign w3170 = ( w246 & w3163 ) | ( w246 & ~w3169 ) | ( w3163 & ~w3169 ) ;
  assign w3171 = w246 & w3170 ;
  assign w3172 = w2941 | w2946 ;
  assign w3173 = w3005 & ~w3172 ;
  assign w3174 = w2944 ^ w3173 ;
  assign w3175 = ( ~w246 & w3163 ) | ( ~w246 & w3169 ) | ( w3163 & w3169 ) ;
  assign w3176 = ~w3163 & w3175 ;
  assign w3177 = w3174 | w3176 ;
  assign w3178 = ( w185 & w3171 ) | ( w185 & ~w3177 ) | ( w3171 & ~w3177 ) ;
  assign w3179 = w185 & w3178 ;
  assign w3180 = w2949 | w2954 ;
  assign w3181 = w3005 & ~w3180 ;
  assign w3182 = w2952 ^ w3181 ;
  assign w3183 = ( ~w185 & w3171 ) | ( ~w185 & w3177 ) | ( w3171 & w3177 ) ;
  assign w3184 = ~w3171 & w3183 ;
  assign w3185 = w3182 | w3184 ;
  assign w3186 = ( w145 & w3179 ) | ( w145 & ~w3185 ) | ( w3179 & ~w3185 ) ;
  assign w3187 = w145 & w3186 ;
  assign w3188 = w2957 | w2962 ;
  assign w3189 = w3005 & ~w3188 ;
  assign w3190 = w2960 ^ w3189 ;
  assign w3191 = ( ~w145 & w3179 ) | ( ~w145 & w3185 ) | ( w3179 & w3185 ) ;
  assign w3192 = ~w3179 & w3191 ;
  assign w3193 = w3190 | w3192 ;
  assign w3194 = ( w132 & w3187 ) | ( w132 & ~w3193 ) | ( w3187 & ~w3193 ) ;
  assign w3195 = w132 & w3194 ;
  assign w3196 = w2965 | w2970 ;
  assign w3197 = w3005 & ~w3196 ;
  assign w3198 = w2968 ^ w3197 ;
  assign w3199 = ( ~w132 & w3187 ) | ( ~w132 & w3193 ) | ( w3187 & w3193 ) ;
  assign w3200 = ~w3187 & w3199 ;
  assign w3201 = w3198 | w3200 ;
  assign w3202 = ~w3195 & w3201 ;
  assign w3203 = w2973 | w2978 ;
  assign w3204 = w3005 & ~w3203 ;
  assign w3205 = w2976 ^ w3204 ;
  assign w3206 = ( ~w2991 & w3202 ) | ( ~w2991 & w3205 ) | ( w3202 & w3205 ) ;
  assign w3207 = w2980 & ~w3206 ;
  assign w3208 = ~w2983 & w3005 ;
  assign w3209 = ( w3206 & ~w3207 ) | ( w3206 & w3208 ) | ( ~w3207 & w3208 ) ;
  assign w3210 = w2991 | w3209 ;
  assign w3211 = ~w129 & w3210 ;
  assign w3212 = ( w3195 & w3201 ) | ( w3195 & w3205 ) | ( w3201 & w3205 ) ;
  assign w3213 = ~w3195 & w3212 ;
  assign w3214 = ( w129 & w2980 ) | ( w129 & w2983 ) | ( w2980 & w2983 ) ;
  assign w3215 = ( w2983 & ~w3005 ) | ( w2983 & w3214 ) | ( ~w3005 & w3214 ) ;
  assign w3216 = w2980 & w3215 ;
  assign w3217 = w3214 ^ w3216 ;
  assign w3218 = ( w2759 & w2764 ) | ( w2759 & w2791 ) | ( w2764 & w2791 ) ;
  assign w3219 = w2791 & ~w3218 ;
  assign w3220 = w2762 ^ w3219 ;
  assign w3221 = ( ~w2995 & w3002 ) | ( ~w2995 & w3220 ) | ( w3002 & w3220 ) ;
  assign w3222 = ~w3002 & w3221 ;
  assign w3223 = ( ~w2989 & w2991 ) | ( ~w2989 & w3222 ) | ( w2991 & w3222 ) ;
  assign w3224 = ~w2991 & w3223 ;
  assign w3225 = w3213 | w3224 ;
  assign w3226 = ( w3211 & ~w3213 ) | ( w3211 & w3217 ) | ( ~w3213 & w3217 ) ;
  assign w3227 = w3225 | w3226 ;
  assign w3228 = ( ~\pi075 & \pi076 ) | ( ~\pi075 & w3005 ) | ( \pi076 & w3005 ) ;
  assign w3229 = ( ~\pi074 & \pi076 ) | ( ~\pi074 & w3228 ) | ( \pi076 & w3228 ) ;
  assign w3230 = ( ~\pi076 & w3005 ) | ( ~\pi076 & w3227 ) | ( w3005 & w3227 ) ;
  assign w3231 = w3229 & w3230 ;
  assign w3232 = ( w2991 & w2995 ) | ( w2991 & ~w3002 ) | ( w2995 & ~w3002 ) ;
  assign w3233 = \pi075 & ~w3232 ;
  assign w3234 = \pi074 | \pi076 ;
  assign w3235 = ( ~w3232 & w3233 ) | ( ~w3232 & w3234 ) | ( w3233 & w3234 ) ;
  assign w3236 = ~w3002 & w3235 ;
  assign w3237 = ~w2989 & w3236 ;
  assign w3238 = ( \pi076 & w3227 ) | ( \pi076 & ~w3236 ) | ( w3227 & ~w3236 ) ;
  assign w3239 = w3237 & ~w3238 ;
  assign w3240 = ~\pi076 & w3227 ;
  assign w3241 = \pi077 ^ w3240 ;
  assign w3242 = w3239 | w3241 ;
  assign w3243 = ( w2791 & w3231 ) | ( w2791 & ~w3242 ) | ( w3231 & ~w3242 ) ;
  assign w3244 = w2791 & w3243 ;
  assign w3245 = ( ~w2791 & w3231 ) | ( ~w2791 & w3242 ) | ( w3231 & w3242 ) ;
  assign w3246 = ~w3231 & w3245 ;
  assign w3247 = w3005 & ~w3224 ;
  assign w3248 = ~w3213 & w3247 ;
  assign w3249 = ~w3226 & w3248 ;
  assign w3250 = \pi077 & w3227 ;
  assign w3251 = ( \pi076 & w3227 ) | ( \pi076 & ~w3250 ) | ( w3227 & ~w3250 ) ;
  assign w3252 = ( ~\pi076 & w3249 ) | ( ~\pi076 & w3251 ) | ( w3249 & w3251 ) ;
  assign w3253 = \pi078 ^ w3252 ;
  assign w3254 = w3246 | w3253 ;
  assign w3255 = ( w2585 & w3244 ) | ( w2585 & ~w3254 ) | ( w3244 & ~w3254 ) ;
  assign w3256 = w2585 & w3255 ;
  assign w3257 = ( w3009 & ~w3017 ) | ( w3009 & w3227 ) | ( ~w3017 & w3227 ) ;
  assign w3258 = ~w3009 & w3257 ;
  assign w3259 = \pi079 ^ w3258 ;
  assign w3260 = w3018 ^ w3259 ;
  assign w3261 = ( ~w2585 & w3244 ) | ( ~w2585 & w3254 ) | ( w3244 & w3254 ) ;
  assign w3262 = ~w3244 & w3261 ;
  assign w3263 = w3260 | w3262 ;
  assign w3264 = ( w2387 & w3256 ) | ( w2387 & ~w3263 ) | ( w3256 & ~w3263 ) ;
  assign w3265 = w2387 & w3264 ;
  assign w3266 = w3022 | w3024 ;
  assign w3267 = w3227 & ~w3266 ;
  assign w3268 = w3031 ^ w3267 ;
  assign w3269 = ( ~w2387 & w3256 ) | ( ~w2387 & w3263 ) | ( w3256 & w3263 ) ;
  assign w3270 = ~w3256 & w3269 ;
  assign w3271 = w3268 | w3270 ;
  assign w3272 = ( w2197 & w3265 ) | ( w2197 & ~w3271 ) | ( w3265 & ~w3271 ) ;
  assign w3273 = w2197 & w3272 ;
  assign w3274 = w3034 | w3040 ;
  assign w3275 = w3227 & ~w3274 ;
  assign w3276 = w3038 ^ w3275 ;
  assign w3277 = ( ~w2197 & w3265 ) | ( ~w2197 & w3271 ) | ( w3265 & w3271 ) ;
  assign w3278 = ~w3265 & w3277 ;
  assign w3279 = w3276 | w3278 ;
  assign w3280 = ( w2015 & w3273 ) | ( w2015 & ~w3279 ) | ( w3273 & ~w3279 ) ;
  assign w3281 = w2015 & w3280 ;
  assign w3282 = w3043 | w3048 ;
  assign w3283 = w3227 & ~w3282 ;
  assign w3284 = w3046 ^ w3283 ;
  assign w3285 = ( ~w2015 & w3273 ) | ( ~w2015 & w3279 ) | ( w3273 & w3279 ) ;
  assign w3286 = ~w3273 & w3285 ;
  assign w3287 = w3284 | w3286 ;
  assign w3288 = ( w1841 & w3281 ) | ( w1841 & ~w3287 ) | ( w3281 & ~w3287 ) ;
  assign w3289 = w1841 & w3288 ;
  assign w3290 = w3051 | w3056 ;
  assign w3291 = w3227 & ~w3290 ;
  assign w3292 = w3054 ^ w3291 ;
  assign w3293 = ( ~w1841 & w3281 ) | ( ~w1841 & w3287 ) | ( w3281 & w3287 ) ;
  assign w3294 = ~w3281 & w3293 ;
  assign w3295 = w3292 | w3294 ;
  assign w3296 = ( w1675 & w3289 ) | ( w1675 & ~w3295 ) | ( w3289 & ~w3295 ) ;
  assign w3297 = w1675 & w3296 ;
  assign w3298 = w3059 | w3064 ;
  assign w3299 = w3227 & ~w3298 ;
  assign w3300 = w3062 ^ w3299 ;
  assign w3301 = ( ~w1675 & w3289 ) | ( ~w1675 & w3295 ) | ( w3289 & w3295 ) ;
  assign w3302 = ~w3289 & w3301 ;
  assign w3303 = w3300 | w3302 ;
  assign w3304 = ( w1517 & w3297 ) | ( w1517 & ~w3303 ) | ( w3297 & ~w3303 ) ;
  assign w3305 = w1517 & w3304 ;
  assign w3306 = w3067 | w3072 ;
  assign w3307 = w3227 & ~w3306 ;
  assign w3308 = w3070 ^ w3307 ;
  assign w3309 = ( ~w1517 & w3297 ) | ( ~w1517 & w3303 ) | ( w3297 & w3303 ) ;
  assign w3310 = ~w3297 & w3309 ;
  assign w3311 = w3308 | w3310 ;
  assign w3312 = ( w1367 & w3305 ) | ( w1367 & ~w3311 ) | ( w3305 & ~w3311 ) ;
  assign w3313 = w1367 & w3312 ;
  assign w3314 = w3075 | w3080 ;
  assign w3315 = w3227 & ~w3314 ;
  assign w3316 = w3078 ^ w3315 ;
  assign w3317 = ( ~w1367 & w3305 ) | ( ~w1367 & w3311 ) | ( w3305 & w3311 ) ;
  assign w3318 = ~w3305 & w3317 ;
  assign w3319 = w3316 | w3318 ;
  assign w3320 = ( w1225 & w3313 ) | ( w1225 & ~w3319 ) | ( w3313 & ~w3319 ) ;
  assign w3321 = w1225 & w3320 ;
  assign w3322 = w3083 | w3088 ;
  assign w3323 = w3227 & ~w3322 ;
  assign w3324 = w3086 ^ w3323 ;
  assign w3325 = ( ~w1225 & w3313 ) | ( ~w1225 & w3319 ) | ( w3313 & w3319 ) ;
  assign w3326 = ~w3313 & w3325 ;
  assign w3327 = w3324 | w3326 ;
  assign w3328 = ( w1091 & w3321 ) | ( w1091 & ~w3327 ) | ( w3321 & ~w3327 ) ;
  assign w3329 = w1091 & w3328 ;
  assign w3330 = w3091 | w3096 ;
  assign w3331 = w3227 & ~w3330 ;
  assign w3332 = w3094 ^ w3331 ;
  assign w3333 = ( ~w1091 & w3321 ) | ( ~w1091 & w3327 ) | ( w3321 & w3327 ) ;
  assign w3334 = ~w3321 & w3333 ;
  assign w3335 = w3332 | w3334 ;
  assign w3336 = ( w965 & w3329 ) | ( w965 & ~w3335 ) | ( w3329 & ~w3335 ) ;
  assign w3337 = w965 & w3336 ;
  assign w3338 = w3099 | w3104 ;
  assign w3339 = w3227 & ~w3338 ;
  assign w3340 = w3102 ^ w3339 ;
  assign w3341 = ( ~w965 & w3329 ) | ( ~w965 & w3335 ) | ( w3329 & w3335 ) ;
  assign w3342 = ~w3329 & w3341 ;
  assign w3343 = w3340 | w3342 ;
  assign w3344 = ( w847 & w3337 ) | ( w847 & ~w3343 ) | ( w3337 & ~w3343 ) ;
  assign w3345 = w847 & w3344 ;
  assign w3346 = w3107 | w3112 ;
  assign w3347 = w3227 & ~w3346 ;
  assign w3348 = w3110 ^ w3347 ;
  assign w3349 = ( ~w847 & w3337 ) | ( ~w847 & w3343 ) | ( w3337 & w3343 ) ;
  assign w3350 = ~w3337 & w3349 ;
  assign w3351 = w3348 | w3350 ;
  assign w3352 = ( w737 & w3345 ) | ( w737 & ~w3351 ) | ( w3345 & ~w3351 ) ;
  assign w3353 = w737 & w3352 ;
  assign w3354 = w3115 | w3120 ;
  assign w3355 = w3227 & ~w3354 ;
  assign w3356 = w3118 ^ w3355 ;
  assign w3357 = ( ~w737 & w3345 ) | ( ~w737 & w3351 ) | ( w3345 & w3351 ) ;
  assign w3358 = ~w3345 & w3357 ;
  assign w3359 = w3356 | w3358 ;
  assign w3360 = ( w635 & w3353 ) | ( w635 & ~w3359 ) | ( w3353 & ~w3359 ) ;
  assign w3361 = w635 & w3360 ;
  assign w3362 = w3123 | w3128 ;
  assign w3363 = w3227 & ~w3362 ;
  assign w3364 = w3126 ^ w3363 ;
  assign w3365 = ( ~w635 & w3353 ) | ( ~w635 & w3359 ) | ( w3353 & w3359 ) ;
  assign w3366 = ~w3353 & w3365 ;
  assign w3367 = w3364 | w3366 ;
  assign w3368 = ( w541 & w3361 ) | ( w541 & ~w3367 ) | ( w3361 & ~w3367 ) ;
  assign w3369 = w541 & w3368 ;
  assign w3370 = w3131 | w3136 ;
  assign w3371 = w3227 & ~w3370 ;
  assign w3372 = w3134 ^ w3371 ;
  assign w3373 = ( ~w541 & w3361 ) | ( ~w541 & w3367 ) | ( w3361 & w3367 ) ;
  assign w3374 = ~w3361 & w3373 ;
  assign w3375 = w3372 | w3374 ;
  assign w3376 = ( w455 & w3369 ) | ( w455 & ~w3375 ) | ( w3369 & ~w3375 ) ;
  assign w3377 = w455 & w3376 ;
  assign w3378 = w3139 | w3144 ;
  assign w3379 = w3227 & ~w3378 ;
  assign w3380 = w3142 ^ w3379 ;
  assign w3381 = ( ~w455 & w3369 ) | ( ~w455 & w3375 ) | ( w3369 & w3375 ) ;
  assign w3382 = ~w3369 & w3381 ;
  assign w3383 = w3380 | w3382 ;
  assign w3384 = ( w377 & w3377 ) | ( w377 & ~w3383 ) | ( w3377 & ~w3383 ) ;
  assign w3385 = w377 & w3384 ;
  assign w3386 = w3147 | w3152 ;
  assign w3387 = w3227 & ~w3386 ;
  assign w3388 = w3150 ^ w3387 ;
  assign w3389 = ( ~w377 & w3377 ) | ( ~w377 & w3383 ) | ( w3377 & w3383 ) ;
  assign w3390 = ~w3377 & w3389 ;
  assign w3391 = w3388 | w3390 ;
  assign w3392 = ( w307 & w3385 ) | ( w307 & ~w3391 ) | ( w3385 & ~w3391 ) ;
  assign w3393 = w307 & w3392 ;
  assign w3394 = w3155 | w3160 ;
  assign w3395 = w3227 & ~w3394 ;
  assign w3396 = w3158 ^ w3395 ;
  assign w3397 = ( ~w307 & w3385 ) | ( ~w307 & w3391 ) | ( w3385 & w3391 ) ;
  assign w3398 = ~w3385 & w3397 ;
  assign w3399 = w3396 | w3398 ;
  assign w3400 = ( w246 & w3393 ) | ( w246 & ~w3399 ) | ( w3393 & ~w3399 ) ;
  assign w3401 = w246 & w3400 ;
  assign w3402 = ( ~w246 & w3393 ) | ( ~w246 & w3399 ) | ( w3393 & w3399 ) ;
  assign w3403 = ~w3393 & w3402 ;
  assign w3404 = w3163 | w3165 ;
  assign w3405 = w3227 & ~w3404 ;
  assign w3406 = w3168 ^ w3405 ;
  assign w3407 = w3403 | w3406 ;
  assign w3408 = ( w185 & w3401 ) | ( w185 & ~w3407 ) | ( w3401 & ~w3407 ) ;
  assign w3409 = w185 & w3408 ;
  assign w3410 = w3171 | w3176 ;
  assign w3411 = w3227 & ~w3410 ;
  assign w3412 = w3174 ^ w3411 ;
  assign w3413 = ( ~w185 & w3401 ) | ( ~w185 & w3407 ) | ( w3401 & w3407 ) ;
  assign w3414 = ~w3401 & w3413 ;
  assign w3415 = w3412 | w3414 ;
  assign w3416 = ( w145 & w3409 ) | ( w145 & ~w3415 ) | ( w3409 & ~w3415 ) ;
  assign w3417 = w145 & w3416 ;
  assign w3418 = w3179 | w3184 ;
  assign w3419 = w3227 & ~w3418 ;
  assign w3420 = w3182 ^ w3419 ;
  assign w3421 = ( ~w145 & w3409 ) | ( ~w145 & w3415 ) | ( w3409 & w3415 ) ;
  assign w3422 = ~w3409 & w3421 ;
  assign w3423 = w3420 | w3422 ;
  assign w3424 = ( w132 & w3417 ) | ( w132 & ~w3423 ) | ( w3417 & ~w3423 ) ;
  assign w3425 = w132 & w3424 ;
  assign w3426 = w3187 | w3192 ;
  assign w3427 = w3227 & ~w3426 ;
  assign w3428 = w3190 ^ w3427 ;
  assign w3429 = ( ~w132 & w3417 ) | ( ~w132 & w3423 ) | ( w3417 & w3423 ) ;
  assign w3430 = ~w3417 & w3429 ;
  assign w3431 = w3428 | w3430 ;
  assign w3432 = ~w3425 & w3431 ;
  assign w3433 = w3195 | w3200 ;
  assign w3434 = w3227 & ~w3433 ;
  assign w3435 = w3198 ^ w3434 ;
  assign w3436 = ( ~w3213 & w3432 ) | ( ~w3213 & w3435 ) | ( w3432 & w3435 ) ;
  assign w3437 = w3202 & ~w3436 ;
  assign w3438 = ~w3205 & w3227 ;
  assign w3439 = ( w3436 & ~w3437 ) | ( w3436 & w3438 ) | ( ~w3437 & w3438 ) ;
  assign w3440 = w3213 | w3439 ;
  assign w3441 = ~w129 & w3440 ;
  assign w3442 = ( w3425 & w3431 ) | ( w3425 & w3435 ) | ( w3431 & w3435 ) ;
  assign w3443 = ~w3425 & w3442 ;
  assign w3444 = ( w129 & w3202 ) | ( w129 & w3205 ) | ( w3202 & w3205 ) ;
  assign w3445 = ( w3205 & ~w3227 ) | ( w3205 & w3444 ) | ( ~w3227 & w3444 ) ;
  assign w3446 = w3202 & w3445 ;
  assign w3447 = w3444 ^ w3446 ;
  assign w3448 = ( w2973 & w2978 ) | ( w2973 & w3005 ) | ( w2978 & w3005 ) ;
  assign w3449 = w3005 & ~w3448 ;
  assign w3450 = w2976 ^ w3449 ;
  assign w3451 = ( ~w3217 & w3224 ) | ( ~w3217 & w3450 ) | ( w3224 & w3450 ) ;
  assign w3452 = ~w3224 & w3451 ;
  assign w3453 = ( ~w3211 & w3213 ) | ( ~w3211 & w3452 ) | ( w3213 & w3452 ) ;
  assign w3454 = ~w3213 & w3453 ;
  assign w3455 = w3443 | w3454 ;
  assign w3456 = ( w3441 & ~w3443 ) | ( w3441 & w3447 ) | ( ~w3443 & w3447 ) ;
  assign w3457 = w3455 | w3456 ;
  assign w3458 = ( ~\pi073 & \pi074 ) | ( ~\pi073 & w3227 ) | ( \pi074 & w3227 ) ;
  assign w3459 = ( ~\pi072 & \pi074 ) | ( ~\pi072 & w3458 ) | ( \pi074 & w3458 ) ;
  assign w3460 = ( ~\pi074 & w3227 ) | ( ~\pi074 & w3457 ) | ( w3227 & w3457 ) ;
  assign w3461 = w3459 & w3460 ;
  assign w3462 = ( w3213 & w3217 ) | ( w3213 & ~w3224 ) | ( w3217 & ~w3224 ) ;
  assign w3463 = \pi073 & ~w3462 ;
  assign w3464 = \pi072 | \pi074 ;
  assign w3465 = ( ~w3462 & w3463 ) | ( ~w3462 & w3464 ) | ( w3463 & w3464 ) ;
  assign w3466 = ~w3224 & w3465 ;
  assign w3467 = ~w3211 & w3466 ;
  assign w3468 = ( \pi074 & w3457 ) | ( \pi074 & ~w3466 ) | ( w3457 & ~w3466 ) ;
  assign w3469 = w3467 & ~w3468 ;
  assign w3470 = ~\pi074 & w3457 ;
  assign w3471 = \pi075 ^ w3470 ;
  assign w3472 = w3469 | w3471 ;
  assign w3473 = ( w3005 & w3461 ) | ( w3005 & ~w3472 ) | ( w3461 & ~w3472 ) ;
  assign w3474 = w3005 & w3473 ;
  assign w3475 = ( ~w3005 & w3461 ) | ( ~w3005 & w3472 ) | ( w3461 & w3472 ) ;
  assign w3476 = ~w3461 & w3475 ;
  assign w3477 = w3227 & ~w3454 ;
  assign w3478 = ~w3443 & w3477 ;
  assign w3479 = ~w3456 & w3478 ;
  assign w3480 = \pi075 & w3457 ;
  assign w3481 = ( \pi074 & w3457 ) | ( \pi074 & ~w3480 ) | ( w3457 & ~w3480 ) ;
  assign w3482 = ( ~\pi074 & w3479 ) | ( ~\pi074 & w3481 ) | ( w3479 & w3481 ) ;
  assign w3483 = \pi076 ^ w3482 ;
  assign w3484 = w3476 | w3483 ;
  assign w3485 = ( w2791 & w3474 ) | ( w2791 & ~w3484 ) | ( w3474 & ~w3484 ) ;
  assign w3486 = w2791 & w3485 ;
  assign w3487 = ( w3231 & ~w3239 ) | ( w3231 & w3457 ) | ( ~w3239 & w3457 ) ;
  assign w3488 = ~w3231 & w3487 ;
  assign w3489 = \pi077 ^ w3488 ;
  assign w3490 = w3240 ^ w3489 ;
  assign w3491 = ( ~w2791 & w3474 ) | ( ~w2791 & w3484 ) | ( w3474 & w3484 ) ;
  assign w3492 = ~w3474 & w3491 ;
  assign w3493 = w3490 | w3492 ;
  assign w3494 = ( w2585 & w3486 ) | ( w2585 & ~w3493 ) | ( w3486 & ~w3493 ) ;
  assign w3495 = w2585 & w3494 ;
  assign w3496 = w3244 | w3246 ;
  assign w3497 = w3457 & ~w3496 ;
  assign w3498 = w3253 ^ w3497 ;
  assign w3499 = ( ~w2585 & w3486 ) | ( ~w2585 & w3493 ) | ( w3486 & w3493 ) ;
  assign w3500 = ~w3486 & w3499 ;
  assign w3501 = w3498 | w3500 ;
  assign w3502 = ( w2387 & w3495 ) | ( w2387 & ~w3501 ) | ( w3495 & ~w3501 ) ;
  assign w3503 = w2387 & w3502 ;
  assign w3504 = w3256 | w3262 ;
  assign w3505 = w3457 & ~w3504 ;
  assign w3506 = w3260 ^ w3505 ;
  assign w3507 = ( ~w2387 & w3495 ) | ( ~w2387 & w3501 ) | ( w3495 & w3501 ) ;
  assign w3508 = ~w3495 & w3507 ;
  assign w3509 = w3506 | w3508 ;
  assign w3510 = ( w2197 & w3503 ) | ( w2197 & ~w3509 ) | ( w3503 & ~w3509 ) ;
  assign w3511 = w2197 & w3510 ;
  assign w3512 = w3265 | w3270 ;
  assign w3513 = w3457 & ~w3512 ;
  assign w3514 = w3268 ^ w3513 ;
  assign w3515 = ( ~w2197 & w3503 ) | ( ~w2197 & w3509 ) | ( w3503 & w3509 ) ;
  assign w3516 = ~w3503 & w3515 ;
  assign w3517 = w3514 | w3516 ;
  assign w3518 = ( w2015 & w3511 ) | ( w2015 & ~w3517 ) | ( w3511 & ~w3517 ) ;
  assign w3519 = w2015 & w3518 ;
  assign w3520 = w3273 | w3278 ;
  assign w3521 = w3457 & ~w3520 ;
  assign w3522 = w3276 ^ w3521 ;
  assign w3523 = ( ~w2015 & w3511 ) | ( ~w2015 & w3517 ) | ( w3511 & w3517 ) ;
  assign w3524 = ~w3511 & w3523 ;
  assign w3525 = w3522 | w3524 ;
  assign w3526 = ( w1841 & w3519 ) | ( w1841 & ~w3525 ) | ( w3519 & ~w3525 ) ;
  assign w3527 = w1841 & w3526 ;
  assign w3528 = w3281 | w3286 ;
  assign w3529 = w3457 & ~w3528 ;
  assign w3530 = w3284 ^ w3529 ;
  assign w3531 = ( ~w1841 & w3519 ) | ( ~w1841 & w3525 ) | ( w3519 & w3525 ) ;
  assign w3532 = ~w3519 & w3531 ;
  assign w3533 = w3530 | w3532 ;
  assign w3534 = ( w1675 & w3527 ) | ( w1675 & ~w3533 ) | ( w3527 & ~w3533 ) ;
  assign w3535 = w1675 & w3534 ;
  assign w3536 = w3289 | w3294 ;
  assign w3537 = w3457 & ~w3536 ;
  assign w3538 = w3292 ^ w3537 ;
  assign w3539 = ( ~w1675 & w3527 ) | ( ~w1675 & w3533 ) | ( w3527 & w3533 ) ;
  assign w3540 = ~w3527 & w3539 ;
  assign w3541 = w3538 | w3540 ;
  assign w3542 = ( w1517 & w3535 ) | ( w1517 & ~w3541 ) | ( w3535 & ~w3541 ) ;
  assign w3543 = w1517 & w3542 ;
  assign w3544 = w3297 | w3302 ;
  assign w3545 = w3457 & ~w3544 ;
  assign w3546 = w3300 ^ w3545 ;
  assign w3547 = ( ~w1517 & w3535 ) | ( ~w1517 & w3541 ) | ( w3535 & w3541 ) ;
  assign w3548 = ~w3535 & w3547 ;
  assign w3549 = w3546 | w3548 ;
  assign w3550 = ( w1367 & w3543 ) | ( w1367 & ~w3549 ) | ( w3543 & ~w3549 ) ;
  assign w3551 = w1367 & w3550 ;
  assign w3552 = w3305 | w3310 ;
  assign w3553 = w3457 & ~w3552 ;
  assign w3554 = w3308 ^ w3553 ;
  assign w3555 = ( ~w1367 & w3543 ) | ( ~w1367 & w3549 ) | ( w3543 & w3549 ) ;
  assign w3556 = ~w3543 & w3555 ;
  assign w3557 = w3554 | w3556 ;
  assign w3558 = ( w1225 & w3551 ) | ( w1225 & ~w3557 ) | ( w3551 & ~w3557 ) ;
  assign w3559 = w1225 & w3558 ;
  assign w3560 = w3313 | w3318 ;
  assign w3561 = w3457 & ~w3560 ;
  assign w3562 = w3316 ^ w3561 ;
  assign w3563 = ( ~w1225 & w3551 ) | ( ~w1225 & w3557 ) | ( w3551 & w3557 ) ;
  assign w3564 = ~w3551 & w3563 ;
  assign w3565 = w3562 | w3564 ;
  assign w3566 = ( w1091 & w3559 ) | ( w1091 & ~w3565 ) | ( w3559 & ~w3565 ) ;
  assign w3567 = w1091 & w3566 ;
  assign w3568 = w3321 | w3326 ;
  assign w3569 = w3457 & ~w3568 ;
  assign w3570 = w3324 ^ w3569 ;
  assign w3571 = ( ~w1091 & w3559 ) | ( ~w1091 & w3565 ) | ( w3559 & w3565 ) ;
  assign w3572 = ~w3559 & w3571 ;
  assign w3573 = w3570 | w3572 ;
  assign w3574 = ( w965 & w3567 ) | ( w965 & ~w3573 ) | ( w3567 & ~w3573 ) ;
  assign w3575 = w965 & w3574 ;
  assign w3576 = w3329 | w3334 ;
  assign w3577 = w3457 & ~w3576 ;
  assign w3578 = w3332 ^ w3577 ;
  assign w3579 = ( ~w965 & w3567 ) | ( ~w965 & w3573 ) | ( w3567 & w3573 ) ;
  assign w3580 = ~w3567 & w3579 ;
  assign w3581 = w3578 | w3580 ;
  assign w3582 = ( w847 & w3575 ) | ( w847 & ~w3581 ) | ( w3575 & ~w3581 ) ;
  assign w3583 = w847 & w3582 ;
  assign w3584 = w3337 | w3342 ;
  assign w3585 = w3457 & ~w3584 ;
  assign w3586 = w3340 ^ w3585 ;
  assign w3587 = ( ~w847 & w3575 ) | ( ~w847 & w3581 ) | ( w3575 & w3581 ) ;
  assign w3588 = ~w3575 & w3587 ;
  assign w3589 = w3586 | w3588 ;
  assign w3590 = ( w737 & w3583 ) | ( w737 & ~w3589 ) | ( w3583 & ~w3589 ) ;
  assign w3591 = w737 & w3590 ;
  assign w3592 = w3345 | w3350 ;
  assign w3593 = w3457 & ~w3592 ;
  assign w3594 = w3348 ^ w3593 ;
  assign w3595 = ( ~w737 & w3583 ) | ( ~w737 & w3589 ) | ( w3583 & w3589 ) ;
  assign w3596 = ~w3583 & w3595 ;
  assign w3597 = w3594 | w3596 ;
  assign w3598 = ( w635 & w3591 ) | ( w635 & ~w3597 ) | ( w3591 & ~w3597 ) ;
  assign w3599 = w635 & w3598 ;
  assign w3600 = w3353 | w3358 ;
  assign w3601 = w3457 & ~w3600 ;
  assign w3602 = w3356 ^ w3601 ;
  assign w3603 = ( ~w635 & w3591 ) | ( ~w635 & w3597 ) | ( w3591 & w3597 ) ;
  assign w3604 = ~w3591 & w3603 ;
  assign w3605 = w3602 | w3604 ;
  assign w3606 = ( w541 & w3599 ) | ( w541 & ~w3605 ) | ( w3599 & ~w3605 ) ;
  assign w3607 = w541 & w3606 ;
  assign w3608 = w3361 | w3366 ;
  assign w3609 = w3457 & ~w3608 ;
  assign w3610 = w3364 ^ w3609 ;
  assign w3611 = ( ~w541 & w3599 ) | ( ~w541 & w3605 ) | ( w3599 & w3605 ) ;
  assign w3612 = ~w3599 & w3611 ;
  assign w3613 = w3610 | w3612 ;
  assign w3614 = ( w455 & w3607 ) | ( w455 & ~w3613 ) | ( w3607 & ~w3613 ) ;
  assign w3615 = w455 & w3614 ;
  assign w3616 = w3369 | w3374 ;
  assign w3617 = w3457 & ~w3616 ;
  assign w3618 = w3372 ^ w3617 ;
  assign w3619 = ( ~w455 & w3607 ) | ( ~w455 & w3613 ) | ( w3607 & w3613 ) ;
  assign w3620 = ~w3607 & w3619 ;
  assign w3621 = w3618 | w3620 ;
  assign w3622 = ( w377 & w3615 ) | ( w377 & ~w3621 ) | ( w3615 & ~w3621 ) ;
  assign w3623 = w377 & w3622 ;
  assign w3624 = w3377 | w3382 ;
  assign w3625 = w3457 & ~w3624 ;
  assign w3626 = w3380 ^ w3625 ;
  assign w3627 = ( ~w377 & w3615 ) | ( ~w377 & w3621 ) | ( w3615 & w3621 ) ;
  assign w3628 = ~w3615 & w3627 ;
  assign w3629 = w3626 | w3628 ;
  assign w3630 = ( w307 & w3623 ) | ( w307 & ~w3629 ) | ( w3623 & ~w3629 ) ;
  assign w3631 = w307 & w3630 ;
  assign w3632 = w3385 | w3390 ;
  assign w3633 = w3457 & ~w3632 ;
  assign w3634 = w3388 ^ w3633 ;
  assign w3635 = ( ~w307 & w3623 ) | ( ~w307 & w3629 ) | ( w3623 & w3629 ) ;
  assign w3636 = ~w3623 & w3635 ;
  assign w3637 = w3634 | w3636 ;
  assign w3638 = ( w246 & w3631 ) | ( w246 & ~w3637 ) | ( w3631 & ~w3637 ) ;
  assign w3639 = w246 & w3638 ;
  assign w3640 = w3393 | w3398 ;
  assign w3641 = w3457 & ~w3640 ;
  assign w3642 = w3396 ^ w3641 ;
  assign w3643 = ( ~w246 & w3631 ) | ( ~w246 & w3637 ) | ( w3631 & w3637 ) ;
  assign w3644 = ~w3631 & w3643 ;
  assign w3645 = w3642 | w3644 ;
  assign w3646 = ( w185 & w3639 ) | ( w185 & ~w3645 ) | ( w3639 & ~w3645 ) ;
  assign w3647 = w185 & w3646 ;
  assign w3648 = ( ~w185 & w3639 ) | ( ~w185 & w3645 ) | ( w3639 & w3645 ) ;
  assign w3649 = ~w3639 & w3648 ;
  assign w3650 = w3401 | w3403 ;
  assign w3651 = w3457 & ~w3650 ;
  assign w3652 = w3406 ^ w3651 ;
  assign w3653 = w3649 | w3652 ;
  assign w3654 = ( w145 & w3647 ) | ( w145 & ~w3653 ) | ( w3647 & ~w3653 ) ;
  assign w3655 = w145 & w3654 ;
  assign w3656 = w3409 | w3414 ;
  assign w3657 = w3457 & ~w3656 ;
  assign w3658 = w3412 ^ w3657 ;
  assign w3659 = ( ~w145 & w3647 ) | ( ~w145 & w3653 ) | ( w3647 & w3653 ) ;
  assign w3660 = ~w3647 & w3659 ;
  assign w3661 = w3658 | w3660 ;
  assign w3662 = ( w132 & w3655 ) | ( w132 & ~w3661 ) | ( w3655 & ~w3661 ) ;
  assign w3663 = w132 & w3662 ;
  assign w3664 = w3417 | w3422 ;
  assign w3665 = w3457 & ~w3664 ;
  assign w3666 = w3420 ^ w3665 ;
  assign w3667 = ( ~w132 & w3655 ) | ( ~w132 & w3661 ) | ( w3655 & w3661 ) ;
  assign w3668 = ~w3655 & w3667 ;
  assign w3669 = w3666 | w3668 ;
  assign w3670 = ~w3663 & w3669 ;
  assign w3671 = w3425 | w3430 ;
  assign w3672 = w3457 & ~w3671 ;
  assign w3673 = w3428 ^ w3672 ;
  assign w3674 = ( ~w3443 & w3670 ) | ( ~w3443 & w3673 ) | ( w3670 & w3673 ) ;
  assign w3675 = w3432 & ~w3674 ;
  assign w3676 = ~w3435 & w3457 ;
  assign w3677 = ( w3674 & ~w3675 ) | ( w3674 & w3676 ) | ( ~w3675 & w3676 ) ;
  assign w3678 = w3443 | w3677 ;
  assign w3679 = ~w129 & w3678 ;
  assign w3680 = ( w3663 & w3669 ) | ( w3663 & w3673 ) | ( w3669 & w3673 ) ;
  assign w3681 = ~w3663 & w3680 ;
  assign w3682 = ( w129 & w3432 ) | ( w129 & w3435 ) | ( w3432 & w3435 ) ;
  assign w3683 = ( w3435 & ~w3457 ) | ( w3435 & w3682 ) | ( ~w3457 & w3682 ) ;
  assign w3684 = w3432 & w3683 ;
  assign w3685 = w3682 ^ w3684 ;
  assign w3686 = ( w3195 & w3200 ) | ( w3195 & w3227 ) | ( w3200 & w3227 ) ;
  assign w3687 = w3227 & ~w3686 ;
  assign w3688 = w3198 ^ w3687 ;
  assign w3689 = ( ~w3447 & w3454 ) | ( ~w3447 & w3688 ) | ( w3454 & w3688 ) ;
  assign w3690 = ~w3454 & w3689 ;
  assign w3691 = ( ~w3441 & w3443 ) | ( ~w3441 & w3690 ) | ( w3443 & w3690 ) ;
  assign w3692 = ~w3443 & w3691 ;
  assign w3693 = w3681 | w3692 ;
  assign w3694 = ( w3679 & ~w3681 ) | ( w3679 & w3685 ) | ( ~w3681 & w3685 ) ;
  assign w3695 = w3693 | w3694 ;
  assign w3696 = ( ~\pi071 & \pi072 ) | ( ~\pi071 & w3457 ) | ( \pi072 & w3457 ) ;
  assign w3697 = ( ~\pi070 & \pi072 ) | ( ~\pi070 & w3696 ) | ( \pi072 & w3696 ) ;
  assign w3698 = ( ~\pi072 & w3457 ) | ( ~\pi072 & w3695 ) | ( w3457 & w3695 ) ;
  assign w3699 = w3697 & w3698 ;
  assign w3700 = ( w3443 & w3447 ) | ( w3443 & ~w3454 ) | ( w3447 & ~w3454 ) ;
  assign w3701 = \pi071 & ~w3700 ;
  assign w3702 = \pi070 | \pi072 ;
  assign w3703 = ( ~w3700 & w3701 ) | ( ~w3700 & w3702 ) | ( w3701 & w3702 ) ;
  assign w3704 = ~w3454 & w3703 ;
  assign w3705 = ~w3441 & w3704 ;
  assign w3706 = ( \pi072 & w3695 ) | ( \pi072 & ~w3704 ) | ( w3695 & ~w3704 ) ;
  assign w3707 = w3705 & ~w3706 ;
  assign w3708 = ~\pi072 & w3695 ;
  assign w3709 = \pi073 ^ w3708 ;
  assign w3710 = w3707 | w3709 ;
  assign w3711 = ( w3227 & w3699 ) | ( w3227 & ~w3710 ) | ( w3699 & ~w3710 ) ;
  assign w3712 = w3227 & w3711 ;
  assign w3713 = ( ~w3227 & w3699 ) | ( ~w3227 & w3710 ) | ( w3699 & w3710 ) ;
  assign w3714 = ~w3699 & w3713 ;
  assign w3715 = w3457 & ~w3692 ;
  assign w3716 = ~w3681 & w3715 ;
  assign w3717 = ~w3694 & w3716 ;
  assign w3718 = \pi073 & w3695 ;
  assign w3719 = ( \pi072 & w3695 ) | ( \pi072 & ~w3718 ) | ( w3695 & ~w3718 ) ;
  assign w3720 = ( ~\pi072 & w3717 ) | ( ~\pi072 & w3719 ) | ( w3717 & w3719 ) ;
  assign w3721 = \pi074 ^ w3720 ;
  assign w3722 = w3714 | w3721 ;
  assign w3723 = ( w3005 & w3712 ) | ( w3005 & ~w3722 ) | ( w3712 & ~w3722 ) ;
  assign w3724 = w3005 & w3723 ;
  assign w3725 = ( w3461 & ~w3469 ) | ( w3461 & w3695 ) | ( ~w3469 & w3695 ) ;
  assign w3726 = ~w3461 & w3725 ;
  assign w3727 = \pi075 ^ w3726 ;
  assign w3728 = w3470 ^ w3727 ;
  assign w3729 = ( ~w3005 & w3712 ) | ( ~w3005 & w3722 ) | ( w3712 & w3722 ) ;
  assign w3730 = ~w3712 & w3729 ;
  assign w3731 = w3728 | w3730 ;
  assign w3732 = ( w2791 & w3724 ) | ( w2791 & ~w3731 ) | ( w3724 & ~w3731 ) ;
  assign w3733 = w2791 & w3732 ;
  assign w3734 = w3474 | w3476 ;
  assign w3735 = w3695 & ~w3734 ;
  assign w3736 = w3483 ^ w3735 ;
  assign w3737 = ( ~w2791 & w3724 ) | ( ~w2791 & w3731 ) | ( w3724 & w3731 ) ;
  assign w3738 = ~w3724 & w3737 ;
  assign w3739 = w3736 | w3738 ;
  assign w3740 = ( w2585 & w3733 ) | ( w2585 & ~w3739 ) | ( w3733 & ~w3739 ) ;
  assign w3741 = w2585 & w3740 ;
  assign w3742 = w3486 | w3492 ;
  assign w3743 = w3695 & ~w3742 ;
  assign w3744 = w3490 ^ w3743 ;
  assign w3745 = ( ~w2585 & w3733 ) | ( ~w2585 & w3739 ) | ( w3733 & w3739 ) ;
  assign w3746 = ~w3733 & w3745 ;
  assign w3747 = w3744 | w3746 ;
  assign w3748 = ( w2387 & w3741 ) | ( w2387 & ~w3747 ) | ( w3741 & ~w3747 ) ;
  assign w3749 = w2387 & w3748 ;
  assign w3750 = w3495 | w3500 ;
  assign w3751 = w3695 & ~w3750 ;
  assign w3752 = w3498 ^ w3751 ;
  assign w3753 = ( ~w2387 & w3741 ) | ( ~w2387 & w3747 ) | ( w3741 & w3747 ) ;
  assign w3754 = ~w3741 & w3753 ;
  assign w3755 = w3752 | w3754 ;
  assign w3756 = ( w2197 & w3749 ) | ( w2197 & ~w3755 ) | ( w3749 & ~w3755 ) ;
  assign w3757 = w2197 & w3756 ;
  assign w3758 = w3503 | w3508 ;
  assign w3759 = w3695 & ~w3758 ;
  assign w3760 = w3506 ^ w3759 ;
  assign w3761 = ( ~w2197 & w3749 ) | ( ~w2197 & w3755 ) | ( w3749 & w3755 ) ;
  assign w3762 = ~w3749 & w3761 ;
  assign w3763 = w3760 | w3762 ;
  assign w3764 = ( w2015 & w3757 ) | ( w2015 & ~w3763 ) | ( w3757 & ~w3763 ) ;
  assign w3765 = w2015 & w3764 ;
  assign w3766 = w3511 | w3516 ;
  assign w3767 = w3695 & ~w3766 ;
  assign w3768 = w3514 ^ w3767 ;
  assign w3769 = ( ~w2015 & w3757 ) | ( ~w2015 & w3763 ) | ( w3757 & w3763 ) ;
  assign w3770 = ~w3757 & w3769 ;
  assign w3771 = w3768 | w3770 ;
  assign w3772 = ( w1841 & w3765 ) | ( w1841 & ~w3771 ) | ( w3765 & ~w3771 ) ;
  assign w3773 = w1841 & w3772 ;
  assign w3774 = w3519 | w3524 ;
  assign w3775 = w3695 & ~w3774 ;
  assign w3776 = w3522 ^ w3775 ;
  assign w3777 = ( ~w1841 & w3765 ) | ( ~w1841 & w3771 ) | ( w3765 & w3771 ) ;
  assign w3778 = ~w3765 & w3777 ;
  assign w3779 = w3776 | w3778 ;
  assign w3780 = ( w1675 & w3773 ) | ( w1675 & ~w3779 ) | ( w3773 & ~w3779 ) ;
  assign w3781 = w1675 & w3780 ;
  assign w3782 = w3527 | w3532 ;
  assign w3783 = w3695 & ~w3782 ;
  assign w3784 = w3530 ^ w3783 ;
  assign w3785 = ( ~w1675 & w3773 ) | ( ~w1675 & w3779 ) | ( w3773 & w3779 ) ;
  assign w3786 = ~w3773 & w3785 ;
  assign w3787 = w3784 | w3786 ;
  assign w3788 = ( w1517 & w3781 ) | ( w1517 & ~w3787 ) | ( w3781 & ~w3787 ) ;
  assign w3789 = w1517 & w3788 ;
  assign w3790 = w3535 | w3540 ;
  assign w3791 = w3695 & ~w3790 ;
  assign w3792 = w3538 ^ w3791 ;
  assign w3793 = ( ~w1517 & w3781 ) | ( ~w1517 & w3787 ) | ( w3781 & w3787 ) ;
  assign w3794 = ~w3781 & w3793 ;
  assign w3795 = w3792 | w3794 ;
  assign w3796 = ( w1367 & w3789 ) | ( w1367 & ~w3795 ) | ( w3789 & ~w3795 ) ;
  assign w3797 = w1367 & w3796 ;
  assign w3798 = w3543 | w3548 ;
  assign w3799 = w3695 & ~w3798 ;
  assign w3800 = w3546 ^ w3799 ;
  assign w3801 = ( ~w1367 & w3789 ) | ( ~w1367 & w3795 ) | ( w3789 & w3795 ) ;
  assign w3802 = ~w3789 & w3801 ;
  assign w3803 = w3800 | w3802 ;
  assign w3804 = ( w1225 & w3797 ) | ( w1225 & ~w3803 ) | ( w3797 & ~w3803 ) ;
  assign w3805 = w1225 & w3804 ;
  assign w3806 = w3551 | w3556 ;
  assign w3807 = w3695 & ~w3806 ;
  assign w3808 = w3554 ^ w3807 ;
  assign w3809 = ( ~w1225 & w3797 ) | ( ~w1225 & w3803 ) | ( w3797 & w3803 ) ;
  assign w3810 = ~w3797 & w3809 ;
  assign w3811 = w3808 | w3810 ;
  assign w3812 = ( w1091 & w3805 ) | ( w1091 & ~w3811 ) | ( w3805 & ~w3811 ) ;
  assign w3813 = w1091 & w3812 ;
  assign w3814 = w3559 | w3564 ;
  assign w3815 = w3695 & ~w3814 ;
  assign w3816 = w3562 ^ w3815 ;
  assign w3817 = ( ~w1091 & w3805 ) | ( ~w1091 & w3811 ) | ( w3805 & w3811 ) ;
  assign w3818 = ~w3805 & w3817 ;
  assign w3819 = w3816 | w3818 ;
  assign w3820 = ( w965 & w3813 ) | ( w965 & ~w3819 ) | ( w3813 & ~w3819 ) ;
  assign w3821 = w965 & w3820 ;
  assign w3822 = w3567 | w3572 ;
  assign w3823 = w3695 & ~w3822 ;
  assign w3824 = w3570 ^ w3823 ;
  assign w3825 = ( ~w965 & w3813 ) | ( ~w965 & w3819 ) | ( w3813 & w3819 ) ;
  assign w3826 = ~w3813 & w3825 ;
  assign w3827 = w3824 | w3826 ;
  assign w3828 = ( w847 & w3821 ) | ( w847 & ~w3827 ) | ( w3821 & ~w3827 ) ;
  assign w3829 = w847 & w3828 ;
  assign w3830 = w3575 | w3580 ;
  assign w3831 = w3695 & ~w3830 ;
  assign w3832 = w3578 ^ w3831 ;
  assign w3833 = ( ~w847 & w3821 ) | ( ~w847 & w3827 ) | ( w3821 & w3827 ) ;
  assign w3834 = ~w3821 & w3833 ;
  assign w3835 = w3832 | w3834 ;
  assign w3836 = ( w737 & w3829 ) | ( w737 & ~w3835 ) | ( w3829 & ~w3835 ) ;
  assign w3837 = w737 & w3836 ;
  assign w3838 = w3583 | w3588 ;
  assign w3839 = w3695 & ~w3838 ;
  assign w3840 = w3586 ^ w3839 ;
  assign w3841 = ( ~w737 & w3829 ) | ( ~w737 & w3835 ) | ( w3829 & w3835 ) ;
  assign w3842 = ~w3829 & w3841 ;
  assign w3843 = w3840 | w3842 ;
  assign w3844 = ( w635 & w3837 ) | ( w635 & ~w3843 ) | ( w3837 & ~w3843 ) ;
  assign w3845 = w635 & w3844 ;
  assign w3846 = w3591 | w3596 ;
  assign w3847 = w3695 & ~w3846 ;
  assign w3848 = w3594 ^ w3847 ;
  assign w3849 = ( ~w635 & w3837 ) | ( ~w635 & w3843 ) | ( w3837 & w3843 ) ;
  assign w3850 = ~w3837 & w3849 ;
  assign w3851 = w3848 | w3850 ;
  assign w3852 = ( w541 & w3845 ) | ( w541 & ~w3851 ) | ( w3845 & ~w3851 ) ;
  assign w3853 = w541 & w3852 ;
  assign w3854 = w3599 | w3604 ;
  assign w3855 = w3695 & ~w3854 ;
  assign w3856 = w3602 ^ w3855 ;
  assign w3857 = ( ~w541 & w3845 ) | ( ~w541 & w3851 ) | ( w3845 & w3851 ) ;
  assign w3858 = ~w3845 & w3857 ;
  assign w3859 = w3856 | w3858 ;
  assign w3860 = ( w455 & w3853 ) | ( w455 & ~w3859 ) | ( w3853 & ~w3859 ) ;
  assign w3861 = w455 & w3860 ;
  assign w3862 = w3607 | w3612 ;
  assign w3863 = w3695 & ~w3862 ;
  assign w3864 = w3610 ^ w3863 ;
  assign w3865 = ( ~w455 & w3853 ) | ( ~w455 & w3859 ) | ( w3853 & w3859 ) ;
  assign w3866 = ~w3853 & w3865 ;
  assign w3867 = w3864 | w3866 ;
  assign w3868 = ( w377 & w3861 ) | ( w377 & ~w3867 ) | ( w3861 & ~w3867 ) ;
  assign w3869 = w377 & w3868 ;
  assign w3870 = w3615 | w3620 ;
  assign w3871 = w3695 & ~w3870 ;
  assign w3872 = w3618 ^ w3871 ;
  assign w3873 = ( ~w377 & w3861 ) | ( ~w377 & w3867 ) | ( w3861 & w3867 ) ;
  assign w3874 = ~w3861 & w3873 ;
  assign w3875 = w3872 | w3874 ;
  assign w3876 = ( w307 & w3869 ) | ( w307 & ~w3875 ) | ( w3869 & ~w3875 ) ;
  assign w3877 = w307 & w3876 ;
  assign w3878 = w3623 | w3628 ;
  assign w3879 = w3695 & ~w3878 ;
  assign w3880 = w3626 ^ w3879 ;
  assign w3881 = ( ~w307 & w3869 ) | ( ~w307 & w3875 ) | ( w3869 & w3875 ) ;
  assign w3882 = ~w3869 & w3881 ;
  assign w3883 = w3880 | w3882 ;
  assign w3884 = ( w246 & w3877 ) | ( w246 & ~w3883 ) | ( w3877 & ~w3883 ) ;
  assign w3885 = w246 & w3884 ;
  assign w3886 = w3631 | w3636 ;
  assign w3887 = w3695 & ~w3886 ;
  assign w3888 = w3634 ^ w3887 ;
  assign w3889 = ( ~w246 & w3877 ) | ( ~w246 & w3883 ) | ( w3877 & w3883 ) ;
  assign w3890 = ~w3877 & w3889 ;
  assign w3891 = w3888 | w3890 ;
  assign w3892 = ( w185 & w3885 ) | ( w185 & ~w3891 ) | ( w3885 & ~w3891 ) ;
  assign w3893 = w185 & w3892 ;
  assign w3894 = w3639 | w3644 ;
  assign w3895 = w3695 & ~w3894 ;
  assign w3896 = w3642 ^ w3895 ;
  assign w3897 = ( ~w185 & w3885 ) | ( ~w185 & w3891 ) | ( w3885 & w3891 ) ;
  assign w3898 = ~w3885 & w3897 ;
  assign w3899 = w3896 | w3898 ;
  assign w3900 = ( w145 & w3893 ) | ( w145 & ~w3899 ) | ( w3893 & ~w3899 ) ;
  assign w3901 = w145 & w3900 ;
  assign w3902 = ( ~w145 & w3893 ) | ( ~w145 & w3899 ) | ( w3893 & w3899 ) ;
  assign w3903 = ~w3893 & w3902 ;
  assign w3904 = w3647 | w3649 ;
  assign w3905 = w3695 & ~w3904 ;
  assign w3906 = w3652 ^ w3905 ;
  assign w3907 = w3903 | w3906 ;
  assign w3908 = ( w132 & w3901 ) | ( w132 & ~w3907 ) | ( w3901 & ~w3907 ) ;
  assign w3909 = w132 & w3908 ;
  assign w3910 = w3655 | w3660 ;
  assign w3911 = w3695 & ~w3910 ;
  assign w3912 = w3658 ^ w3911 ;
  assign w3913 = ( ~w132 & w3901 ) | ( ~w132 & w3907 ) | ( w3901 & w3907 ) ;
  assign w3914 = ~w3901 & w3913 ;
  assign w3915 = w3912 | w3914 ;
  assign w3916 = ~w3909 & w3915 ;
  assign w3917 = w3663 | w3668 ;
  assign w3918 = w3695 & ~w3917 ;
  assign w3919 = w3666 ^ w3918 ;
  assign w3920 = ( ~w3681 & w3916 ) | ( ~w3681 & w3919 ) | ( w3916 & w3919 ) ;
  assign w3921 = w3670 & ~w3920 ;
  assign w3922 = ~w3673 & w3695 ;
  assign w3923 = ( w3920 & ~w3921 ) | ( w3920 & w3922 ) | ( ~w3921 & w3922 ) ;
  assign w3924 = w3681 | w3923 ;
  assign w3925 = ~w129 & w3924 ;
  assign w3926 = ( w3909 & w3915 ) | ( w3909 & w3919 ) | ( w3915 & w3919 ) ;
  assign w3927 = ~w3909 & w3926 ;
  assign w3928 = ( w129 & w3670 ) | ( w129 & w3673 ) | ( w3670 & w3673 ) ;
  assign w3929 = ( w3673 & ~w3695 ) | ( w3673 & w3928 ) | ( ~w3695 & w3928 ) ;
  assign w3930 = w3670 & w3929 ;
  assign w3931 = w3928 ^ w3930 ;
  assign w3932 = ( w3425 & w3430 ) | ( w3425 & w3457 ) | ( w3430 & w3457 ) ;
  assign w3933 = w3457 & ~w3932 ;
  assign w3934 = w3428 ^ w3933 ;
  assign w3935 = ( ~w3685 & w3692 ) | ( ~w3685 & w3934 ) | ( w3692 & w3934 ) ;
  assign w3936 = ~w3692 & w3935 ;
  assign w3937 = ( ~w3679 & w3681 ) | ( ~w3679 & w3936 ) | ( w3681 & w3936 ) ;
  assign w3938 = ~w3681 & w3937 ;
  assign w3939 = w3927 | w3938 ;
  assign w3940 = ( w3925 & ~w3927 ) | ( w3925 & w3931 ) | ( ~w3927 & w3931 ) ;
  assign w3941 = w3939 | w3940 ;
  assign w3942 = ( ~\pi069 & \pi070 ) | ( ~\pi069 & w3695 ) | ( \pi070 & w3695 ) ;
  assign w3943 = ( ~\pi068 & \pi070 ) | ( ~\pi068 & w3942 ) | ( \pi070 & w3942 ) ;
  assign w3944 = ( ~\pi070 & w3695 ) | ( ~\pi070 & w3941 ) | ( w3695 & w3941 ) ;
  assign w3945 = w3943 & w3944 ;
  assign w3946 = ( w3681 & w3685 ) | ( w3681 & ~w3692 ) | ( w3685 & ~w3692 ) ;
  assign w3947 = \pi069 & ~w3946 ;
  assign w3948 = \pi068 | \pi070 ;
  assign w3949 = ( ~w3946 & w3947 ) | ( ~w3946 & w3948 ) | ( w3947 & w3948 ) ;
  assign w3950 = ~w3692 & w3949 ;
  assign w3951 = ~w3679 & w3950 ;
  assign w3952 = ( \pi070 & w3941 ) | ( \pi070 & ~w3950 ) | ( w3941 & ~w3950 ) ;
  assign w3953 = w3951 & ~w3952 ;
  assign w3954 = ~\pi070 & w3941 ;
  assign w3955 = \pi071 ^ w3954 ;
  assign w3956 = w3953 | w3955 ;
  assign w3957 = ( w3457 & w3945 ) | ( w3457 & ~w3956 ) | ( w3945 & ~w3956 ) ;
  assign w3958 = w3457 & w3957 ;
  assign w3959 = ( ~w3457 & w3945 ) | ( ~w3457 & w3956 ) | ( w3945 & w3956 ) ;
  assign w3960 = ~w3945 & w3959 ;
  assign w3961 = w3695 & ~w3938 ;
  assign w3962 = ~w3927 & w3961 ;
  assign w3963 = ~w3940 & w3962 ;
  assign w3964 = \pi071 & w3941 ;
  assign w3965 = ( \pi070 & w3941 ) | ( \pi070 & ~w3964 ) | ( w3941 & ~w3964 ) ;
  assign w3966 = ( ~\pi070 & w3963 ) | ( ~\pi070 & w3965 ) | ( w3963 & w3965 ) ;
  assign w3967 = \pi072 ^ w3966 ;
  assign w3968 = w3960 | w3967 ;
  assign w3969 = ( w3227 & w3958 ) | ( w3227 & ~w3968 ) | ( w3958 & ~w3968 ) ;
  assign w3970 = w3227 & w3969 ;
  assign w3971 = ( w3699 & ~w3707 ) | ( w3699 & w3941 ) | ( ~w3707 & w3941 ) ;
  assign w3972 = ~w3699 & w3971 ;
  assign w3973 = \pi073 ^ w3972 ;
  assign w3974 = w3708 ^ w3973 ;
  assign w3975 = ( ~w3227 & w3958 ) | ( ~w3227 & w3968 ) | ( w3958 & w3968 ) ;
  assign w3976 = ~w3958 & w3975 ;
  assign w3977 = w3974 | w3976 ;
  assign w3978 = ( w3005 & w3970 ) | ( w3005 & ~w3977 ) | ( w3970 & ~w3977 ) ;
  assign w3979 = w3005 & w3978 ;
  assign w3980 = w3712 | w3714 ;
  assign w3981 = w3941 & ~w3980 ;
  assign w3982 = w3721 ^ w3981 ;
  assign w3983 = ( ~w3005 & w3970 ) | ( ~w3005 & w3977 ) | ( w3970 & w3977 ) ;
  assign w3984 = ~w3970 & w3983 ;
  assign w3985 = w3982 | w3984 ;
  assign w3986 = ( w2791 & w3979 ) | ( w2791 & ~w3985 ) | ( w3979 & ~w3985 ) ;
  assign w3987 = w2791 & w3986 ;
  assign w3988 = w3724 | w3730 ;
  assign w3989 = w3941 & ~w3988 ;
  assign w3990 = w3728 ^ w3989 ;
  assign w3991 = ( ~w2791 & w3979 ) | ( ~w2791 & w3985 ) | ( w3979 & w3985 ) ;
  assign w3992 = ~w3979 & w3991 ;
  assign w3993 = w3990 | w3992 ;
  assign w3994 = ( w2585 & w3987 ) | ( w2585 & ~w3993 ) | ( w3987 & ~w3993 ) ;
  assign w3995 = w2585 & w3994 ;
  assign w3996 = w3733 | w3738 ;
  assign w3997 = w3941 & ~w3996 ;
  assign w3998 = w3736 ^ w3997 ;
  assign w3999 = ( ~w2585 & w3987 ) | ( ~w2585 & w3993 ) | ( w3987 & w3993 ) ;
  assign w4000 = ~w3987 & w3999 ;
  assign w4001 = w3998 | w4000 ;
  assign w4002 = ( w2387 & w3995 ) | ( w2387 & ~w4001 ) | ( w3995 & ~w4001 ) ;
  assign w4003 = w2387 & w4002 ;
  assign w4004 = w3741 | w3746 ;
  assign w4005 = w3941 & ~w4004 ;
  assign w4006 = w3744 ^ w4005 ;
  assign w4007 = ( ~w2387 & w3995 ) | ( ~w2387 & w4001 ) | ( w3995 & w4001 ) ;
  assign w4008 = ~w3995 & w4007 ;
  assign w4009 = w4006 | w4008 ;
  assign w4010 = ( w2197 & w4003 ) | ( w2197 & ~w4009 ) | ( w4003 & ~w4009 ) ;
  assign w4011 = w2197 & w4010 ;
  assign w4012 = w3749 | w3754 ;
  assign w4013 = w3941 & ~w4012 ;
  assign w4014 = w3752 ^ w4013 ;
  assign w4015 = ( ~w2197 & w4003 ) | ( ~w2197 & w4009 ) | ( w4003 & w4009 ) ;
  assign w4016 = ~w4003 & w4015 ;
  assign w4017 = w4014 | w4016 ;
  assign w4018 = ( w2015 & w4011 ) | ( w2015 & ~w4017 ) | ( w4011 & ~w4017 ) ;
  assign w4019 = w2015 & w4018 ;
  assign w4020 = w3757 | w3762 ;
  assign w4021 = w3941 & ~w4020 ;
  assign w4022 = w3760 ^ w4021 ;
  assign w4023 = ( ~w2015 & w4011 ) | ( ~w2015 & w4017 ) | ( w4011 & w4017 ) ;
  assign w4024 = ~w4011 & w4023 ;
  assign w4025 = w4022 | w4024 ;
  assign w4026 = ( w1841 & w4019 ) | ( w1841 & ~w4025 ) | ( w4019 & ~w4025 ) ;
  assign w4027 = w1841 & w4026 ;
  assign w4028 = w3765 | w3770 ;
  assign w4029 = w3941 & ~w4028 ;
  assign w4030 = w3768 ^ w4029 ;
  assign w4031 = ( ~w1841 & w4019 ) | ( ~w1841 & w4025 ) | ( w4019 & w4025 ) ;
  assign w4032 = ~w4019 & w4031 ;
  assign w4033 = w4030 | w4032 ;
  assign w4034 = ( w1675 & w4027 ) | ( w1675 & ~w4033 ) | ( w4027 & ~w4033 ) ;
  assign w4035 = w1675 & w4034 ;
  assign w4036 = w3773 | w3778 ;
  assign w4037 = w3941 & ~w4036 ;
  assign w4038 = w3776 ^ w4037 ;
  assign w4039 = ( ~w1675 & w4027 ) | ( ~w1675 & w4033 ) | ( w4027 & w4033 ) ;
  assign w4040 = ~w4027 & w4039 ;
  assign w4041 = w4038 | w4040 ;
  assign w4042 = ( w1517 & w4035 ) | ( w1517 & ~w4041 ) | ( w4035 & ~w4041 ) ;
  assign w4043 = w1517 & w4042 ;
  assign w4044 = w3781 | w3786 ;
  assign w4045 = w3941 & ~w4044 ;
  assign w4046 = w3784 ^ w4045 ;
  assign w4047 = ( ~w1517 & w4035 ) | ( ~w1517 & w4041 ) | ( w4035 & w4041 ) ;
  assign w4048 = ~w4035 & w4047 ;
  assign w4049 = w4046 | w4048 ;
  assign w4050 = ( w1367 & w4043 ) | ( w1367 & ~w4049 ) | ( w4043 & ~w4049 ) ;
  assign w4051 = w1367 & w4050 ;
  assign w4052 = w3789 | w3794 ;
  assign w4053 = w3941 & ~w4052 ;
  assign w4054 = w3792 ^ w4053 ;
  assign w4055 = ( ~w1367 & w4043 ) | ( ~w1367 & w4049 ) | ( w4043 & w4049 ) ;
  assign w4056 = ~w4043 & w4055 ;
  assign w4057 = w4054 | w4056 ;
  assign w4058 = ( w1225 & w4051 ) | ( w1225 & ~w4057 ) | ( w4051 & ~w4057 ) ;
  assign w4059 = w1225 & w4058 ;
  assign w4060 = w3797 | w3802 ;
  assign w4061 = w3941 & ~w4060 ;
  assign w4062 = w3800 ^ w4061 ;
  assign w4063 = ( ~w1225 & w4051 ) | ( ~w1225 & w4057 ) | ( w4051 & w4057 ) ;
  assign w4064 = ~w4051 & w4063 ;
  assign w4065 = w4062 | w4064 ;
  assign w4066 = ( w1091 & w4059 ) | ( w1091 & ~w4065 ) | ( w4059 & ~w4065 ) ;
  assign w4067 = w1091 & w4066 ;
  assign w4068 = w3805 | w3810 ;
  assign w4069 = w3941 & ~w4068 ;
  assign w4070 = w3808 ^ w4069 ;
  assign w4071 = ( ~w1091 & w4059 ) | ( ~w1091 & w4065 ) | ( w4059 & w4065 ) ;
  assign w4072 = ~w4059 & w4071 ;
  assign w4073 = w4070 | w4072 ;
  assign w4074 = ( w965 & w4067 ) | ( w965 & ~w4073 ) | ( w4067 & ~w4073 ) ;
  assign w4075 = w965 & w4074 ;
  assign w4076 = w3813 | w3818 ;
  assign w4077 = w3941 & ~w4076 ;
  assign w4078 = w3816 ^ w4077 ;
  assign w4079 = ( ~w965 & w4067 ) | ( ~w965 & w4073 ) | ( w4067 & w4073 ) ;
  assign w4080 = ~w4067 & w4079 ;
  assign w4081 = w4078 | w4080 ;
  assign w4082 = ( w847 & w4075 ) | ( w847 & ~w4081 ) | ( w4075 & ~w4081 ) ;
  assign w4083 = w847 & w4082 ;
  assign w4084 = w3821 | w3826 ;
  assign w4085 = w3941 & ~w4084 ;
  assign w4086 = w3824 ^ w4085 ;
  assign w4087 = ( ~w847 & w4075 ) | ( ~w847 & w4081 ) | ( w4075 & w4081 ) ;
  assign w4088 = ~w4075 & w4087 ;
  assign w4089 = w4086 | w4088 ;
  assign w4090 = ( w737 & w4083 ) | ( w737 & ~w4089 ) | ( w4083 & ~w4089 ) ;
  assign w4091 = w737 & w4090 ;
  assign w4092 = w3829 | w3834 ;
  assign w4093 = w3941 & ~w4092 ;
  assign w4094 = w3832 ^ w4093 ;
  assign w4095 = ( ~w737 & w4083 ) | ( ~w737 & w4089 ) | ( w4083 & w4089 ) ;
  assign w4096 = ~w4083 & w4095 ;
  assign w4097 = w4094 | w4096 ;
  assign w4098 = ( w635 & w4091 ) | ( w635 & ~w4097 ) | ( w4091 & ~w4097 ) ;
  assign w4099 = w635 & w4098 ;
  assign w4100 = w3837 | w3842 ;
  assign w4101 = w3941 & ~w4100 ;
  assign w4102 = w3840 ^ w4101 ;
  assign w4103 = ( ~w635 & w4091 ) | ( ~w635 & w4097 ) | ( w4091 & w4097 ) ;
  assign w4104 = ~w4091 & w4103 ;
  assign w4105 = w4102 | w4104 ;
  assign w4106 = ( w541 & w4099 ) | ( w541 & ~w4105 ) | ( w4099 & ~w4105 ) ;
  assign w4107 = w541 & w4106 ;
  assign w4108 = w3845 | w3850 ;
  assign w4109 = w3941 & ~w4108 ;
  assign w4110 = w3848 ^ w4109 ;
  assign w4111 = ( ~w541 & w4099 ) | ( ~w541 & w4105 ) | ( w4099 & w4105 ) ;
  assign w4112 = ~w4099 & w4111 ;
  assign w4113 = w4110 | w4112 ;
  assign w4114 = ( w455 & w4107 ) | ( w455 & ~w4113 ) | ( w4107 & ~w4113 ) ;
  assign w4115 = w455 & w4114 ;
  assign w4116 = w3853 | w3858 ;
  assign w4117 = w3941 & ~w4116 ;
  assign w4118 = w3856 ^ w4117 ;
  assign w4119 = ( ~w455 & w4107 ) | ( ~w455 & w4113 ) | ( w4107 & w4113 ) ;
  assign w4120 = ~w4107 & w4119 ;
  assign w4121 = w4118 | w4120 ;
  assign w4122 = ( w377 & w4115 ) | ( w377 & ~w4121 ) | ( w4115 & ~w4121 ) ;
  assign w4123 = w377 & w4122 ;
  assign w4124 = w3861 | w3866 ;
  assign w4125 = w3941 & ~w4124 ;
  assign w4126 = w3864 ^ w4125 ;
  assign w4127 = ( ~w377 & w4115 ) | ( ~w377 & w4121 ) | ( w4115 & w4121 ) ;
  assign w4128 = ~w4115 & w4127 ;
  assign w4129 = w4126 | w4128 ;
  assign w4130 = ( w307 & w4123 ) | ( w307 & ~w4129 ) | ( w4123 & ~w4129 ) ;
  assign w4131 = w307 & w4130 ;
  assign w4132 = w3869 | w3874 ;
  assign w4133 = w3941 & ~w4132 ;
  assign w4134 = w3872 ^ w4133 ;
  assign w4135 = ( ~w307 & w4123 ) | ( ~w307 & w4129 ) | ( w4123 & w4129 ) ;
  assign w4136 = ~w4123 & w4135 ;
  assign w4137 = w4134 | w4136 ;
  assign w4138 = ( w246 & w4131 ) | ( w246 & ~w4137 ) | ( w4131 & ~w4137 ) ;
  assign w4139 = w246 & w4138 ;
  assign w4140 = w3877 | w3882 ;
  assign w4141 = w3941 & ~w4140 ;
  assign w4142 = w3880 ^ w4141 ;
  assign w4143 = ( ~w246 & w4131 ) | ( ~w246 & w4137 ) | ( w4131 & w4137 ) ;
  assign w4144 = ~w4131 & w4143 ;
  assign w4145 = w4142 | w4144 ;
  assign w4146 = ( w185 & w4139 ) | ( w185 & ~w4145 ) | ( w4139 & ~w4145 ) ;
  assign w4147 = w185 & w4146 ;
  assign w4148 = w3885 | w3890 ;
  assign w4149 = w3941 & ~w4148 ;
  assign w4150 = w3888 ^ w4149 ;
  assign w4151 = ( ~w185 & w4139 ) | ( ~w185 & w4145 ) | ( w4139 & w4145 ) ;
  assign w4152 = ~w4139 & w4151 ;
  assign w4153 = w4150 | w4152 ;
  assign w4154 = ( w145 & w4147 ) | ( w145 & ~w4153 ) | ( w4147 & ~w4153 ) ;
  assign w4155 = w145 & w4154 ;
  assign w4156 = w3893 | w3898 ;
  assign w4157 = w3941 & ~w4156 ;
  assign w4158 = w3896 ^ w4157 ;
  assign w4159 = ( ~w145 & w4147 ) | ( ~w145 & w4153 ) | ( w4147 & w4153 ) ;
  assign w4160 = ~w4147 & w4159 ;
  assign w4161 = w4158 | w4160 ;
  assign w4162 = ( w132 & w4155 ) | ( w132 & ~w4161 ) | ( w4155 & ~w4161 ) ;
  assign w4163 = w132 & w4162 ;
  assign w4164 = ( ~w132 & w4155 ) | ( ~w132 & w4161 ) | ( w4155 & w4161 ) ;
  assign w4165 = ~w4155 & w4164 ;
  assign w4166 = w3901 | w3903 ;
  assign w4167 = w3941 & ~w4166 ;
  assign w4168 = w3906 ^ w4167 ;
  assign w4169 = w4165 | w4168 ;
  assign w4170 = ~w4163 & w4169 ;
  assign w4171 = w3909 | w3914 ;
  assign w4172 = w3941 & ~w4171 ;
  assign w4173 = w3912 ^ w4172 ;
  assign w4174 = ( ~w3927 & w4170 ) | ( ~w3927 & w4173 ) | ( w4170 & w4173 ) ;
  assign w4175 = w3916 & ~w4174 ;
  assign w4176 = ~w3919 & w3941 ;
  assign w4177 = ( w4174 & ~w4175 ) | ( w4174 & w4176 ) | ( ~w4175 & w4176 ) ;
  assign w4178 = w3927 | w4177 ;
  assign w4179 = ~w129 & w4178 ;
  assign w4180 = ( w4163 & w4169 ) | ( w4163 & w4173 ) | ( w4169 & w4173 ) ;
  assign w4181 = ~w4163 & w4180 ;
  assign w4182 = ( w129 & w3916 ) | ( w129 & w3919 ) | ( w3916 & w3919 ) ;
  assign w4183 = ( w3919 & ~w3941 ) | ( w3919 & w4182 ) | ( ~w3941 & w4182 ) ;
  assign w4184 = w3916 & w4183 ;
  assign w4185 = w4182 ^ w4184 ;
  assign w4186 = ( w3663 & w3668 ) | ( w3663 & w3695 ) | ( w3668 & w3695 ) ;
  assign w4187 = w3695 & ~w4186 ;
  assign w4188 = w3666 ^ w4187 ;
  assign w4189 = ( ~w3931 & w3938 ) | ( ~w3931 & w4188 ) | ( w3938 & w4188 ) ;
  assign w4190 = ~w3938 & w4189 ;
  assign w4191 = ( ~w3925 & w3927 ) | ( ~w3925 & w4190 ) | ( w3927 & w4190 ) ;
  assign w4192 = ~w3927 & w4191 ;
  assign w4193 = w4181 | w4192 ;
  assign w4194 = ( w4179 & ~w4181 ) | ( w4179 & w4185 ) | ( ~w4181 & w4185 ) ;
  assign w4195 = w4193 | w4194 ;
  assign w4196 = ( ~\pi067 & \pi068 ) | ( ~\pi067 & w3941 ) | ( \pi068 & w3941 ) ;
  assign w4197 = ( ~\pi066 & \pi068 ) | ( ~\pi066 & w4196 ) | ( \pi068 & w4196 ) ;
  assign w4198 = ( ~\pi068 & w3941 ) | ( ~\pi068 & w4195 ) | ( w3941 & w4195 ) ;
  assign w4199 = w4197 & w4198 ;
  assign w4200 = ( w3927 & w3931 ) | ( w3927 & ~w3938 ) | ( w3931 & ~w3938 ) ;
  assign w4201 = \pi067 & ~w4200 ;
  assign w4202 = \pi066 | \pi068 ;
  assign w4203 = ( ~w4200 & w4201 ) | ( ~w4200 & w4202 ) | ( w4201 & w4202 ) ;
  assign w4204 = ~w3938 & w4203 ;
  assign w4205 = ~w3925 & w4204 ;
  assign w4206 = ( \pi068 & w4195 ) | ( \pi068 & ~w4204 ) | ( w4195 & ~w4204 ) ;
  assign w4207 = w4205 & ~w4206 ;
  assign w4208 = ~\pi068 & w4195 ;
  assign w4209 = \pi069 ^ w4208 ;
  assign w4210 = w4207 | w4209 ;
  assign w4211 = ( w3695 & w4199 ) | ( w3695 & ~w4210 ) | ( w4199 & ~w4210 ) ;
  assign w4212 = w3695 & w4211 ;
  assign w4213 = ( ~w3695 & w4199 ) | ( ~w3695 & w4210 ) | ( w4199 & w4210 ) ;
  assign w4214 = ~w4199 & w4213 ;
  assign w4215 = w3941 & ~w4192 ;
  assign w4216 = ~w4181 & w4215 ;
  assign w4217 = ~w4194 & w4216 ;
  assign w4218 = \pi069 & w4195 ;
  assign w4219 = ( \pi068 & w4195 ) | ( \pi068 & ~w4218 ) | ( w4195 & ~w4218 ) ;
  assign w4220 = ( ~\pi068 & w4217 ) | ( ~\pi068 & w4219 ) | ( w4217 & w4219 ) ;
  assign w4221 = \pi070 ^ w4220 ;
  assign w4222 = w4214 | w4221 ;
  assign w4223 = ( w3457 & w4212 ) | ( w3457 & ~w4222 ) | ( w4212 & ~w4222 ) ;
  assign w4224 = w3457 & w4223 ;
  assign w4225 = ( w3945 & ~w3953 ) | ( w3945 & w4195 ) | ( ~w3953 & w4195 ) ;
  assign w4226 = ~w3945 & w4225 ;
  assign w4227 = \pi071 ^ w4226 ;
  assign w4228 = w3954 ^ w4227 ;
  assign w4229 = ( ~w3457 & w4212 ) | ( ~w3457 & w4222 ) | ( w4212 & w4222 ) ;
  assign w4230 = ~w4212 & w4229 ;
  assign w4231 = w4228 | w4230 ;
  assign w4232 = ( w3227 & w4224 ) | ( w3227 & ~w4231 ) | ( w4224 & ~w4231 ) ;
  assign w4233 = w3227 & w4232 ;
  assign w4234 = w3958 | w3960 ;
  assign w4235 = w4195 & ~w4234 ;
  assign w4236 = w3967 ^ w4235 ;
  assign w4237 = ( ~w3227 & w4224 ) | ( ~w3227 & w4231 ) | ( w4224 & w4231 ) ;
  assign w4238 = ~w4224 & w4237 ;
  assign w4239 = w4236 | w4238 ;
  assign w4240 = ( w3005 & w4233 ) | ( w3005 & ~w4239 ) | ( w4233 & ~w4239 ) ;
  assign w4241 = w3005 & w4240 ;
  assign w4242 = w3970 | w3976 ;
  assign w4243 = w4195 & ~w4242 ;
  assign w4244 = w3974 ^ w4243 ;
  assign w4245 = ( ~w3005 & w4233 ) | ( ~w3005 & w4239 ) | ( w4233 & w4239 ) ;
  assign w4246 = ~w4233 & w4245 ;
  assign w4247 = w4244 | w4246 ;
  assign w4248 = ( w2791 & w4241 ) | ( w2791 & ~w4247 ) | ( w4241 & ~w4247 ) ;
  assign w4249 = w2791 & w4248 ;
  assign w4250 = w3979 | w3984 ;
  assign w4251 = w4195 & ~w4250 ;
  assign w4252 = w3982 ^ w4251 ;
  assign w4253 = ( ~w2791 & w4241 ) | ( ~w2791 & w4247 ) | ( w4241 & w4247 ) ;
  assign w4254 = ~w4241 & w4253 ;
  assign w4255 = w4252 | w4254 ;
  assign w4256 = ( w2585 & w4249 ) | ( w2585 & ~w4255 ) | ( w4249 & ~w4255 ) ;
  assign w4257 = w2585 & w4256 ;
  assign w4258 = w3987 | w3992 ;
  assign w4259 = w4195 & ~w4258 ;
  assign w4260 = w3990 ^ w4259 ;
  assign w4261 = ( ~w2585 & w4249 ) | ( ~w2585 & w4255 ) | ( w4249 & w4255 ) ;
  assign w4262 = ~w4249 & w4261 ;
  assign w4263 = w4260 | w4262 ;
  assign w4264 = ( w2387 & w4257 ) | ( w2387 & ~w4263 ) | ( w4257 & ~w4263 ) ;
  assign w4265 = w2387 & w4264 ;
  assign w4266 = w3995 | w4000 ;
  assign w4267 = w4195 & ~w4266 ;
  assign w4268 = w3998 ^ w4267 ;
  assign w4269 = ( ~w2387 & w4257 ) | ( ~w2387 & w4263 ) | ( w4257 & w4263 ) ;
  assign w4270 = ~w4257 & w4269 ;
  assign w4271 = w4268 | w4270 ;
  assign w4272 = ( w2197 & w4265 ) | ( w2197 & ~w4271 ) | ( w4265 & ~w4271 ) ;
  assign w4273 = w2197 & w4272 ;
  assign w4274 = w4003 | w4008 ;
  assign w4275 = w4195 & ~w4274 ;
  assign w4276 = w4006 ^ w4275 ;
  assign w4277 = ( ~w2197 & w4265 ) | ( ~w2197 & w4271 ) | ( w4265 & w4271 ) ;
  assign w4278 = ~w4265 & w4277 ;
  assign w4279 = w4276 | w4278 ;
  assign w4280 = ( w2015 & w4273 ) | ( w2015 & ~w4279 ) | ( w4273 & ~w4279 ) ;
  assign w4281 = w2015 & w4280 ;
  assign w4282 = w4011 | w4016 ;
  assign w4283 = w4195 & ~w4282 ;
  assign w4284 = w4014 ^ w4283 ;
  assign w4285 = ( ~w2015 & w4273 ) | ( ~w2015 & w4279 ) | ( w4273 & w4279 ) ;
  assign w4286 = ~w4273 & w4285 ;
  assign w4287 = w4284 | w4286 ;
  assign w4288 = ( w1841 & w4281 ) | ( w1841 & ~w4287 ) | ( w4281 & ~w4287 ) ;
  assign w4289 = w1841 & w4288 ;
  assign w4290 = w4019 | w4024 ;
  assign w4291 = w4195 & ~w4290 ;
  assign w4292 = w4022 ^ w4291 ;
  assign w4293 = ( ~w1841 & w4281 ) | ( ~w1841 & w4287 ) | ( w4281 & w4287 ) ;
  assign w4294 = ~w4281 & w4293 ;
  assign w4295 = w4292 | w4294 ;
  assign w4296 = ( w1675 & w4289 ) | ( w1675 & ~w4295 ) | ( w4289 & ~w4295 ) ;
  assign w4297 = w1675 & w4296 ;
  assign w4298 = w4027 | w4032 ;
  assign w4299 = w4195 & ~w4298 ;
  assign w4300 = w4030 ^ w4299 ;
  assign w4301 = ( ~w1675 & w4289 ) | ( ~w1675 & w4295 ) | ( w4289 & w4295 ) ;
  assign w4302 = ~w4289 & w4301 ;
  assign w4303 = w4300 | w4302 ;
  assign w4304 = ( w1517 & w4297 ) | ( w1517 & ~w4303 ) | ( w4297 & ~w4303 ) ;
  assign w4305 = w1517 & w4304 ;
  assign w4306 = w4035 | w4040 ;
  assign w4307 = w4195 & ~w4306 ;
  assign w4308 = w4038 ^ w4307 ;
  assign w4309 = ( ~w1517 & w4297 ) | ( ~w1517 & w4303 ) | ( w4297 & w4303 ) ;
  assign w4310 = ~w4297 & w4309 ;
  assign w4311 = w4308 | w4310 ;
  assign w4312 = ( w1367 & w4305 ) | ( w1367 & ~w4311 ) | ( w4305 & ~w4311 ) ;
  assign w4313 = w1367 & w4312 ;
  assign w4314 = w4043 | w4048 ;
  assign w4315 = w4195 & ~w4314 ;
  assign w4316 = w4046 ^ w4315 ;
  assign w4317 = ( ~w1367 & w4305 ) | ( ~w1367 & w4311 ) | ( w4305 & w4311 ) ;
  assign w4318 = ~w4305 & w4317 ;
  assign w4319 = w4316 | w4318 ;
  assign w4320 = ( w1225 & w4313 ) | ( w1225 & ~w4319 ) | ( w4313 & ~w4319 ) ;
  assign w4321 = w1225 & w4320 ;
  assign w4322 = w4051 | w4056 ;
  assign w4323 = w4195 & ~w4322 ;
  assign w4324 = w4054 ^ w4323 ;
  assign w4325 = ( ~w1225 & w4313 ) | ( ~w1225 & w4319 ) | ( w4313 & w4319 ) ;
  assign w4326 = ~w4313 & w4325 ;
  assign w4327 = w4324 | w4326 ;
  assign w4328 = ( w1091 & w4321 ) | ( w1091 & ~w4327 ) | ( w4321 & ~w4327 ) ;
  assign w4329 = w1091 & w4328 ;
  assign w4330 = w4059 | w4064 ;
  assign w4331 = w4195 & ~w4330 ;
  assign w4332 = w4062 ^ w4331 ;
  assign w4333 = ( ~w1091 & w4321 ) | ( ~w1091 & w4327 ) | ( w4321 & w4327 ) ;
  assign w4334 = ~w4321 & w4333 ;
  assign w4335 = w4332 | w4334 ;
  assign w4336 = ( w965 & w4329 ) | ( w965 & ~w4335 ) | ( w4329 & ~w4335 ) ;
  assign w4337 = w965 & w4336 ;
  assign w4338 = w4067 | w4072 ;
  assign w4339 = w4195 & ~w4338 ;
  assign w4340 = w4070 ^ w4339 ;
  assign w4341 = ( ~w965 & w4329 ) | ( ~w965 & w4335 ) | ( w4329 & w4335 ) ;
  assign w4342 = ~w4329 & w4341 ;
  assign w4343 = w4340 | w4342 ;
  assign w4344 = ( w847 & w4337 ) | ( w847 & ~w4343 ) | ( w4337 & ~w4343 ) ;
  assign w4345 = w847 & w4344 ;
  assign w4346 = w4075 | w4080 ;
  assign w4347 = w4195 & ~w4346 ;
  assign w4348 = w4078 ^ w4347 ;
  assign w4349 = ( ~w847 & w4337 ) | ( ~w847 & w4343 ) | ( w4337 & w4343 ) ;
  assign w4350 = ~w4337 & w4349 ;
  assign w4351 = w4348 | w4350 ;
  assign w4352 = ( w737 & w4345 ) | ( w737 & ~w4351 ) | ( w4345 & ~w4351 ) ;
  assign w4353 = w737 & w4352 ;
  assign w4354 = w4083 | w4088 ;
  assign w4355 = w4195 & ~w4354 ;
  assign w4356 = w4086 ^ w4355 ;
  assign w4357 = ( ~w737 & w4345 ) | ( ~w737 & w4351 ) | ( w4345 & w4351 ) ;
  assign w4358 = ~w4345 & w4357 ;
  assign w4359 = w4356 | w4358 ;
  assign w4360 = ( w635 & w4353 ) | ( w635 & ~w4359 ) | ( w4353 & ~w4359 ) ;
  assign w4361 = w635 & w4360 ;
  assign w4362 = w4091 | w4096 ;
  assign w4363 = w4195 & ~w4362 ;
  assign w4364 = w4094 ^ w4363 ;
  assign w4365 = ( ~w635 & w4353 ) | ( ~w635 & w4359 ) | ( w4353 & w4359 ) ;
  assign w4366 = ~w4353 & w4365 ;
  assign w4367 = w4364 | w4366 ;
  assign w4368 = ( w541 & w4361 ) | ( w541 & ~w4367 ) | ( w4361 & ~w4367 ) ;
  assign w4369 = w541 & w4368 ;
  assign w4370 = w4099 | w4104 ;
  assign w4371 = w4195 & ~w4370 ;
  assign w4372 = w4102 ^ w4371 ;
  assign w4373 = ( ~w541 & w4361 ) | ( ~w541 & w4367 ) | ( w4361 & w4367 ) ;
  assign w4374 = ~w4361 & w4373 ;
  assign w4375 = w4372 | w4374 ;
  assign w4376 = ( w455 & w4369 ) | ( w455 & ~w4375 ) | ( w4369 & ~w4375 ) ;
  assign w4377 = w455 & w4376 ;
  assign w4378 = w4107 | w4112 ;
  assign w4379 = w4195 & ~w4378 ;
  assign w4380 = w4110 ^ w4379 ;
  assign w4381 = ( ~w455 & w4369 ) | ( ~w455 & w4375 ) | ( w4369 & w4375 ) ;
  assign w4382 = ~w4369 & w4381 ;
  assign w4383 = w4380 | w4382 ;
  assign w4384 = ( w377 & w4377 ) | ( w377 & ~w4383 ) | ( w4377 & ~w4383 ) ;
  assign w4385 = w377 & w4384 ;
  assign w4386 = w4115 | w4120 ;
  assign w4387 = w4195 & ~w4386 ;
  assign w4388 = w4118 ^ w4387 ;
  assign w4389 = ( ~w377 & w4377 ) | ( ~w377 & w4383 ) | ( w4377 & w4383 ) ;
  assign w4390 = ~w4377 & w4389 ;
  assign w4391 = w4388 | w4390 ;
  assign w4392 = ( w307 & w4385 ) | ( w307 & ~w4391 ) | ( w4385 & ~w4391 ) ;
  assign w4393 = w307 & w4392 ;
  assign w4394 = w4123 | w4128 ;
  assign w4395 = w4195 & ~w4394 ;
  assign w4396 = w4126 ^ w4395 ;
  assign w4397 = ( ~w307 & w4385 ) | ( ~w307 & w4391 ) | ( w4385 & w4391 ) ;
  assign w4398 = ~w4385 & w4397 ;
  assign w4399 = w4396 | w4398 ;
  assign w4400 = ( w246 & w4393 ) | ( w246 & ~w4399 ) | ( w4393 & ~w4399 ) ;
  assign w4401 = w246 & w4400 ;
  assign w4402 = w4131 | w4136 ;
  assign w4403 = w4195 & ~w4402 ;
  assign w4404 = w4134 ^ w4403 ;
  assign w4405 = ( ~w246 & w4393 ) | ( ~w246 & w4399 ) | ( w4393 & w4399 ) ;
  assign w4406 = ~w4393 & w4405 ;
  assign w4407 = w4404 | w4406 ;
  assign w4408 = ( w185 & w4401 ) | ( w185 & ~w4407 ) | ( w4401 & ~w4407 ) ;
  assign w4409 = w185 & w4408 ;
  assign w4410 = w4139 | w4144 ;
  assign w4411 = w4195 & ~w4410 ;
  assign w4412 = w4142 ^ w4411 ;
  assign w4413 = ( ~w185 & w4401 ) | ( ~w185 & w4407 ) | ( w4401 & w4407 ) ;
  assign w4414 = ~w4401 & w4413 ;
  assign w4415 = w4412 | w4414 ;
  assign w4416 = ( w145 & w4409 ) | ( w145 & ~w4415 ) | ( w4409 & ~w4415 ) ;
  assign w4417 = w145 & w4416 ;
  assign w4418 = w4147 | w4152 ;
  assign w4419 = w4195 & ~w4418 ;
  assign w4420 = w4150 ^ w4419 ;
  assign w4421 = ( ~w145 & w4409 ) | ( ~w145 & w4415 ) | ( w4409 & w4415 ) ;
  assign w4422 = ~w4409 & w4421 ;
  assign w4423 = w4420 | w4422 ;
  assign w4424 = ( w132 & w4417 ) | ( w132 & ~w4423 ) | ( w4417 & ~w4423 ) ;
  assign w4425 = w132 & w4424 ;
  assign w4426 = w4155 | w4160 ;
  assign w4427 = w4195 & ~w4426 ;
  assign w4428 = w4158 ^ w4427 ;
  assign w4429 = ( ~w132 & w4417 ) | ( ~w132 & w4423 ) | ( w4417 & w4423 ) ;
  assign w4430 = ~w4417 & w4429 ;
  assign w4431 = w4428 | w4430 ;
  assign w4432 = ~w4425 & w4431 ;
  assign w4433 = w4163 | w4165 ;
  assign w4434 = w4195 & ~w4433 ;
  assign w4435 = w4168 ^ w4434 ;
  assign w4436 = ( ~w4181 & w4432 ) | ( ~w4181 & w4435 ) | ( w4432 & w4435 ) ;
  assign w4437 = w4170 & ~w4436 ;
  assign w4438 = ~w4173 & w4195 ;
  assign w4439 = ( w4436 & ~w4437 ) | ( w4436 & w4438 ) | ( ~w4437 & w4438 ) ;
  assign w4440 = w4181 | w4439 ;
  assign w4441 = ~w129 & w4440 ;
  assign w4442 = ( w4425 & w4431 ) | ( w4425 & w4435 ) | ( w4431 & w4435 ) ;
  assign w4443 = ~w4425 & w4442 ;
  assign w4444 = ( w129 & w4170 ) | ( w129 & w4173 ) | ( w4170 & w4173 ) ;
  assign w4445 = ( w4173 & ~w4195 ) | ( w4173 & w4444 ) | ( ~w4195 & w4444 ) ;
  assign w4446 = w4170 & w4445 ;
  assign w4447 = w4444 ^ w4446 ;
  assign w4448 = ( w3909 & w3914 ) | ( w3909 & w3941 ) | ( w3914 & w3941 ) ;
  assign w4449 = w3941 & ~w4448 ;
  assign w4450 = w3912 ^ w4449 ;
  assign w4451 = ( ~w4185 & w4192 ) | ( ~w4185 & w4450 ) | ( w4192 & w4450 ) ;
  assign w4452 = ~w4192 & w4451 ;
  assign w4453 = ( ~w4179 & w4181 ) | ( ~w4179 & w4452 ) | ( w4181 & w4452 ) ;
  assign w4454 = ~w4181 & w4453 ;
  assign w4455 = w4443 | w4454 ;
  assign w4456 = ( w4441 & ~w4443 ) | ( w4441 & w4447 ) | ( ~w4443 & w4447 ) ;
  assign w4457 = w4455 | w4456 ;
  assign w4458 = ( ~\pi065 & \pi066 ) | ( ~\pi065 & w4195 ) | ( \pi066 & w4195 ) ;
  assign w4459 = ( ~\pi064 & \pi066 ) | ( ~\pi064 & w4458 ) | ( \pi066 & w4458 ) ;
  assign w4460 = ( ~\pi066 & w4195 ) | ( ~\pi066 & w4457 ) | ( w4195 & w4457 ) ;
  assign w4461 = w4459 & w4460 ;
  assign w4462 = ( w4181 & w4185 ) | ( w4181 & ~w4192 ) | ( w4185 & ~w4192 ) ;
  assign w4463 = \pi065 & ~w4462 ;
  assign w4464 = \pi064 | \pi066 ;
  assign w4465 = ( ~w4462 & w4463 ) | ( ~w4462 & w4464 ) | ( w4463 & w4464 ) ;
  assign w4466 = ~w4192 & w4465 ;
  assign w4467 = ~w4179 & w4466 ;
  assign w4468 = ( \pi066 & w4457 ) | ( \pi066 & ~w4466 ) | ( w4457 & ~w4466 ) ;
  assign w4469 = w4467 & ~w4468 ;
  assign w4470 = ~\pi066 & w4457 ;
  assign w4471 = \pi067 ^ w4470 ;
  assign w4472 = w4469 | w4471 ;
  assign w4473 = ( w3941 & w4461 ) | ( w3941 & ~w4472 ) | ( w4461 & ~w4472 ) ;
  assign w4474 = w3941 & w4473 ;
  assign w4475 = ( ~w3941 & w4461 ) | ( ~w3941 & w4472 ) | ( w4461 & w4472 ) ;
  assign w4476 = ~w4461 & w4475 ;
  assign w4477 = w4195 & ~w4454 ;
  assign w4478 = ~w4443 & w4477 ;
  assign w4479 = ~w4456 & w4478 ;
  assign w4480 = \pi067 & w4457 ;
  assign w4481 = ( \pi066 & w4457 ) | ( \pi066 & ~w4480 ) | ( w4457 & ~w4480 ) ;
  assign w4482 = ( ~\pi066 & w4479 ) | ( ~\pi066 & w4481 ) | ( w4479 & w4481 ) ;
  assign w4483 = \pi068 ^ w4482 ;
  assign w4484 = w4476 | w4483 ;
  assign w4485 = ( w3695 & w4474 ) | ( w3695 & ~w4484 ) | ( w4474 & ~w4484 ) ;
  assign w4486 = w3695 & w4485 ;
  assign w4487 = ( w4199 & ~w4207 ) | ( w4199 & w4457 ) | ( ~w4207 & w4457 ) ;
  assign w4488 = ~w4199 & w4487 ;
  assign w4489 = \pi069 ^ w4488 ;
  assign w4490 = w4208 ^ w4489 ;
  assign w4491 = ( ~w3695 & w4474 ) | ( ~w3695 & w4484 ) | ( w4474 & w4484 ) ;
  assign w4492 = ~w4474 & w4491 ;
  assign w4493 = w4490 | w4492 ;
  assign w4494 = ( w3457 & w4486 ) | ( w3457 & ~w4493 ) | ( w4486 & ~w4493 ) ;
  assign w4495 = w3457 & w4494 ;
  assign w4496 = w4212 | w4214 ;
  assign w4497 = w4457 & ~w4496 ;
  assign w4498 = w4221 ^ w4497 ;
  assign w4499 = ( ~w3457 & w4486 ) | ( ~w3457 & w4493 ) | ( w4486 & w4493 ) ;
  assign w4500 = ~w4486 & w4499 ;
  assign w4501 = w4498 | w4500 ;
  assign w4502 = ( w3227 & w4495 ) | ( w3227 & ~w4501 ) | ( w4495 & ~w4501 ) ;
  assign w4503 = w3227 & w4502 ;
  assign w4504 = w4224 | w4230 ;
  assign w4505 = w4457 & ~w4504 ;
  assign w4506 = w4228 ^ w4505 ;
  assign w4507 = ( ~w3227 & w4495 ) | ( ~w3227 & w4501 ) | ( w4495 & w4501 ) ;
  assign w4508 = ~w4495 & w4507 ;
  assign w4509 = w4506 | w4508 ;
  assign w4510 = ( w3005 & w4503 ) | ( w3005 & ~w4509 ) | ( w4503 & ~w4509 ) ;
  assign w4511 = w3005 & w4510 ;
  assign w4512 = w4233 | w4238 ;
  assign w4513 = w4457 & ~w4512 ;
  assign w4514 = w4236 ^ w4513 ;
  assign w4515 = ( ~w3005 & w4503 ) | ( ~w3005 & w4509 ) | ( w4503 & w4509 ) ;
  assign w4516 = ~w4503 & w4515 ;
  assign w4517 = w4514 | w4516 ;
  assign w4518 = ( w2791 & w4511 ) | ( w2791 & ~w4517 ) | ( w4511 & ~w4517 ) ;
  assign w4519 = w2791 & w4518 ;
  assign w4520 = w4241 | w4246 ;
  assign w4521 = w4457 & ~w4520 ;
  assign w4522 = w4244 ^ w4521 ;
  assign w4523 = ( ~w2791 & w4511 ) | ( ~w2791 & w4517 ) | ( w4511 & w4517 ) ;
  assign w4524 = ~w4511 & w4523 ;
  assign w4525 = w4522 | w4524 ;
  assign w4526 = ( w2585 & w4519 ) | ( w2585 & ~w4525 ) | ( w4519 & ~w4525 ) ;
  assign w4527 = w2585 & w4526 ;
  assign w4528 = w4249 | w4254 ;
  assign w4529 = w4457 & ~w4528 ;
  assign w4530 = w4252 ^ w4529 ;
  assign w4531 = ( ~w2585 & w4519 ) | ( ~w2585 & w4525 ) | ( w4519 & w4525 ) ;
  assign w4532 = ~w4519 & w4531 ;
  assign w4533 = w4530 | w4532 ;
  assign w4534 = ( w2387 & w4527 ) | ( w2387 & ~w4533 ) | ( w4527 & ~w4533 ) ;
  assign w4535 = w2387 & w4534 ;
  assign w4536 = w4257 | w4262 ;
  assign w4537 = w4457 & ~w4536 ;
  assign w4538 = w4260 ^ w4537 ;
  assign w4539 = ( ~w2387 & w4527 ) | ( ~w2387 & w4533 ) | ( w4527 & w4533 ) ;
  assign w4540 = ~w4527 & w4539 ;
  assign w4541 = w4538 | w4540 ;
  assign w4542 = ( w2197 & w4535 ) | ( w2197 & ~w4541 ) | ( w4535 & ~w4541 ) ;
  assign w4543 = w2197 & w4542 ;
  assign w4544 = w4265 | w4270 ;
  assign w4545 = w4457 & ~w4544 ;
  assign w4546 = w4268 ^ w4545 ;
  assign w4547 = ( ~w2197 & w4535 ) | ( ~w2197 & w4541 ) | ( w4535 & w4541 ) ;
  assign w4548 = ~w4535 & w4547 ;
  assign w4549 = w4546 | w4548 ;
  assign w4550 = ( w2015 & w4543 ) | ( w2015 & ~w4549 ) | ( w4543 & ~w4549 ) ;
  assign w4551 = w2015 & w4550 ;
  assign w4552 = w4273 | w4278 ;
  assign w4553 = w4457 & ~w4552 ;
  assign w4554 = w4276 ^ w4553 ;
  assign w4555 = ( ~w2015 & w4543 ) | ( ~w2015 & w4549 ) | ( w4543 & w4549 ) ;
  assign w4556 = ~w4543 & w4555 ;
  assign w4557 = w4554 | w4556 ;
  assign w4558 = ( w1841 & w4551 ) | ( w1841 & ~w4557 ) | ( w4551 & ~w4557 ) ;
  assign w4559 = w1841 & w4558 ;
  assign w4560 = w4281 | w4286 ;
  assign w4561 = w4457 & ~w4560 ;
  assign w4562 = w4284 ^ w4561 ;
  assign w4563 = ( ~w1841 & w4551 ) | ( ~w1841 & w4557 ) | ( w4551 & w4557 ) ;
  assign w4564 = ~w4551 & w4563 ;
  assign w4565 = w4562 | w4564 ;
  assign w4566 = ( w1675 & w4559 ) | ( w1675 & ~w4565 ) | ( w4559 & ~w4565 ) ;
  assign w4567 = w1675 & w4566 ;
  assign w4568 = w4289 | w4294 ;
  assign w4569 = w4457 & ~w4568 ;
  assign w4570 = w4292 ^ w4569 ;
  assign w4571 = ( ~w1675 & w4559 ) | ( ~w1675 & w4565 ) | ( w4559 & w4565 ) ;
  assign w4572 = ~w4559 & w4571 ;
  assign w4573 = w4570 | w4572 ;
  assign w4574 = ( w1517 & w4567 ) | ( w1517 & ~w4573 ) | ( w4567 & ~w4573 ) ;
  assign w4575 = w1517 & w4574 ;
  assign w4576 = w4297 | w4302 ;
  assign w4577 = w4457 & ~w4576 ;
  assign w4578 = w4300 ^ w4577 ;
  assign w4579 = ( ~w1517 & w4567 ) | ( ~w1517 & w4573 ) | ( w4567 & w4573 ) ;
  assign w4580 = ~w4567 & w4579 ;
  assign w4581 = w4578 | w4580 ;
  assign w4582 = ( w1367 & w4575 ) | ( w1367 & ~w4581 ) | ( w4575 & ~w4581 ) ;
  assign w4583 = w1367 & w4582 ;
  assign w4584 = w4305 | w4310 ;
  assign w4585 = w4457 & ~w4584 ;
  assign w4586 = w4308 ^ w4585 ;
  assign w4587 = ( ~w1367 & w4575 ) | ( ~w1367 & w4581 ) | ( w4575 & w4581 ) ;
  assign w4588 = ~w4575 & w4587 ;
  assign w4589 = w4586 | w4588 ;
  assign w4590 = ( w1225 & w4583 ) | ( w1225 & ~w4589 ) | ( w4583 & ~w4589 ) ;
  assign w4591 = w1225 & w4590 ;
  assign w4592 = w4313 | w4318 ;
  assign w4593 = w4457 & ~w4592 ;
  assign w4594 = w4316 ^ w4593 ;
  assign w4595 = ( ~w1225 & w4583 ) | ( ~w1225 & w4589 ) | ( w4583 & w4589 ) ;
  assign w4596 = ~w4583 & w4595 ;
  assign w4597 = w4594 | w4596 ;
  assign w4598 = ( w1091 & w4591 ) | ( w1091 & ~w4597 ) | ( w4591 & ~w4597 ) ;
  assign w4599 = w1091 & w4598 ;
  assign w4600 = w4321 | w4326 ;
  assign w4601 = w4457 & ~w4600 ;
  assign w4602 = w4324 ^ w4601 ;
  assign w4603 = ( ~w1091 & w4591 ) | ( ~w1091 & w4597 ) | ( w4591 & w4597 ) ;
  assign w4604 = ~w4591 & w4603 ;
  assign w4605 = w4602 | w4604 ;
  assign w4606 = ( w965 & w4599 ) | ( w965 & ~w4605 ) | ( w4599 & ~w4605 ) ;
  assign w4607 = w965 & w4606 ;
  assign w4608 = w4329 | w4334 ;
  assign w4609 = w4457 & ~w4608 ;
  assign w4610 = w4332 ^ w4609 ;
  assign w4611 = ( ~w965 & w4599 ) | ( ~w965 & w4605 ) | ( w4599 & w4605 ) ;
  assign w4612 = ~w4599 & w4611 ;
  assign w4613 = w4610 | w4612 ;
  assign w4614 = ( w847 & w4607 ) | ( w847 & ~w4613 ) | ( w4607 & ~w4613 ) ;
  assign w4615 = w847 & w4614 ;
  assign w4616 = w4337 | w4342 ;
  assign w4617 = w4457 & ~w4616 ;
  assign w4618 = w4340 ^ w4617 ;
  assign w4619 = ( ~w847 & w4607 ) | ( ~w847 & w4613 ) | ( w4607 & w4613 ) ;
  assign w4620 = ~w4607 & w4619 ;
  assign w4621 = w4618 | w4620 ;
  assign w4622 = ( w737 & w4615 ) | ( w737 & ~w4621 ) | ( w4615 & ~w4621 ) ;
  assign w4623 = w737 & w4622 ;
  assign w4624 = w4345 | w4350 ;
  assign w4625 = w4457 & ~w4624 ;
  assign w4626 = w4348 ^ w4625 ;
  assign w4627 = ( ~w737 & w4615 ) | ( ~w737 & w4621 ) | ( w4615 & w4621 ) ;
  assign w4628 = ~w4615 & w4627 ;
  assign w4629 = w4626 | w4628 ;
  assign w4630 = ( w635 & w4623 ) | ( w635 & ~w4629 ) | ( w4623 & ~w4629 ) ;
  assign w4631 = w635 & w4630 ;
  assign w4632 = w4353 | w4358 ;
  assign w4633 = w4457 & ~w4632 ;
  assign w4634 = w4356 ^ w4633 ;
  assign w4635 = ( ~w635 & w4623 ) | ( ~w635 & w4629 ) | ( w4623 & w4629 ) ;
  assign w4636 = ~w4623 & w4635 ;
  assign w4637 = w4634 | w4636 ;
  assign w4638 = ( w541 & w4631 ) | ( w541 & ~w4637 ) | ( w4631 & ~w4637 ) ;
  assign w4639 = w541 & w4638 ;
  assign w4640 = w4361 | w4366 ;
  assign w4641 = w4457 & ~w4640 ;
  assign w4642 = w4364 ^ w4641 ;
  assign w4643 = ( ~w541 & w4631 ) | ( ~w541 & w4637 ) | ( w4631 & w4637 ) ;
  assign w4644 = ~w4631 & w4643 ;
  assign w4645 = w4642 | w4644 ;
  assign w4646 = ( w455 & w4639 ) | ( w455 & ~w4645 ) | ( w4639 & ~w4645 ) ;
  assign w4647 = w455 & w4646 ;
  assign w4648 = w4369 | w4374 ;
  assign w4649 = w4457 & ~w4648 ;
  assign w4650 = w4372 ^ w4649 ;
  assign w4651 = ( ~w455 & w4639 ) | ( ~w455 & w4645 ) | ( w4639 & w4645 ) ;
  assign w4652 = ~w4639 & w4651 ;
  assign w4653 = w4650 | w4652 ;
  assign w4654 = ( w377 & w4647 ) | ( w377 & ~w4653 ) | ( w4647 & ~w4653 ) ;
  assign w4655 = w377 & w4654 ;
  assign w4656 = w4377 | w4382 ;
  assign w4657 = w4457 & ~w4656 ;
  assign w4658 = w4380 ^ w4657 ;
  assign w4659 = ( ~w377 & w4647 ) | ( ~w377 & w4653 ) | ( w4647 & w4653 ) ;
  assign w4660 = ~w4647 & w4659 ;
  assign w4661 = w4658 | w4660 ;
  assign w4662 = ( w307 & w4655 ) | ( w307 & ~w4661 ) | ( w4655 & ~w4661 ) ;
  assign w4663 = w307 & w4662 ;
  assign w4664 = w4385 | w4390 ;
  assign w4665 = w4457 & ~w4664 ;
  assign w4666 = w4388 ^ w4665 ;
  assign w4667 = ( ~w307 & w4655 ) | ( ~w307 & w4661 ) | ( w4655 & w4661 ) ;
  assign w4668 = ~w4655 & w4667 ;
  assign w4669 = w4666 | w4668 ;
  assign w4670 = ( w246 & w4663 ) | ( w246 & ~w4669 ) | ( w4663 & ~w4669 ) ;
  assign w4671 = w246 & w4670 ;
  assign w4672 = w4393 | w4398 ;
  assign w4673 = w4457 & ~w4672 ;
  assign w4674 = w4396 ^ w4673 ;
  assign w4675 = ( ~w246 & w4663 ) | ( ~w246 & w4669 ) | ( w4663 & w4669 ) ;
  assign w4676 = ~w4663 & w4675 ;
  assign w4677 = w4674 | w4676 ;
  assign w4678 = ( w185 & w4671 ) | ( w185 & ~w4677 ) | ( w4671 & ~w4677 ) ;
  assign w4679 = w185 & w4678 ;
  assign w4680 = w4401 | w4406 ;
  assign w4681 = w4457 & ~w4680 ;
  assign w4682 = w4404 ^ w4681 ;
  assign w4683 = ( ~w185 & w4671 ) | ( ~w185 & w4677 ) | ( w4671 & w4677 ) ;
  assign w4684 = ~w4671 & w4683 ;
  assign w4685 = w4682 | w4684 ;
  assign w4686 = ( w145 & w4679 ) | ( w145 & ~w4685 ) | ( w4679 & ~w4685 ) ;
  assign w4687 = w145 & w4686 ;
  assign w4688 = w4409 | w4414 ;
  assign w4689 = w4457 & ~w4688 ;
  assign w4690 = w4412 ^ w4689 ;
  assign w4691 = ( ~w145 & w4679 ) | ( ~w145 & w4685 ) | ( w4679 & w4685 ) ;
  assign w4692 = ~w4679 & w4691 ;
  assign w4693 = w4690 | w4692 ;
  assign w4694 = ( w132 & w4687 ) | ( w132 & ~w4693 ) | ( w4687 & ~w4693 ) ;
  assign w4695 = w132 & w4694 ;
  assign w4696 = w4417 | w4422 ;
  assign w4697 = w4457 & ~w4696 ;
  assign w4698 = w4420 ^ w4697 ;
  assign w4699 = ( ~w132 & w4687 ) | ( ~w132 & w4693 ) | ( w4687 & w4693 ) ;
  assign w4700 = ~w4687 & w4699 ;
  assign w4701 = w4698 | w4700 ;
  assign w4702 = ~w4695 & w4701 ;
  assign w4703 = w4425 | w4430 ;
  assign w4704 = w4457 & ~w4703 ;
  assign w4705 = w4428 ^ w4704 ;
  assign w4706 = ( ~w4443 & w4702 ) | ( ~w4443 & w4705 ) | ( w4702 & w4705 ) ;
  assign w4707 = w4432 & ~w4706 ;
  assign w4708 = ~w4435 & w4457 ;
  assign w4709 = ( w4706 & ~w4707 ) | ( w4706 & w4708 ) | ( ~w4707 & w4708 ) ;
  assign w4710 = w4443 | w4709 ;
  assign w4711 = ~w129 & w4710 ;
  assign w4712 = ( w4695 & w4701 ) | ( w4695 & w4705 ) | ( w4701 & w4705 ) ;
  assign w4713 = ~w4695 & w4712 ;
  assign w4714 = ( w129 & w4432 ) | ( w129 & w4435 ) | ( w4432 & w4435 ) ;
  assign w4715 = ( w4435 & ~w4457 ) | ( w4435 & w4714 ) | ( ~w4457 & w4714 ) ;
  assign w4716 = w4432 & w4715 ;
  assign w4717 = w4714 ^ w4716 ;
  assign w4718 = ( w4163 & w4165 ) | ( w4163 & w4195 ) | ( w4165 & w4195 ) ;
  assign w4719 = w4195 & ~w4718 ;
  assign w4720 = w4168 ^ w4719 ;
  assign w4721 = ( ~w4447 & w4454 ) | ( ~w4447 & w4720 ) | ( w4454 & w4720 ) ;
  assign w4722 = ~w4454 & w4721 ;
  assign w4723 = ( ~w4441 & w4443 ) | ( ~w4441 & w4722 ) | ( w4443 & w4722 ) ;
  assign w4724 = ~w4443 & w4723 ;
  assign w4725 = w4713 | w4724 ;
  assign w4726 = ( w4711 & ~w4713 ) | ( w4711 & w4717 ) | ( ~w4713 & w4717 ) ;
  assign w4727 = w4725 | w4726 ;
  assign w4728 = ( ~\pi063 & \pi064 ) | ( ~\pi063 & w4457 ) | ( \pi064 & w4457 ) ;
  assign w4729 = ( ~\pi062 & \pi064 ) | ( ~\pi062 & w4728 ) | ( \pi064 & w4728 ) ;
  assign w4730 = ( ~\pi064 & w4457 ) | ( ~\pi064 & w4727 ) | ( w4457 & w4727 ) ;
  assign w4731 = w4729 & w4730 ;
  assign w4732 = ( w4443 & w4447 ) | ( w4443 & ~w4454 ) | ( w4447 & ~w4454 ) ;
  assign w4733 = \pi063 & ~w4732 ;
  assign w4734 = \pi062 | \pi064 ;
  assign w4735 = ( ~w4732 & w4733 ) | ( ~w4732 & w4734 ) | ( w4733 & w4734 ) ;
  assign w4736 = ~w4454 & w4735 ;
  assign w4737 = ~w4441 & w4736 ;
  assign w4738 = ( \pi064 & w4727 ) | ( \pi064 & ~w4736 ) | ( w4727 & ~w4736 ) ;
  assign w4739 = w4737 & ~w4738 ;
  assign w4740 = ~\pi064 & w4727 ;
  assign w4741 = \pi065 ^ w4740 ;
  assign w4742 = w4739 | w4741 ;
  assign w4743 = ( w4195 & w4731 ) | ( w4195 & ~w4742 ) | ( w4731 & ~w4742 ) ;
  assign w4744 = w4195 & w4743 ;
  assign w4745 = ( ~w4195 & w4731 ) | ( ~w4195 & w4742 ) | ( w4731 & w4742 ) ;
  assign w4746 = ~w4731 & w4745 ;
  assign w4747 = w4457 & ~w4724 ;
  assign w4748 = ~w4713 & w4747 ;
  assign w4749 = ~w4726 & w4748 ;
  assign w4750 = \pi065 & w4727 ;
  assign w4751 = ( \pi064 & w4727 ) | ( \pi064 & ~w4750 ) | ( w4727 & ~w4750 ) ;
  assign w4752 = ( ~\pi064 & w4749 ) | ( ~\pi064 & w4751 ) | ( w4749 & w4751 ) ;
  assign w4753 = \pi066 ^ w4752 ;
  assign w4754 = w4746 | w4753 ;
  assign w4755 = ( w3941 & w4744 ) | ( w3941 & ~w4754 ) | ( w4744 & ~w4754 ) ;
  assign w4756 = w3941 & w4755 ;
  assign w4757 = ( w4461 & ~w4469 ) | ( w4461 & w4727 ) | ( ~w4469 & w4727 ) ;
  assign w4758 = ~w4461 & w4757 ;
  assign w4759 = \pi067 ^ w4758 ;
  assign w4760 = w4470 ^ w4759 ;
  assign w4761 = ( ~w3941 & w4744 ) | ( ~w3941 & w4754 ) | ( w4744 & w4754 ) ;
  assign w4762 = ~w4744 & w4761 ;
  assign w4763 = w4760 | w4762 ;
  assign w4764 = ( w3695 & w4756 ) | ( w3695 & ~w4763 ) | ( w4756 & ~w4763 ) ;
  assign w4765 = w3695 & w4764 ;
  assign w4766 = w4474 | w4476 ;
  assign w4767 = w4727 & ~w4766 ;
  assign w4768 = w4483 ^ w4767 ;
  assign w4769 = ( ~w3695 & w4756 ) | ( ~w3695 & w4763 ) | ( w4756 & w4763 ) ;
  assign w4770 = ~w4756 & w4769 ;
  assign w4771 = w4768 | w4770 ;
  assign w4772 = ( w3457 & w4765 ) | ( w3457 & ~w4771 ) | ( w4765 & ~w4771 ) ;
  assign w4773 = w3457 & w4772 ;
  assign w4774 = w4486 | w4492 ;
  assign w4775 = w4727 & ~w4774 ;
  assign w4776 = w4490 ^ w4775 ;
  assign w4777 = ( ~w3457 & w4765 ) | ( ~w3457 & w4771 ) | ( w4765 & w4771 ) ;
  assign w4778 = ~w4765 & w4777 ;
  assign w4779 = w4776 | w4778 ;
  assign w4780 = ( w3227 & w4773 ) | ( w3227 & ~w4779 ) | ( w4773 & ~w4779 ) ;
  assign w4781 = w3227 & w4780 ;
  assign w4782 = w4495 | w4500 ;
  assign w4783 = w4727 & ~w4782 ;
  assign w4784 = w4498 ^ w4783 ;
  assign w4785 = ( ~w3227 & w4773 ) | ( ~w3227 & w4779 ) | ( w4773 & w4779 ) ;
  assign w4786 = ~w4773 & w4785 ;
  assign w4787 = w4784 | w4786 ;
  assign w4788 = ( w3005 & w4781 ) | ( w3005 & ~w4787 ) | ( w4781 & ~w4787 ) ;
  assign w4789 = w3005 & w4788 ;
  assign w4790 = w4503 | w4508 ;
  assign w4791 = w4727 & ~w4790 ;
  assign w4792 = w4506 ^ w4791 ;
  assign w4793 = ( ~w3005 & w4781 ) | ( ~w3005 & w4787 ) | ( w4781 & w4787 ) ;
  assign w4794 = ~w4781 & w4793 ;
  assign w4795 = w4792 | w4794 ;
  assign w4796 = ( w2791 & w4789 ) | ( w2791 & ~w4795 ) | ( w4789 & ~w4795 ) ;
  assign w4797 = w2791 & w4796 ;
  assign w4798 = w4511 | w4516 ;
  assign w4799 = w4727 & ~w4798 ;
  assign w4800 = w4514 ^ w4799 ;
  assign w4801 = ( ~w2791 & w4789 ) | ( ~w2791 & w4795 ) | ( w4789 & w4795 ) ;
  assign w4802 = ~w4789 & w4801 ;
  assign w4803 = w4800 | w4802 ;
  assign w4804 = ( w2585 & w4797 ) | ( w2585 & ~w4803 ) | ( w4797 & ~w4803 ) ;
  assign w4805 = w2585 & w4804 ;
  assign w4806 = w4519 | w4524 ;
  assign w4807 = w4727 & ~w4806 ;
  assign w4808 = w4522 ^ w4807 ;
  assign w4809 = ( ~w2585 & w4797 ) | ( ~w2585 & w4803 ) | ( w4797 & w4803 ) ;
  assign w4810 = ~w4797 & w4809 ;
  assign w4811 = w4808 | w4810 ;
  assign w4812 = ( w2387 & w4805 ) | ( w2387 & ~w4811 ) | ( w4805 & ~w4811 ) ;
  assign w4813 = w2387 & w4812 ;
  assign w4814 = w4527 | w4532 ;
  assign w4815 = w4727 & ~w4814 ;
  assign w4816 = w4530 ^ w4815 ;
  assign w4817 = ( ~w2387 & w4805 ) | ( ~w2387 & w4811 ) | ( w4805 & w4811 ) ;
  assign w4818 = ~w4805 & w4817 ;
  assign w4819 = w4816 | w4818 ;
  assign w4820 = ( w2197 & w4813 ) | ( w2197 & ~w4819 ) | ( w4813 & ~w4819 ) ;
  assign w4821 = w2197 & w4820 ;
  assign w4822 = w4535 | w4540 ;
  assign w4823 = w4727 & ~w4822 ;
  assign w4824 = w4538 ^ w4823 ;
  assign w4825 = ( ~w2197 & w4813 ) | ( ~w2197 & w4819 ) | ( w4813 & w4819 ) ;
  assign w4826 = ~w4813 & w4825 ;
  assign w4827 = w4824 | w4826 ;
  assign w4828 = ( w2015 & w4821 ) | ( w2015 & ~w4827 ) | ( w4821 & ~w4827 ) ;
  assign w4829 = w2015 & w4828 ;
  assign w4830 = w4543 | w4548 ;
  assign w4831 = w4727 & ~w4830 ;
  assign w4832 = w4546 ^ w4831 ;
  assign w4833 = ( ~w2015 & w4821 ) | ( ~w2015 & w4827 ) | ( w4821 & w4827 ) ;
  assign w4834 = ~w4821 & w4833 ;
  assign w4835 = w4832 | w4834 ;
  assign w4836 = ( w1841 & w4829 ) | ( w1841 & ~w4835 ) | ( w4829 & ~w4835 ) ;
  assign w4837 = w1841 & w4836 ;
  assign w4838 = w4551 | w4556 ;
  assign w4839 = w4727 & ~w4838 ;
  assign w4840 = w4554 ^ w4839 ;
  assign w4841 = ( ~w1841 & w4829 ) | ( ~w1841 & w4835 ) | ( w4829 & w4835 ) ;
  assign w4842 = ~w4829 & w4841 ;
  assign w4843 = w4840 | w4842 ;
  assign w4844 = ( w1675 & w4837 ) | ( w1675 & ~w4843 ) | ( w4837 & ~w4843 ) ;
  assign w4845 = w1675 & w4844 ;
  assign w4846 = w4559 | w4564 ;
  assign w4847 = w4727 & ~w4846 ;
  assign w4848 = w4562 ^ w4847 ;
  assign w4849 = ( ~w1675 & w4837 ) | ( ~w1675 & w4843 ) | ( w4837 & w4843 ) ;
  assign w4850 = ~w4837 & w4849 ;
  assign w4851 = w4848 | w4850 ;
  assign w4852 = ( w1517 & w4845 ) | ( w1517 & ~w4851 ) | ( w4845 & ~w4851 ) ;
  assign w4853 = w1517 & w4852 ;
  assign w4854 = w4567 | w4572 ;
  assign w4855 = w4727 & ~w4854 ;
  assign w4856 = w4570 ^ w4855 ;
  assign w4857 = ( ~w1517 & w4845 ) | ( ~w1517 & w4851 ) | ( w4845 & w4851 ) ;
  assign w4858 = ~w4845 & w4857 ;
  assign w4859 = w4856 | w4858 ;
  assign w4860 = ( w1367 & w4853 ) | ( w1367 & ~w4859 ) | ( w4853 & ~w4859 ) ;
  assign w4861 = w1367 & w4860 ;
  assign w4862 = w4575 | w4580 ;
  assign w4863 = w4727 & ~w4862 ;
  assign w4864 = w4578 ^ w4863 ;
  assign w4865 = ( ~w1367 & w4853 ) | ( ~w1367 & w4859 ) | ( w4853 & w4859 ) ;
  assign w4866 = ~w4853 & w4865 ;
  assign w4867 = w4864 | w4866 ;
  assign w4868 = ( w1225 & w4861 ) | ( w1225 & ~w4867 ) | ( w4861 & ~w4867 ) ;
  assign w4869 = w1225 & w4868 ;
  assign w4870 = w4583 | w4588 ;
  assign w4871 = w4727 & ~w4870 ;
  assign w4872 = w4586 ^ w4871 ;
  assign w4873 = ( ~w1225 & w4861 ) | ( ~w1225 & w4867 ) | ( w4861 & w4867 ) ;
  assign w4874 = ~w4861 & w4873 ;
  assign w4875 = w4872 | w4874 ;
  assign w4876 = ( w1091 & w4869 ) | ( w1091 & ~w4875 ) | ( w4869 & ~w4875 ) ;
  assign w4877 = w1091 & w4876 ;
  assign w4878 = w4591 | w4596 ;
  assign w4879 = w4727 & ~w4878 ;
  assign w4880 = w4594 ^ w4879 ;
  assign w4881 = ( ~w1091 & w4869 ) | ( ~w1091 & w4875 ) | ( w4869 & w4875 ) ;
  assign w4882 = ~w4869 & w4881 ;
  assign w4883 = w4880 | w4882 ;
  assign w4884 = ( w965 & w4877 ) | ( w965 & ~w4883 ) | ( w4877 & ~w4883 ) ;
  assign w4885 = w965 & w4884 ;
  assign w4886 = w4599 | w4604 ;
  assign w4887 = w4727 & ~w4886 ;
  assign w4888 = w4602 ^ w4887 ;
  assign w4889 = ( ~w965 & w4877 ) | ( ~w965 & w4883 ) | ( w4877 & w4883 ) ;
  assign w4890 = ~w4877 & w4889 ;
  assign w4891 = w4888 | w4890 ;
  assign w4892 = ( w847 & w4885 ) | ( w847 & ~w4891 ) | ( w4885 & ~w4891 ) ;
  assign w4893 = w847 & w4892 ;
  assign w4894 = w4607 | w4612 ;
  assign w4895 = w4727 & ~w4894 ;
  assign w4896 = w4610 ^ w4895 ;
  assign w4897 = ( ~w847 & w4885 ) | ( ~w847 & w4891 ) | ( w4885 & w4891 ) ;
  assign w4898 = ~w4885 & w4897 ;
  assign w4899 = w4896 | w4898 ;
  assign w4900 = ( w737 & w4893 ) | ( w737 & ~w4899 ) | ( w4893 & ~w4899 ) ;
  assign w4901 = w737 & w4900 ;
  assign w4902 = w4615 | w4620 ;
  assign w4903 = w4727 & ~w4902 ;
  assign w4904 = w4618 ^ w4903 ;
  assign w4905 = ( ~w737 & w4893 ) | ( ~w737 & w4899 ) | ( w4893 & w4899 ) ;
  assign w4906 = ~w4893 & w4905 ;
  assign w4907 = w4904 | w4906 ;
  assign w4908 = ( w635 & w4901 ) | ( w635 & ~w4907 ) | ( w4901 & ~w4907 ) ;
  assign w4909 = w635 & w4908 ;
  assign w4910 = w4623 | w4628 ;
  assign w4911 = w4727 & ~w4910 ;
  assign w4912 = w4626 ^ w4911 ;
  assign w4913 = ( ~w635 & w4901 ) | ( ~w635 & w4907 ) | ( w4901 & w4907 ) ;
  assign w4914 = ~w4901 & w4913 ;
  assign w4915 = w4912 | w4914 ;
  assign w4916 = ( w541 & w4909 ) | ( w541 & ~w4915 ) | ( w4909 & ~w4915 ) ;
  assign w4917 = w541 & w4916 ;
  assign w4918 = w4631 | w4636 ;
  assign w4919 = w4727 & ~w4918 ;
  assign w4920 = w4634 ^ w4919 ;
  assign w4921 = ( ~w541 & w4909 ) | ( ~w541 & w4915 ) | ( w4909 & w4915 ) ;
  assign w4922 = ~w4909 & w4921 ;
  assign w4923 = w4920 | w4922 ;
  assign w4924 = ( w455 & w4917 ) | ( w455 & ~w4923 ) | ( w4917 & ~w4923 ) ;
  assign w4925 = w455 & w4924 ;
  assign w4926 = w4639 | w4644 ;
  assign w4927 = w4727 & ~w4926 ;
  assign w4928 = w4642 ^ w4927 ;
  assign w4929 = ( ~w455 & w4917 ) | ( ~w455 & w4923 ) | ( w4917 & w4923 ) ;
  assign w4930 = ~w4917 & w4929 ;
  assign w4931 = w4928 | w4930 ;
  assign w4932 = ( w377 & w4925 ) | ( w377 & ~w4931 ) | ( w4925 & ~w4931 ) ;
  assign w4933 = w377 & w4932 ;
  assign w4934 = w4647 | w4652 ;
  assign w4935 = w4727 & ~w4934 ;
  assign w4936 = w4650 ^ w4935 ;
  assign w4937 = ( ~w377 & w4925 ) | ( ~w377 & w4931 ) | ( w4925 & w4931 ) ;
  assign w4938 = ~w4925 & w4937 ;
  assign w4939 = w4936 | w4938 ;
  assign w4940 = ( w307 & w4933 ) | ( w307 & ~w4939 ) | ( w4933 & ~w4939 ) ;
  assign w4941 = w307 & w4940 ;
  assign w4942 = w4655 | w4660 ;
  assign w4943 = w4727 & ~w4942 ;
  assign w4944 = w4658 ^ w4943 ;
  assign w4945 = ( ~w307 & w4933 ) | ( ~w307 & w4939 ) | ( w4933 & w4939 ) ;
  assign w4946 = ~w4933 & w4945 ;
  assign w4947 = w4944 | w4946 ;
  assign w4948 = ( w246 & w4941 ) | ( w246 & ~w4947 ) | ( w4941 & ~w4947 ) ;
  assign w4949 = w246 & w4948 ;
  assign w4950 = w4663 | w4668 ;
  assign w4951 = w4727 & ~w4950 ;
  assign w4952 = w4666 ^ w4951 ;
  assign w4953 = ( ~w246 & w4941 ) | ( ~w246 & w4947 ) | ( w4941 & w4947 ) ;
  assign w4954 = ~w4941 & w4953 ;
  assign w4955 = w4952 | w4954 ;
  assign w4956 = ( w185 & w4949 ) | ( w185 & ~w4955 ) | ( w4949 & ~w4955 ) ;
  assign w4957 = w185 & w4956 ;
  assign w4958 = w4671 | w4676 ;
  assign w4959 = w4727 & ~w4958 ;
  assign w4960 = w4674 ^ w4959 ;
  assign w4961 = ( ~w185 & w4949 ) | ( ~w185 & w4955 ) | ( w4949 & w4955 ) ;
  assign w4962 = ~w4949 & w4961 ;
  assign w4963 = w4960 | w4962 ;
  assign w4964 = ( w145 & w4957 ) | ( w145 & ~w4963 ) | ( w4957 & ~w4963 ) ;
  assign w4965 = w145 & w4964 ;
  assign w4966 = w4679 | w4684 ;
  assign w4967 = w4727 & ~w4966 ;
  assign w4968 = w4682 ^ w4967 ;
  assign w4969 = ( ~w145 & w4957 ) | ( ~w145 & w4963 ) | ( w4957 & w4963 ) ;
  assign w4970 = ~w4957 & w4969 ;
  assign w4971 = w4968 | w4970 ;
  assign w4972 = ( w132 & w4965 ) | ( w132 & ~w4971 ) | ( w4965 & ~w4971 ) ;
  assign w4973 = w132 & w4972 ;
  assign w4974 = w4687 | w4692 ;
  assign w4975 = w4727 & ~w4974 ;
  assign w4976 = w4690 ^ w4975 ;
  assign w4977 = ( ~w132 & w4965 ) | ( ~w132 & w4971 ) | ( w4965 & w4971 ) ;
  assign w4978 = ~w4965 & w4977 ;
  assign w4979 = w4976 | w4978 ;
  assign w4980 = ~w4973 & w4979 ;
  assign w4981 = w4695 | w4700 ;
  assign w4982 = w4727 & ~w4981 ;
  assign w4983 = w4698 ^ w4982 ;
  assign w4984 = ( ~w4713 & w4980 ) | ( ~w4713 & w4983 ) | ( w4980 & w4983 ) ;
  assign w4985 = w4702 & ~w4984 ;
  assign w4986 = ~w4705 & w4727 ;
  assign w4987 = ( w4984 & ~w4985 ) | ( w4984 & w4986 ) | ( ~w4985 & w4986 ) ;
  assign w4988 = w4713 | w4987 ;
  assign w4989 = ~w129 & w4988 ;
  assign w4990 = ( w4973 & w4979 ) | ( w4973 & w4983 ) | ( w4979 & w4983 ) ;
  assign w4991 = ~w4973 & w4990 ;
  assign w4992 = ( w129 & w4702 ) | ( w129 & w4705 ) | ( w4702 & w4705 ) ;
  assign w4993 = ( w4705 & ~w4727 ) | ( w4705 & w4992 ) | ( ~w4727 & w4992 ) ;
  assign w4994 = w4702 & w4993 ;
  assign w4995 = w4992 ^ w4994 ;
  assign w4996 = ( w4425 & w4430 ) | ( w4425 & w4457 ) | ( w4430 & w4457 ) ;
  assign w4997 = w4457 & ~w4996 ;
  assign w4998 = w4428 ^ w4997 ;
  assign w4999 = ( ~w4717 & w4724 ) | ( ~w4717 & w4998 ) | ( w4724 & w4998 ) ;
  assign w5000 = ~w4724 & w4999 ;
  assign w5001 = ( ~w4711 & w4713 ) | ( ~w4711 & w5000 ) | ( w4713 & w5000 ) ;
  assign w5002 = ~w4713 & w5001 ;
  assign w5003 = w4991 | w5002 ;
  assign w5004 = ( w4989 & ~w4991 ) | ( w4989 & w4995 ) | ( ~w4991 & w4995 ) ;
  assign w5005 = w5003 | w5004 ;
  assign w5006 = ( ~\pi061 & \pi062 ) | ( ~\pi061 & w4727 ) | ( \pi062 & w4727 ) ;
  assign w5007 = ( ~\pi060 & \pi062 ) | ( ~\pi060 & w5006 ) | ( \pi062 & w5006 ) ;
  assign w5008 = ( ~\pi062 & w4727 ) | ( ~\pi062 & w5005 ) | ( w4727 & w5005 ) ;
  assign w5009 = w5007 & w5008 ;
  assign w5010 = ( w4713 & w4717 ) | ( w4713 & ~w4724 ) | ( w4717 & ~w4724 ) ;
  assign w5011 = \pi061 & ~w5010 ;
  assign w5012 = \pi060 | \pi062 ;
  assign w5013 = ( ~w5010 & w5011 ) | ( ~w5010 & w5012 ) | ( w5011 & w5012 ) ;
  assign w5014 = ~w4724 & w5013 ;
  assign w5015 = ~w4711 & w5014 ;
  assign w5016 = ( \pi062 & w5005 ) | ( \pi062 & ~w5014 ) | ( w5005 & ~w5014 ) ;
  assign w5017 = w5015 & ~w5016 ;
  assign w5018 = ~\pi062 & w5005 ;
  assign w5019 = \pi063 ^ w5018 ;
  assign w5020 = w5017 | w5019 ;
  assign w5021 = ( w4457 & w5009 ) | ( w4457 & ~w5020 ) | ( w5009 & ~w5020 ) ;
  assign w5022 = w4457 & w5021 ;
  assign w5023 = ( ~w4457 & w5009 ) | ( ~w4457 & w5020 ) | ( w5009 & w5020 ) ;
  assign w5024 = ~w5009 & w5023 ;
  assign w5025 = w4727 & ~w5002 ;
  assign w5026 = ~w4991 & w5025 ;
  assign w5027 = ~w5004 & w5026 ;
  assign w5028 = \pi063 & w5005 ;
  assign w5029 = ( \pi062 & w5005 ) | ( \pi062 & ~w5028 ) | ( w5005 & ~w5028 ) ;
  assign w5030 = ( ~\pi062 & w5027 ) | ( ~\pi062 & w5029 ) | ( w5027 & w5029 ) ;
  assign w5031 = \pi064 ^ w5030 ;
  assign w5032 = w5024 | w5031 ;
  assign w5033 = ( w4195 & w5022 ) | ( w4195 & ~w5032 ) | ( w5022 & ~w5032 ) ;
  assign w5034 = w4195 & w5033 ;
  assign w5035 = ( ~w4195 & w5022 ) | ( ~w4195 & w5032 ) | ( w5022 & w5032 ) ;
  assign w5036 = ~w5022 & w5035 ;
  assign w5037 = ( w4731 & ~w4739 ) | ( w4731 & w5005 ) | ( ~w4739 & w5005 ) ;
  assign w5038 = ~w4731 & w5037 ;
  assign w5039 = \pi065 ^ w5038 ;
  assign w5040 = w4740 ^ w5039 ;
  assign w5041 = w5036 | w5040 ;
  assign w5042 = ( w3941 & w5034 ) | ( w3941 & ~w5041 ) | ( w5034 & ~w5041 ) ;
  assign w5043 = w3941 & w5042 ;
  assign w5044 = w4744 | w4746 ;
  assign w5045 = w5005 & ~w5044 ;
  assign w5046 = w4753 ^ w5045 ;
  assign w5047 = ( ~w3941 & w5034 ) | ( ~w3941 & w5041 ) | ( w5034 & w5041 ) ;
  assign w5048 = ~w5034 & w5047 ;
  assign w5049 = w5046 | w5048 ;
  assign w5050 = ( w3695 & w5043 ) | ( w3695 & ~w5049 ) | ( w5043 & ~w5049 ) ;
  assign w5051 = w3695 & w5050 ;
  assign w5052 = w4756 | w4762 ;
  assign w5053 = w5005 & ~w5052 ;
  assign w5054 = w4760 ^ w5053 ;
  assign w5055 = ( ~w3695 & w5043 ) | ( ~w3695 & w5049 ) | ( w5043 & w5049 ) ;
  assign w5056 = ~w5043 & w5055 ;
  assign w5057 = w5054 | w5056 ;
  assign w5058 = ( w3457 & w5051 ) | ( w3457 & ~w5057 ) | ( w5051 & ~w5057 ) ;
  assign w5059 = w3457 & w5058 ;
  assign w5060 = w4765 | w4770 ;
  assign w5061 = w5005 & ~w5060 ;
  assign w5062 = w4768 ^ w5061 ;
  assign w5063 = ( ~w3457 & w5051 ) | ( ~w3457 & w5057 ) | ( w5051 & w5057 ) ;
  assign w5064 = ~w5051 & w5063 ;
  assign w5065 = w5062 | w5064 ;
  assign w5066 = ( w3227 & w5059 ) | ( w3227 & ~w5065 ) | ( w5059 & ~w5065 ) ;
  assign w5067 = w3227 & w5066 ;
  assign w5068 = w4773 | w4778 ;
  assign w5069 = w5005 & ~w5068 ;
  assign w5070 = w4776 ^ w5069 ;
  assign w5071 = ( ~w3227 & w5059 ) | ( ~w3227 & w5065 ) | ( w5059 & w5065 ) ;
  assign w5072 = ~w5059 & w5071 ;
  assign w5073 = w5070 | w5072 ;
  assign w5074 = ( w3005 & w5067 ) | ( w3005 & ~w5073 ) | ( w5067 & ~w5073 ) ;
  assign w5075 = w3005 & w5074 ;
  assign w5076 = w4781 | w4786 ;
  assign w5077 = w5005 & ~w5076 ;
  assign w5078 = w4784 ^ w5077 ;
  assign w5079 = ( ~w3005 & w5067 ) | ( ~w3005 & w5073 ) | ( w5067 & w5073 ) ;
  assign w5080 = ~w5067 & w5079 ;
  assign w5081 = w5078 | w5080 ;
  assign w5082 = ( w2791 & w5075 ) | ( w2791 & ~w5081 ) | ( w5075 & ~w5081 ) ;
  assign w5083 = w2791 & w5082 ;
  assign w5084 = w4789 | w4794 ;
  assign w5085 = w5005 & ~w5084 ;
  assign w5086 = w4792 ^ w5085 ;
  assign w5087 = ( ~w2791 & w5075 ) | ( ~w2791 & w5081 ) | ( w5075 & w5081 ) ;
  assign w5088 = ~w5075 & w5087 ;
  assign w5089 = w5086 | w5088 ;
  assign w5090 = ( w2585 & w5083 ) | ( w2585 & ~w5089 ) | ( w5083 & ~w5089 ) ;
  assign w5091 = w2585 & w5090 ;
  assign w5092 = w4797 | w4802 ;
  assign w5093 = w5005 & ~w5092 ;
  assign w5094 = w4800 ^ w5093 ;
  assign w5095 = ( ~w2585 & w5083 ) | ( ~w2585 & w5089 ) | ( w5083 & w5089 ) ;
  assign w5096 = ~w5083 & w5095 ;
  assign w5097 = w5094 | w5096 ;
  assign w5098 = ( w2387 & w5091 ) | ( w2387 & ~w5097 ) | ( w5091 & ~w5097 ) ;
  assign w5099 = w2387 & w5098 ;
  assign w5100 = w4805 | w4810 ;
  assign w5101 = w5005 & ~w5100 ;
  assign w5102 = w4808 ^ w5101 ;
  assign w5103 = ( ~w2387 & w5091 ) | ( ~w2387 & w5097 ) | ( w5091 & w5097 ) ;
  assign w5104 = ~w5091 & w5103 ;
  assign w5105 = w5102 | w5104 ;
  assign w5106 = ( w2197 & w5099 ) | ( w2197 & ~w5105 ) | ( w5099 & ~w5105 ) ;
  assign w5107 = w2197 & w5106 ;
  assign w5108 = w4813 | w4818 ;
  assign w5109 = w5005 & ~w5108 ;
  assign w5110 = w4816 ^ w5109 ;
  assign w5111 = ( ~w2197 & w5099 ) | ( ~w2197 & w5105 ) | ( w5099 & w5105 ) ;
  assign w5112 = ~w5099 & w5111 ;
  assign w5113 = w5110 | w5112 ;
  assign w5114 = ( w2015 & w5107 ) | ( w2015 & ~w5113 ) | ( w5107 & ~w5113 ) ;
  assign w5115 = w2015 & w5114 ;
  assign w5116 = w4821 | w4826 ;
  assign w5117 = w5005 & ~w5116 ;
  assign w5118 = w4824 ^ w5117 ;
  assign w5119 = ( ~w2015 & w5107 ) | ( ~w2015 & w5113 ) | ( w5107 & w5113 ) ;
  assign w5120 = ~w5107 & w5119 ;
  assign w5121 = w5118 | w5120 ;
  assign w5122 = ( w1841 & w5115 ) | ( w1841 & ~w5121 ) | ( w5115 & ~w5121 ) ;
  assign w5123 = w1841 & w5122 ;
  assign w5124 = w4829 | w4834 ;
  assign w5125 = w5005 & ~w5124 ;
  assign w5126 = w4832 ^ w5125 ;
  assign w5127 = ( ~w1841 & w5115 ) | ( ~w1841 & w5121 ) | ( w5115 & w5121 ) ;
  assign w5128 = ~w5115 & w5127 ;
  assign w5129 = w5126 | w5128 ;
  assign w5130 = ( w1675 & w5123 ) | ( w1675 & ~w5129 ) | ( w5123 & ~w5129 ) ;
  assign w5131 = w1675 & w5130 ;
  assign w5132 = w4837 | w4842 ;
  assign w5133 = w5005 & ~w5132 ;
  assign w5134 = w4840 ^ w5133 ;
  assign w5135 = ( ~w1675 & w5123 ) | ( ~w1675 & w5129 ) | ( w5123 & w5129 ) ;
  assign w5136 = ~w5123 & w5135 ;
  assign w5137 = w5134 | w5136 ;
  assign w5138 = ( w1517 & w5131 ) | ( w1517 & ~w5137 ) | ( w5131 & ~w5137 ) ;
  assign w5139 = w1517 & w5138 ;
  assign w5140 = w4845 | w4850 ;
  assign w5141 = w5005 & ~w5140 ;
  assign w5142 = w4848 ^ w5141 ;
  assign w5143 = ( ~w1517 & w5131 ) | ( ~w1517 & w5137 ) | ( w5131 & w5137 ) ;
  assign w5144 = ~w5131 & w5143 ;
  assign w5145 = w5142 | w5144 ;
  assign w5146 = ( w1367 & w5139 ) | ( w1367 & ~w5145 ) | ( w5139 & ~w5145 ) ;
  assign w5147 = w1367 & w5146 ;
  assign w5148 = w4853 | w4858 ;
  assign w5149 = w5005 & ~w5148 ;
  assign w5150 = w4856 ^ w5149 ;
  assign w5151 = ( ~w1367 & w5139 ) | ( ~w1367 & w5145 ) | ( w5139 & w5145 ) ;
  assign w5152 = ~w5139 & w5151 ;
  assign w5153 = w5150 | w5152 ;
  assign w5154 = ( w1225 & w5147 ) | ( w1225 & ~w5153 ) | ( w5147 & ~w5153 ) ;
  assign w5155 = w1225 & w5154 ;
  assign w5156 = w4861 | w4866 ;
  assign w5157 = w5005 & ~w5156 ;
  assign w5158 = w4864 ^ w5157 ;
  assign w5159 = ( ~w1225 & w5147 ) | ( ~w1225 & w5153 ) | ( w5147 & w5153 ) ;
  assign w5160 = ~w5147 & w5159 ;
  assign w5161 = w5158 | w5160 ;
  assign w5162 = ( w1091 & w5155 ) | ( w1091 & ~w5161 ) | ( w5155 & ~w5161 ) ;
  assign w5163 = w1091 & w5162 ;
  assign w5164 = w4869 | w4874 ;
  assign w5165 = w5005 & ~w5164 ;
  assign w5166 = w4872 ^ w5165 ;
  assign w5167 = ( ~w1091 & w5155 ) | ( ~w1091 & w5161 ) | ( w5155 & w5161 ) ;
  assign w5168 = ~w5155 & w5167 ;
  assign w5169 = w5166 | w5168 ;
  assign w5170 = ( w965 & w5163 ) | ( w965 & ~w5169 ) | ( w5163 & ~w5169 ) ;
  assign w5171 = w965 & w5170 ;
  assign w5172 = w4877 | w4882 ;
  assign w5173 = w5005 & ~w5172 ;
  assign w5174 = w4880 ^ w5173 ;
  assign w5175 = ( ~w965 & w5163 ) | ( ~w965 & w5169 ) | ( w5163 & w5169 ) ;
  assign w5176 = ~w5163 & w5175 ;
  assign w5177 = w5174 | w5176 ;
  assign w5178 = ( w847 & w5171 ) | ( w847 & ~w5177 ) | ( w5171 & ~w5177 ) ;
  assign w5179 = w847 & w5178 ;
  assign w5180 = w4885 | w4890 ;
  assign w5181 = w5005 & ~w5180 ;
  assign w5182 = w4888 ^ w5181 ;
  assign w5183 = ( ~w847 & w5171 ) | ( ~w847 & w5177 ) | ( w5171 & w5177 ) ;
  assign w5184 = ~w5171 & w5183 ;
  assign w5185 = w5182 | w5184 ;
  assign w5186 = ( w737 & w5179 ) | ( w737 & ~w5185 ) | ( w5179 & ~w5185 ) ;
  assign w5187 = w737 & w5186 ;
  assign w5188 = w4893 | w4898 ;
  assign w5189 = w5005 & ~w5188 ;
  assign w5190 = w4896 ^ w5189 ;
  assign w5191 = ( ~w737 & w5179 ) | ( ~w737 & w5185 ) | ( w5179 & w5185 ) ;
  assign w5192 = ~w5179 & w5191 ;
  assign w5193 = w5190 | w5192 ;
  assign w5194 = ( w635 & w5187 ) | ( w635 & ~w5193 ) | ( w5187 & ~w5193 ) ;
  assign w5195 = w635 & w5194 ;
  assign w5196 = w4901 | w4906 ;
  assign w5197 = w5005 & ~w5196 ;
  assign w5198 = w4904 ^ w5197 ;
  assign w5199 = ( ~w635 & w5187 ) | ( ~w635 & w5193 ) | ( w5187 & w5193 ) ;
  assign w5200 = ~w5187 & w5199 ;
  assign w5201 = w5198 | w5200 ;
  assign w5202 = ( w541 & w5195 ) | ( w541 & ~w5201 ) | ( w5195 & ~w5201 ) ;
  assign w5203 = w541 & w5202 ;
  assign w5204 = w4909 | w4914 ;
  assign w5205 = w5005 & ~w5204 ;
  assign w5206 = w4912 ^ w5205 ;
  assign w5207 = ( ~w541 & w5195 ) | ( ~w541 & w5201 ) | ( w5195 & w5201 ) ;
  assign w5208 = ~w5195 & w5207 ;
  assign w5209 = w5206 | w5208 ;
  assign w5210 = ( w455 & w5203 ) | ( w455 & ~w5209 ) | ( w5203 & ~w5209 ) ;
  assign w5211 = w455 & w5210 ;
  assign w5212 = w4917 | w4922 ;
  assign w5213 = w5005 & ~w5212 ;
  assign w5214 = w4920 ^ w5213 ;
  assign w5215 = ( ~w455 & w5203 ) | ( ~w455 & w5209 ) | ( w5203 & w5209 ) ;
  assign w5216 = ~w5203 & w5215 ;
  assign w5217 = w5214 | w5216 ;
  assign w5218 = ( w377 & w5211 ) | ( w377 & ~w5217 ) | ( w5211 & ~w5217 ) ;
  assign w5219 = w377 & w5218 ;
  assign w5220 = w4925 | w4930 ;
  assign w5221 = w5005 & ~w5220 ;
  assign w5222 = w4928 ^ w5221 ;
  assign w5223 = ( ~w377 & w5211 ) | ( ~w377 & w5217 ) | ( w5211 & w5217 ) ;
  assign w5224 = ~w5211 & w5223 ;
  assign w5225 = w5222 | w5224 ;
  assign w5226 = ( w307 & w5219 ) | ( w307 & ~w5225 ) | ( w5219 & ~w5225 ) ;
  assign w5227 = w307 & w5226 ;
  assign w5228 = w4933 | w4938 ;
  assign w5229 = w5005 & ~w5228 ;
  assign w5230 = w4936 ^ w5229 ;
  assign w5231 = ( ~w307 & w5219 ) | ( ~w307 & w5225 ) | ( w5219 & w5225 ) ;
  assign w5232 = ~w5219 & w5231 ;
  assign w5233 = w5230 | w5232 ;
  assign w5234 = ( w246 & w5227 ) | ( w246 & ~w5233 ) | ( w5227 & ~w5233 ) ;
  assign w5235 = w246 & w5234 ;
  assign w5236 = w4941 | w4946 ;
  assign w5237 = w5005 & ~w5236 ;
  assign w5238 = w4944 ^ w5237 ;
  assign w5239 = ( ~w246 & w5227 ) | ( ~w246 & w5233 ) | ( w5227 & w5233 ) ;
  assign w5240 = ~w5227 & w5239 ;
  assign w5241 = w5238 | w5240 ;
  assign w5242 = ( w185 & w5235 ) | ( w185 & ~w5241 ) | ( w5235 & ~w5241 ) ;
  assign w5243 = w185 & w5242 ;
  assign w5244 = w4949 | w4954 ;
  assign w5245 = w5005 & ~w5244 ;
  assign w5246 = w4952 ^ w5245 ;
  assign w5247 = ( ~w185 & w5235 ) | ( ~w185 & w5241 ) | ( w5235 & w5241 ) ;
  assign w5248 = ~w5235 & w5247 ;
  assign w5249 = w5246 | w5248 ;
  assign w5250 = ( w145 & w5243 ) | ( w145 & ~w5249 ) | ( w5243 & ~w5249 ) ;
  assign w5251 = w145 & w5250 ;
  assign w5252 = w4957 | w4962 ;
  assign w5253 = w5005 & ~w5252 ;
  assign w5254 = w4960 ^ w5253 ;
  assign w5255 = ( ~w145 & w5243 ) | ( ~w145 & w5249 ) | ( w5243 & w5249 ) ;
  assign w5256 = ~w5243 & w5255 ;
  assign w5257 = w5254 | w5256 ;
  assign w5258 = ( w132 & w5251 ) | ( w132 & ~w5257 ) | ( w5251 & ~w5257 ) ;
  assign w5259 = w132 & w5258 ;
  assign w5260 = w4965 | w4970 ;
  assign w5261 = w5005 & ~w5260 ;
  assign w5262 = w4968 ^ w5261 ;
  assign w5263 = ( ~w132 & w5251 ) | ( ~w132 & w5257 ) | ( w5251 & w5257 ) ;
  assign w5264 = ~w5251 & w5263 ;
  assign w5265 = w5262 | w5264 ;
  assign w5266 = ~w5259 & w5265 ;
  assign w5267 = w4973 | w4978 ;
  assign w5268 = w5005 & ~w5267 ;
  assign w5269 = w4976 ^ w5268 ;
  assign w5270 = ( ~w4991 & w5266 ) | ( ~w4991 & w5269 ) | ( w5266 & w5269 ) ;
  assign w5271 = w4980 & ~w5270 ;
  assign w5272 = ~w4983 & w5005 ;
  assign w5273 = ( w5270 & ~w5271 ) | ( w5270 & w5272 ) | ( ~w5271 & w5272 ) ;
  assign w5274 = w4991 | w5273 ;
  assign w5275 = ~w129 & w5274 ;
  assign w5276 = ( w5259 & w5265 ) | ( w5259 & w5269 ) | ( w5265 & w5269 ) ;
  assign w5277 = ~w5259 & w5276 ;
  assign w5278 = ( w129 & w4980 ) | ( w129 & w4983 ) | ( w4980 & w4983 ) ;
  assign w5279 = ( w4983 & ~w5005 ) | ( w4983 & w5278 ) | ( ~w5005 & w5278 ) ;
  assign w5280 = w4980 & w5279 ;
  assign w5281 = w5278 ^ w5280 ;
  assign w5282 = ( w4695 & w4700 ) | ( w4695 & w4727 ) | ( w4700 & w4727 ) ;
  assign w5283 = w4727 & ~w5282 ;
  assign w5284 = w4698 ^ w5283 ;
  assign w5285 = ( ~w4995 & w5002 ) | ( ~w4995 & w5284 ) | ( w5002 & w5284 ) ;
  assign w5286 = ~w5002 & w5285 ;
  assign w5287 = ( ~w4989 & w4991 ) | ( ~w4989 & w5286 ) | ( w4991 & w5286 ) ;
  assign w5288 = ~w4991 & w5287 ;
  assign w5289 = w5277 | w5288 ;
  assign w5290 = ( w5275 & ~w5277 ) | ( w5275 & w5281 ) | ( ~w5277 & w5281 ) ;
  assign w5291 = w5289 | w5290 ;
  assign w5292 = ( ~\pi059 & \pi060 ) | ( ~\pi059 & w5005 ) | ( \pi060 & w5005 ) ;
  assign w5293 = ( ~\pi058 & \pi060 ) | ( ~\pi058 & w5292 ) | ( \pi060 & w5292 ) ;
  assign w5294 = ( ~\pi060 & w5005 ) | ( ~\pi060 & w5291 ) | ( w5005 & w5291 ) ;
  assign w5295 = w5293 & w5294 ;
  assign w5296 = ( w4991 & w4995 ) | ( w4991 & ~w5002 ) | ( w4995 & ~w5002 ) ;
  assign w5297 = \pi059 & ~w5296 ;
  assign w5298 = \pi058 | \pi060 ;
  assign w5299 = ( ~w5296 & w5297 ) | ( ~w5296 & w5298 ) | ( w5297 & w5298 ) ;
  assign w5300 = ~w5002 & w5299 ;
  assign w5301 = ~w4989 & w5300 ;
  assign w5302 = ( \pi060 & w5291 ) | ( \pi060 & ~w5300 ) | ( w5291 & ~w5300 ) ;
  assign w5303 = w5301 & ~w5302 ;
  assign w5304 = ~\pi060 & w5291 ;
  assign w5305 = \pi061 ^ w5304 ;
  assign w5306 = w5303 | w5305 ;
  assign w5307 = ( w4727 & w5295 ) | ( w4727 & ~w5306 ) | ( w5295 & ~w5306 ) ;
  assign w5308 = w4727 & w5307 ;
  assign w5309 = ( ~w4727 & w5295 ) | ( ~w4727 & w5306 ) | ( w5295 & w5306 ) ;
  assign w5310 = ~w5295 & w5309 ;
  assign w5311 = w5005 & ~w5288 ;
  assign w5312 = ~w5277 & w5311 ;
  assign w5313 = ~w5290 & w5312 ;
  assign w5314 = \pi061 & w5291 ;
  assign w5315 = ( \pi060 & w5291 ) | ( \pi060 & ~w5314 ) | ( w5291 & ~w5314 ) ;
  assign w5316 = ( ~\pi060 & w5313 ) | ( ~\pi060 & w5315 ) | ( w5313 & w5315 ) ;
  assign w5317 = \pi062 ^ w5316 ;
  assign w5318 = w5310 | w5317 ;
  assign w5319 = ( w4457 & w5308 ) | ( w4457 & ~w5318 ) | ( w5308 & ~w5318 ) ;
  assign w5320 = w4457 & w5319 ;
  assign w5321 = ( w5009 & ~w5017 ) | ( w5009 & w5291 ) | ( ~w5017 & w5291 ) ;
  assign w5322 = ~w5009 & w5321 ;
  assign w5323 = \pi063 ^ w5322 ;
  assign w5324 = w5018 ^ w5323 ;
  assign w5325 = ( ~w4457 & w5308 ) | ( ~w4457 & w5318 ) | ( w5308 & w5318 ) ;
  assign w5326 = ~w5308 & w5325 ;
  assign w5327 = w5324 | w5326 ;
  assign w5328 = ( w4195 & w5320 ) | ( w4195 & ~w5327 ) | ( w5320 & ~w5327 ) ;
  assign w5329 = w4195 & w5328 ;
  assign w5330 = w5022 | w5024 ;
  assign w5331 = w5291 & ~w5330 ;
  assign w5332 = w5031 ^ w5331 ;
  assign w5333 = ( ~w4195 & w5320 ) | ( ~w4195 & w5327 ) | ( w5320 & w5327 ) ;
  assign w5334 = ~w5320 & w5333 ;
  assign w5335 = w5332 | w5334 ;
  assign w5336 = ( w3941 & w5329 ) | ( w3941 & ~w5335 ) | ( w5329 & ~w5335 ) ;
  assign w5337 = w3941 & w5336 ;
  assign w5338 = ( ~w3941 & w5329 ) | ( ~w3941 & w5335 ) | ( w5329 & w5335 ) ;
  assign w5339 = ~w5329 & w5338 ;
  assign w5340 = w5034 | w5036 ;
  assign w5341 = w5291 & ~w5340 ;
  assign w5342 = w5040 ^ w5341 ;
  assign w5343 = w5339 | w5342 ;
  assign w5344 = ( w3695 & w5337 ) | ( w3695 & ~w5343 ) | ( w5337 & ~w5343 ) ;
  assign w5345 = w3695 & w5344 ;
  assign w5346 = w5043 | w5048 ;
  assign w5347 = w5291 & ~w5346 ;
  assign w5348 = w5046 ^ w5347 ;
  assign w5349 = ( ~w3695 & w5337 ) | ( ~w3695 & w5343 ) | ( w5337 & w5343 ) ;
  assign w5350 = ~w5337 & w5349 ;
  assign w5351 = w5348 | w5350 ;
  assign w5352 = ( w3457 & w5345 ) | ( w3457 & ~w5351 ) | ( w5345 & ~w5351 ) ;
  assign w5353 = w3457 & w5352 ;
  assign w5354 = w5051 | w5056 ;
  assign w5355 = w5291 & ~w5354 ;
  assign w5356 = w5054 ^ w5355 ;
  assign w5357 = ( ~w3457 & w5345 ) | ( ~w3457 & w5351 ) | ( w5345 & w5351 ) ;
  assign w5358 = ~w5345 & w5357 ;
  assign w5359 = w5356 | w5358 ;
  assign w5360 = ( w3227 & w5353 ) | ( w3227 & ~w5359 ) | ( w5353 & ~w5359 ) ;
  assign w5361 = w3227 & w5360 ;
  assign w5362 = w5059 | w5064 ;
  assign w5363 = w5291 & ~w5362 ;
  assign w5364 = w5062 ^ w5363 ;
  assign w5365 = ( ~w3227 & w5353 ) | ( ~w3227 & w5359 ) | ( w5353 & w5359 ) ;
  assign w5366 = ~w5353 & w5365 ;
  assign w5367 = w5364 | w5366 ;
  assign w5368 = ( w3005 & w5361 ) | ( w3005 & ~w5367 ) | ( w5361 & ~w5367 ) ;
  assign w5369 = w3005 & w5368 ;
  assign w5370 = w5067 | w5072 ;
  assign w5371 = w5291 & ~w5370 ;
  assign w5372 = w5070 ^ w5371 ;
  assign w5373 = ( ~w3005 & w5361 ) | ( ~w3005 & w5367 ) | ( w5361 & w5367 ) ;
  assign w5374 = ~w5361 & w5373 ;
  assign w5375 = w5372 | w5374 ;
  assign w5376 = ( w2791 & w5369 ) | ( w2791 & ~w5375 ) | ( w5369 & ~w5375 ) ;
  assign w5377 = w2791 & w5376 ;
  assign w5378 = w5075 | w5080 ;
  assign w5379 = w5291 & ~w5378 ;
  assign w5380 = w5078 ^ w5379 ;
  assign w5381 = ( ~w2791 & w5369 ) | ( ~w2791 & w5375 ) | ( w5369 & w5375 ) ;
  assign w5382 = ~w5369 & w5381 ;
  assign w5383 = w5380 | w5382 ;
  assign w5384 = ( w2585 & w5377 ) | ( w2585 & ~w5383 ) | ( w5377 & ~w5383 ) ;
  assign w5385 = w2585 & w5384 ;
  assign w5386 = w5083 | w5088 ;
  assign w5387 = w5291 & ~w5386 ;
  assign w5388 = w5086 ^ w5387 ;
  assign w5389 = ( ~w2585 & w5377 ) | ( ~w2585 & w5383 ) | ( w5377 & w5383 ) ;
  assign w5390 = ~w5377 & w5389 ;
  assign w5391 = w5388 | w5390 ;
  assign w5392 = ( w2387 & w5385 ) | ( w2387 & ~w5391 ) | ( w5385 & ~w5391 ) ;
  assign w5393 = w2387 & w5392 ;
  assign w5394 = w5091 | w5096 ;
  assign w5395 = w5291 & ~w5394 ;
  assign w5396 = w5094 ^ w5395 ;
  assign w5397 = ( ~w2387 & w5385 ) | ( ~w2387 & w5391 ) | ( w5385 & w5391 ) ;
  assign w5398 = ~w5385 & w5397 ;
  assign w5399 = w5396 | w5398 ;
  assign w5400 = ( w2197 & w5393 ) | ( w2197 & ~w5399 ) | ( w5393 & ~w5399 ) ;
  assign w5401 = w2197 & w5400 ;
  assign w5402 = w5099 | w5104 ;
  assign w5403 = w5291 & ~w5402 ;
  assign w5404 = w5102 ^ w5403 ;
  assign w5405 = ( ~w2197 & w5393 ) | ( ~w2197 & w5399 ) | ( w5393 & w5399 ) ;
  assign w5406 = ~w5393 & w5405 ;
  assign w5407 = w5404 | w5406 ;
  assign w5408 = ( w2015 & w5401 ) | ( w2015 & ~w5407 ) | ( w5401 & ~w5407 ) ;
  assign w5409 = w2015 & w5408 ;
  assign w5410 = w5107 | w5112 ;
  assign w5411 = w5291 & ~w5410 ;
  assign w5412 = w5110 ^ w5411 ;
  assign w5413 = ( ~w2015 & w5401 ) | ( ~w2015 & w5407 ) | ( w5401 & w5407 ) ;
  assign w5414 = ~w5401 & w5413 ;
  assign w5415 = w5412 | w5414 ;
  assign w5416 = ( w1841 & w5409 ) | ( w1841 & ~w5415 ) | ( w5409 & ~w5415 ) ;
  assign w5417 = w1841 & w5416 ;
  assign w5418 = w5115 | w5120 ;
  assign w5419 = w5291 & ~w5418 ;
  assign w5420 = w5118 ^ w5419 ;
  assign w5421 = ( ~w1841 & w5409 ) | ( ~w1841 & w5415 ) | ( w5409 & w5415 ) ;
  assign w5422 = ~w5409 & w5421 ;
  assign w5423 = w5420 | w5422 ;
  assign w5424 = ( w1675 & w5417 ) | ( w1675 & ~w5423 ) | ( w5417 & ~w5423 ) ;
  assign w5425 = w1675 & w5424 ;
  assign w5426 = w5123 | w5128 ;
  assign w5427 = w5291 & ~w5426 ;
  assign w5428 = w5126 ^ w5427 ;
  assign w5429 = ( ~w1675 & w5417 ) | ( ~w1675 & w5423 ) | ( w5417 & w5423 ) ;
  assign w5430 = ~w5417 & w5429 ;
  assign w5431 = w5428 | w5430 ;
  assign w5432 = ( w1517 & w5425 ) | ( w1517 & ~w5431 ) | ( w5425 & ~w5431 ) ;
  assign w5433 = w1517 & w5432 ;
  assign w5434 = w5131 | w5136 ;
  assign w5435 = w5291 & ~w5434 ;
  assign w5436 = w5134 ^ w5435 ;
  assign w5437 = ( ~w1517 & w5425 ) | ( ~w1517 & w5431 ) | ( w5425 & w5431 ) ;
  assign w5438 = ~w5425 & w5437 ;
  assign w5439 = w5436 | w5438 ;
  assign w5440 = ( w1367 & w5433 ) | ( w1367 & ~w5439 ) | ( w5433 & ~w5439 ) ;
  assign w5441 = w1367 & w5440 ;
  assign w5442 = w5139 | w5144 ;
  assign w5443 = w5291 & ~w5442 ;
  assign w5444 = w5142 ^ w5443 ;
  assign w5445 = ( ~w1367 & w5433 ) | ( ~w1367 & w5439 ) | ( w5433 & w5439 ) ;
  assign w5446 = ~w5433 & w5445 ;
  assign w5447 = w5444 | w5446 ;
  assign w5448 = ( w1225 & w5441 ) | ( w1225 & ~w5447 ) | ( w5441 & ~w5447 ) ;
  assign w5449 = w1225 & w5448 ;
  assign w5450 = w5147 | w5152 ;
  assign w5451 = w5291 & ~w5450 ;
  assign w5452 = w5150 ^ w5451 ;
  assign w5453 = ( ~w1225 & w5441 ) | ( ~w1225 & w5447 ) | ( w5441 & w5447 ) ;
  assign w5454 = ~w5441 & w5453 ;
  assign w5455 = w5452 | w5454 ;
  assign w5456 = ( w1091 & w5449 ) | ( w1091 & ~w5455 ) | ( w5449 & ~w5455 ) ;
  assign w5457 = w1091 & w5456 ;
  assign w5458 = w5155 | w5160 ;
  assign w5459 = w5291 & ~w5458 ;
  assign w5460 = w5158 ^ w5459 ;
  assign w5461 = ( ~w1091 & w5449 ) | ( ~w1091 & w5455 ) | ( w5449 & w5455 ) ;
  assign w5462 = ~w5449 & w5461 ;
  assign w5463 = w5460 | w5462 ;
  assign w5464 = ( w965 & w5457 ) | ( w965 & ~w5463 ) | ( w5457 & ~w5463 ) ;
  assign w5465 = w965 & w5464 ;
  assign w5466 = w5163 | w5168 ;
  assign w5467 = w5291 & ~w5466 ;
  assign w5468 = w5166 ^ w5467 ;
  assign w5469 = ( ~w965 & w5457 ) | ( ~w965 & w5463 ) | ( w5457 & w5463 ) ;
  assign w5470 = ~w5457 & w5469 ;
  assign w5471 = w5468 | w5470 ;
  assign w5472 = ( w847 & w5465 ) | ( w847 & ~w5471 ) | ( w5465 & ~w5471 ) ;
  assign w5473 = w847 & w5472 ;
  assign w5474 = w5171 | w5176 ;
  assign w5475 = w5291 & ~w5474 ;
  assign w5476 = w5174 ^ w5475 ;
  assign w5477 = ( ~w847 & w5465 ) | ( ~w847 & w5471 ) | ( w5465 & w5471 ) ;
  assign w5478 = ~w5465 & w5477 ;
  assign w5479 = w5476 | w5478 ;
  assign w5480 = ( w737 & w5473 ) | ( w737 & ~w5479 ) | ( w5473 & ~w5479 ) ;
  assign w5481 = w737 & w5480 ;
  assign w5482 = w5179 | w5184 ;
  assign w5483 = w5291 & ~w5482 ;
  assign w5484 = w5182 ^ w5483 ;
  assign w5485 = ( ~w737 & w5473 ) | ( ~w737 & w5479 ) | ( w5473 & w5479 ) ;
  assign w5486 = ~w5473 & w5485 ;
  assign w5487 = w5484 | w5486 ;
  assign w5488 = ( w635 & w5481 ) | ( w635 & ~w5487 ) | ( w5481 & ~w5487 ) ;
  assign w5489 = w635 & w5488 ;
  assign w5490 = w5187 | w5192 ;
  assign w5491 = w5291 & ~w5490 ;
  assign w5492 = w5190 ^ w5491 ;
  assign w5493 = ( ~w635 & w5481 ) | ( ~w635 & w5487 ) | ( w5481 & w5487 ) ;
  assign w5494 = ~w5481 & w5493 ;
  assign w5495 = w5492 | w5494 ;
  assign w5496 = ( w541 & w5489 ) | ( w541 & ~w5495 ) | ( w5489 & ~w5495 ) ;
  assign w5497 = w541 & w5496 ;
  assign w5498 = w5195 | w5200 ;
  assign w5499 = w5291 & ~w5498 ;
  assign w5500 = w5198 ^ w5499 ;
  assign w5501 = ( ~w541 & w5489 ) | ( ~w541 & w5495 ) | ( w5489 & w5495 ) ;
  assign w5502 = ~w5489 & w5501 ;
  assign w5503 = w5500 | w5502 ;
  assign w5504 = ( w455 & w5497 ) | ( w455 & ~w5503 ) | ( w5497 & ~w5503 ) ;
  assign w5505 = w455 & w5504 ;
  assign w5506 = w5203 | w5208 ;
  assign w5507 = w5291 & ~w5506 ;
  assign w5508 = w5206 ^ w5507 ;
  assign w5509 = ( ~w455 & w5497 ) | ( ~w455 & w5503 ) | ( w5497 & w5503 ) ;
  assign w5510 = ~w5497 & w5509 ;
  assign w5511 = w5508 | w5510 ;
  assign w5512 = ( w377 & w5505 ) | ( w377 & ~w5511 ) | ( w5505 & ~w5511 ) ;
  assign w5513 = w377 & w5512 ;
  assign w5514 = w5211 | w5216 ;
  assign w5515 = w5291 & ~w5514 ;
  assign w5516 = w5214 ^ w5515 ;
  assign w5517 = ( ~w377 & w5505 ) | ( ~w377 & w5511 ) | ( w5505 & w5511 ) ;
  assign w5518 = ~w5505 & w5517 ;
  assign w5519 = w5516 | w5518 ;
  assign w5520 = ( w307 & w5513 ) | ( w307 & ~w5519 ) | ( w5513 & ~w5519 ) ;
  assign w5521 = w307 & w5520 ;
  assign w5522 = w5219 | w5224 ;
  assign w5523 = w5291 & ~w5522 ;
  assign w5524 = w5222 ^ w5523 ;
  assign w5525 = ( ~w307 & w5513 ) | ( ~w307 & w5519 ) | ( w5513 & w5519 ) ;
  assign w5526 = ~w5513 & w5525 ;
  assign w5527 = w5524 | w5526 ;
  assign w5528 = ( w246 & w5521 ) | ( w246 & ~w5527 ) | ( w5521 & ~w5527 ) ;
  assign w5529 = w246 & w5528 ;
  assign w5530 = w5227 | w5232 ;
  assign w5531 = w5291 & ~w5530 ;
  assign w5532 = w5230 ^ w5531 ;
  assign w5533 = ( ~w246 & w5521 ) | ( ~w246 & w5527 ) | ( w5521 & w5527 ) ;
  assign w5534 = ~w5521 & w5533 ;
  assign w5535 = w5532 | w5534 ;
  assign w5536 = ( w185 & w5529 ) | ( w185 & ~w5535 ) | ( w5529 & ~w5535 ) ;
  assign w5537 = w185 & w5536 ;
  assign w5538 = w5235 | w5240 ;
  assign w5539 = w5291 & ~w5538 ;
  assign w5540 = w5238 ^ w5539 ;
  assign w5541 = ( ~w185 & w5529 ) | ( ~w185 & w5535 ) | ( w5529 & w5535 ) ;
  assign w5542 = ~w5529 & w5541 ;
  assign w5543 = w5540 | w5542 ;
  assign w5544 = ( w145 & w5537 ) | ( w145 & ~w5543 ) | ( w5537 & ~w5543 ) ;
  assign w5545 = w145 & w5544 ;
  assign w5546 = w5243 | w5248 ;
  assign w5547 = w5291 & ~w5546 ;
  assign w5548 = w5246 ^ w5547 ;
  assign w5549 = ( ~w145 & w5537 ) | ( ~w145 & w5543 ) | ( w5537 & w5543 ) ;
  assign w5550 = ~w5537 & w5549 ;
  assign w5551 = w5548 | w5550 ;
  assign w5552 = ( w132 & w5545 ) | ( w132 & ~w5551 ) | ( w5545 & ~w5551 ) ;
  assign w5553 = w132 & w5552 ;
  assign w5554 = w5251 | w5256 ;
  assign w5555 = w5291 & ~w5554 ;
  assign w5556 = w5254 ^ w5555 ;
  assign w5557 = ( ~w132 & w5545 ) | ( ~w132 & w5551 ) | ( w5545 & w5551 ) ;
  assign w5558 = ~w5545 & w5557 ;
  assign w5559 = w5556 | w5558 ;
  assign w5560 = ~w5553 & w5559 ;
  assign w5561 = w5259 | w5264 ;
  assign w5562 = w5291 & ~w5561 ;
  assign w5563 = w5262 ^ w5562 ;
  assign w5564 = ( ~w5277 & w5560 ) | ( ~w5277 & w5563 ) | ( w5560 & w5563 ) ;
  assign w5565 = w5266 & ~w5564 ;
  assign w5566 = ~w5269 & w5291 ;
  assign w5567 = ( w5564 & ~w5565 ) | ( w5564 & w5566 ) | ( ~w5565 & w5566 ) ;
  assign w5568 = w5277 | w5567 ;
  assign w5569 = ~w129 & w5568 ;
  assign w5570 = ( w5553 & w5559 ) | ( w5553 & w5563 ) | ( w5559 & w5563 ) ;
  assign w5571 = ~w5553 & w5570 ;
  assign w5572 = ( w129 & w5266 ) | ( w129 & w5269 ) | ( w5266 & w5269 ) ;
  assign w5573 = ( w5269 & ~w5291 ) | ( w5269 & w5572 ) | ( ~w5291 & w5572 ) ;
  assign w5574 = w5266 & w5573 ;
  assign w5575 = w5572 ^ w5574 ;
  assign w5576 = ( w4973 & w4978 ) | ( w4973 & w5005 ) | ( w4978 & w5005 ) ;
  assign w5577 = w5005 & ~w5576 ;
  assign w5578 = w4976 ^ w5577 ;
  assign w5579 = ( ~w5281 & w5288 ) | ( ~w5281 & w5578 ) | ( w5288 & w5578 ) ;
  assign w5580 = ~w5288 & w5579 ;
  assign w5581 = ( ~w5275 & w5277 ) | ( ~w5275 & w5580 ) | ( w5277 & w5580 ) ;
  assign w5582 = ~w5277 & w5581 ;
  assign w5583 = w5571 | w5582 ;
  assign w5584 = ( w5569 & ~w5571 ) | ( w5569 & w5575 ) | ( ~w5571 & w5575 ) ;
  assign w5585 = w5583 | w5584 ;
  assign w5586 = ( ~\pi057 & \pi058 ) | ( ~\pi057 & w5291 ) | ( \pi058 & w5291 ) ;
  assign w5587 = ( ~\pi056 & \pi058 ) | ( ~\pi056 & w5586 ) | ( \pi058 & w5586 ) ;
  assign w5588 = ( ~\pi058 & w5291 ) | ( ~\pi058 & w5585 ) | ( w5291 & w5585 ) ;
  assign w5589 = w5587 & w5588 ;
  assign w5590 = ( w5277 & w5281 ) | ( w5277 & ~w5288 ) | ( w5281 & ~w5288 ) ;
  assign w5591 = \pi057 & ~w5590 ;
  assign w5592 = \pi056 | \pi058 ;
  assign w5593 = ( ~w5590 & w5591 ) | ( ~w5590 & w5592 ) | ( w5591 & w5592 ) ;
  assign w5594 = ~w5288 & w5593 ;
  assign w5595 = ~w5275 & w5594 ;
  assign w5596 = ( \pi058 & w5585 ) | ( \pi058 & ~w5594 ) | ( w5585 & ~w5594 ) ;
  assign w5597 = w5595 & ~w5596 ;
  assign w5598 = ~\pi058 & w5585 ;
  assign w5599 = \pi059 ^ w5598 ;
  assign w5600 = w5597 | w5599 ;
  assign w5601 = ( w5005 & w5589 ) | ( w5005 & ~w5600 ) | ( w5589 & ~w5600 ) ;
  assign w5602 = w5005 & w5601 ;
  assign w5603 = ( ~w5005 & w5589 ) | ( ~w5005 & w5600 ) | ( w5589 & w5600 ) ;
  assign w5604 = ~w5589 & w5603 ;
  assign w5605 = w5291 & ~w5582 ;
  assign w5606 = ~w5571 & w5605 ;
  assign w5607 = ~w5584 & w5606 ;
  assign w5608 = \pi059 & w5585 ;
  assign w5609 = ( \pi058 & w5585 ) | ( \pi058 & ~w5608 ) | ( w5585 & ~w5608 ) ;
  assign w5610 = ( ~\pi058 & w5607 ) | ( ~\pi058 & w5609 ) | ( w5607 & w5609 ) ;
  assign w5611 = \pi060 ^ w5610 ;
  assign w5612 = w5604 | w5611 ;
  assign w5613 = ( w4727 & w5602 ) | ( w4727 & ~w5612 ) | ( w5602 & ~w5612 ) ;
  assign w5614 = w4727 & w5613 ;
  assign w5615 = ( w5295 & ~w5303 ) | ( w5295 & w5585 ) | ( ~w5303 & w5585 ) ;
  assign w5616 = ~w5295 & w5615 ;
  assign w5617 = \pi061 ^ w5616 ;
  assign w5618 = w5304 ^ w5617 ;
  assign w5619 = ( ~w4727 & w5602 ) | ( ~w4727 & w5612 ) | ( w5602 & w5612 ) ;
  assign w5620 = ~w5602 & w5619 ;
  assign w5621 = w5618 | w5620 ;
  assign w5622 = ( w4457 & w5614 ) | ( w4457 & ~w5621 ) | ( w5614 & ~w5621 ) ;
  assign w5623 = w4457 & w5622 ;
  assign w5624 = w5308 | w5310 ;
  assign w5625 = w5585 & ~w5624 ;
  assign w5626 = w5317 ^ w5625 ;
  assign w5627 = ( ~w4457 & w5614 ) | ( ~w4457 & w5621 ) | ( w5614 & w5621 ) ;
  assign w5628 = ~w5614 & w5627 ;
  assign w5629 = w5626 | w5628 ;
  assign w5630 = ( w4195 & w5623 ) | ( w4195 & ~w5629 ) | ( w5623 & ~w5629 ) ;
  assign w5631 = w4195 & w5630 ;
  assign w5632 = w5320 | w5326 ;
  assign w5633 = w5585 & ~w5632 ;
  assign w5634 = w5324 ^ w5633 ;
  assign w5635 = ( ~w4195 & w5623 ) | ( ~w4195 & w5629 ) | ( w5623 & w5629 ) ;
  assign w5636 = ~w5623 & w5635 ;
  assign w5637 = w5634 | w5636 ;
  assign w5638 = ( w3941 & w5631 ) | ( w3941 & ~w5637 ) | ( w5631 & ~w5637 ) ;
  assign w5639 = w3941 & w5638 ;
  assign w5640 = w5329 | w5334 ;
  assign w5641 = w5585 & ~w5640 ;
  assign w5642 = w5332 ^ w5641 ;
  assign w5643 = ( ~w3941 & w5631 ) | ( ~w3941 & w5637 ) | ( w5631 & w5637 ) ;
  assign w5644 = ~w5631 & w5643 ;
  assign w5645 = w5642 | w5644 ;
  assign w5646 = ( w3695 & w5639 ) | ( w3695 & ~w5645 ) | ( w5639 & ~w5645 ) ;
  assign w5647 = w3695 & w5646 ;
  assign w5648 = ( ~w3695 & w5639 ) | ( ~w3695 & w5645 ) | ( w5639 & w5645 ) ;
  assign w5649 = ~w5639 & w5648 ;
  assign w5650 = w5337 | w5339 ;
  assign w5651 = w5585 & ~w5650 ;
  assign w5652 = w5342 ^ w5651 ;
  assign w5653 = w5649 | w5652 ;
  assign w5654 = ( w3457 & w5647 ) | ( w3457 & ~w5653 ) | ( w5647 & ~w5653 ) ;
  assign w5655 = w3457 & w5654 ;
  assign w5656 = w5345 | w5350 ;
  assign w5657 = w5585 & ~w5656 ;
  assign w5658 = w5348 ^ w5657 ;
  assign w5659 = ( ~w3457 & w5647 ) | ( ~w3457 & w5653 ) | ( w5647 & w5653 ) ;
  assign w5660 = ~w5647 & w5659 ;
  assign w5661 = w5658 | w5660 ;
  assign w5662 = ( w3227 & w5655 ) | ( w3227 & ~w5661 ) | ( w5655 & ~w5661 ) ;
  assign w5663 = w3227 & w5662 ;
  assign w5664 = w5353 | w5358 ;
  assign w5665 = w5585 & ~w5664 ;
  assign w5666 = w5356 ^ w5665 ;
  assign w5667 = ( ~w3227 & w5655 ) | ( ~w3227 & w5661 ) | ( w5655 & w5661 ) ;
  assign w5668 = ~w5655 & w5667 ;
  assign w5669 = w5666 | w5668 ;
  assign w5670 = ( w3005 & w5663 ) | ( w3005 & ~w5669 ) | ( w5663 & ~w5669 ) ;
  assign w5671 = w3005 & w5670 ;
  assign w5672 = w5361 | w5366 ;
  assign w5673 = w5585 & ~w5672 ;
  assign w5674 = w5364 ^ w5673 ;
  assign w5675 = ( ~w3005 & w5663 ) | ( ~w3005 & w5669 ) | ( w5663 & w5669 ) ;
  assign w5676 = ~w5663 & w5675 ;
  assign w5677 = w5674 | w5676 ;
  assign w5678 = ( w2791 & w5671 ) | ( w2791 & ~w5677 ) | ( w5671 & ~w5677 ) ;
  assign w5679 = w2791 & w5678 ;
  assign w5680 = w5369 | w5374 ;
  assign w5681 = w5585 & ~w5680 ;
  assign w5682 = w5372 ^ w5681 ;
  assign w5683 = ( ~w2791 & w5671 ) | ( ~w2791 & w5677 ) | ( w5671 & w5677 ) ;
  assign w5684 = ~w5671 & w5683 ;
  assign w5685 = w5682 | w5684 ;
  assign w5686 = ( w2585 & w5679 ) | ( w2585 & ~w5685 ) | ( w5679 & ~w5685 ) ;
  assign w5687 = w2585 & w5686 ;
  assign w5688 = w5377 | w5382 ;
  assign w5689 = w5585 & ~w5688 ;
  assign w5690 = w5380 ^ w5689 ;
  assign w5691 = ( ~w2585 & w5679 ) | ( ~w2585 & w5685 ) | ( w5679 & w5685 ) ;
  assign w5692 = ~w5679 & w5691 ;
  assign w5693 = w5690 | w5692 ;
  assign w5694 = ( w2387 & w5687 ) | ( w2387 & ~w5693 ) | ( w5687 & ~w5693 ) ;
  assign w5695 = w2387 & w5694 ;
  assign w5696 = w5385 | w5390 ;
  assign w5697 = w5585 & ~w5696 ;
  assign w5698 = w5388 ^ w5697 ;
  assign w5699 = ( ~w2387 & w5687 ) | ( ~w2387 & w5693 ) | ( w5687 & w5693 ) ;
  assign w5700 = ~w5687 & w5699 ;
  assign w5701 = w5698 | w5700 ;
  assign w5702 = ( w2197 & w5695 ) | ( w2197 & ~w5701 ) | ( w5695 & ~w5701 ) ;
  assign w5703 = w2197 & w5702 ;
  assign w5704 = w5393 | w5398 ;
  assign w5705 = w5585 & ~w5704 ;
  assign w5706 = w5396 ^ w5705 ;
  assign w5707 = ( ~w2197 & w5695 ) | ( ~w2197 & w5701 ) | ( w5695 & w5701 ) ;
  assign w5708 = ~w5695 & w5707 ;
  assign w5709 = w5706 | w5708 ;
  assign w5710 = ( w2015 & w5703 ) | ( w2015 & ~w5709 ) | ( w5703 & ~w5709 ) ;
  assign w5711 = w2015 & w5710 ;
  assign w5712 = w5401 | w5406 ;
  assign w5713 = w5585 & ~w5712 ;
  assign w5714 = w5404 ^ w5713 ;
  assign w5715 = ( ~w2015 & w5703 ) | ( ~w2015 & w5709 ) | ( w5703 & w5709 ) ;
  assign w5716 = ~w5703 & w5715 ;
  assign w5717 = w5714 | w5716 ;
  assign w5718 = ( w1841 & w5711 ) | ( w1841 & ~w5717 ) | ( w5711 & ~w5717 ) ;
  assign w5719 = w1841 & w5718 ;
  assign w5720 = w5409 | w5414 ;
  assign w5721 = w5585 & ~w5720 ;
  assign w5722 = w5412 ^ w5721 ;
  assign w5723 = ( ~w1841 & w5711 ) | ( ~w1841 & w5717 ) | ( w5711 & w5717 ) ;
  assign w5724 = ~w5711 & w5723 ;
  assign w5725 = w5722 | w5724 ;
  assign w5726 = ( w1675 & w5719 ) | ( w1675 & ~w5725 ) | ( w5719 & ~w5725 ) ;
  assign w5727 = w1675 & w5726 ;
  assign w5728 = w5417 | w5422 ;
  assign w5729 = w5585 & ~w5728 ;
  assign w5730 = w5420 ^ w5729 ;
  assign w5731 = ( ~w1675 & w5719 ) | ( ~w1675 & w5725 ) | ( w5719 & w5725 ) ;
  assign w5732 = ~w5719 & w5731 ;
  assign w5733 = w5730 | w5732 ;
  assign w5734 = ( w1517 & w5727 ) | ( w1517 & ~w5733 ) | ( w5727 & ~w5733 ) ;
  assign w5735 = w1517 & w5734 ;
  assign w5736 = w5425 | w5430 ;
  assign w5737 = w5585 & ~w5736 ;
  assign w5738 = w5428 ^ w5737 ;
  assign w5739 = ( ~w1517 & w5727 ) | ( ~w1517 & w5733 ) | ( w5727 & w5733 ) ;
  assign w5740 = ~w5727 & w5739 ;
  assign w5741 = w5738 | w5740 ;
  assign w5742 = ( w1367 & w5735 ) | ( w1367 & ~w5741 ) | ( w5735 & ~w5741 ) ;
  assign w5743 = w1367 & w5742 ;
  assign w5744 = w5433 | w5438 ;
  assign w5745 = w5585 & ~w5744 ;
  assign w5746 = w5436 ^ w5745 ;
  assign w5747 = ( ~w1367 & w5735 ) | ( ~w1367 & w5741 ) | ( w5735 & w5741 ) ;
  assign w5748 = ~w5735 & w5747 ;
  assign w5749 = w5746 | w5748 ;
  assign w5750 = ( w1225 & w5743 ) | ( w1225 & ~w5749 ) | ( w5743 & ~w5749 ) ;
  assign w5751 = w1225 & w5750 ;
  assign w5752 = w5441 | w5446 ;
  assign w5753 = w5585 & ~w5752 ;
  assign w5754 = w5444 ^ w5753 ;
  assign w5755 = ( ~w1225 & w5743 ) | ( ~w1225 & w5749 ) | ( w5743 & w5749 ) ;
  assign w5756 = ~w5743 & w5755 ;
  assign w5757 = w5754 | w5756 ;
  assign w5758 = ( w1091 & w5751 ) | ( w1091 & ~w5757 ) | ( w5751 & ~w5757 ) ;
  assign w5759 = w1091 & w5758 ;
  assign w5760 = w5449 | w5454 ;
  assign w5761 = w5585 & ~w5760 ;
  assign w5762 = w5452 ^ w5761 ;
  assign w5763 = ( ~w1091 & w5751 ) | ( ~w1091 & w5757 ) | ( w5751 & w5757 ) ;
  assign w5764 = ~w5751 & w5763 ;
  assign w5765 = w5762 | w5764 ;
  assign w5766 = ( w965 & w5759 ) | ( w965 & ~w5765 ) | ( w5759 & ~w5765 ) ;
  assign w5767 = w965 & w5766 ;
  assign w5768 = w5457 | w5462 ;
  assign w5769 = w5585 & ~w5768 ;
  assign w5770 = w5460 ^ w5769 ;
  assign w5771 = ( ~w965 & w5759 ) | ( ~w965 & w5765 ) | ( w5759 & w5765 ) ;
  assign w5772 = ~w5759 & w5771 ;
  assign w5773 = w5770 | w5772 ;
  assign w5774 = ( w847 & w5767 ) | ( w847 & ~w5773 ) | ( w5767 & ~w5773 ) ;
  assign w5775 = w847 & w5774 ;
  assign w5776 = w5465 | w5470 ;
  assign w5777 = w5585 & ~w5776 ;
  assign w5778 = w5468 ^ w5777 ;
  assign w5779 = ( ~w847 & w5767 ) | ( ~w847 & w5773 ) | ( w5767 & w5773 ) ;
  assign w5780 = ~w5767 & w5779 ;
  assign w5781 = w5778 | w5780 ;
  assign w5782 = ( w737 & w5775 ) | ( w737 & ~w5781 ) | ( w5775 & ~w5781 ) ;
  assign w5783 = w737 & w5782 ;
  assign w5784 = w5473 | w5478 ;
  assign w5785 = w5585 & ~w5784 ;
  assign w5786 = w5476 ^ w5785 ;
  assign w5787 = ( ~w737 & w5775 ) | ( ~w737 & w5781 ) | ( w5775 & w5781 ) ;
  assign w5788 = ~w5775 & w5787 ;
  assign w5789 = w5786 | w5788 ;
  assign w5790 = ( w635 & w5783 ) | ( w635 & ~w5789 ) | ( w5783 & ~w5789 ) ;
  assign w5791 = w635 & w5790 ;
  assign w5792 = w5481 | w5486 ;
  assign w5793 = w5585 & ~w5792 ;
  assign w5794 = w5484 ^ w5793 ;
  assign w5795 = ( ~w635 & w5783 ) | ( ~w635 & w5789 ) | ( w5783 & w5789 ) ;
  assign w5796 = ~w5783 & w5795 ;
  assign w5797 = w5794 | w5796 ;
  assign w5798 = ( w541 & w5791 ) | ( w541 & ~w5797 ) | ( w5791 & ~w5797 ) ;
  assign w5799 = w541 & w5798 ;
  assign w5800 = w5489 | w5494 ;
  assign w5801 = w5585 & ~w5800 ;
  assign w5802 = w5492 ^ w5801 ;
  assign w5803 = ( ~w541 & w5791 ) | ( ~w541 & w5797 ) | ( w5791 & w5797 ) ;
  assign w5804 = ~w5791 & w5803 ;
  assign w5805 = w5802 | w5804 ;
  assign w5806 = ( w455 & w5799 ) | ( w455 & ~w5805 ) | ( w5799 & ~w5805 ) ;
  assign w5807 = w455 & w5806 ;
  assign w5808 = w5497 | w5502 ;
  assign w5809 = w5585 & ~w5808 ;
  assign w5810 = w5500 ^ w5809 ;
  assign w5811 = ( ~w455 & w5799 ) | ( ~w455 & w5805 ) | ( w5799 & w5805 ) ;
  assign w5812 = ~w5799 & w5811 ;
  assign w5813 = w5810 | w5812 ;
  assign w5814 = ( w377 & w5807 ) | ( w377 & ~w5813 ) | ( w5807 & ~w5813 ) ;
  assign w5815 = w377 & w5814 ;
  assign w5816 = w5505 | w5510 ;
  assign w5817 = w5585 & ~w5816 ;
  assign w5818 = w5508 ^ w5817 ;
  assign w5819 = ( ~w377 & w5807 ) | ( ~w377 & w5813 ) | ( w5807 & w5813 ) ;
  assign w5820 = ~w5807 & w5819 ;
  assign w5821 = w5818 | w5820 ;
  assign w5822 = ( w307 & w5815 ) | ( w307 & ~w5821 ) | ( w5815 & ~w5821 ) ;
  assign w5823 = w307 & w5822 ;
  assign w5824 = w5513 | w5518 ;
  assign w5825 = w5585 & ~w5824 ;
  assign w5826 = w5516 ^ w5825 ;
  assign w5827 = ( ~w307 & w5815 ) | ( ~w307 & w5821 ) | ( w5815 & w5821 ) ;
  assign w5828 = ~w5815 & w5827 ;
  assign w5829 = w5826 | w5828 ;
  assign w5830 = ( w246 & w5823 ) | ( w246 & ~w5829 ) | ( w5823 & ~w5829 ) ;
  assign w5831 = w246 & w5830 ;
  assign w5832 = w5521 | w5526 ;
  assign w5833 = w5585 & ~w5832 ;
  assign w5834 = w5524 ^ w5833 ;
  assign w5835 = ( ~w246 & w5823 ) | ( ~w246 & w5829 ) | ( w5823 & w5829 ) ;
  assign w5836 = ~w5823 & w5835 ;
  assign w5837 = w5834 | w5836 ;
  assign w5838 = ( w185 & w5831 ) | ( w185 & ~w5837 ) | ( w5831 & ~w5837 ) ;
  assign w5839 = w185 & w5838 ;
  assign w5840 = w5529 | w5534 ;
  assign w5841 = w5585 & ~w5840 ;
  assign w5842 = w5532 ^ w5841 ;
  assign w5843 = ( ~w185 & w5831 ) | ( ~w185 & w5837 ) | ( w5831 & w5837 ) ;
  assign w5844 = ~w5831 & w5843 ;
  assign w5845 = w5842 | w5844 ;
  assign w5846 = ( w145 & w5839 ) | ( w145 & ~w5845 ) | ( w5839 & ~w5845 ) ;
  assign w5847 = w145 & w5846 ;
  assign w5848 = w5537 | w5542 ;
  assign w5849 = w5585 & ~w5848 ;
  assign w5850 = w5540 ^ w5849 ;
  assign w5851 = ( ~w145 & w5839 ) | ( ~w145 & w5845 ) | ( w5839 & w5845 ) ;
  assign w5852 = ~w5839 & w5851 ;
  assign w5853 = w5850 | w5852 ;
  assign w5854 = ( w132 & w5847 ) | ( w132 & ~w5853 ) | ( w5847 & ~w5853 ) ;
  assign w5855 = w132 & w5854 ;
  assign w5856 = w5545 | w5550 ;
  assign w5857 = w5585 & ~w5856 ;
  assign w5858 = w5548 ^ w5857 ;
  assign w5859 = ( ~w132 & w5847 ) | ( ~w132 & w5853 ) | ( w5847 & w5853 ) ;
  assign w5860 = ~w5847 & w5859 ;
  assign w5861 = w5858 | w5860 ;
  assign w5862 = ~w5855 & w5861 ;
  assign w5863 = w5553 | w5558 ;
  assign w5864 = w5585 & ~w5863 ;
  assign w5865 = w5556 ^ w5864 ;
  assign w5866 = ( ~w5571 & w5862 ) | ( ~w5571 & w5865 ) | ( w5862 & w5865 ) ;
  assign w5867 = w5560 & ~w5866 ;
  assign w5868 = ~w5563 & w5585 ;
  assign w5869 = ( w5866 & ~w5867 ) | ( w5866 & w5868 ) | ( ~w5867 & w5868 ) ;
  assign w5870 = w5571 | w5869 ;
  assign w5871 = ~w129 & w5870 ;
  assign w5872 = ( w5855 & w5861 ) | ( w5855 & w5865 ) | ( w5861 & w5865 ) ;
  assign w5873 = ~w5855 & w5872 ;
  assign w5874 = ( w129 & w5560 ) | ( w129 & w5563 ) | ( w5560 & w5563 ) ;
  assign w5875 = ( w5563 & ~w5585 ) | ( w5563 & w5874 ) | ( ~w5585 & w5874 ) ;
  assign w5876 = w5560 & w5875 ;
  assign w5877 = w5874 ^ w5876 ;
  assign w5878 = ( w5259 & w5264 ) | ( w5259 & w5291 ) | ( w5264 & w5291 ) ;
  assign w5879 = w5291 & ~w5878 ;
  assign w5880 = w5262 ^ w5879 ;
  assign w5881 = ( ~w5575 & w5582 ) | ( ~w5575 & w5880 ) | ( w5582 & w5880 ) ;
  assign w5882 = ~w5582 & w5881 ;
  assign w5883 = ( ~w5569 & w5571 ) | ( ~w5569 & w5882 ) | ( w5571 & w5882 ) ;
  assign w5884 = ~w5571 & w5883 ;
  assign w5885 = w5873 | w5884 ;
  assign w5886 = ( w5871 & ~w5873 ) | ( w5871 & w5877 ) | ( ~w5873 & w5877 ) ;
  assign w5887 = w5885 | w5886 ;
  assign w5888 = ( ~\pi055 & \pi056 ) | ( ~\pi055 & w5585 ) | ( \pi056 & w5585 ) ;
  assign w5889 = ( ~\pi054 & \pi056 ) | ( ~\pi054 & w5888 ) | ( \pi056 & w5888 ) ;
  assign w5890 = ( ~\pi056 & w5585 ) | ( ~\pi056 & w5887 ) | ( w5585 & w5887 ) ;
  assign w5891 = w5889 & w5890 ;
  assign w5892 = ( w5571 & w5575 ) | ( w5571 & ~w5582 ) | ( w5575 & ~w5582 ) ;
  assign w5893 = \pi055 & ~w5892 ;
  assign w5894 = \pi054 | \pi056 ;
  assign w5895 = ( ~w5892 & w5893 ) | ( ~w5892 & w5894 ) | ( w5893 & w5894 ) ;
  assign w5896 = ~w5582 & w5895 ;
  assign w5897 = ~w5569 & w5896 ;
  assign w5898 = ( \pi056 & w5887 ) | ( \pi056 & ~w5896 ) | ( w5887 & ~w5896 ) ;
  assign w5899 = w5897 & ~w5898 ;
  assign w5900 = ~\pi056 & w5887 ;
  assign w5901 = \pi057 ^ w5900 ;
  assign w5902 = w5899 | w5901 ;
  assign w5903 = ( w5291 & w5891 ) | ( w5291 & ~w5902 ) | ( w5891 & ~w5902 ) ;
  assign w5904 = w5291 & w5903 ;
  assign w5905 = ( ~w5291 & w5891 ) | ( ~w5291 & w5902 ) | ( w5891 & w5902 ) ;
  assign w5906 = ~w5891 & w5905 ;
  assign w5907 = w5585 & ~w5884 ;
  assign w5908 = ~w5873 & w5907 ;
  assign w5909 = ~w5886 & w5908 ;
  assign w5910 = \pi057 & w5887 ;
  assign w5911 = ( \pi056 & w5887 ) | ( \pi056 & ~w5910 ) | ( w5887 & ~w5910 ) ;
  assign w5912 = ( ~\pi056 & w5909 ) | ( ~\pi056 & w5911 ) | ( w5909 & w5911 ) ;
  assign w5913 = \pi058 ^ w5912 ;
  assign w5914 = w5906 | w5913 ;
  assign w5915 = ( w5005 & w5904 ) | ( w5005 & ~w5914 ) | ( w5904 & ~w5914 ) ;
  assign w5916 = w5005 & w5915 ;
  assign w5917 = ( w5589 & ~w5597 ) | ( w5589 & w5887 ) | ( ~w5597 & w5887 ) ;
  assign w5918 = ~w5589 & w5917 ;
  assign w5919 = \pi059 ^ w5918 ;
  assign w5920 = w5598 ^ w5919 ;
  assign w5921 = ( ~w5005 & w5904 ) | ( ~w5005 & w5914 ) | ( w5904 & w5914 ) ;
  assign w5922 = ~w5904 & w5921 ;
  assign w5923 = w5920 | w5922 ;
  assign w5924 = ( w4727 & w5916 ) | ( w4727 & ~w5923 ) | ( w5916 & ~w5923 ) ;
  assign w5925 = w4727 & w5924 ;
  assign w5926 = w5602 | w5604 ;
  assign w5927 = w5887 & ~w5926 ;
  assign w5928 = w5611 ^ w5927 ;
  assign w5929 = ( ~w4727 & w5916 ) | ( ~w4727 & w5923 ) | ( w5916 & w5923 ) ;
  assign w5930 = ~w5916 & w5929 ;
  assign w5931 = w5928 | w5930 ;
  assign w5932 = ( w4457 & w5925 ) | ( w4457 & ~w5931 ) | ( w5925 & ~w5931 ) ;
  assign w5933 = w4457 & w5932 ;
  assign w5934 = w5614 | w5620 ;
  assign w5935 = w5887 & ~w5934 ;
  assign w5936 = w5618 ^ w5935 ;
  assign w5937 = ( ~w4457 & w5925 ) | ( ~w4457 & w5931 ) | ( w5925 & w5931 ) ;
  assign w5938 = ~w5925 & w5937 ;
  assign w5939 = w5936 | w5938 ;
  assign w5940 = ( w4195 & w5933 ) | ( w4195 & ~w5939 ) | ( w5933 & ~w5939 ) ;
  assign w5941 = w4195 & w5940 ;
  assign w5942 = w5623 | w5628 ;
  assign w5943 = w5887 & ~w5942 ;
  assign w5944 = w5626 ^ w5943 ;
  assign w5945 = ( ~w4195 & w5933 ) | ( ~w4195 & w5939 ) | ( w5933 & w5939 ) ;
  assign w5946 = ~w5933 & w5945 ;
  assign w5947 = w5944 | w5946 ;
  assign w5948 = ( w3941 & w5941 ) | ( w3941 & ~w5947 ) | ( w5941 & ~w5947 ) ;
  assign w5949 = w3941 & w5948 ;
  assign w5950 = w5631 | w5636 ;
  assign w5951 = w5887 & ~w5950 ;
  assign w5952 = w5634 ^ w5951 ;
  assign w5953 = ( ~w3941 & w5941 ) | ( ~w3941 & w5947 ) | ( w5941 & w5947 ) ;
  assign w5954 = ~w5941 & w5953 ;
  assign w5955 = w5952 | w5954 ;
  assign w5956 = ( w3695 & w5949 ) | ( w3695 & ~w5955 ) | ( w5949 & ~w5955 ) ;
  assign w5957 = w3695 & w5956 ;
  assign w5958 = w5639 | w5644 ;
  assign w5959 = w5887 & ~w5958 ;
  assign w5960 = w5642 ^ w5959 ;
  assign w5961 = ( ~w3695 & w5949 ) | ( ~w3695 & w5955 ) | ( w5949 & w5955 ) ;
  assign w5962 = ~w5949 & w5961 ;
  assign w5963 = w5960 | w5962 ;
  assign w5964 = ( w3457 & w5957 ) | ( w3457 & ~w5963 ) | ( w5957 & ~w5963 ) ;
  assign w5965 = w3457 & w5964 ;
  assign w5966 = ( ~w3457 & w5957 ) | ( ~w3457 & w5963 ) | ( w5957 & w5963 ) ;
  assign w5967 = ~w5957 & w5966 ;
  assign w5968 = w5647 | w5649 ;
  assign w5969 = w5887 & ~w5968 ;
  assign w5970 = w5652 ^ w5969 ;
  assign w5971 = w5967 | w5970 ;
  assign w5972 = ( w3227 & w5965 ) | ( w3227 & ~w5971 ) | ( w5965 & ~w5971 ) ;
  assign w5973 = w3227 & w5972 ;
  assign w5974 = w5655 | w5660 ;
  assign w5975 = w5887 & ~w5974 ;
  assign w5976 = w5658 ^ w5975 ;
  assign w5977 = ( ~w3227 & w5965 ) | ( ~w3227 & w5971 ) | ( w5965 & w5971 ) ;
  assign w5978 = ~w5965 & w5977 ;
  assign w5979 = w5976 | w5978 ;
  assign w5980 = ( w3005 & w5973 ) | ( w3005 & ~w5979 ) | ( w5973 & ~w5979 ) ;
  assign w5981 = w3005 & w5980 ;
  assign w5982 = w5663 | w5668 ;
  assign w5983 = w5887 & ~w5982 ;
  assign w5984 = w5666 ^ w5983 ;
  assign w5985 = ( ~w3005 & w5973 ) | ( ~w3005 & w5979 ) | ( w5973 & w5979 ) ;
  assign w5986 = ~w5973 & w5985 ;
  assign w5987 = w5984 | w5986 ;
  assign w5988 = ( w2791 & w5981 ) | ( w2791 & ~w5987 ) | ( w5981 & ~w5987 ) ;
  assign w5989 = w2791 & w5988 ;
  assign w5990 = w5671 | w5676 ;
  assign w5991 = w5887 & ~w5990 ;
  assign w5992 = w5674 ^ w5991 ;
  assign w5993 = ( ~w2791 & w5981 ) | ( ~w2791 & w5987 ) | ( w5981 & w5987 ) ;
  assign w5994 = ~w5981 & w5993 ;
  assign w5995 = w5992 | w5994 ;
  assign w5996 = ( w2585 & w5989 ) | ( w2585 & ~w5995 ) | ( w5989 & ~w5995 ) ;
  assign w5997 = w2585 & w5996 ;
  assign w5998 = w5679 | w5684 ;
  assign w5999 = w5887 & ~w5998 ;
  assign w6000 = w5682 ^ w5999 ;
  assign w6001 = ( ~w2585 & w5989 ) | ( ~w2585 & w5995 ) | ( w5989 & w5995 ) ;
  assign w6002 = ~w5989 & w6001 ;
  assign w6003 = w6000 | w6002 ;
  assign w6004 = ( w2387 & w5997 ) | ( w2387 & ~w6003 ) | ( w5997 & ~w6003 ) ;
  assign w6005 = w2387 & w6004 ;
  assign w6006 = w5687 | w5692 ;
  assign w6007 = w5887 & ~w6006 ;
  assign w6008 = w5690 ^ w6007 ;
  assign w6009 = ( ~w2387 & w5997 ) | ( ~w2387 & w6003 ) | ( w5997 & w6003 ) ;
  assign w6010 = ~w5997 & w6009 ;
  assign w6011 = w6008 | w6010 ;
  assign w6012 = ( w2197 & w6005 ) | ( w2197 & ~w6011 ) | ( w6005 & ~w6011 ) ;
  assign w6013 = w2197 & w6012 ;
  assign w6014 = w5695 | w5700 ;
  assign w6015 = w5887 & ~w6014 ;
  assign w6016 = w5698 ^ w6015 ;
  assign w6017 = ( ~w2197 & w6005 ) | ( ~w2197 & w6011 ) | ( w6005 & w6011 ) ;
  assign w6018 = ~w6005 & w6017 ;
  assign w6019 = w6016 | w6018 ;
  assign w6020 = ( w2015 & w6013 ) | ( w2015 & ~w6019 ) | ( w6013 & ~w6019 ) ;
  assign w6021 = w2015 & w6020 ;
  assign w6022 = w5703 | w5708 ;
  assign w6023 = w5887 & ~w6022 ;
  assign w6024 = w5706 ^ w6023 ;
  assign w6025 = ( ~w2015 & w6013 ) | ( ~w2015 & w6019 ) | ( w6013 & w6019 ) ;
  assign w6026 = ~w6013 & w6025 ;
  assign w6027 = w6024 | w6026 ;
  assign w6028 = ( w1841 & w6021 ) | ( w1841 & ~w6027 ) | ( w6021 & ~w6027 ) ;
  assign w6029 = w1841 & w6028 ;
  assign w6030 = w5711 | w5716 ;
  assign w6031 = w5887 & ~w6030 ;
  assign w6032 = w5714 ^ w6031 ;
  assign w6033 = ( ~w1841 & w6021 ) | ( ~w1841 & w6027 ) | ( w6021 & w6027 ) ;
  assign w6034 = ~w6021 & w6033 ;
  assign w6035 = w6032 | w6034 ;
  assign w6036 = ( w1675 & w6029 ) | ( w1675 & ~w6035 ) | ( w6029 & ~w6035 ) ;
  assign w6037 = w1675 & w6036 ;
  assign w6038 = w5719 | w5724 ;
  assign w6039 = w5887 & ~w6038 ;
  assign w6040 = w5722 ^ w6039 ;
  assign w6041 = ( ~w1675 & w6029 ) | ( ~w1675 & w6035 ) | ( w6029 & w6035 ) ;
  assign w6042 = ~w6029 & w6041 ;
  assign w6043 = w6040 | w6042 ;
  assign w6044 = ( w1517 & w6037 ) | ( w1517 & ~w6043 ) | ( w6037 & ~w6043 ) ;
  assign w6045 = w1517 & w6044 ;
  assign w6046 = w5727 | w5732 ;
  assign w6047 = w5887 & ~w6046 ;
  assign w6048 = w5730 ^ w6047 ;
  assign w6049 = ( ~w1517 & w6037 ) | ( ~w1517 & w6043 ) | ( w6037 & w6043 ) ;
  assign w6050 = ~w6037 & w6049 ;
  assign w6051 = w6048 | w6050 ;
  assign w6052 = ( w1367 & w6045 ) | ( w1367 & ~w6051 ) | ( w6045 & ~w6051 ) ;
  assign w6053 = w1367 & w6052 ;
  assign w6054 = w5735 | w5740 ;
  assign w6055 = w5887 & ~w6054 ;
  assign w6056 = w5738 ^ w6055 ;
  assign w6057 = ( ~w1367 & w6045 ) | ( ~w1367 & w6051 ) | ( w6045 & w6051 ) ;
  assign w6058 = ~w6045 & w6057 ;
  assign w6059 = w6056 | w6058 ;
  assign w6060 = ( w1225 & w6053 ) | ( w1225 & ~w6059 ) | ( w6053 & ~w6059 ) ;
  assign w6061 = w1225 & w6060 ;
  assign w6062 = w5743 | w5748 ;
  assign w6063 = w5887 & ~w6062 ;
  assign w6064 = w5746 ^ w6063 ;
  assign w6065 = ( ~w1225 & w6053 ) | ( ~w1225 & w6059 ) | ( w6053 & w6059 ) ;
  assign w6066 = ~w6053 & w6065 ;
  assign w6067 = w6064 | w6066 ;
  assign w6068 = ( w1091 & w6061 ) | ( w1091 & ~w6067 ) | ( w6061 & ~w6067 ) ;
  assign w6069 = w1091 & w6068 ;
  assign w6070 = w5751 | w5756 ;
  assign w6071 = w5887 & ~w6070 ;
  assign w6072 = w5754 ^ w6071 ;
  assign w6073 = ( ~w1091 & w6061 ) | ( ~w1091 & w6067 ) | ( w6061 & w6067 ) ;
  assign w6074 = ~w6061 & w6073 ;
  assign w6075 = w6072 | w6074 ;
  assign w6076 = ( w965 & w6069 ) | ( w965 & ~w6075 ) | ( w6069 & ~w6075 ) ;
  assign w6077 = w965 & w6076 ;
  assign w6078 = w5759 | w5764 ;
  assign w6079 = w5887 & ~w6078 ;
  assign w6080 = w5762 ^ w6079 ;
  assign w6081 = ( ~w965 & w6069 ) | ( ~w965 & w6075 ) | ( w6069 & w6075 ) ;
  assign w6082 = ~w6069 & w6081 ;
  assign w6083 = w6080 | w6082 ;
  assign w6084 = ( w847 & w6077 ) | ( w847 & ~w6083 ) | ( w6077 & ~w6083 ) ;
  assign w6085 = w847 & w6084 ;
  assign w6086 = w5767 | w5772 ;
  assign w6087 = w5887 & ~w6086 ;
  assign w6088 = w5770 ^ w6087 ;
  assign w6089 = ( ~w847 & w6077 ) | ( ~w847 & w6083 ) | ( w6077 & w6083 ) ;
  assign w6090 = ~w6077 & w6089 ;
  assign w6091 = w6088 | w6090 ;
  assign w6092 = ( w737 & w6085 ) | ( w737 & ~w6091 ) | ( w6085 & ~w6091 ) ;
  assign w6093 = w737 & w6092 ;
  assign w6094 = w5775 | w5780 ;
  assign w6095 = w5887 & ~w6094 ;
  assign w6096 = w5778 ^ w6095 ;
  assign w6097 = ( ~w737 & w6085 ) | ( ~w737 & w6091 ) | ( w6085 & w6091 ) ;
  assign w6098 = ~w6085 & w6097 ;
  assign w6099 = w6096 | w6098 ;
  assign w6100 = ( w635 & w6093 ) | ( w635 & ~w6099 ) | ( w6093 & ~w6099 ) ;
  assign w6101 = w635 & w6100 ;
  assign w6102 = w5783 | w5788 ;
  assign w6103 = w5887 & ~w6102 ;
  assign w6104 = w5786 ^ w6103 ;
  assign w6105 = ( ~w635 & w6093 ) | ( ~w635 & w6099 ) | ( w6093 & w6099 ) ;
  assign w6106 = ~w6093 & w6105 ;
  assign w6107 = w6104 | w6106 ;
  assign w6108 = ( w541 & w6101 ) | ( w541 & ~w6107 ) | ( w6101 & ~w6107 ) ;
  assign w6109 = w541 & w6108 ;
  assign w6110 = w5791 | w5796 ;
  assign w6111 = w5887 & ~w6110 ;
  assign w6112 = w5794 ^ w6111 ;
  assign w6113 = ( ~w541 & w6101 ) | ( ~w541 & w6107 ) | ( w6101 & w6107 ) ;
  assign w6114 = ~w6101 & w6113 ;
  assign w6115 = w6112 | w6114 ;
  assign w6116 = ( w455 & w6109 ) | ( w455 & ~w6115 ) | ( w6109 & ~w6115 ) ;
  assign w6117 = w455 & w6116 ;
  assign w6118 = w5799 | w5804 ;
  assign w6119 = w5887 & ~w6118 ;
  assign w6120 = w5802 ^ w6119 ;
  assign w6121 = ( ~w455 & w6109 ) | ( ~w455 & w6115 ) | ( w6109 & w6115 ) ;
  assign w6122 = ~w6109 & w6121 ;
  assign w6123 = w6120 | w6122 ;
  assign w6124 = ( w377 & w6117 ) | ( w377 & ~w6123 ) | ( w6117 & ~w6123 ) ;
  assign w6125 = w377 & w6124 ;
  assign w6126 = w5807 | w5812 ;
  assign w6127 = w5887 & ~w6126 ;
  assign w6128 = w5810 ^ w6127 ;
  assign w6129 = ( ~w377 & w6117 ) | ( ~w377 & w6123 ) | ( w6117 & w6123 ) ;
  assign w6130 = ~w6117 & w6129 ;
  assign w6131 = w6128 | w6130 ;
  assign w6132 = ( w307 & w6125 ) | ( w307 & ~w6131 ) | ( w6125 & ~w6131 ) ;
  assign w6133 = w307 & w6132 ;
  assign w6134 = w5815 | w5820 ;
  assign w6135 = w5887 & ~w6134 ;
  assign w6136 = w5818 ^ w6135 ;
  assign w6137 = ( ~w307 & w6125 ) | ( ~w307 & w6131 ) | ( w6125 & w6131 ) ;
  assign w6138 = ~w6125 & w6137 ;
  assign w6139 = w6136 | w6138 ;
  assign w6140 = ( w246 & w6133 ) | ( w246 & ~w6139 ) | ( w6133 & ~w6139 ) ;
  assign w6141 = w246 & w6140 ;
  assign w6142 = w5823 | w5828 ;
  assign w6143 = w5887 & ~w6142 ;
  assign w6144 = w5826 ^ w6143 ;
  assign w6145 = ( ~w246 & w6133 ) | ( ~w246 & w6139 ) | ( w6133 & w6139 ) ;
  assign w6146 = ~w6133 & w6145 ;
  assign w6147 = w6144 | w6146 ;
  assign w6148 = ( w185 & w6141 ) | ( w185 & ~w6147 ) | ( w6141 & ~w6147 ) ;
  assign w6149 = w185 & w6148 ;
  assign w6150 = w5831 | w5836 ;
  assign w6151 = w5887 & ~w6150 ;
  assign w6152 = w5834 ^ w6151 ;
  assign w6153 = ( ~w185 & w6141 ) | ( ~w185 & w6147 ) | ( w6141 & w6147 ) ;
  assign w6154 = ~w6141 & w6153 ;
  assign w6155 = w6152 | w6154 ;
  assign w6156 = ( w145 & w6149 ) | ( w145 & ~w6155 ) | ( w6149 & ~w6155 ) ;
  assign w6157 = w145 & w6156 ;
  assign w6158 = w5839 | w5844 ;
  assign w6159 = w5887 & ~w6158 ;
  assign w6160 = w5842 ^ w6159 ;
  assign w6161 = ( ~w145 & w6149 ) | ( ~w145 & w6155 ) | ( w6149 & w6155 ) ;
  assign w6162 = ~w6149 & w6161 ;
  assign w6163 = w6160 | w6162 ;
  assign w6164 = ( w132 & w6157 ) | ( w132 & ~w6163 ) | ( w6157 & ~w6163 ) ;
  assign w6165 = w132 & w6164 ;
  assign w6166 = w5847 | w5852 ;
  assign w6167 = w5887 & ~w6166 ;
  assign w6168 = w5850 ^ w6167 ;
  assign w6169 = ( ~w132 & w6157 ) | ( ~w132 & w6163 ) | ( w6157 & w6163 ) ;
  assign w6170 = ~w6157 & w6169 ;
  assign w6171 = w6168 | w6170 ;
  assign w6172 = ~w6165 & w6171 ;
  assign w6173 = w5855 | w5860 ;
  assign w6174 = w5887 & ~w6173 ;
  assign w6175 = w5858 ^ w6174 ;
  assign w6176 = ( ~w5873 & w6172 ) | ( ~w5873 & w6175 ) | ( w6172 & w6175 ) ;
  assign w6177 = w5862 & ~w6176 ;
  assign w6178 = ~w5865 & w5887 ;
  assign w6179 = ( w6176 & ~w6177 ) | ( w6176 & w6178 ) | ( ~w6177 & w6178 ) ;
  assign w6180 = w5873 | w6179 ;
  assign w6181 = ~w129 & w6180 ;
  assign w6182 = ( w6165 & w6171 ) | ( w6165 & w6175 ) | ( w6171 & w6175 ) ;
  assign w6183 = ~w6165 & w6182 ;
  assign w6184 = ( w129 & w5862 ) | ( w129 & w5865 ) | ( w5862 & w5865 ) ;
  assign w6185 = ( w5865 & ~w5887 ) | ( w5865 & w6184 ) | ( ~w5887 & w6184 ) ;
  assign w6186 = w5862 & w6185 ;
  assign w6187 = w6184 ^ w6186 ;
  assign w6188 = ( w5553 & w5558 ) | ( w5553 & w5585 ) | ( w5558 & w5585 ) ;
  assign w6189 = w5585 & ~w6188 ;
  assign w6190 = w5556 ^ w6189 ;
  assign w6191 = ( ~w5877 & w5884 ) | ( ~w5877 & w6190 ) | ( w5884 & w6190 ) ;
  assign w6192 = ~w5884 & w6191 ;
  assign w6193 = ( ~w5871 & w5873 ) | ( ~w5871 & w6192 ) | ( w5873 & w6192 ) ;
  assign w6194 = ~w5873 & w6193 ;
  assign w6195 = w6183 | w6194 ;
  assign w6196 = ( w6181 & ~w6183 ) | ( w6181 & w6187 ) | ( ~w6183 & w6187 ) ;
  assign w6197 = w6195 | w6196 ;
  assign w6198 = ( ~\pi053 & \pi054 ) | ( ~\pi053 & w5887 ) | ( \pi054 & w5887 ) ;
  assign w6199 = ( ~\pi052 & \pi054 ) | ( ~\pi052 & w6198 ) | ( \pi054 & w6198 ) ;
  assign w6200 = ( ~\pi054 & w5887 ) | ( ~\pi054 & w6197 ) | ( w5887 & w6197 ) ;
  assign w6201 = w6199 & w6200 ;
  assign w6202 = ( w5873 & w5877 ) | ( w5873 & ~w5884 ) | ( w5877 & ~w5884 ) ;
  assign w6203 = \pi053 & ~w6202 ;
  assign w6204 = \pi052 | \pi054 ;
  assign w6205 = ( ~w6202 & w6203 ) | ( ~w6202 & w6204 ) | ( w6203 & w6204 ) ;
  assign w6206 = ~w5884 & w6205 ;
  assign w6207 = ~w5871 & w6206 ;
  assign w6208 = ( \pi054 & w6197 ) | ( \pi054 & ~w6206 ) | ( w6197 & ~w6206 ) ;
  assign w6209 = w6207 & ~w6208 ;
  assign w6210 = ~\pi054 & w6197 ;
  assign w6211 = \pi055 ^ w6210 ;
  assign w6212 = w6209 | w6211 ;
  assign w6213 = ( w5585 & w6201 ) | ( w5585 & ~w6212 ) | ( w6201 & ~w6212 ) ;
  assign w6214 = w5585 & w6213 ;
  assign w6215 = ( ~w5585 & w6201 ) | ( ~w5585 & w6212 ) | ( w6201 & w6212 ) ;
  assign w6216 = ~w6201 & w6215 ;
  assign w6217 = w5887 & ~w6194 ;
  assign w6218 = ~w6183 & w6217 ;
  assign w6219 = ~w6196 & w6218 ;
  assign w6220 = \pi055 & w6197 ;
  assign w6221 = ( \pi054 & w6197 ) | ( \pi054 & ~w6220 ) | ( w6197 & ~w6220 ) ;
  assign w6222 = ( ~\pi054 & w6219 ) | ( ~\pi054 & w6221 ) | ( w6219 & w6221 ) ;
  assign w6223 = \pi056 ^ w6222 ;
  assign w6224 = w6216 | w6223 ;
  assign w6225 = ( w5291 & w6214 ) | ( w5291 & ~w6224 ) | ( w6214 & ~w6224 ) ;
  assign w6226 = w5291 & w6225 ;
  assign w6227 = ( w5891 & ~w5899 ) | ( w5891 & w6197 ) | ( ~w5899 & w6197 ) ;
  assign w6228 = ~w5891 & w6227 ;
  assign w6229 = \pi057 ^ w6228 ;
  assign w6230 = w5900 ^ w6229 ;
  assign w6231 = ( ~w5291 & w6214 ) | ( ~w5291 & w6224 ) | ( w6214 & w6224 ) ;
  assign w6232 = ~w6214 & w6231 ;
  assign w6233 = w6230 | w6232 ;
  assign w6234 = ( w5005 & w6226 ) | ( w5005 & ~w6233 ) | ( w6226 & ~w6233 ) ;
  assign w6235 = w5005 & w6234 ;
  assign w6236 = w5904 | w5906 ;
  assign w6237 = w6197 & ~w6236 ;
  assign w6238 = w5913 ^ w6237 ;
  assign w6239 = ( ~w5005 & w6226 ) | ( ~w5005 & w6233 ) | ( w6226 & w6233 ) ;
  assign w6240 = ~w6226 & w6239 ;
  assign w6241 = w6238 | w6240 ;
  assign w6242 = ( w4727 & w6235 ) | ( w4727 & ~w6241 ) | ( w6235 & ~w6241 ) ;
  assign w6243 = w4727 & w6242 ;
  assign w6244 = w5916 | w5922 ;
  assign w6245 = w6197 & ~w6244 ;
  assign w6246 = w5920 ^ w6245 ;
  assign w6247 = ( ~w4727 & w6235 ) | ( ~w4727 & w6241 ) | ( w6235 & w6241 ) ;
  assign w6248 = ~w6235 & w6247 ;
  assign w6249 = w6246 | w6248 ;
  assign w6250 = ( w4457 & w6243 ) | ( w4457 & ~w6249 ) | ( w6243 & ~w6249 ) ;
  assign w6251 = w4457 & w6250 ;
  assign w6252 = w5925 | w5930 ;
  assign w6253 = w6197 & ~w6252 ;
  assign w6254 = w5928 ^ w6253 ;
  assign w6255 = ( ~w4457 & w6243 ) | ( ~w4457 & w6249 ) | ( w6243 & w6249 ) ;
  assign w6256 = ~w6243 & w6255 ;
  assign w6257 = w6254 | w6256 ;
  assign w6258 = ( w4195 & w6251 ) | ( w4195 & ~w6257 ) | ( w6251 & ~w6257 ) ;
  assign w6259 = w4195 & w6258 ;
  assign w6260 = w5933 | w5938 ;
  assign w6261 = w6197 & ~w6260 ;
  assign w6262 = w5936 ^ w6261 ;
  assign w6263 = ( ~w4195 & w6251 ) | ( ~w4195 & w6257 ) | ( w6251 & w6257 ) ;
  assign w6264 = ~w6251 & w6263 ;
  assign w6265 = w6262 | w6264 ;
  assign w6266 = ( w3941 & w6259 ) | ( w3941 & ~w6265 ) | ( w6259 & ~w6265 ) ;
  assign w6267 = w3941 & w6266 ;
  assign w6268 = w5941 | w5946 ;
  assign w6269 = w6197 & ~w6268 ;
  assign w6270 = w5944 ^ w6269 ;
  assign w6271 = ( ~w3941 & w6259 ) | ( ~w3941 & w6265 ) | ( w6259 & w6265 ) ;
  assign w6272 = ~w6259 & w6271 ;
  assign w6273 = w6270 | w6272 ;
  assign w6274 = ( w3695 & w6267 ) | ( w3695 & ~w6273 ) | ( w6267 & ~w6273 ) ;
  assign w6275 = w3695 & w6274 ;
  assign w6276 = w5949 | w5954 ;
  assign w6277 = w6197 & ~w6276 ;
  assign w6278 = w5952 ^ w6277 ;
  assign w6279 = ( ~w3695 & w6267 ) | ( ~w3695 & w6273 ) | ( w6267 & w6273 ) ;
  assign w6280 = ~w6267 & w6279 ;
  assign w6281 = w6278 | w6280 ;
  assign w6282 = ( w3457 & w6275 ) | ( w3457 & ~w6281 ) | ( w6275 & ~w6281 ) ;
  assign w6283 = w3457 & w6282 ;
  assign w6284 = w5957 | w5962 ;
  assign w6285 = w6197 & ~w6284 ;
  assign w6286 = w5960 ^ w6285 ;
  assign w6287 = ( ~w3457 & w6275 ) | ( ~w3457 & w6281 ) | ( w6275 & w6281 ) ;
  assign w6288 = ~w6275 & w6287 ;
  assign w6289 = w6286 | w6288 ;
  assign w6290 = ( w3227 & w6283 ) | ( w3227 & ~w6289 ) | ( w6283 & ~w6289 ) ;
  assign w6291 = w3227 & w6290 ;
  assign w6292 = ( ~w3227 & w6283 ) | ( ~w3227 & w6289 ) | ( w6283 & w6289 ) ;
  assign w6293 = ~w6283 & w6292 ;
  assign w6294 = w5965 | w5967 ;
  assign w6295 = w6197 & ~w6294 ;
  assign w6296 = w5970 ^ w6295 ;
  assign w6297 = w6293 | w6296 ;
  assign w6298 = ( w3005 & w6291 ) | ( w3005 & ~w6297 ) | ( w6291 & ~w6297 ) ;
  assign w6299 = w3005 & w6298 ;
  assign w6300 = w5973 | w5978 ;
  assign w6301 = w6197 & ~w6300 ;
  assign w6302 = w5976 ^ w6301 ;
  assign w6303 = ( ~w3005 & w6291 ) | ( ~w3005 & w6297 ) | ( w6291 & w6297 ) ;
  assign w6304 = ~w6291 & w6303 ;
  assign w6305 = w6302 | w6304 ;
  assign w6306 = ( w2791 & w6299 ) | ( w2791 & ~w6305 ) | ( w6299 & ~w6305 ) ;
  assign w6307 = w2791 & w6306 ;
  assign w6308 = w5981 | w5986 ;
  assign w6309 = w6197 & ~w6308 ;
  assign w6310 = w5984 ^ w6309 ;
  assign w6311 = ( ~w2791 & w6299 ) | ( ~w2791 & w6305 ) | ( w6299 & w6305 ) ;
  assign w6312 = ~w6299 & w6311 ;
  assign w6313 = w6310 | w6312 ;
  assign w6314 = ( w2585 & w6307 ) | ( w2585 & ~w6313 ) | ( w6307 & ~w6313 ) ;
  assign w6315 = w2585 & w6314 ;
  assign w6316 = w5989 | w5994 ;
  assign w6317 = w6197 & ~w6316 ;
  assign w6318 = w5992 ^ w6317 ;
  assign w6319 = ( ~w2585 & w6307 ) | ( ~w2585 & w6313 ) | ( w6307 & w6313 ) ;
  assign w6320 = ~w6307 & w6319 ;
  assign w6321 = w6318 | w6320 ;
  assign w6322 = ( w2387 & w6315 ) | ( w2387 & ~w6321 ) | ( w6315 & ~w6321 ) ;
  assign w6323 = w2387 & w6322 ;
  assign w6324 = w5997 | w6002 ;
  assign w6325 = w6197 & ~w6324 ;
  assign w6326 = w6000 ^ w6325 ;
  assign w6327 = ( ~w2387 & w6315 ) | ( ~w2387 & w6321 ) | ( w6315 & w6321 ) ;
  assign w6328 = ~w6315 & w6327 ;
  assign w6329 = w6326 | w6328 ;
  assign w6330 = ( w2197 & w6323 ) | ( w2197 & ~w6329 ) | ( w6323 & ~w6329 ) ;
  assign w6331 = w2197 & w6330 ;
  assign w6332 = w6005 | w6010 ;
  assign w6333 = w6197 & ~w6332 ;
  assign w6334 = w6008 ^ w6333 ;
  assign w6335 = ( ~w2197 & w6323 ) | ( ~w2197 & w6329 ) | ( w6323 & w6329 ) ;
  assign w6336 = ~w6323 & w6335 ;
  assign w6337 = w6334 | w6336 ;
  assign w6338 = ( w2015 & w6331 ) | ( w2015 & ~w6337 ) | ( w6331 & ~w6337 ) ;
  assign w6339 = w2015 & w6338 ;
  assign w6340 = w6013 | w6018 ;
  assign w6341 = w6197 & ~w6340 ;
  assign w6342 = w6016 ^ w6341 ;
  assign w6343 = ( ~w2015 & w6331 ) | ( ~w2015 & w6337 ) | ( w6331 & w6337 ) ;
  assign w6344 = ~w6331 & w6343 ;
  assign w6345 = w6342 | w6344 ;
  assign w6346 = ( w1841 & w6339 ) | ( w1841 & ~w6345 ) | ( w6339 & ~w6345 ) ;
  assign w6347 = w1841 & w6346 ;
  assign w6348 = w6021 | w6026 ;
  assign w6349 = w6197 & ~w6348 ;
  assign w6350 = w6024 ^ w6349 ;
  assign w6351 = ( ~w1841 & w6339 ) | ( ~w1841 & w6345 ) | ( w6339 & w6345 ) ;
  assign w6352 = ~w6339 & w6351 ;
  assign w6353 = w6350 | w6352 ;
  assign w6354 = ( w1675 & w6347 ) | ( w1675 & ~w6353 ) | ( w6347 & ~w6353 ) ;
  assign w6355 = w1675 & w6354 ;
  assign w6356 = w6029 | w6034 ;
  assign w6357 = w6197 & ~w6356 ;
  assign w6358 = w6032 ^ w6357 ;
  assign w6359 = ( ~w1675 & w6347 ) | ( ~w1675 & w6353 ) | ( w6347 & w6353 ) ;
  assign w6360 = ~w6347 & w6359 ;
  assign w6361 = w6358 | w6360 ;
  assign w6362 = ( w1517 & w6355 ) | ( w1517 & ~w6361 ) | ( w6355 & ~w6361 ) ;
  assign w6363 = w1517 & w6362 ;
  assign w6364 = w6037 | w6042 ;
  assign w6365 = w6197 & ~w6364 ;
  assign w6366 = w6040 ^ w6365 ;
  assign w6367 = ( ~w1517 & w6355 ) | ( ~w1517 & w6361 ) | ( w6355 & w6361 ) ;
  assign w6368 = ~w6355 & w6367 ;
  assign w6369 = w6366 | w6368 ;
  assign w6370 = ( w1367 & w6363 ) | ( w1367 & ~w6369 ) | ( w6363 & ~w6369 ) ;
  assign w6371 = w1367 & w6370 ;
  assign w6372 = w6045 | w6050 ;
  assign w6373 = w6197 & ~w6372 ;
  assign w6374 = w6048 ^ w6373 ;
  assign w6375 = ( ~w1367 & w6363 ) | ( ~w1367 & w6369 ) | ( w6363 & w6369 ) ;
  assign w6376 = ~w6363 & w6375 ;
  assign w6377 = w6374 | w6376 ;
  assign w6378 = ( w1225 & w6371 ) | ( w1225 & ~w6377 ) | ( w6371 & ~w6377 ) ;
  assign w6379 = w1225 & w6378 ;
  assign w6380 = w6053 | w6058 ;
  assign w6381 = w6197 & ~w6380 ;
  assign w6382 = w6056 ^ w6381 ;
  assign w6383 = ( ~w1225 & w6371 ) | ( ~w1225 & w6377 ) | ( w6371 & w6377 ) ;
  assign w6384 = ~w6371 & w6383 ;
  assign w6385 = w6382 | w6384 ;
  assign w6386 = ( w1091 & w6379 ) | ( w1091 & ~w6385 ) | ( w6379 & ~w6385 ) ;
  assign w6387 = w1091 & w6386 ;
  assign w6388 = w6061 | w6066 ;
  assign w6389 = w6197 & ~w6388 ;
  assign w6390 = w6064 ^ w6389 ;
  assign w6391 = ( ~w1091 & w6379 ) | ( ~w1091 & w6385 ) | ( w6379 & w6385 ) ;
  assign w6392 = ~w6379 & w6391 ;
  assign w6393 = w6390 | w6392 ;
  assign w6394 = ( w965 & w6387 ) | ( w965 & ~w6393 ) | ( w6387 & ~w6393 ) ;
  assign w6395 = w965 & w6394 ;
  assign w6396 = w6069 | w6074 ;
  assign w6397 = w6197 & ~w6396 ;
  assign w6398 = w6072 ^ w6397 ;
  assign w6399 = ( ~w965 & w6387 ) | ( ~w965 & w6393 ) | ( w6387 & w6393 ) ;
  assign w6400 = ~w6387 & w6399 ;
  assign w6401 = w6398 | w6400 ;
  assign w6402 = ( w847 & w6395 ) | ( w847 & ~w6401 ) | ( w6395 & ~w6401 ) ;
  assign w6403 = w847 & w6402 ;
  assign w6404 = w6077 | w6082 ;
  assign w6405 = w6197 & ~w6404 ;
  assign w6406 = w6080 ^ w6405 ;
  assign w6407 = ( ~w847 & w6395 ) | ( ~w847 & w6401 ) | ( w6395 & w6401 ) ;
  assign w6408 = ~w6395 & w6407 ;
  assign w6409 = w6406 | w6408 ;
  assign w6410 = ( w737 & w6403 ) | ( w737 & ~w6409 ) | ( w6403 & ~w6409 ) ;
  assign w6411 = w737 & w6410 ;
  assign w6412 = w6085 | w6090 ;
  assign w6413 = w6197 & ~w6412 ;
  assign w6414 = w6088 ^ w6413 ;
  assign w6415 = ( ~w737 & w6403 ) | ( ~w737 & w6409 ) | ( w6403 & w6409 ) ;
  assign w6416 = ~w6403 & w6415 ;
  assign w6417 = w6414 | w6416 ;
  assign w6418 = ( w635 & w6411 ) | ( w635 & ~w6417 ) | ( w6411 & ~w6417 ) ;
  assign w6419 = w635 & w6418 ;
  assign w6420 = w6093 | w6098 ;
  assign w6421 = w6197 & ~w6420 ;
  assign w6422 = w6096 ^ w6421 ;
  assign w6423 = ( ~w635 & w6411 ) | ( ~w635 & w6417 ) | ( w6411 & w6417 ) ;
  assign w6424 = ~w6411 & w6423 ;
  assign w6425 = w6422 | w6424 ;
  assign w6426 = ( w541 & w6419 ) | ( w541 & ~w6425 ) | ( w6419 & ~w6425 ) ;
  assign w6427 = w541 & w6426 ;
  assign w6428 = w6101 | w6106 ;
  assign w6429 = w6197 & ~w6428 ;
  assign w6430 = w6104 ^ w6429 ;
  assign w6431 = ( ~w541 & w6419 ) | ( ~w541 & w6425 ) | ( w6419 & w6425 ) ;
  assign w6432 = ~w6419 & w6431 ;
  assign w6433 = w6430 | w6432 ;
  assign w6434 = ( w455 & w6427 ) | ( w455 & ~w6433 ) | ( w6427 & ~w6433 ) ;
  assign w6435 = w455 & w6434 ;
  assign w6436 = w6109 | w6114 ;
  assign w6437 = w6197 & ~w6436 ;
  assign w6438 = w6112 ^ w6437 ;
  assign w6439 = ( ~w455 & w6427 ) | ( ~w455 & w6433 ) | ( w6427 & w6433 ) ;
  assign w6440 = ~w6427 & w6439 ;
  assign w6441 = w6438 | w6440 ;
  assign w6442 = ( w377 & w6435 ) | ( w377 & ~w6441 ) | ( w6435 & ~w6441 ) ;
  assign w6443 = w377 & w6442 ;
  assign w6444 = w6117 | w6122 ;
  assign w6445 = w6197 & ~w6444 ;
  assign w6446 = w6120 ^ w6445 ;
  assign w6447 = ( ~w377 & w6435 ) | ( ~w377 & w6441 ) | ( w6435 & w6441 ) ;
  assign w6448 = ~w6435 & w6447 ;
  assign w6449 = w6446 | w6448 ;
  assign w6450 = ( w307 & w6443 ) | ( w307 & ~w6449 ) | ( w6443 & ~w6449 ) ;
  assign w6451 = w307 & w6450 ;
  assign w6452 = w6125 | w6130 ;
  assign w6453 = w6197 & ~w6452 ;
  assign w6454 = w6128 ^ w6453 ;
  assign w6455 = ( ~w307 & w6443 ) | ( ~w307 & w6449 ) | ( w6443 & w6449 ) ;
  assign w6456 = ~w6443 & w6455 ;
  assign w6457 = w6454 | w6456 ;
  assign w6458 = ( w246 & w6451 ) | ( w246 & ~w6457 ) | ( w6451 & ~w6457 ) ;
  assign w6459 = w246 & w6458 ;
  assign w6460 = w6133 | w6138 ;
  assign w6461 = w6197 & ~w6460 ;
  assign w6462 = w6136 ^ w6461 ;
  assign w6463 = ( ~w246 & w6451 ) | ( ~w246 & w6457 ) | ( w6451 & w6457 ) ;
  assign w6464 = ~w6451 & w6463 ;
  assign w6465 = w6462 | w6464 ;
  assign w6466 = ( w185 & w6459 ) | ( w185 & ~w6465 ) | ( w6459 & ~w6465 ) ;
  assign w6467 = w185 & w6466 ;
  assign w6468 = w6141 | w6146 ;
  assign w6469 = w6197 & ~w6468 ;
  assign w6470 = w6144 ^ w6469 ;
  assign w6471 = ( ~w185 & w6459 ) | ( ~w185 & w6465 ) | ( w6459 & w6465 ) ;
  assign w6472 = ~w6459 & w6471 ;
  assign w6473 = w6470 | w6472 ;
  assign w6474 = ( w145 & w6467 ) | ( w145 & ~w6473 ) | ( w6467 & ~w6473 ) ;
  assign w6475 = w145 & w6474 ;
  assign w6476 = w6149 | w6154 ;
  assign w6477 = w6197 & ~w6476 ;
  assign w6478 = w6152 ^ w6477 ;
  assign w6479 = ( ~w145 & w6467 ) | ( ~w145 & w6473 ) | ( w6467 & w6473 ) ;
  assign w6480 = ~w6467 & w6479 ;
  assign w6481 = w6478 | w6480 ;
  assign w6482 = ( w132 & w6475 ) | ( w132 & ~w6481 ) | ( w6475 & ~w6481 ) ;
  assign w6483 = w132 & w6482 ;
  assign w6484 = w6157 | w6162 ;
  assign w6485 = w6197 & ~w6484 ;
  assign w6486 = w6160 ^ w6485 ;
  assign w6487 = ( ~w132 & w6475 ) | ( ~w132 & w6481 ) | ( w6475 & w6481 ) ;
  assign w6488 = ~w6475 & w6487 ;
  assign w6489 = w6486 | w6488 ;
  assign w6490 = ~w6483 & w6489 ;
  assign w6491 = w6165 | w6170 ;
  assign w6492 = w6197 & ~w6491 ;
  assign w6493 = w6168 ^ w6492 ;
  assign w6494 = ( ~w6183 & w6490 ) | ( ~w6183 & w6493 ) | ( w6490 & w6493 ) ;
  assign w6495 = w6172 & ~w6494 ;
  assign w6496 = ~w6175 & w6197 ;
  assign w6497 = ( w6494 & ~w6495 ) | ( w6494 & w6496 ) | ( ~w6495 & w6496 ) ;
  assign w6498 = w6183 | w6497 ;
  assign w6499 = ~w129 & w6498 ;
  assign w6500 = ( w6483 & w6489 ) | ( w6483 & w6493 ) | ( w6489 & w6493 ) ;
  assign w6501 = ~w6483 & w6500 ;
  assign w6502 = ( w129 & w6172 ) | ( w129 & w6175 ) | ( w6172 & w6175 ) ;
  assign w6503 = ( w6175 & ~w6197 ) | ( w6175 & w6502 ) | ( ~w6197 & w6502 ) ;
  assign w6504 = w6172 & w6503 ;
  assign w6505 = w6502 ^ w6504 ;
  assign w6506 = ( w5855 & w5860 ) | ( w5855 & w5887 ) | ( w5860 & w5887 ) ;
  assign w6507 = w5887 & ~w6506 ;
  assign w6508 = w5858 ^ w6507 ;
  assign w6509 = ( ~w6187 & w6194 ) | ( ~w6187 & w6508 ) | ( w6194 & w6508 ) ;
  assign w6510 = ~w6194 & w6509 ;
  assign w6511 = ( ~w6181 & w6183 ) | ( ~w6181 & w6510 ) | ( w6183 & w6510 ) ;
  assign w6512 = ~w6183 & w6511 ;
  assign w6513 = w6501 | w6512 ;
  assign w6514 = ( w6499 & ~w6501 ) | ( w6499 & w6505 ) | ( ~w6501 & w6505 ) ;
  assign w6515 = w6513 | w6514 ;
  assign w6516 = ( ~\pi051 & \pi052 ) | ( ~\pi051 & w6197 ) | ( \pi052 & w6197 ) ;
  assign w6517 = ( ~\pi050 & \pi052 ) | ( ~\pi050 & w6516 ) | ( \pi052 & w6516 ) ;
  assign w6518 = ( ~\pi052 & w6197 ) | ( ~\pi052 & w6515 ) | ( w6197 & w6515 ) ;
  assign w6519 = w6517 & w6518 ;
  assign w6520 = ( w6183 & w6187 ) | ( w6183 & ~w6194 ) | ( w6187 & ~w6194 ) ;
  assign w6521 = \pi051 & ~w6520 ;
  assign w6522 = \pi050 | \pi052 ;
  assign w6523 = ( ~w6520 & w6521 ) | ( ~w6520 & w6522 ) | ( w6521 & w6522 ) ;
  assign w6524 = ~w6194 & w6523 ;
  assign w6525 = ~w6181 & w6524 ;
  assign w6526 = ( \pi052 & w6515 ) | ( \pi052 & ~w6524 ) | ( w6515 & ~w6524 ) ;
  assign w6527 = w6525 & ~w6526 ;
  assign w6528 = ~\pi052 & w6515 ;
  assign w6529 = \pi053 ^ w6528 ;
  assign w6530 = w6527 | w6529 ;
  assign w6531 = ( w5887 & w6519 ) | ( w5887 & ~w6530 ) | ( w6519 & ~w6530 ) ;
  assign w6532 = w5887 & w6531 ;
  assign w6533 = ( ~w5887 & w6519 ) | ( ~w5887 & w6530 ) | ( w6519 & w6530 ) ;
  assign w6534 = ~w6519 & w6533 ;
  assign w6535 = w6197 & ~w6512 ;
  assign w6536 = ~w6501 & w6535 ;
  assign w6537 = ~w6514 & w6536 ;
  assign w6538 = \pi053 & w6515 ;
  assign w6539 = ( \pi052 & w6515 ) | ( \pi052 & ~w6538 ) | ( w6515 & ~w6538 ) ;
  assign w6540 = ( ~\pi052 & w6537 ) | ( ~\pi052 & w6539 ) | ( w6537 & w6539 ) ;
  assign w6541 = \pi054 ^ w6540 ;
  assign w6542 = w6534 | w6541 ;
  assign w6543 = ( w5585 & w6532 ) | ( w5585 & ~w6542 ) | ( w6532 & ~w6542 ) ;
  assign w6544 = w5585 & w6543 ;
  assign w6545 = ( w6201 & ~w6209 ) | ( w6201 & w6515 ) | ( ~w6209 & w6515 ) ;
  assign w6546 = ~w6201 & w6545 ;
  assign w6547 = \pi055 ^ w6546 ;
  assign w6548 = w6210 ^ w6547 ;
  assign w6549 = ( ~w5585 & w6532 ) | ( ~w5585 & w6542 ) | ( w6532 & w6542 ) ;
  assign w6550 = ~w6532 & w6549 ;
  assign w6551 = w6548 | w6550 ;
  assign w6552 = ( w5291 & w6544 ) | ( w5291 & ~w6551 ) | ( w6544 & ~w6551 ) ;
  assign w6553 = w5291 & w6552 ;
  assign w6554 = w6214 | w6216 ;
  assign w6555 = w6515 & ~w6554 ;
  assign w6556 = w6223 ^ w6555 ;
  assign w6557 = ( ~w5291 & w6544 ) | ( ~w5291 & w6551 ) | ( w6544 & w6551 ) ;
  assign w6558 = ~w6544 & w6557 ;
  assign w6559 = w6556 | w6558 ;
  assign w6560 = ( w5005 & w6553 ) | ( w5005 & ~w6559 ) | ( w6553 & ~w6559 ) ;
  assign w6561 = w5005 & w6560 ;
  assign w6562 = w6226 | w6232 ;
  assign w6563 = w6515 & ~w6562 ;
  assign w6564 = w6230 ^ w6563 ;
  assign w6565 = ( ~w5005 & w6553 ) | ( ~w5005 & w6559 ) | ( w6553 & w6559 ) ;
  assign w6566 = ~w6553 & w6565 ;
  assign w6567 = w6564 | w6566 ;
  assign w6568 = ( w4727 & w6561 ) | ( w4727 & ~w6567 ) | ( w6561 & ~w6567 ) ;
  assign w6569 = w4727 & w6568 ;
  assign w6570 = w6235 | w6240 ;
  assign w6571 = w6515 & ~w6570 ;
  assign w6572 = w6238 ^ w6571 ;
  assign w6573 = ( ~w4727 & w6561 ) | ( ~w4727 & w6567 ) | ( w6561 & w6567 ) ;
  assign w6574 = ~w6561 & w6573 ;
  assign w6575 = w6572 | w6574 ;
  assign w6576 = ( w4457 & w6569 ) | ( w4457 & ~w6575 ) | ( w6569 & ~w6575 ) ;
  assign w6577 = w4457 & w6576 ;
  assign w6578 = w6243 | w6248 ;
  assign w6579 = w6515 & ~w6578 ;
  assign w6580 = w6246 ^ w6579 ;
  assign w6581 = ( ~w4457 & w6569 ) | ( ~w4457 & w6575 ) | ( w6569 & w6575 ) ;
  assign w6582 = ~w6569 & w6581 ;
  assign w6583 = w6580 | w6582 ;
  assign w6584 = ( w4195 & w6577 ) | ( w4195 & ~w6583 ) | ( w6577 & ~w6583 ) ;
  assign w6585 = w4195 & w6584 ;
  assign w6586 = w6251 | w6256 ;
  assign w6587 = w6515 & ~w6586 ;
  assign w6588 = w6254 ^ w6587 ;
  assign w6589 = ( ~w4195 & w6577 ) | ( ~w4195 & w6583 ) | ( w6577 & w6583 ) ;
  assign w6590 = ~w6577 & w6589 ;
  assign w6591 = w6588 | w6590 ;
  assign w6592 = ( w3941 & w6585 ) | ( w3941 & ~w6591 ) | ( w6585 & ~w6591 ) ;
  assign w6593 = w3941 & w6592 ;
  assign w6594 = w6259 | w6264 ;
  assign w6595 = w6515 & ~w6594 ;
  assign w6596 = w6262 ^ w6595 ;
  assign w6597 = ( ~w3941 & w6585 ) | ( ~w3941 & w6591 ) | ( w6585 & w6591 ) ;
  assign w6598 = ~w6585 & w6597 ;
  assign w6599 = w6596 | w6598 ;
  assign w6600 = ( w3695 & w6593 ) | ( w3695 & ~w6599 ) | ( w6593 & ~w6599 ) ;
  assign w6601 = w3695 & w6600 ;
  assign w6602 = w6267 | w6272 ;
  assign w6603 = w6515 & ~w6602 ;
  assign w6604 = w6270 ^ w6603 ;
  assign w6605 = ( ~w3695 & w6593 ) | ( ~w3695 & w6599 ) | ( w6593 & w6599 ) ;
  assign w6606 = ~w6593 & w6605 ;
  assign w6607 = w6604 | w6606 ;
  assign w6608 = ( w3457 & w6601 ) | ( w3457 & ~w6607 ) | ( w6601 & ~w6607 ) ;
  assign w6609 = w3457 & w6608 ;
  assign w6610 = w6275 | w6280 ;
  assign w6611 = w6515 & ~w6610 ;
  assign w6612 = w6278 ^ w6611 ;
  assign w6613 = ( ~w3457 & w6601 ) | ( ~w3457 & w6607 ) | ( w6601 & w6607 ) ;
  assign w6614 = ~w6601 & w6613 ;
  assign w6615 = w6612 | w6614 ;
  assign w6616 = ( w3227 & w6609 ) | ( w3227 & ~w6615 ) | ( w6609 & ~w6615 ) ;
  assign w6617 = w3227 & w6616 ;
  assign w6618 = w6283 | w6288 ;
  assign w6619 = w6515 & ~w6618 ;
  assign w6620 = w6286 ^ w6619 ;
  assign w6621 = ( ~w3227 & w6609 ) | ( ~w3227 & w6615 ) | ( w6609 & w6615 ) ;
  assign w6622 = ~w6609 & w6621 ;
  assign w6623 = w6620 | w6622 ;
  assign w6624 = ( w3005 & w6617 ) | ( w3005 & ~w6623 ) | ( w6617 & ~w6623 ) ;
  assign w6625 = w3005 & w6624 ;
  assign w6626 = ( ~w3005 & w6617 ) | ( ~w3005 & w6623 ) | ( w6617 & w6623 ) ;
  assign w6627 = ~w6617 & w6626 ;
  assign w6628 = w6291 | w6293 ;
  assign w6629 = w6515 & ~w6628 ;
  assign w6630 = w6296 ^ w6629 ;
  assign w6631 = w6627 | w6630 ;
  assign w6632 = ( w2791 & w6625 ) | ( w2791 & ~w6631 ) | ( w6625 & ~w6631 ) ;
  assign w6633 = w2791 & w6632 ;
  assign w6634 = w6299 | w6304 ;
  assign w6635 = w6515 & ~w6634 ;
  assign w6636 = w6302 ^ w6635 ;
  assign w6637 = ( ~w2791 & w6625 ) | ( ~w2791 & w6631 ) | ( w6625 & w6631 ) ;
  assign w6638 = ~w6625 & w6637 ;
  assign w6639 = w6636 | w6638 ;
  assign w6640 = ( w2585 & w6633 ) | ( w2585 & ~w6639 ) | ( w6633 & ~w6639 ) ;
  assign w6641 = w2585 & w6640 ;
  assign w6642 = w6307 | w6312 ;
  assign w6643 = w6515 & ~w6642 ;
  assign w6644 = w6310 ^ w6643 ;
  assign w6645 = ( ~w2585 & w6633 ) | ( ~w2585 & w6639 ) | ( w6633 & w6639 ) ;
  assign w6646 = ~w6633 & w6645 ;
  assign w6647 = w6644 | w6646 ;
  assign w6648 = ( w2387 & w6641 ) | ( w2387 & ~w6647 ) | ( w6641 & ~w6647 ) ;
  assign w6649 = w2387 & w6648 ;
  assign w6650 = w6315 | w6320 ;
  assign w6651 = w6515 & ~w6650 ;
  assign w6652 = w6318 ^ w6651 ;
  assign w6653 = ( ~w2387 & w6641 ) | ( ~w2387 & w6647 ) | ( w6641 & w6647 ) ;
  assign w6654 = ~w6641 & w6653 ;
  assign w6655 = w6652 | w6654 ;
  assign w6656 = ( w2197 & w6649 ) | ( w2197 & ~w6655 ) | ( w6649 & ~w6655 ) ;
  assign w6657 = w2197 & w6656 ;
  assign w6658 = w6323 | w6328 ;
  assign w6659 = w6515 & ~w6658 ;
  assign w6660 = w6326 ^ w6659 ;
  assign w6661 = ( ~w2197 & w6649 ) | ( ~w2197 & w6655 ) | ( w6649 & w6655 ) ;
  assign w6662 = ~w6649 & w6661 ;
  assign w6663 = w6660 | w6662 ;
  assign w6664 = ( w2015 & w6657 ) | ( w2015 & ~w6663 ) | ( w6657 & ~w6663 ) ;
  assign w6665 = w2015 & w6664 ;
  assign w6666 = w6331 | w6336 ;
  assign w6667 = w6515 & ~w6666 ;
  assign w6668 = w6334 ^ w6667 ;
  assign w6669 = ( ~w2015 & w6657 ) | ( ~w2015 & w6663 ) | ( w6657 & w6663 ) ;
  assign w6670 = ~w6657 & w6669 ;
  assign w6671 = w6668 | w6670 ;
  assign w6672 = ( w1841 & w6665 ) | ( w1841 & ~w6671 ) | ( w6665 & ~w6671 ) ;
  assign w6673 = w1841 & w6672 ;
  assign w6674 = w6339 | w6344 ;
  assign w6675 = w6515 & ~w6674 ;
  assign w6676 = w6342 ^ w6675 ;
  assign w6677 = ( ~w1841 & w6665 ) | ( ~w1841 & w6671 ) | ( w6665 & w6671 ) ;
  assign w6678 = ~w6665 & w6677 ;
  assign w6679 = w6676 | w6678 ;
  assign w6680 = ( w1675 & w6673 ) | ( w1675 & ~w6679 ) | ( w6673 & ~w6679 ) ;
  assign w6681 = w1675 & w6680 ;
  assign w6682 = w6347 | w6352 ;
  assign w6683 = w6515 & ~w6682 ;
  assign w6684 = w6350 ^ w6683 ;
  assign w6685 = ( ~w1675 & w6673 ) | ( ~w1675 & w6679 ) | ( w6673 & w6679 ) ;
  assign w6686 = ~w6673 & w6685 ;
  assign w6687 = w6684 | w6686 ;
  assign w6688 = ( w1517 & w6681 ) | ( w1517 & ~w6687 ) | ( w6681 & ~w6687 ) ;
  assign w6689 = w1517 & w6688 ;
  assign w6690 = w6355 | w6360 ;
  assign w6691 = w6515 & ~w6690 ;
  assign w6692 = w6358 ^ w6691 ;
  assign w6693 = ( ~w1517 & w6681 ) | ( ~w1517 & w6687 ) | ( w6681 & w6687 ) ;
  assign w6694 = ~w6681 & w6693 ;
  assign w6695 = w6692 | w6694 ;
  assign w6696 = ( w1367 & w6689 ) | ( w1367 & ~w6695 ) | ( w6689 & ~w6695 ) ;
  assign w6697 = w1367 & w6696 ;
  assign w6698 = w6363 | w6368 ;
  assign w6699 = w6515 & ~w6698 ;
  assign w6700 = w6366 ^ w6699 ;
  assign w6701 = ( ~w1367 & w6689 ) | ( ~w1367 & w6695 ) | ( w6689 & w6695 ) ;
  assign w6702 = ~w6689 & w6701 ;
  assign w6703 = w6700 | w6702 ;
  assign w6704 = ( w1225 & w6697 ) | ( w1225 & ~w6703 ) | ( w6697 & ~w6703 ) ;
  assign w6705 = w1225 & w6704 ;
  assign w6706 = w6371 | w6376 ;
  assign w6707 = w6515 & ~w6706 ;
  assign w6708 = w6374 ^ w6707 ;
  assign w6709 = ( ~w1225 & w6697 ) | ( ~w1225 & w6703 ) | ( w6697 & w6703 ) ;
  assign w6710 = ~w6697 & w6709 ;
  assign w6711 = w6708 | w6710 ;
  assign w6712 = ( w1091 & w6705 ) | ( w1091 & ~w6711 ) | ( w6705 & ~w6711 ) ;
  assign w6713 = w1091 & w6712 ;
  assign w6714 = w6379 | w6384 ;
  assign w6715 = w6515 & ~w6714 ;
  assign w6716 = w6382 ^ w6715 ;
  assign w6717 = ( ~w1091 & w6705 ) | ( ~w1091 & w6711 ) | ( w6705 & w6711 ) ;
  assign w6718 = ~w6705 & w6717 ;
  assign w6719 = w6716 | w6718 ;
  assign w6720 = ( w965 & w6713 ) | ( w965 & ~w6719 ) | ( w6713 & ~w6719 ) ;
  assign w6721 = w965 & w6720 ;
  assign w6722 = w6387 | w6392 ;
  assign w6723 = w6515 & ~w6722 ;
  assign w6724 = w6390 ^ w6723 ;
  assign w6725 = ( ~w965 & w6713 ) | ( ~w965 & w6719 ) | ( w6713 & w6719 ) ;
  assign w6726 = ~w6713 & w6725 ;
  assign w6727 = w6724 | w6726 ;
  assign w6728 = ( w847 & w6721 ) | ( w847 & ~w6727 ) | ( w6721 & ~w6727 ) ;
  assign w6729 = w847 & w6728 ;
  assign w6730 = w6395 | w6400 ;
  assign w6731 = w6515 & ~w6730 ;
  assign w6732 = w6398 ^ w6731 ;
  assign w6733 = ( ~w847 & w6721 ) | ( ~w847 & w6727 ) | ( w6721 & w6727 ) ;
  assign w6734 = ~w6721 & w6733 ;
  assign w6735 = w6732 | w6734 ;
  assign w6736 = ( w737 & w6729 ) | ( w737 & ~w6735 ) | ( w6729 & ~w6735 ) ;
  assign w6737 = w737 & w6736 ;
  assign w6738 = w6403 | w6408 ;
  assign w6739 = w6515 & ~w6738 ;
  assign w6740 = w6406 ^ w6739 ;
  assign w6741 = ( ~w737 & w6729 ) | ( ~w737 & w6735 ) | ( w6729 & w6735 ) ;
  assign w6742 = ~w6729 & w6741 ;
  assign w6743 = w6740 | w6742 ;
  assign w6744 = ( w635 & w6737 ) | ( w635 & ~w6743 ) | ( w6737 & ~w6743 ) ;
  assign w6745 = w635 & w6744 ;
  assign w6746 = w6411 | w6416 ;
  assign w6747 = w6515 & ~w6746 ;
  assign w6748 = w6414 ^ w6747 ;
  assign w6749 = ( ~w635 & w6737 ) | ( ~w635 & w6743 ) | ( w6737 & w6743 ) ;
  assign w6750 = ~w6737 & w6749 ;
  assign w6751 = w6748 | w6750 ;
  assign w6752 = ( w541 & w6745 ) | ( w541 & ~w6751 ) | ( w6745 & ~w6751 ) ;
  assign w6753 = w541 & w6752 ;
  assign w6754 = w6419 | w6424 ;
  assign w6755 = w6515 & ~w6754 ;
  assign w6756 = w6422 ^ w6755 ;
  assign w6757 = ( ~w541 & w6745 ) | ( ~w541 & w6751 ) | ( w6745 & w6751 ) ;
  assign w6758 = ~w6745 & w6757 ;
  assign w6759 = w6756 | w6758 ;
  assign w6760 = ( w455 & w6753 ) | ( w455 & ~w6759 ) | ( w6753 & ~w6759 ) ;
  assign w6761 = w455 & w6760 ;
  assign w6762 = w6427 | w6432 ;
  assign w6763 = w6515 & ~w6762 ;
  assign w6764 = w6430 ^ w6763 ;
  assign w6765 = ( ~w455 & w6753 ) | ( ~w455 & w6759 ) | ( w6753 & w6759 ) ;
  assign w6766 = ~w6753 & w6765 ;
  assign w6767 = w6764 | w6766 ;
  assign w6768 = ( w377 & w6761 ) | ( w377 & ~w6767 ) | ( w6761 & ~w6767 ) ;
  assign w6769 = w377 & w6768 ;
  assign w6770 = w6435 | w6440 ;
  assign w6771 = w6515 & ~w6770 ;
  assign w6772 = w6438 ^ w6771 ;
  assign w6773 = ( ~w377 & w6761 ) | ( ~w377 & w6767 ) | ( w6761 & w6767 ) ;
  assign w6774 = ~w6761 & w6773 ;
  assign w6775 = w6772 | w6774 ;
  assign w6776 = ( w307 & w6769 ) | ( w307 & ~w6775 ) | ( w6769 & ~w6775 ) ;
  assign w6777 = w307 & w6776 ;
  assign w6778 = w6443 | w6448 ;
  assign w6779 = w6515 & ~w6778 ;
  assign w6780 = w6446 ^ w6779 ;
  assign w6781 = ( ~w307 & w6769 ) | ( ~w307 & w6775 ) | ( w6769 & w6775 ) ;
  assign w6782 = ~w6769 & w6781 ;
  assign w6783 = w6780 | w6782 ;
  assign w6784 = ( w246 & w6777 ) | ( w246 & ~w6783 ) | ( w6777 & ~w6783 ) ;
  assign w6785 = w246 & w6784 ;
  assign w6786 = w6451 | w6456 ;
  assign w6787 = w6515 & ~w6786 ;
  assign w6788 = w6454 ^ w6787 ;
  assign w6789 = ( ~w246 & w6777 ) | ( ~w246 & w6783 ) | ( w6777 & w6783 ) ;
  assign w6790 = ~w6777 & w6789 ;
  assign w6791 = w6788 | w6790 ;
  assign w6792 = ( w185 & w6785 ) | ( w185 & ~w6791 ) | ( w6785 & ~w6791 ) ;
  assign w6793 = w185 & w6792 ;
  assign w6794 = w6459 | w6464 ;
  assign w6795 = w6515 & ~w6794 ;
  assign w6796 = w6462 ^ w6795 ;
  assign w6797 = ( ~w185 & w6785 ) | ( ~w185 & w6791 ) | ( w6785 & w6791 ) ;
  assign w6798 = ~w6785 & w6797 ;
  assign w6799 = w6796 | w6798 ;
  assign w6800 = ( w145 & w6793 ) | ( w145 & ~w6799 ) | ( w6793 & ~w6799 ) ;
  assign w6801 = w145 & w6800 ;
  assign w6802 = w6467 | w6472 ;
  assign w6803 = w6515 & ~w6802 ;
  assign w6804 = w6470 ^ w6803 ;
  assign w6805 = ( ~w145 & w6793 ) | ( ~w145 & w6799 ) | ( w6793 & w6799 ) ;
  assign w6806 = ~w6793 & w6805 ;
  assign w6807 = w6804 | w6806 ;
  assign w6808 = ( w132 & w6801 ) | ( w132 & ~w6807 ) | ( w6801 & ~w6807 ) ;
  assign w6809 = w132 & w6808 ;
  assign w6810 = w6475 | w6480 ;
  assign w6811 = w6515 & ~w6810 ;
  assign w6812 = w6478 ^ w6811 ;
  assign w6813 = ( ~w132 & w6801 ) | ( ~w132 & w6807 ) | ( w6801 & w6807 ) ;
  assign w6814 = ~w6801 & w6813 ;
  assign w6815 = w6812 | w6814 ;
  assign w6816 = ~w6809 & w6815 ;
  assign w6817 = w6483 | w6488 ;
  assign w6818 = w6515 & ~w6817 ;
  assign w6819 = w6486 ^ w6818 ;
  assign w6820 = ( ~w6501 & w6816 ) | ( ~w6501 & w6819 ) | ( w6816 & w6819 ) ;
  assign w6821 = w6490 & ~w6820 ;
  assign w6822 = ~w6493 & w6515 ;
  assign w6823 = ( w6820 & ~w6821 ) | ( w6820 & w6822 ) | ( ~w6821 & w6822 ) ;
  assign w6824 = w6501 | w6823 ;
  assign w6825 = ~w129 & w6824 ;
  assign w6826 = ( w6809 & w6815 ) | ( w6809 & w6819 ) | ( w6815 & w6819 ) ;
  assign w6827 = ~w6809 & w6826 ;
  assign w6828 = ( w129 & w6490 ) | ( w129 & w6493 ) | ( w6490 & w6493 ) ;
  assign w6829 = ( w6493 & ~w6515 ) | ( w6493 & w6828 ) | ( ~w6515 & w6828 ) ;
  assign w6830 = w6490 & w6829 ;
  assign w6831 = w6828 ^ w6830 ;
  assign w6832 = ( w6165 & w6170 ) | ( w6165 & w6197 ) | ( w6170 & w6197 ) ;
  assign w6833 = w6197 & ~w6832 ;
  assign w6834 = w6168 ^ w6833 ;
  assign w6835 = ( ~w6505 & w6512 ) | ( ~w6505 & w6834 ) | ( w6512 & w6834 ) ;
  assign w6836 = ~w6512 & w6835 ;
  assign w6837 = ( ~w6499 & w6501 ) | ( ~w6499 & w6836 ) | ( w6501 & w6836 ) ;
  assign w6838 = ~w6501 & w6837 ;
  assign w6839 = w6827 | w6838 ;
  assign w6840 = ( w6825 & ~w6827 ) | ( w6825 & w6831 ) | ( ~w6827 & w6831 ) ;
  assign w6841 = w6839 | w6840 ;
  assign w6842 = ( ~\pi049 & \pi050 ) | ( ~\pi049 & w6515 ) | ( \pi050 & w6515 ) ;
  assign w6843 = ( ~\pi048 & \pi050 ) | ( ~\pi048 & w6842 ) | ( \pi050 & w6842 ) ;
  assign w6844 = ( ~\pi050 & w6515 ) | ( ~\pi050 & w6841 ) | ( w6515 & w6841 ) ;
  assign w6845 = w6843 & w6844 ;
  assign w6846 = ( w6501 & w6505 ) | ( w6501 & ~w6512 ) | ( w6505 & ~w6512 ) ;
  assign w6847 = \pi049 & ~w6846 ;
  assign w6848 = \pi048 | \pi050 ;
  assign w6849 = ( ~w6846 & w6847 ) | ( ~w6846 & w6848 ) | ( w6847 & w6848 ) ;
  assign w6850 = ~w6512 & w6849 ;
  assign w6851 = ~w6499 & w6850 ;
  assign w6852 = ( \pi050 & w6841 ) | ( \pi050 & ~w6850 ) | ( w6841 & ~w6850 ) ;
  assign w6853 = w6851 & ~w6852 ;
  assign w6854 = ~\pi050 & w6841 ;
  assign w6855 = \pi051 ^ w6854 ;
  assign w6856 = w6853 | w6855 ;
  assign w6857 = ( w6197 & w6845 ) | ( w6197 & ~w6856 ) | ( w6845 & ~w6856 ) ;
  assign w6858 = w6197 & w6857 ;
  assign w6859 = ( ~w6197 & w6845 ) | ( ~w6197 & w6856 ) | ( w6845 & w6856 ) ;
  assign w6860 = ~w6845 & w6859 ;
  assign w6861 = w6515 & ~w6838 ;
  assign w6862 = ~w6827 & w6861 ;
  assign w6863 = ~w6840 & w6862 ;
  assign w6864 = \pi051 & w6841 ;
  assign w6865 = ( \pi050 & w6841 ) | ( \pi050 & ~w6864 ) | ( w6841 & ~w6864 ) ;
  assign w6866 = ( ~\pi050 & w6863 ) | ( ~\pi050 & w6865 ) | ( w6863 & w6865 ) ;
  assign w6867 = \pi052 ^ w6866 ;
  assign w6868 = w6860 | w6867 ;
  assign w6869 = ( w5887 & w6858 ) | ( w5887 & ~w6868 ) | ( w6858 & ~w6868 ) ;
  assign w6870 = w5887 & w6869 ;
  assign w6871 = ( w6519 & ~w6527 ) | ( w6519 & w6841 ) | ( ~w6527 & w6841 ) ;
  assign w6872 = ~w6519 & w6871 ;
  assign w6873 = \pi053 ^ w6872 ;
  assign w6874 = w6528 ^ w6873 ;
  assign w6875 = ( ~w5887 & w6858 ) | ( ~w5887 & w6868 ) | ( w6858 & w6868 ) ;
  assign w6876 = ~w6858 & w6875 ;
  assign w6877 = w6874 | w6876 ;
  assign w6878 = ( w5585 & w6870 ) | ( w5585 & ~w6877 ) | ( w6870 & ~w6877 ) ;
  assign w6879 = w5585 & w6878 ;
  assign w6880 = w6532 | w6534 ;
  assign w6881 = w6841 & ~w6880 ;
  assign w6882 = w6541 ^ w6881 ;
  assign w6883 = ( ~w5585 & w6870 ) | ( ~w5585 & w6877 ) | ( w6870 & w6877 ) ;
  assign w6884 = ~w6870 & w6883 ;
  assign w6885 = w6882 | w6884 ;
  assign w6886 = ( w5291 & w6879 ) | ( w5291 & ~w6885 ) | ( w6879 & ~w6885 ) ;
  assign w6887 = w5291 & w6886 ;
  assign w6888 = w6544 | w6550 ;
  assign w6889 = w6841 & ~w6888 ;
  assign w6890 = w6548 ^ w6889 ;
  assign w6891 = ( ~w5291 & w6879 ) | ( ~w5291 & w6885 ) | ( w6879 & w6885 ) ;
  assign w6892 = ~w6879 & w6891 ;
  assign w6893 = w6890 | w6892 ;
  assign w6894 = ( w5005 & w6887 ) | ( w5005 & ~w6893 ) | ( w6887 & ~w6893 ) ;
  assign w6895 = w5005 & w6894 ;
  assign w6896 = w6553 | w6558 ;
  assign w6897 = w6841 & ~w6896 ;
  assign w6898 = w6556 ^ w6897 ;
  assign w6899 = ( ~w5005 & w6887 ) | ( ~w5005 & w6893 ) | ( w6887 & w6893 ) ;
  assign w6900 = ~w6887 & w6899 ;
  assign w6901 = w6898 | w6900 ;
  assign w6902 = ( w4727 & w6895 ) | ( w4727 & ~w6901 ) | ( w6895 & ~w6901 ) ;
  assign w6903 = w4727 & w6902 ;
  assign w6904 = w6561 | w6566 ;
  assign w6905 = w6841 & ~w6904 ;
  assign w6906 = w6564 ^ w6905 ;
  assign w6907 = ( ~w4727 & w6895 ) | ( ~w4727 & w6901 ) | ( w6895 & w6901 ) ;
  assign w6908 = ~w6895 & w6907 ;
  assign w6909 = w6906 | w6908 ;
  assign w6910 = ( w4457 & w6903 ) | ( w4457 & ~w6909 ) | ( w6903 & ~w6909 ) ;
  assign w6911 = w4457 & w6910 ;
  assign w6912 = w6569 | w6574 ;
  assign w6913 = w6841 & ~w6912 ;
  assign w6914 = w6572 ^ w6913 ;
  assign w6915 = ( ~w4457 & w6903 ) | ( ~w4457 & w6909 ) | ( w6903 & w6909 ) ;
  assign w6916 = ~w6903 & w6915 ;
  assign w6917 = w6914 | w6916 ;
  assign w6918 = ( w4195 & w6911 ) | ( w4195 & ~w6917 ) | ( w6911 & ~w6917 ) ;
  assign w6919 = w4195 & w6918 ;
  assign w6920 = w6577 | w6582 ;
  assign w6921 = w6841 & ~w6920 ;
  assign w6922 = w6580 ^ w6921 ;
  assign w6923 = ( ~w4195 & w6911 ) | ( ~w4195 & w6917 ) | ( w6911 & w6917 ) ;
  assign w6924 = ~w6911 & w6923 ;
  assign w6925 = w6922 | w6924 ;
  assign w6926 = ( w3941 & w6919 ) | ( w3941 & ~w6925 ) | ( w6919 & ~w6925 ) ;
  assign w6927 = w3941 & w6926 ;
  assign w6928 = w6585 | w6590 ;
  assign w6929 = w6841 & ~w6928 ;
  assign w6930 = w6588 ^ w6929 ;
  assign w6931 = ( ~w3941 & w6919 ) | ( ~w3941 & w6925 ) | ( w6919 & w6925 ) ;
  assign w6932 = ~w6919 & w6931 ;
  assign w6933 = w6930 | w6932 ;
  assign w6934 = ( w3695 & w6927 ) | ( w3695 & ~w6933 ) | ( w6927 & ~w6933 ) ;
  assign w6935 = w3695 & w6934 ;
  assign w6936 = w6593 | w6598 ;
  assign w6937 = w6841 & ~w6936 ;
  assign w6938 = w6596 ^ w6937 ;
  assign w6939 = ( ~w3695 & w6927 ) | ( ~w3695 & w6933 ) | ( w6927 & w6933 ) ;
  assign w6940 = ~w6927 & w6939 ;
  assign w6941 = w6938 | w6940 ;
  assign w6942 = ( w3457 & w6935 ) | ( w3457 & ~w6941 ) | ( w6935 & ~w6941 ) ;
  assign w6943 = w3457 & w6942 ;
  assign w6944 = w6601 | w6606 ;
  assign w6945 = w6841 & ~w6944 ;
  assign w6946 = w6604 ^ w6945 ;
  assign w6947 = ( ~w3457 & w6935 ) | ( ~w3457 & w6941 ) | ( w6935 & w6941 ) ;
  assign w6948 = ~w6935 & w6947 ;
  assign w6949 = w6946 | w6948 ;
  assign w6950 = ( w3227 & w6943 ) | ( w3227 & ~w6949 ) | ( w6943 & ~w6949 ) ;
  assign w6951 = w3227 & w6950 ;
  assign w6952 = w6609 | w6614 ;
  assign w6953 = w6841 & ~w6952 ;
  assign w6954 = w6612 ^ w6953 ;
  assign w6955 = ( ~w3227 & w6943 ) | ( ~w3227 & w6949 ) | ( w6943 & w6949 ) ;
  assign w6956 = ~w6943 & w6955 ;
  assign w6957 = w6954 | w6956 ;
  assign w6958 = ( w3005 & w6951 ) | ( w3005 & ~w6957 ) | ( w6951 & ~w6957 ) ;
  assign w6959 = w3005 & w6958 ;
  assign w6960 = w6617 | w6622 ;
  assign w6961 = w6841 & ~w6960 ;
  assign w6962 = w6620 ^ w6961 ;
  assign w6963 = ( ~w3005 & w6951 ) | ( ~w3005 & w6957 ) | ( w6951 & w6957 ) ;
  assign w6964 = ~w6951 & w6963 ;
  assign w6965 = w6962 | w6964 ;
  assign w6966 = ( w2791 & w6959 ) | ( w2791 & ~w6965 ) | ( w6959 & ~w6965 ) ;
  assign w6967 = w2791 & w6966 ;
  assign w6968 = ( ~w2791 & w6959 ) | ( ~w2791 & w6965 ) | ( w6959 & w6965 ) ;
  assign w6969 = ~w6959 & w6968 ;
  assign w6970 = w6625 | w6627 ;
  assign w6971 = w6841 & ~w6970 ;
  assign w6972 = w6630 ^ w6971 ;
  assign w6973 = w6969 | w6972 ;
  assign w6974 = ( w2585 & w6967 ) | ( w2585 & ~w6973 ) | ( w6967 & ~w6973 ) ;
  assign w6975 = w2585 & w6974 ;
  assign w6976 = w6633 | w6638 ;
  assign w6977 = w6841 & ~w6976 ;
  assign w6978 = w6636 ^ w6977 ;
  assign w6979 = ( ~w2585 & w6967 ) | ( ~w2585 & w6973 ) | ( w6967 & w6973 ) ;
  assign w6980 = ~w6967 & w6979 ;
  assign w6981 = w6978 | w6980 ;
  assign w6982 = ( w2387 & w6975 ) | ( w2387 & ~w6981 ) | ( w6975 & ~w6981 ) ;
  assign w6983 = w2387 & w6982 ;
  assign w6984 = w6641 | w6646 ;
  assign w6985 = w6841 & ~w6984 ;
  assign w6986 = w6644 ^ w6985 ;
  assign w6987 = ( ~w2387 & w6975 ) | ( ~w2387 & w6981 ) | ( w6975 & w6981 ) ;
  assign w6988 = ~w6975 & w6987 ;
  assign w6989 = w6986 | w6988 ;
  assign w6990 = ( w2197 & w6983 ) | ( w2197 & ~w6989 ) | ( w6983 & ~w6989 ) ;
  assign w6991 = w2197 & w6990 ;
  assign w6992 = w6649 | w6654 ;
  assign w6993 = w6841 & ~w6992 ;
  assign w6994 = w6652 ^ w6993 ;
  assign w6995 = ( ~w2197 & w6983 ) | ( ~w2197 & w6989 ) | ( w6983 & w6989 ) ;
  assign w6996 = ~w6983 & w6995 ;
  assign w6997 = w6994 | w6996 ;
  assign w6998 = ( w2015 & w6991 ) | ( w2015 & ~w6997 ) | ( w6991 & ~w6997 ) ;
  assign w6999 = w2015 & w6998 ;
  assign w7000 = w6657 | w6662 ;
  assign w7001 = w6841 & ~w7000 ;
  assign w7002 = w6660 ^ w7001 ;
  assign w7003 = ( ~w2015 & w6991 ) | ( ~w2015 & w6997 ) | ( w6991 & w6997 ) ;
  assign w7004 = ~w6991 & w7003 ;
  assign w7005 = w7002 | w7004 ;
  assign w7006 = ( w1841 & w6999 ) | ( w1841 & ~w7005 ) | ( w6999 & ~w7005 ) ;
  assign w7007 = w1841 & w7006 ;
  assign w7008 = w6665 | w6670 ;
  assign w7009 = w6841 & ~w7008 ;
  assign w7010 = w6668 ^ w7009 ;
  assign w7011 = ( ~w1841 & w6999 ) | ( ~w1841 & w7005 ) | ( w6999 & w7005 ) ;
  assign w7012 = ~w6999 & w7011 ;
  assign w7013 = w7010 | w7012 ;
  assign w7014 = ( w1675 & w7007 ) | ( w1675 & ~w7013 ) | ( w7007 & ~w7013 ) ;
  assign w7015 = w1675 & w7014 ;
  assign w7016 = w6673 | w6678 ;
  assign w7017 = w6841 & ~w7016 ;
  assign w7018 = w6676 ^ w7017 ;
  assign w7019 = ( ~w1675 & w7007 ) | ( ~w1675 & w7013 ) | ( w7007 & w7013 ) ;
  assign w7020 = ~w7007 & w7019 ;
  assign w7021 = w7018 | w7020 ;
  assign w7022 = ( w1517 & w7015 ) | ( w1517 & ~w7021 ) | ( w7015 & ~w7021 ) ;
  assign w7023 = w1517 & w7022 ;
  assign w7024 = w6681 | w6686 ;
  assign w7025 = w6841 & ~w7024 ;
  assign w7026 = w6684 ^ w7025 ;
  assign w7027 = ( ~w1517 & w7015 ) | ( ~w1517 & w7021 ) | ( w7015 & w7021 ) ;
  assign w7028 = ~w7015 & w7027 ;
  assign w7029 = w7026 | w7028 ;
  assign w7030 = ( w1367 & w7023 ) | ( w1367 & ~w7029 ) | ( w7023 & ~w7029 ) ;
  assign w7031 = w1367 & w7030 ;
  assign w7032 = w6689 | w6694 ;
  assign w7033 = w6841 & ~w7032 ;
  assign w7034 = w6692 ^ w7033 ;
  assign w7035 = ( ~w1367 & w7023 ) | ( ~w1367 & w7029 ) | ( w7023 & w7029 ) ;
  assign w7036 = ~w7023 & w7035 ;
  assign w7037 = w7034 | w7036 ;
  assign w7038 = ( w1225 & w7031 ) | ( w1225 & ~w7037 ) | ( w7031 & ~w7037 ) ;
  assign w7039 = w1225 & w7038 ;
  assign w7040 = w6697 | w6702 ;
  assign w7041 = w6841 & ~w7040 ;
  assign w7042 = w6700 ^ w7041 ;
  assign w7043 = ( ~w1225 & w7031 ) | ( ~w1225 & w7037 ) | ( w7031 & w7037 ) ;
  assign w7044 = ~w7031 & w7043 ;
  assign w7045 = w7042 | w7044 ;
  assign w7046 = ( w1091 & w7039 ) | ( w1091 & ~w7045 ) | ( w7039 & ~w7045 ) ;
  assign w7047 = w1091 & w7046 ;
  assign w7048 = w6705 | w6710 ;
  assign w7049 = w6841 & ~w7048 ;
  assign w7050 = w6708 ^ w7049 ;
  assign w7051 = ( ~w1091 & w7039 ) | ( ~w1091 & w7045 ) | ( w7039 & w7045 ) ;
  assign w7052 = ~w7039 & w7051 ;
  assign w7053 = w7050 | w7052 ;
  assign w7054 = ( w965 & w7047 ) | ( w965 & ~w7053 ) | ( w7047 & ~w7053 ) ;
  assign w7055 = w965 & w7054 ;
  assign w7056 = w6713 | w6718 ;
  assign w7057 = w6841 & ~w7056 ;
  assign w7058 = w6716 ^ w7057 ;
  assign w7059 = ( ~w965 & w7047 ) | ( ~w965 & w7053 ) | ( w7047 & w7053 ) ;
  assign w7060 = ~w7047 & w7059 ;
  assign w7061 = w7058 | w7060 ;
  assign w7062 = ( w847 & w7055 ) | ( w847 & ~w7061 ) | ( w7055 & ~w7061 ) ;
  assign w7063 = w847 & w7062 ;
  assign w7064 = w6721 | w6726 ;
  assign w7065 = w6841 & ~w7064 ;
  assign w7066 = w6724 ^ w7065 ;
  assign w7067 = ( ~w847 & w7055 ) | ( ~w847 & w7061 ) | ( w7055 & w7061 ) ;
  assign w7068 = ~w7055 & w7067 ;
  assign w7069 = w7066 | w7068 ;
  assign w7070 = ( w737 & w7063 ) | ( w737 & ~w7069 ) | ( w7063 & ~w7069 ) ;
  assign w7071 = w737 & w7070 ;
  assign w7072 = w6729 | w6734 ;
  assign w7073 = w6841 & ~w7072 ;
  assign w7074 = w6732 ^ w7073 ;
  assign w7075 = ( ~w737 & w7063 ) | ( ~w737 & w7069 ) | ( w7063 & w7069 ) ;
  assign w7076 = ~w7063 & w7075 ;
  assign w7077 = w7074 | w7076 ;
  assign w7078 = ( w635 & w7071 ) | ( w635 & ~w7077 ) | ( w7071 & ~w7077 ) ;
  assign w7079 = w635 & w7078 ;
  assign w7080 = w6737 | w6742 ;
  assign w7081 = w6841 & ~w7080 ;
  assign w7082 = w6740 ^ w7081 ;
  assign w7083 = ( ~w635 & w7071 ) | ( ~w635 & w7077 ) | ( w7071 & w7077 ) ;
  assign w7084 = ~w7071 & w7083 ;
  assign w7085 = w7082 | w7084 ;
  assign w7086 = ( w541 & w7079 ) | ( w541 & ~w7085 ) | ( w7079 & ~w7085 ) ;
  assign w7087 = w541 & w7086 ;
  assign w7088 = w6745 | w6750 ;
  assign w7089 = w6841 & ~w7088 ;
  assign w7090 = w6748 ^ w7089 ;
  assign w7091 = ( ~w541 & w7079 ) | ( ~w541 & w7085 ) | ( w7079 & w7085 ) ;
  assign w7092 = ~w7079 & w7091 ;
  assign w7093 = w7090 | w7092 ;
  assign w7094 = ( w455 & w7087 ) | ( w455 & ~w7093 ) | ( w7087 & ~w7093 ) ;
  assign w7095 = w455 & w7094 ;
  assign w7096 = w6753 | w6758 ;
  assign w7097 = w6841 & ~w7096 ;
  assign w7098 = w6756 ^ w7097 ;
  assign w7099 = ( ~w455 & w7087 ) | ( ~w455 & w7093 ) | ( w7087 & w7093 ) ;
  assign w7100 = ~w7087 & w7099 ;
  assign w7101 = w7098 | w7100 ;
  assign w7102 = ( w377 & w7095 ) | ( w377 & ~w7101 ) | ( w7095 & ~w7101 ) ;
  assign w7103 = w377 & w7102 ;
  assign w7104 = w6761 | w6766 ;
  assign w7105 = w6841 & ~w7104 ;
  assign w7106 = w6764 ^ w7105 ;
  assign w7107 = ( ~w377 & w7095 ) | ( ~w377 & w7101 ) | ( w7095 & w7101 ) ;
  assign w7108 = ~w7095 & w7107 ;
  assign w7109 = w7106 | w7108 ;
  assign w7110 = ( w307 & w7103 ) | ( w307 & ~w7109 ) | ( w7103 & ~w7109 ) ;
  assign w7111 = w307 & w7110 ;
  assign w7112 = w6769 | w6774 ;
  assign w7113 = w6841 & ~w7112 ;
  assign w7114 = w6772 ^ w7113 ;
  assign w7115 = ( ~w307 & w7103 ) | ( ~w307 & w7109 ) | ( w7103 & w7109 ) ;
  assign w7116 = ~w7103 & w7115 ;
  assign w7117 = w7114 | w7116 ;
  assign w7118 = ( w246 & w7111 ) | ( w246 & ~w7117 ) | ( w7111 & ~w7117 ) ;
  assign w7119 = w246 & w7118 ;
  assign w7120 = w6777 | w6782 ;
  assign w7121 = w6841 & ~w7120 ;
  assign w7122 = w6780 ^ w7121 ;
  assign w7123 = ( ~w246 & w7111 ) | ( ~w246 & w7117 ) | ( w7111 & w7117 ) ;
  assign w7124 = ~w7111 & w7123 ;
  assign w7125 = w7122 | w7124 ;
  assign w7126 = ( w185 & w7119 ) | ( w185 & ~w7125 ) | ( w7119 & ~w7125 ) ;
  assign w7127 = w185 & w7126 ;
  assign w7128 = w6785 | w6790 ;
  assign w7129 = w6841 & ~w7128 ;
  assign w7130 = w6788 ^ w7129 ;
  assign w7131 = ( ~w185 & w7119 ) | ( ~w185 & w7125 ) | ( w7119 & w7125 ) ;
  assign w7132 = ~w7119 & w7131 ;
  assign w7133 = w7130 | w7132 ;
  assign w7134 = ( w145 & w7127 ) | ( w145 & ~w7133 ) | ( w7127 & ~w7133 ) ;
  assign w7135 = w145 & w7134 ;
  assign w7136 = w6793 | w6798 ;
  assign w7137 = w6841 & ~w7136 ;
  assign w7138 = w6796 ^ w7137 ;
  assign w7139 = ( ~w145 & w7127 ) | ( ~w145 & w7133 ) | ( w7127 & w7133 ) ;
  assign w7140 = ~w7127 & w7139 ;
  assign w7141 = w7138 | w7140 ;
  assign w7142 = ( w132 & w7135 ) | ( w132 & ~w7141 ) | ( w7135 & ~w7141 ) ;
  assign w7143 = w132 & w7142 ;
  assign w7144 = w6801 | w6806 ;
  assign w7145 = w6841 & ~w7144 ;
  assign w7146 = w6804 ^ w7145 ;
  assign w7147 = ( ~w132 & w7135 ) | ( ~w132 & w7141 ) | ( w7135 & w7141 ) ;
  assign w7148 = ~w7135 & w7147 ;
  assign w7149 = w7146 | w7148 ;
  assign w7150 = ~w7143 & w7149 ;
  assign w7151 = w6809 | w6814 ;
  assign w7152 = w6841 & ~w7151 ;
  assign w7153 = w6812 ^ w7152 ;
  assign w7154 = ( ~w6827 & w7150 ) | ( ~w6827 & w7153 ) | ( w7150 & w7153 ) ;
  assign w7155 = w6816 & ~w7154 ;
  assign w7156 = ~w6819 & w6841 ;
  assign w7157 = ( w7154 & ~w7155 ) | ( w7154 & w7156 ) | ( ~w7155 & w7156 ) ;
  assign w7158 = w6827 | w7157 ;
  assign w7159 = ~w129 & w7158 ;
  assign w7160 = ( w7143 & w7149 ) | ( w7143 & w7153 ) | ( w7149 & w7153 ) ;
  assign w7161 = ~w7143 & w7160 ;
  assign w7162 = ( w129 & w6816 ) | ( w129 & w6819 ) | ( w6816 & w6819 ) ;
  assign w7163 = ( w6819 & ~w6841 ) | ( w6819 & w7162 ) | ( ~w6841 & w7162 ) ;
  assign w7164 = w6816 & w7163 ;
  assign w7165 = w7162 ^ w7164 ;
  assign w7166 = ( w6483 & w6488 ) | ( w6483 & w6515 ) | ( w6488 & w6515 ) ;
  assign w7167 = w6515 & ~w7166 ;
  assign w7168 = w6486 ^ w7167 ;
  assign w7169 = ( ~w6831 & w6838 ) | ( ~w6831 & w7168 ) | ( w6838 & w7168 ) ;
  assign w7170 = ~w6838 & w7169 ;
  assign w7171 = ( ~w6825 & w6827 ) | ( ~w6825 & w7170 ) | ( w6827 & w7170 ) ;
  assign w7172 = ~w6827 & w7171 ;
  assign w7173 = w7161 | w7172 ;
  assign w7174 = ( w7159 & ~w7161 ) | ( w7159 & w7165 ) | ( ~w7161 & w7165 ) ;
  assign w7175 = w7173 | w7174 ;
  assign w7176 = ( ~\pi047 & \pi048 ) | ( ~\pi047 & w6841 ) | ( \pi048 & w6841 ) ;
  assign w7177 = ( ~\pi046 & \pi048 ) | ( ~\pi046 & w7176 ) | ( \pi048 & w7176 ) ;
  assign w7178 = ( ~\pi048 & w6841 ) | ( ~\pi048 & w7175 ) | ( w6841 & w7175 ) ;
  assign w7179 = w7177 & w7178 ;
  assign w7180 = ( w6827 & w6831 ) | ( w6827 & ~w6838 ) | ( w6831 & ~w6838 ) ;
  assign w7181 = \pi047 & ~w7180 ;
  assign w7182 = \pi046 | \pi048 ;
  assign w7183 = ( ~w7180 & w7181 ) | ( ~w7180 & w7182 ) | ( w7181 & w7182 ) ;
  assign w7184 = ~w6838 & w7183 ;
  assign w7185 = ~w6825 & w7184 ;
  assign w7186 = ( \pi048 & w7175 ) | ( \pi048 & ~w7184 ) | ( w7175 & ~w7184 ) ;
  assign w7187 = w7185 & ~w7186 ;
  assign w7188 = ~\pi048 & w7175 ;
  assign w7189 = \pi049 ^ w7188 ;
  assign w7190 = w7187 | w7189 ;
  assign w7191 = ( w6515 & w7179 ) | ( w6515 & ~w7190 ) | ( w7179 & ~w7190 ) ;
  assign w7192 = w6515 & w7191 ;
  assign w7193 = ( ~w6515 & w7179 ) | ( ~w6515 & w7190 ) | ( w7179 & w7190 ) ;
  assign w7194 = ~w7179 & w7193 ;
  assign w7195 = w6841 & ~w7172 ;
  assign w7196 = ~w7161 & w7195 ;
  assign w7197 = ~w7174 & w7196 ;
  assign w7198 = \pi049 & w7175 ;
  assign w7199 = ( \pi048 & w7175 ) | ( \pi048 & ~w7198 ) | ( w7175 & ~w7198 ) ;
  assign w7200 = ( ~\pi048 & w7197 ) | ( ~\pi048 & w7199 ) | ( w7197 & w7199 ) ;
  assign w7201 = \pi050 ^ w7200 ;
  assign w7202 = w7194 | w7201 ;
  assign w7203 = ( w6197 & w7192 ) | ( w6197 & ~w7202 ) | ( w7192 & ~w7202 ) ;
  assign w7204 = w6197 & w7203 ;
  assign w7205 = ( w6845 & ~w6853 ) | ( w6845 & w7175 ) | ( ~w6853 & w7175 ) ;
  assign w7206 = ~w6845 & w7205 ;
  assign w7207 = \pi051 ^ w7206 ;
  assign w7208 = w6854 ^ w7207 ;
  assign w7209 = ( ~w6197 & w7192 ) | ( ~w6197 & w7202 ) | ( w7192 & w7202 ) ;
  assign w7210 = ~w7192 & w7209 ;
  assign w7211 = w7208 | w7210 ;
  assign w7212 = ( w5887 & w7204 ) | ( w5887 & ~w7211 ) | ( w7204 & ~w7211 ) ;
  assign w7213 = w5887 & w7212 ;
  assign w7214 = w6858 | w6860 ;
  assign w7215 = w7175 & ~w7214 ;
  assign w7216 = w6867 ^ w7215 ;
  assign w7217 = ( ~w5887 & w7204 ) | ( ~w5887 & w7211 ) | ( w7204 & w7211 ) ;
  assign w7218 = ~w7204 & w7217 ;
  assign w7219 = w7216 | w7218 ;
  assign w7220 = ( w5585 & w7213 ) | ( w5585 & ~w7219 ) | ( w7213 & ~w7219 ) ;
  assign w7221 = w5585 & w7220 ;
  assign w7222 = w6870 | w6876 ;
  assign w7223 = w7175 & ~w7222 ;
  assign w7224 = w6874 ^ w7223 ;
  assign w7225 = ( ~w5585 & w7213 ) | ( ~w5585 & w7219 ) | ( w7213 & w7219 ) ;
  assign w7226 = ~w7213 & w7225 ;
  assign w7227 = w7224 | w7226 ;
  assign w7228 = ( w5291 & w7221 ) | ( w5291 & ~w7227 ) | ( w7221 & ~w7227 ) ;
  assign w7229 = w5291 & w7228 ;
  assign w7230 = w6879 | w6884 ;
  assign w7231 = w7175 & ~w7230 ;
  assign w7232 = w6882 ^ w7231 ;
  assign w7233 = ( ~w5291 & w7221 ) | ( ~w5291 & w7227 ) | ( w7221 & w7227 ) ;
  assign w7234 = ~w7221 & w7233 ;
  assign w7235 = w7232 | w7234 ;
  assign w7236 = ( w5005 & w7229 ) | ( w5005 & ~w7235 ) | ( w7229 & ~w7235 ) ;
  assign w7237 = w5005 & w7236 ;
  assign w7238 = w6887 | w6892 ;
  assign w7239 = w7175 & ~w7238 ;
  assign w7240 = w6890 ^ w7239 ;
  assign w7241 = ( ~w5005 & w7229 ) | ( ~w5005 & w7235 ) | ( w7229 & w7235 ) ;
  assign w7242 = ~w7229 & w7241 ;
  assign w7243 = w7240 | w7242 ;
  assign w7244 = ( w4727 & w7237 ) | ( w4727 & ~w7243 ) | ( w7237 & ~w7243 ) ;
  assign w7245 = w4727 & w7244 ;
  assign w7246 = w6895 | w6900 ;
  assign w7247 = w7175 & ~w7246 ;
  assign w7248 = w6898 ^ w7247 ;
  assign w7249 = ( ~w4727 & w7237 ) | ( ~w4727 & w7243 ) | ( w7237 & w7243 ) ;
  assign w7250 = ~w7237 & w7249 ;
  assign w7251 = w7248 | w7250 ;
  assign w7252 = ( w4457 & w7245 ) | ( w4457 & ~w7251 ) | ( w7245 & ~w7251 ) ;
  assign w7253 = w4457 & w7252 ;
  assign w7254 = w6903 | w6908 ;
  assign w7255 = w7175 & ~w7254 ;
  assign w7256 = w6906 ^ w7255 ;
  assign w7257 = ( ~w4457 & w7245 ) | ( ~w4457 & w7251 ) | ( w7245 & w7251 ) ;
  assign w7258 = ~w7245 & w7257 ;
  assign w7259 = w7256 | w7258 ;
  assign w7260 = ( w4195 & w7253 ) | ( w4195 & ~w7259 ) | ( w7253 & ~w7259 ) ;
  assign w7261 = w4195 & w7260 ;
  assign w7262 = w6911 | w6916 ;
  assign w7263 = w7175 & ~w7262 ;
  assign w7264 = w6914 ^ w7263 ;
  assign w7265 = ( ~w4195 & w7253 ) | ( ~w4195 & w7259 ) | ( w7253 & w7259 ) ;
  assign w7266 = ~w7253 & w7265 ;
  assign w7267 = w7264 | w7266 ;
  assign w7268 = ( w3941 & w7261 ) | ( w3941 & ~w7267 ) | ( w7261 & ~w7267 ) ;
  assign w7269 = w3941 & w7268 ;
  assign w7270 = w6919 | w6924 ;
  assign w7271 = w7175 & ~w7270 ;
  assign w7272 = w6922 ^ w7271 ;
  assign w7273 = ( ~w3941 & w7261 ) | ( ~w3941 & w7267 ) | ( w7261 & w7267 ) ;
  assign w7274 = ~w7261 & w7273 ;
  assign w7275 = w7272 | w7274 ;
  assign w7276 = ( w3695 & w7269 ) | ( w3695 & ~w7275 ) | ( w7269 & ~w7275 ) ;
  assign w7277 = w3695 & w7276 ;
  assign w7278 = w6927 | w6932 ;
  assign w7279 = w7175 & ~w7278 ;
  assign w7280 = w6930 ^ w7279 ;
  assign w7281 = ( ~w3695 & w7269 ) | ( ~w3695 & w7275 ) | ( w7269 & w7275 ) ;
  assign w7282 = ~w7269 & w7281 ;
  assign w7283 = w7280 | w7282 ;
  assign w7284 = ( w3457 & w7277 ) | ( w3457 & ~w7283 ) | ( w7277 & ~w7283 ) ;
  assign w7285 = w3457 & w7284 ;
  assign w7286 = w6935 | w6940 ;
  assign w7287 = w7175 & ~w7286 ;
  assign w7288 = w6938 ^ w7287 ;
  assign w7289 = ( ~w3457 & w7277 ) | ( ~w3457 & w7283 ) | ( w7277 & w7283 ) ;
  assign w7290 = ~w7277 & w7289 ;
  assign w7291 = w7288 | w7290 ;
  assign w7292 = ( w3227 & w7285 ) | ( w3227 & ~w7291 ) | ( w7285 & ~w7291 ) ;
  assign w7293 = w3227 & w7292 ;
  assign w7294 = w6943 | w6948 ;
  assign w7295 = w7175 & ~w7294 ;
  assign w7296 = w6946 ^ w7295 ;
  assign w7297 = ( ~w3227 & w7285 ) | ( ~w3227 & w7291 ) | ( w7285 & w7291 ) ;
  assign w7298 = ~w7285 & w7297 ;
  assign w7299 = w7296 | w7298 ;
  assign w7300 = ( w3005 & w7293 ) | ( w3005 & ~w7299 ) | ( w7293 & ~w7299 ) ;
  assign w7301 = w3005 & w7300 ;
  assign w7302 = w6951 | w6956 ;
  assign w7303 = w7175 & ~w7302 ;
  assign w7304 = w6954 ^ w7303 ;
  assign w7305 = ( ~w3005 & w7293 ) | ( ~w3005 & w7299 ) | ( w7293 & w7299 ) ;
  assign w7306 = ~w7293 & w7305 ;
  assign w7307 = w7304 | w7306 ;
  assign w7308 = ( w2791 & w7301 ) | ( w2791 & ~w7307 ) | ( w7301 & ~w7307 ) ;
  assign w7309 = w2791 & w7308 ;
  assign w7310 = w6959 | w6964 ;
  assign w7311 = w7175 & ~w7310 ;
  assign w7312 = w6962 ^ w7311 ;
  assign w7313 = ( ~w2791 & w7301 ) | ( ~w2791 & w7307 ) | ( w7301 & w7307 ) ;
  assign w7314 = ~w7301 & w7313 ;
  assign w7315 = w7312 | w7314 ;
  assign w7316 = ( w2585 & w7309 ) | ( w2585 & ~w7315 ) | ( w7309 & ~w7315 ) ;
  assign w7317 = w2585 & w7316 ;
  assign w7318 = ( ~w2585 & w7309 ) | ( ~w2585 & w7315 ) | ( w7309 & w7315 ) ;
  assign w7319 = ~w7309 & w7318 ;
  assign w7320 = w6967 | w6969 ;
  assign w7321 = w7175 & ~w7320 ;
  assign w7322 = w6972 ^ w7321 ;
  assign w7323 = w7319 | w7322 ;
  assign w7324 = ( w2387 & w7317 ) | ( w2387 & ~w7323 ) | ( w7317 & ~w7323 ) ;
  assign w7325 = w2387 & w7324 ;
  assign w7326 = w6975 | w6980 ;
  assign w7327 = w7175 & ~w7326 ;
  assign w7328 = w6978 ^ w7327 ;
  assign w7329 = ( ~w2387 & w7317 ) | ( ~w2387 & w7323 ) | ( w7317 & w7323 ) ;
  assign w7330 = ~w7317 & w7329 ;
  assign w7331 = w7328 | w7330 ;
  assign w7332 = ( w2197 & w7325 ) | ( w2197 & ~w7331 ) | ( w7325 & ~w7331 ) ;
  assign w7333 = w2197 & w7332 ;
  assign w7334 = w6983 | w6988 ;
  assign w7335 = w7175 & ~w7334 ;
  assign w7336 = w6986 ^ w7335 ;
  assign w7337 = ( ~w2197 & w7325 ) | ( ~w2197 & w7331 ) | ( w7325 & w7331 ) ;
  assign w7338 = ~w7325 & w7337 ;
  assign w7339 = w7336 | w7338 ;
  assign w7340 = ( w2015 & w7333 ) | ( w2015 & ~w7339 ) | ( w7333 & ~w7339 ) ;
  assign w7341 = w2015 & w7340 ;
  assign w7342 = w6991 | w6996 ;
  assign w7343 = w7175 & ~w7342 ;
  assign w7344 = w6994 ^ w7343 ;
  assign w7345 = ( ~w2015 & w7333 ) | ( ~w2015 & w7339 ) | ( w7333 & w7339 ) ;
  assign w7346 = ~w7333 & w7345 ;
  assign w7347 = w7344 | w7346 ;
  assign w7348 = ( w1841 & w7341 ) | ( w1841 & ~w7347 ) | ( w7341 & ~w7347 ) ;
  assign w7349 = w1841 & w7348 ;
  assign w7350 = w6999 | w7004 ;
  assign w7351 = w7175 & ~w7350 ;
  assign w7352 = w7002 ^ w7351 ;
  assign w7353 = ( ~w1841 & w7341 ) | ( ~w1841 & w7347 ) | ( w7341 & w7347 ) ;
  assign w7354 = ~w7341 & w7353 ;
  assign w7355 = w7352 | w7354 ;
  assign w7356 = ( w1675 & w7349 ) | ( w1675 & ~w7355 ) | ( w7349 & ~w7355 ) ;
  assign w7357 = w1675 & w7356 ;
  assign w7358 = w7007 | w7012 ;
  assign w7359 = w7175 & ~w7358 ;
  assign w7360 = w7010 ^ w7359 ;
  assign w7361 = ( ~w1675 & w7349 ) | ( ~w1675 & w7355 ) | ( w7349 & w7355 ) ;
  assign w7362 = ~w7349 & w7361 ;
  assign w7363 = w7360 | w7362 ;
  assign w7364 = ( w1517 & w7357 ) | ( w1517 & ~w7363 ) | ( w7357 & ~w7363 ) ;
  assign w7365 = w1517 & w7364 ;
  assign w7366 = w7015 | w7020 ;
  assign w7367 = w7175 & ~w7366 ;
  assign w7368 = w7018 ^ w7367 ;
  assign w7369 = ( ~w1517 & w7357 ) | ( ~w1517 & w7363 ) | ( w7357 & w7363 ) ;
  assign w7370 = ~w7357 & w7369 ;
  assign w7371 = w7368 | w7370 ;
  assign w7372 = ( w1367 & w7365 ) | ( w1367 & ~w7371 ) | ( w7365 & ~w7371 ) ;
  assign w7373 = w1367 & w7372 ;
  assign w7374 = w7023 | w7028 ;
  assign w7375 = w7175 & ~w7374 ;
  assign w7376 = w7026 ^ w7375 ;
  assign w7377 = ( ~w1367 & w7365 ) | ( ~w1367 & w7371 ) | ( w7365 & w7371 ) ;
  assign w7378 = ~w7365 & w7377 ;
  assign w7379 = w7376 | w7378 ;
  assign w7380 = ( w1225 & w7373 ) | ( w1225 & ~w7379 ) | ( w7373 & ~w7379 ) ;
  assign w7381 = w1225 & w7380 ;
  assign w7382 = w7031 | w7036 ;
  assign w7383 = w7175 & ~w7382 ;
  assign w7384 = w7034 ^ w7383 ;
  assign w7385 = ( ~w1225 & w7373 ) | ( ~w1225 & w7379 ) | ( w7373 & w7379 ) ;
  assign w7386 = ~w7373 & w7385 ;
  assign w7387 = w7384 | w7386 ;
  assign w7388 = ( w1091 & w7381 ) | ( w1091 & ~w7387 ) | ( w7381 & ~w7387 ) ;
  assign w7389 = w1091 & w7388 ;
  assign w7390 = w7039 | w7044 ;
  assign w7391 = w7175 & ~w7390 ;
  assign w7392 = w7042 ^ w7391 ;
  assign w7393 = ( ~w1091 & w7381 ) | ( ~w1091 & w7387 ) | ( w7381 & w7387 ) ;
  assign w7394 = ~w7381 & w7393 ;
  assign w7395 = w7392 | w7394 ;
  assign w7396 = ( w965 & w7389 ) | ( w965 & ~w7395 ) | ( w7389 & ~w7395 ) ;
  assign w7397 = w965 & w7396 ;
  assign w7398 = w7047 | w7052 ;
  assign w7399 = w7175 & ~w7398 ;
  assign w7400 = w7050 ^ w7399 ;
  assign w7401 = ( ~w965 & w7389 ) | ( ~w965 & w7395 ) | ( w7389 & w7395 ) ;
  assign w7402 = ~w7389 & w7401 ;
  assign w7403 = w7400 | w7402 ;
  assign w7404 = ( w847 & w7397 ) | ( w847 & ~w7403 ) | ( w7397 & ~w7403 ) ;
  assign w7405 = w847 & w7404 ;
  assign w7406 = w7055 | w7060 ;
  assign w7407 = w7175 & ~w7406 ;
  assign w7408 = w7058 ^ w7407 ;
  assign w7409 = ( ~w847 & w7397 ) | ( ~w847 & w7403 ) | ( w7397 & w7403 ) ;
  assign w7410 = ~w7397 & w7409 ;
  assign w7411 = w7408 | w7410 ;
  assign w7412 = ( w737 & w7405 ) | ( w737 & ~w7411 ) | ( w7405 & ~w7411 ) ;
  assign w7413 = w737 & w7412 ;
  assign w7414 = w7063 | w7068 ;
  assign w7415 = w7175 & ~w7414 ;
  assign w7416 = w7066 ^ w7415 ;
  assign w7417 = ( ~w737 & w7405 ) | ( ~w737 & w7411 ) | ( w7405 & w7411 ) ;
  assign w7418 = ~w7405 & w7417 ;
  assign w7419 = w7416 | w7418 ;
  assign w7420 = ( w635 & w7413 ) | ( w635 & ~w7419 ) | ( w7413 & ~w7419 ) ;
  assign w7421 = w635 & w7420 ;
  assign w7422 = w7071 | w7076 ;
  assign w7423 = w7175 & ~w7422 ;
  assign w7424 = w7074 ^ w7423 ;
  assign w7425 = ( ~w635 & w7413 ) | ( ~w635 & w7419 ) | ( w7413 & w7419 ) ;
  assign w7426 = ~w7413 & w7425 ;
  assign w7427 = w7424 | w7426 ;
  assign w7428 = ( w541 & w7421 ) | ( w541 & ~w7427 ) | ( w7421 & ~w7427 ) ;
  assign w7429 = w541 & w7428 ;
  assign w7430 = w7079 | w7084 ;
  assign w7431 = w7175 & ~w7430 ;
  assign w7432 = w7082 ^ w7431 ;
  assign w7433 = ( ~w541 & w7421 ) | ( ~w541 & w7427 ) | ( w7421 & w7427 ) ;
  assign w7434 = ~w7421 & w7433 ;
  assign w7435 = w7432 | w7434 ;
  assign w7436 = ( w455 & w7429 ) | ( w455 & ~w7435 ) | ( w7429 & ~w7435 ) ;
  assign w7437 = w455 & w7436 ;
  assign w7438 = w7087 | w7092 ;
  assign w7439 = w7175 & ~w7438 ;
  assign w7440 = w7090 ^ w7439 ;
  assign w7441 = ( ~w455 & w7429 ) | ( ~w455 & w7435 ) | ( w7429 & w7435 ) ;
  assign w7442 = ~w7429 & w7441 ;
  assign w7443 = w7440 | w7442 ;
  assign w7444 = ( w377 & w7437 ) | ( w377 & ~w7443 ) | ( w7437 & ~w7443 ) ;
  assign w7445 = w377 & w7444 ;
  assign w7446 = w7095 | w7100 ;
  assign w7447 = w7175 & ~w7446 ;
  assign w7448 = w7098 ^ w7447 ;
  assign w7449 = ( ~w377 & w7437 ) | ( ~w377 & w7443 ) | ( w7437 & w7443 ) ;
  assign w7450 = ~w7437 & w7449 ;
  assign w7451 = w7448 | w7450 ;
  assign w7452 = ( w307 & w7445 ) | ( w307 & ~w7451 ) | ( w7445 & ~w7451 ) ;
  assign w7453 = w307 & w7452 ;
  assign w7454 = w7103 | w7108 ;
  assign w7455 = w7175 & ~w7454 ;
  assign w7456 = w7106 ^ w7455 ;
  assign w7457 = ( ~w307 & w7445 ) | ( ~w307 & w7451 ) | ( w7445 & w7451 ) ;
  assign w7458 = ~w7445 & w7457 ;
  assign w7459 = w7456 | w7458 ;
  assign w7460 = ( w246 & w7453 ) | ( w246 & ~w7459 ) | ( w7453 & ~w7459 ) ;
  assign w7461 = w246 & w7460 ;
  assign w7462 = w7111 | w7116 ;
  assign w7463 = w7175 & ~w7462 ;
  assign w7464 = w7114 ^ w7463 ;
  assign w7465 = ( ~w246 & w7453 ) | ( ~w246 & w7459 ) | ( w7453 & w7459 ) ;
  assign w7466 = ~w7453 & w7465 ;
  assign w7467 = w7464 | w7466 ;
  assign w7468 = ( w185 & w7461 ) | ( w185 & ~w7467 ) | ( w7461 & ~w7467 ) ;
  assign w7469 = w185 & w7468 ;
  assign w7470 = w7119 | w7124 ;
  assign w7471 = w7175 & ~w7470 ;
  assign w7472 = w7122 ^ w7471 ;
  assign w7473 = ( ~w185 & w7461 ) | ( ~w185 & w7467 ) | ( w7461 & w7467 ) ;
  assign w7474 = ~w7461 & w7473 ;
  assign w7475 = w7472 | w7474 ;
  assign w7476 = ( w145 & w7469 ) | ( w145 & ~w7475 ) | ( w7469 & ~w7475 ) ;
  assign w7477 = w145 & w7476 ;
  assign w7478 = w7127 | w7132 ;
  assign w7479 = w7175 & ~w7478 ;
  assign w7480 = w7130 ^ w7479 ;
  assign w7481 = ( ~w145 & w7469 ) | ( ~w145 & w7475 ) | ( w7469 & w7475 ) ;
  assign w7482 = ~w7469 & w7481 ;
  assign w7483 = w7480 | w7482 ;
  assign w7484 = ( w132 & w7477 ) | ( w132 & ~w7483 ) | ( w7477 & ~w7483 ) ;
  assign w7485 = w132 & w7484 ;
  assign w7486 = w7135 | w7140 ;
  assign w7487 = w7175 & ~w7486 ;
  assign w7488 = w7138 ^ w7487 ;
  assign w7489 = ( ~w132 & w7477 ) | ( ~w132 & w7483 ) | ( w7477 & w7483 ) ;
  assign w7490 = ~w7477 & w7489 ;
  assign w7491 = w7488 | w7490 ;
  assign w7492 = ~w7485 & w7491 ;
  assign w7493 = w7143 | w7148 ;
  assign w7494 = w7175 & ~w7493 ;
  assign w7495 = w7146 ^ w7494 ;
  assign w7496 = ( ~w7161 & w7492 ) | ( ~w7161 & w7495 ) | ( w7492 & w7495 ) ;
  assign w7497 = w7150 & ~w7496 ;
  assign w7498 = ~w7153 & w7175 ;
  assign w7499 = ( w7496 & ~w7497 ) | ( w7496 & w7498 ) | ( ~w7497 & w7498 ) ;
  assign w7500 = w7161 | w7499 ;
  assign w7501 = ~w129 & w7500 ;
  assign w7502 = ( w7485 & w7491 ) | ( w7485 & w7495 ) | ( w7491 & w7495 ) ;
  assign w7503 = ~w7485 & w7502 ;
  assign w7504 = ( w129 & w7150 ) | ( w129 & w7153 ) | ( w7150 & w7153 ) ;
  assign w7505 = ( w7153 & ~w7175 ) | ( w7153 & w7504 ) | ( ~w7175 & w7504 ) ;
  assign w7506 = w7150 & w7505 ;
  assign w7507 = w7504 ^ w7506 ;
  assign w7508 = ( w6809 & w6814 ) | ( w6809 & w6841 ) | ( w6814 & w6841 ) ;
  assign w7509 = w6841 & ~w7508 ;
  assign w7510 = w6812 ^ w7509 ;
  assign w7511 = ( ~w7165 & w7172 ) | ( ~w7165 & w7510 ) | ( w7172 & w7510 ) ;
  assign w7512 = ~w7172 & w7511 ;
  assign w7513 = ( ~w7159 & w7161 ) | ( ~w7159 & w7512 ) | ( w7161 & w7512 ) ;
  assign w7514 = ~w7161 & w7513 ;
  assign w7515 = w7503 | w7514 ;
  assign w7516 = ( w7501 & ~w7503 ) | ( w7501 & w7507 ) | ( ~w7503 & w7507 ) ;
  assign w7517 = w7515 | w7516 ;
  assign w7518 = ( ~\pi045 & \pi046 ) | ( ~\pi045 & w7175 ) | ( \pi046 & w7175 ) ;
  assign w7519 = ( ~\pi044 & \pi046 ) | ( ~\pi044 & w7518 ) | ( \pi046 & w7518 ) ;
  assign w7520 = ( ~\pi046 & w7175 ) | ( ~\pi046 & w7517 ) | ( w7175 & w7517 ) ;
  assign w7521 = w7519 & w7520 ;
  assign w7522 = ( w7161 & w7165 ) | ( w7161 & ~w7172 ) | ( w7165 & ~w7172 ) ;
  assign w7523 = \pi045 & ~w7522 ;
  assign w7524 = \pi044 | \pi046 ;
  assign w7525 = ( ~w7522 & w7523 ) | ( ~w7522 & w7524 ) | ( w7523 & w7524 ) ;
  assign w7526 = ~w7172 & w7525 ;
  assign w7527 = ~w7159 & w7526 ;
  assign w7528 = ( \pi046 & w7517 ) | ( \pi046 & ~w7526 ) | ( w7517 & ~w7526 ) ;
  assign w7529 = w7527 & ~w7528 ;
  assign w7530 = ~\pi046 & w7517 ;
  assign w7531 = \pi047 ^ w7530 ;
  assign w7532 = w7529 | w7531 ;
  assign w7533 = ( w6841 & w7521 ) | ( w6841 & ~w7532 ) | ( w7521 & ~w7532 ) ;
  assign w7534 = w6841 & w7533 ;
  assign w7535 = ( ~w6841 & w7521 ) | ( ~w6841 & w7532 ) | ( w7521 & w7532 ) ;
  assign w7536 = ~w7521 & w7535 ;
  assign w7537 = w7175 & ~w7514 ;
  assign w7538 = ~w7503 & w7537 ;
  assign w7539 = ~w7516 & w7538 ;
  assign w7540 = \pi047 & w7517 ;
  assign w7541 = ( \pi046 & w7517 ) | ( \pi046 & ~w7540 ) | ( w7517 & ~w7540 ) ;
  assign w7542 = ( ~\pi046 & w7539 ) | ( ~\pi046 & w7541 ) | ( w7539 & w7541 ) ;
  assign w7543 = \pi048 ^ w7542 ;
  assign w7544 = w7536 | w7543 ;
  assign w7545 = ( w6515 & w7534 ) | ( w6515 & ~w7544 ) | ( w7534 & ~w7544 ) ;
  assign w7546 = w6515 & w7545 ;
  assign w7547 = ( w7179 & ~w7187 ) | ( w7179 & w7517 ) | ( ~w7187 & w7517 ) ;
  assign w7548 = ~w7179 & w7547 ;
  assign w7549 = \pi049 ^ w7548 ;
  assign w7550 = w7188 ^ w7549 ;
  assign w7551 = ( ~w6515 & w7534 ) | ( ~w6515 & w7544 ) | ( w7534 & w7544 ) ;
  assign w7552 = ~w7534 & w7551 ;
  assign w7553 = w7550 | w7552 ;
  assign w7554 = ( w6197 & w7546 ) | ( w6197 & ~w7553 ) | ( w7546 & ~w7553 ) ;
  assign w7555 = w6197 & w7554 ;
  assign w7556 = w7192 | w7194 ;
  assign w7557 = w7517 & ~w7556 ;
  assign w7558 = w7201 ^ w7557 ;
  assign w7559 = ( ~w6197 & w7546 ) | ( ~w6197 & w7553 ) | ( w7546 & w7553 ) ;
  assign w7560 = ~w7546 & w7559 ;
  assign w7561 = w7558 | w7560 ;
  assign w7562 = ( w5887 & w7555 ) | ( w5887 & ~w7561 ) | ( w7555 & ~w7561 ) ;
  assign w7563 = w5887 & w7562 ;
  assign w7564 = w7204 | w7210 ;
  assign w7565 = w7517 & ~w7564 ;
  assign w7566 = w7208 ^ w7565 ;
  assign w7567 = ( ~w5887 & w7555 ) | ( ~w5887 & w7561 ) | ( w7555 & w7561 ) ;
  assign w7568 = ~w7555 & w7567 ;
  assign w7569 = w7566 | w7568 ;
  assign w7570 = ( w5585 & w7563 ) | ( w5585 & ~w7569 ) | ( w7563 & ~w7569 ) ;
  assign w7571 = w5585 & w7570 ;
  assign w7572 = w7213 | w7218 ;
  assign w7573 = w7517 & ~w7572 ;
  assign w7574 = w7216 ^ w7573 ;
  assign w7575 = ( ~w5585 & w7563 ) | ( ~w5585 & w7569 ) | ( w7563 & w7569 ) ;
  assign w7576 = ~w7563 & w7575 ;
  assign w7577 = w7574 | w7576 ;
  assign w7578 = ( w5291 & w7571 ) | ( w5291 & ~w7577 ) | ( w7571 & ~w7577 ) ;
  assign w7579 = w5291 & w7578 ;
  assign w7580 = w7221 | w7226 ;
  assign w7581 = w7517 & ~w7580 ;
  assign w7582 = w7224 ^ w7581 ;
  assign w7583 = ( ~w5291 & w7571 ) | ( ~w5291 & w7577 ) | ( w7571 & w7577 ) ;
  assign w7584 = ~w7571 & w7583 ;
  assign w7585 = w7582 | w7584 ;
  assign w7586 = ( w5005 & w7579 ) | ( w5005 & ~w7585 ) | ( w7579 & ~w7585 ) ;
  assign w7587 = w5005 & w7586 ;
  assign w7588 = w7229 | w7234 ;
  assign w7589 = w7517 & ~w7588 ;
  assign w7590 = w7232 ^ w7589 ;
  assign w7591 = ( ~w5005 & w7579 ) | ( ~w5005 & w7585 ) | ( w7579 & w7585 ) ;
  assign w7592 = ~w7579 & w7591 ;
  assign w7593 = w7590 | w7592 ;
  assign w7594 = ( w4727 & w7587 ) | ( w4727 & ~w7593 ) | ( w7587 & ~w7593 ) ;
  assign w7595 = w4727 & w7594 ;
  assign w7596 = w7237 | w7242 ;
  assign w7597 = w7517 & ~w7596 ;
  assign w7598 = w7240 ^ w7597 ;
  assign w7599 = ( ~w4727 & w7587 ) | ( ~w4727 & w7593 ) | ( w7587 & w7593 ) ;
  assign w7600 = ~w7587 & w7599 ;
  assign w7601 = w7598 | w7600 ;
  assign w7602 = ( w4457 & w7595 ) | ( w4457 & ~w7601 ) | ( w7595 & ~w7601 ) ;
  assign w7603 = w4457 & w7602 ;
  assign w7604 = w7245 | w7250 ;
  assign w7605 = w7517 & ~w7604 ;
  assign w7606 = w7248 ^ w7605 ;
  assign w7607 = ( ~w4457 & w7595 ) | ( ~w4457 & w7601 ) | ( w7595 & w7601 ) ;
  assign w7608 = ~w7595 & w7607 ;
  assign w7609 = w7606 | w7608 ;
  assign w7610 = ( w4195 & w7603 ) | ( w4195 & ~w7609 ) | ( w7603 & ~w7609 ) ;
  assign w7611 = w4195 & w7610 ;
  assign w7612 = w7253 | w7258 ;
  assign w7613 = w7517 & ~w7612 ;
  assign w7614 = w7256 ^ w7613 ;
  assign w7615 = ( ~w4195 & w7603 ) | ( ~w4195 & w7609 ) | ( w7603 & w7609 ) ;
  assign w7616 = ~w7603 & w7615 ;
  assign w7617 = w7614 | w7616 ;
  assign w7618 = ( w3941 & w7611 ) | ( w3941 & ~w7617 ) | ( w7611 & ~w7617 ) ;
  assign w7619 = w3941 & w7618 ;
  assign w7620 = w7261 | w7266 ;
  assign w7621 = w7517 & ~w7620 ;
  assign w7622 = w7264 ^ w7621 ;
  assign w7623 = ( ~w3941 & w7611 ) | ( ~w3941 & w7617 ) | ( w7611 & w7617 ) ;
  assign w7624 = ~w7611 & w7623 ;
  assign w7625 = w7622 | w7624 ;
  assign w7626 = ( w3695 & w7619 ) | ( w3695 & ~w7625 ) | ( w7619 & ~w7625 ) ;
  assign w7627 = w3695 & w7626 ;
  assign w7628 = w7269 | w7274 ;
  assign w7629 = w7517 & ~w7628 ;
  assign w7630 = w7272 ^ w7629 ;
  assign w7631 = ( ~w3695 & w7619 ) | ( ~w3695 & w7625 ) | ( w7619 & w7625 ) ;
  assign w7632 = ~w7619 & w7631 ;
  assign w7633 = w7630 | w7632 ;
  assign w7634 = ( w3457 & w7627 ) | ( w3457 & ~w7633 ) | ( w7627 & ~w7633 ) ;
  assign w7635 = w3457 & w7634 ;
  assign w7636 = w7277 | w7282 ;
  assign w7637 = w7517 & ~w7636 ;
  assign w7638 = w7280 ^ w7637 ;
  assign w7639 = ( ~w3457 & w7627 ) | ( ~w3457 & w7633 ) | ( w7627 & w7633 ) ;
  assign w7640 = ~w7627 & w7639 ;
  assign w7641 = w7638 | w7640 ;
  assign w7642 = ( w3227 & w7635 ) | ( w3227 & ~w7641 ) | ( w7635 & ~w7641 ) ;
  assign w7643 = w3227 & w7642 ;
  assign w7644 = w7285 | w7290 ;
  assign w7645 = w7517 & ~w7644 ;
  assign w7646 = w7288 ^ w7645 ;
  assign w7647 = ( ~w3227 & w7635 ) | ( ~w3227 & w7641 ) | ( w7635 & w7641 ) ;
  assign w7648 = ~w7635 & w7647 ;
  assign w7649 = w7646 | w7648 ;
  assign w7650 = ( w3005 & w7643 ) | ( w3005 & ~w7649 ) | ( w7643 & ~w7649 ) ;
  assign w7651 = w3005 & w7650 ;
  assign w7652 = w7293 | w7298 ;
  assign w7653 = w7517 & ~w7652 ;
  assign w7654 = w7296 ^ w7653 ;
  assign w7655 = ( ~w3005 & w7643 ) | ( ~w3005 & w7649 ) | ( w7643 & w7649 ) ;
  assign w7656 = ~w7643 & w7655 ;
  assign w7657 = w7654 | w7656 ;
  assign w7658 = ( w2791 & w7651 ) | ( w2791 & ~w7657 ) | ( w7651 & ~w7657 ) ;
  assign w7659 = w2791 & w7658 ;
  assign w7660 = w7301 | w7306 ;
  assign w7661 = w7517 & ~w7660 ;
  assign w7662 = w7304 ^ w7661 ;
  assign w7663 = ( ~w2791 & w7651 ) | ( ~w2791 & w7657 ) | ( w7651 & w7657 ) ;
  assign w7664 = ~w7651 & w7663 ;
  assign w7665 = w7662 | w7664 ;
  assign w7666 = ( w2585 & w7659 ) | ( w2585 & ~w7665 ) | ( w7659 & ~w7665 ) ;
  assign w7667 = w2585 & w7666 ;
  assign w7668 = w7309 | w7314 ;
  assign w7669 = w7517 & ~w7668 ;
  assign w7670 = w7312 ^ w7669 ;
  assign w7671 = ( ~w2585 & w7659 ) | ( ~w2585 & w7665 ) | ( w7659 & w7665 ) ;
  assign w7672 = ~w7659 & w7671 ;
  assign w7673 = w7670 | w7672 ;
  assign w7674 = ( w2387 & w7667 ) | ( w2387 & ~w7673 ) | ( w7667 & ~w7673 ) ;
  assign w7675 = w2387 & w7674 ;
  assign w7676 = ( ~w2387 & w7667 ) | ( ~w2387 & w7673 ) | ( w7667 & w7673 ) ;
  assign w7677 = ~w7667 & w7676 ;
  assign w7678 = w7317 | w7319 ;
  assign w7679 = w7517 & ~w7678 ;
  assign w7680 = w7322 ^ w7679 ;
  assign w7681 = w7677 | w7680 ;
  assign w7682 = ( w2197 & w7675 ) | ( w2197 & ~w7681 ) | ( w7675 & ~w7681 ) ;
  assign w7683 = w2197 & w7682 ;
  assign w7684 = w7325 | w7330 ;
  assign w7685 = w7517 & ~w7684 ;
  assign w7686 = w7328 ^ w7685 ;
  assign w7687 = ( ~w2197 & w7675 ) | ( ~w2197 & w7681 ) | ( w7675 & w7681 ) ;
  assign w7688 = ~w7675 & w7687 ;
  assign w7689 = w7686 | w7688 ;
  assign w7690 = ( w2015 & w7683 ) | ( w2015 & ~w7689 ) | ( w7683 & ~w7689 ) ;
  assign w7691 = w2015 & w7690 ;
  assign w7692 = w7333 | w7338 ;
  assign w7693 = w7517 & ~w7692 ;
  assign w7694 = w7336 ^ w7693 ;
  assign w7695 = ( ~w2015 & w7683 ) | ( ~w2015 & w7689 ) | ( w7683 & w7689 ) ;
  assign w7696 = ~w7683 & w7695 ;
  assign w7697 = w7694 | w7696 ;
  assign w7698 = ( w1841 & w7691 ) | ( w1841 & ~w7697 ) | ( w7691 & ~w7697 ) ;
  assign w7699 = w1841 & w7698 ;
  assign w7700 = w7341 | w7346 ;
  assign w7701 = w7517 & ~w7700 ;
  assign w7702 = w7344 ^ w7701 ;
  assign w7703 = ( ~w1841 & w7691 ) | ( ~w1841 & w7697 ) | ( w7691 & w7697 ) ;
  assign w7704 = ~w7691 & w7703 ;
  assign w7705 = w7702 | w7704 ;
  assign w7706 = ( w1675 & w7699 ) | ( w1675 & ~w7705 ) | ( w7699 & ~w7705 ) ;
  assign w7707 = w1675 & w7706 ;
  assign w7708 = w7349 | w7354 ;
  assign w7709 = w7517 & ~w7708 ;
  assign w7710 = w7352 ^ w7709 ;
  assign w7711 = ( ~w1675 & w7699 ) | ( ~w1675 & w7705 ) | ( w7699 & w7705 ) ;
  assign w7712 = ~w7699 & w7711 ;
  assign w7713 = w7710 | w7712 ;
  assign w7714 = ( w1517 & w7707 ) | ( w1517 & ~w7713 ) | ( w7707 & ~w7713 ) ;
  assign w7715 = w1517 & w7714 ;
  assign w7716 = w7357 | w7362 ;
  assign w7717 = w7517 & ~w7716 ;
  assign w7718 = w7360 ^ w7717 ;
  assign w7719 = ( ~w1517 & w7707 ) | ( ~w1517 & w7713 ) | ( w7707 & w7713 ) ;
  assign w7720 = ~w7707 & w7719 ;
  assign w7721 = w7718 | w7720 ;
  assign w7722 = ( w1367 & w7715 ) | ( w1367 & ~w7721 ) | ( w7715 & ~w7721 ) ;
  assign w7723 = w1367 & w7722 ;
  assign w7724 = w7365 | w7370 ;
  assign w7725 = w7517 & ~w7724 ;
  assign w7726 = w7368 ^ w7725 ;
  assign w7727 = ( ~w1367 & w7715 ) | ( ~w1367 & w7721 ) | ( w7715 & w7721 ) ;
  assign w7728 = ~w7715 & w7727 ;
  assign w7729 = w7726 | w7728 ;
  assign w7730 = ( w1225 & w7723 ) | ( w1225 & ~w7729 ) | ( w7723 & ~w7729 ) ;
  assign w7731 = w1225 & w7730 ;
  assign w7732 = w7373 | w7378 ;
  assign w7733 = w7517 & ~w7732 ;
  assign w7734 = w7376 ^ w7733 ;
  assign w7735 = ( ~w1225 & w7723 ) | ( ~w1225 & w7729 ) | ( w7723 & w7729 ) ;
  assign w7736 = ~w7723 & w7735 ;
  assign w7737 = w7734 | w7736 ;
  assign w7738 = ( w1091 & w7731 ) | ( w1091 & ~w7737 ) | ( w7731 & ~w7737 ) ;
  assign w7739 = w1091 & w7738 ;
  assign w7740 = w7381 | w7386 ;
  assign w7741 = w7517 & ~w7740 ;
  assign w7742 = w7384 ^ w7741 ;
  assign w7743 = ( ~w1091 & w7731 ) | ( ~w1091 & w7737 ) | ( w7731 & w7737 ) ;
  assign w7744 = ~w7731 & w7743 ;
  assign w7745 = w7742 | w7744 ;
  assign w7746 = ( w965 & w7739 ) | ( w965 & ~w7745 ) | ( w7739 & ~w7745 ) ;
  assign w7747 = w965 & w7746 ;
  assign w7748 = w7389 | w7394 ;
  assign w7749 = w7517 & ~w7748 ;
  assign w7750 = w7392 ^ w7749 ;
  assign w7751 = ( ~w965 & w7739 ) | ( ~w965 & w7745 ) | ( w7739 & w7745 ) ;
  assign w7752 = ~w7739 & w7751 ;
  assign w7753 = w7750 | w7752 ;
  assign w7754 = ( w847 & w7747 ) | ( w847 & ~w7753 ) | ( w7747 & ~w7753 ) ;
  assign w7755 = w847 & w7754 ;
  assign w7756 = w7397 | w7402 ;
  assign w7757 = w7517 & ~w7756 ;
  assign w7758 = w7400 ^ w7757 ;
  assign w7759 = ( ~w847 & w7747 ) | ( ~w847 & w7753 ) | ( w7747 & w7753 ) ;
  assign w7760 = ~w7747 & w7759 ;
  assign w7761 = w7758 | w7760 ;
  assign w7762 = ( w737 & w7755 ) | ( w737 & ~w7761 ) | ( w7755 & ~w7761 ) ;
  assign w7763 = w737 & w7762 ;
  assign w7764 = w7405 | w7410 ;
  assign w7765 = w7517 & ~w7764 ;
  assign w7766 = w7408 ^ w7765 ;
  assign w7767 = ( ~w737 & w7755 ) | ( ~w737 & w7761 ) | ( w7755 & w7761 ) ;
  assign w7768 = ~w7755 & w7767 ;
  assign w7769 = w7766 | w7768 ;
  assign w7770 = ( w635 & w7763 ) | ( w635 & ~w7769 ) | ( w7763 & ~w7769 ) ;
  assign w7771 = w635 & w7770 ;
  assign w7772 = w7413 | w7418 ;
  assign w7773 = w7517 & ~w7772 ;
  assign w7774 = w7416 ^ w7773 ;
  assign w7775 = ( ~w635 & w7763 ) | ( ~w635 & w7769 ) | ( w7763 & w7769 ) ;
  assign w7776 = ~w7763 & w7775 ;
  assign w7777 = w7774 | w7776 ;
  assign w7778 = ( w541 & w7771 ) | ( w541 & ~w7777 ) | ( w7771 & ~w7777 ) ;
  assign w7779 = w541 & w7778 ;
  assign w7780 = w7421 | w7426 ;
  assign w7781 = w7517 & ~w7780 ;
  assign w7782 = w7424 ^ w7781 ;
  assign w7783 = ( ~w541 & w7771 ) | ( ~w541 & w7777 ) | ( w7771 & w7777 ) ;
  assign w7784 = ~w7771 & w7783 ;
  assign w7785 = w7782 | w7784 ;
  assign w7786 = ( w455 & w7779 ) | ( w455 & ~w7785 ) | ( w7779 & ~w7785 ) ;
  assign w7787 = w455 & w7786 ;
  assign w7788 = w7429 | w7434 ;
  assign w7789 = w7517 & ~w7788 ;
  assign w7790 = w7432 ^ w7789 ;
  assign w7791 = ( ~w455 & w7779 ) | ( ~w455 & w7785 ) | ( w7779 & w7785 ) ;
  assign w7792 = ~w7779 & w7791 ;
  assign w7793 = w7790 | w7792 ;
  assign w7794 = ( w377 & w7787 ) | ( w377 & ~w7793 ) | ( w7787 & ~w7793 ) ;
  assign w7795 = w377 & w7794 ;
  assign w7796 = w7437 | w7442 ;
  assign w7797 = w7517 & ~w7796 ;
  assign w7798 = w7440 ^ w7797 ;
  assign w7799 = ( ~w377 & w7787 ) | ( ~w377 & w7793 ) | ( w7787 & w7793 ) ;
  assign w7800 = ~w7787 & w7799 ;
  assign w7801 = w7798 | w7800 ;
  assign w7802 = ( w307 & w7795 ) | ( w307 & ~w7801 ) | ( w7795 & ~w7801 ) ;
  assign w7803 = w307 & w7802 ;
  assign w7804 = w7445 | w7450 ;
  assign w7805 = w7517 & ~w7804 ;
  assign w7806 = w7448 ^ w7805 ;
  assign w7807 = ( ~w307 & w7795 ) | ( ~w307 & w7801 ) | ( w7795 & w7801 ) ;
  assign w7808 = ~w7795 & w7807 ;
  assign w7809 = w7806 | w7808 ;
  assign w7810 = ( w246 & w7803 ) | ( w246 & ~w7809 ) | ( w7803 & ~w7809 ) ;
  assign w7811 = w246 & w7810 ;
  assign w7812 = w7453 | w7458 ;
  assign w7813 = w7517 & ~w7812 ;
  assign w7814 = w7456 ^ w7813 ;
  assign w7815 = ( ~w246 & w7803 ) | ( ~w246 & w7809 ) | ( w7803 & w7809 ) ;
  assign w7816 = ~w7803 & w7815 ;
  assign w7817 = w7814 | w7816 ;
  assign w7818 = ( w185 & w7811 ) | ( w185 & ~w7817 ) | ( w7811 & ~w7817 ) ;
  assign w7819 = w185 & w7818 ;
  assign w7820 = w7461 | w7466 ;
  assign w7821 = w7517 & ~w7820 ;
  assign w7822 = w7464 ^ w7821 ;
  assign w7823 = ( ~w185 & w7811 ) | ( ~w185 & w7817 ) | ( w7811 & w7817 ) ;
  assign w7824 = ~w7811 & w7823 ;
  assign w7825 = w7822 | w7824 ;
  assign w7826 = ( w145 & w7819 ) | ( w145 & ~w7825 ) | ( w7819 & ~w7825 ) ;
  assign w7827 = w145 & w7826 ;
  assign w7828 = w7469 | w7474 ;
  assign w7829 = w7517 & ~w7828 ;
  assign w7830 = w7472 ^ w7829 ;
  assign w7831 = ( ~w145 & w7819 ) | ( ~w145 & w7825 ) | ( w7819 & w7825 ) ;
  assign w7832 = ~w7819 & w7831 ;
  assign w7833 = w7830 | w7832 ;
  assign w7834 = ( w132 & w7827 ) | ( w132 & ~w7833 ) | ( w7827 & ~w7833 ) ;
  assign w7835 = w132 & w7834 ;
  assign w7836 = w7477 | w7482 ;
  assign w7837 = w7517 & ~w7836 ;
  assign w7838 = w7480 ^ w7837 ;
  assign w7839 = ( ~w132 & w7827 ) | ( ~w132 & w7833 ) | ( w7827 & w7833 ) ;
  assign w7840 = ~w7827 & w7839 ;
  assign w7841 = w7838 | w7840 ;
  assign w7842 = ~w7835 & w7841 ;
  assign w7843 = w7485 | w7490 ;
  assign w7844 = w7517 & ~w7843 ;
  assign w7845 = w7488 ^ w7844 ;
  assign w7846 = ( ~w7503 & w7842 ) | ( ~w7503 & w7845 ) | ( w7842 & w7845 ) ;
  assign w7847 = w7492 & ~w7846 ;
  assign w7848 = ~w7495 & w7517 ;
  assign w7849 = ( w7846 & ~w7847 ) | ( w7846 & w7848 ) | ( ~w7847 & w7848 ) ;
  assign w7850 = w7503 | w7849 ;
  assign w7851 = ~w129 & w7850 ;
  assign w7852 = ( w7835 & w7841 ) | ( w7835 & w7845 ) | ( w7841 & w7845 ) ;
  assign w7853 = ~w7835 & w7852 ;
  assign w7854 = ( w129 & w7492 ) | ( w129 & w7495 ) | ( w7492 & w7495 ) ;
  assign w7855 = ( w7495 & ~w7517 ) | ( w7495 & w7854 ) | ( ~w7517 & w7854 ) ;
  assign w7856 = w7492 & w7855 ;
  assign w7857 = w7854 ^ w7856 ;
  assign w7858 = ( w7143 & w7148 ) | ( w7143 & w7175 ) | ( w7148 & w7175 ) ;
  assign w7859 = w7175 & ~w7858 ;
  assign w7860 = w7146 ^ w7859 ;
  assign w7861 = ( ~w7507 & w7514 ) | ( ~w7507 & w7860 ) | ( w7514 & w7860 ) ;
  assign w7862 = ~w7514 & w7861 ;
  assign w7863 = ( ~w7501 & w7503 ) | ( ~w7501 & w7862 ) | ( w7503 & w7862 ) ;
  assign w7864 = ~w7503 & w7863 ;
  assign w7865 = w7853 | w7864 ;
  assign w7866 = ( w7851 & ~w7853 ) | ( w7851 & w7857 ) | ( ~w7853 & w7857 ) ;
  assign w7867 = w7865 | w7866 ;
  assign w7868 = ( ~\pi043 & \pi044 ) | ( ~\pi043 & w7517 ) | ( \pi044 & w7517 ) ;
  assign w7869 = ( ~\pi042 & \pi044 ) | ( ~\pi042 & w7868 ) | ( \pi044 & w7868 ) ;
  assign w7870 = ( ~\pi044 & w7517 ) | ( ~\pi044 & w7867 ) | ( w7517 & w7867 ) ;
  assign w7871 = w7869 & w7870 ;
  assign w7872 = ( w7503 & w7507 ) | ( w7503 & ~w7514 ) | ( w7507 & ~w7514 ) ;
  assign w7873 = \pi043 & ~w7872 ;
  assign w7874 = \pi042 | \pi044 ;
  assign w7875 = ( ~w7872 & w7873 ) | ( ~w7872 & w7874 ) | ( w7873 & w7874 ) ;
  assign w7876 = ~w7514 & w7875 ;
  assign w7877 = ~w7501 & w7876 ;
  assign w7878 = ( \pi044 & w7867 ) | ( \pi044 & ~w7876 ) | ( w7867 & ~w7876 ) ;
  assign w7879 = w7877 & ~w7878 ;
  assign w7880 = ~\pi044 & w7867 ;
  assign w7881 = \pi045 ^ w7880 ;
  assign w7882 = w7879 | w7881 ;
  assign w7883 = ( w7175 & w7871 ) | ( w7175 & ~w7882 ) | ( w7871 & ~w7882 ) ;
  assign w7884 = w7175 & w7883 ;
  assign w7885 = ( ~w7175 & w7871 ) | ( ~w7175 & w7882 ) | ( w7871 & w7882 ) ;
  assign w7886 = ~w7871 & w7885 ;
  assign w7887 = w7517 & ~w7864 ;
  assign w7888 = ~w7853 & w7887 ;
  assign w7889 = ~w7866 & w7888 ;
  assign w7890 = \pi045 & w7867 ;
  assign w7891 = ( \pi044 & w7867 ) | ( \pi044 & ~w7890 ) | ( w7867 & ~w7890 ) ;
  assign w7892 = ( ~\pi044 & w7889 ) | ( ~\pi044 & w7891 ) | ( w7889 & w7891 ) ;
  assign w7893 = \pi046 ^ w7892 ;
  assign w7894 = w7886 | w7893 ;
  assign w7895 = ( w6841 & w7884 ) | ( w6841 & ~w7894 ) | ( w7884 & ~w7894 ) ;
  assign w7896 = w6841 & w7895 ;
  assign w7897 = ( w7521 & ~w7529 ) | ( w7521 & w7867 ) | ( ~w7529 & w7867 ) ;
  assign w7898 = ~w7521 & w7897 ;
  assign w7899 = \pi047 ^ w7898 ;
  assign w7900 = w7530 ^ w7899 ;
  assign w7901 = ( ~w6841 & w7884 ) | ( ~w6841 & w7894 ) | ( w7884 & w7894 ) ;
  assign w7902 = ~w7884 & w7901 ;
  assign w7903 = w7900 | w7902 ;
  assign w7904 = ( w6515 & w7896 ) | ( w6515 & ~w7903 ) | ( w7896 & ~w7903 ) ;
  assign w7905 = w6515 & w7904 ;
  assign w7906 = w7534 | w7536 ;
  assign w7907 = w7867 & ~w7906 ;
  assign w7908 = w7543 ^ w7907 ;
  assign w7909 = ( ~w6515 & w7896 ) | ( ~w6515 & w7903 ) | ( w7896 & w7903 ) ;
  assign w7910 = ~w7896 & w7909 ;
  assign w7911 = w7908 | w7910 ;
  assign w7912 = ( w6197 & w7905 ) | ( w6197 & ~w7911 ) | ( w7905 & ~w7911 ) ;
  assign w7913 = w6197 & w7912 ;
  assign w7914 = w7546 | w7552 ;
  assign w7915 = w7867 & ~w7914 ;
  assign w7916 = w7550 ^ w7915 ;
  assign w7917 = ( ~w6197 & w7905 ) | ( ~w6197 & w7911 ) | ( w7905 & w7911 ) ;
  assign w7918 = ~w7905 & w7917 ;
  assign w7919 = w7916 | w7918 ;
  assign w7920 = ( w5887 & w7913 ) | ( w5887 & ~w7919 ) | ( w7913 & ~w7919 ) ;
  assign w7921 = w5887 & w7920 ;
  assign w7922 = w7555 | w7560 ;
  assign w7923 = w7867 & ~w7922 ;
  assign w7924 = w7558 ^ w7923 ;
  assign w7925 = ( ~w5887 & w7913 ) | ( ~w5887 & w7919 ) | ( w7913 & w7919 ) ;
  assign w7926 = ~w7913 & w7925 ;
  assign w7927 = w7924 | w7926 ;
  assign w7928 = ( w5585 & w7921 ) | ( w5585 & ~w7927 ) | ( w7921 & ~w7927 ) ;
  assign w7929 = w5585 & w7928 ;
  assign w7930 = w7563 | w7568 ;
  assign w7931 = w7867 & ~w7930 ;
  assign w7932 = w7566 ^ w7931 ;
  assign w7933 = ( ~w5585 & w7921 ) | ( ~w5585 & w7927 ) | ( w7921 & w7927 ) ;
  assign w7934 = ~w7921 & w7933 ;
  assign w7935 = w7932 | w7934 ;
  assign w7936 = ( w5291 & w7929 ) | ( w5291 & ~w7935 ) | ( w7929 & ~w7935 ) ;
  assign w7937 = w5291 & w7936 ;
  assign w7938 = w7571 | w7576 ;
  assign w7939 = w7867 & ~w7938 ;
  assign w7940 = w7574 ^ w7939 ;
  assign w7941 = ( ~w5291 & w7929 ) | ( ~w5291 & w7935 ) | ( w7929 & w7935 ) ;
  assign w7942 = ~w7929 & w7941 ;
  assign w7943 = w7940 | w7942 ;
  assign w7944 = ( w5005 & w7937 ) | ( w5005 & ~w7943 ) | ( w7937 & ~w7943 ) ;
  assign w7945 = w5005 & w7944 ;
  assign w7946 = w7579 | w7584 ;
  assign w7947 = w7867 & ~w7946 ;
  assign w7948 = w7582 ^ w7947 ;
  assign w7949 = ( ~w5005 & w7937 ) | ( ~w5005 & w7943 ) | ( w7937 & w7943 ) ;
  assign w7950 = ~w7937 & w7949 ;
  assign w7951 = w7948 | w7950 ;
  assign w7952 = ( w4727 & w7945 ) | ( w4727 & ~w7951 ) | ( w7945 & ~w7951 ) ;
  assign w7953 = w4727 & w7952 ;
  assign w7954 = w7587 | w7592 ;
  assign w7955 = w7867 & ~w7954 ;
  assign w7956 = w7590 ^ w7955 ;
  assign w7957 = ( ~w4727 & w7945 ) | ( ~w4727 & w7951 ) | ( w7945 & w7951 ) ;
  assign w7958 = ~w7945 & w7957 ;
  assign w7959 = w7956 | w7958 ;
  assign w7960 = ( w4457 & w7953 ) | ( w4457 & ~w7959 ) | ( w7953 & ~w7959 ) ;
  assign w7961 = w4457 & w7960 ;
  assign w7962 = w7595 | w7600 ;
  assign w7963 = w7867 & ~w7962 ;
  assign w7964 = w7598 ^ w7963 ;
  assign w7965 = ( ~w4457 & w7953 ) | ( ~w4457 & w7959 ) | ( w7953 & w7959 ) ;
  assign w7966 = ~w7953 & w7965 ;
  assign w7967 = w7964 | w7966 ;
  assign w7968 = ( w4195 & w7961 ) | ( w4195 & ~w7967 ) | ( w7961 & ~w7967 ) ;
  assign w7969 = w4195 & w7968 ;
  assign w7970 = w7603 | w7608 ;
  assign w7971 = w7867 & ~w7970 ;
  assign w7972 = w7606 ^ w7971 ;
  assign w7973 = ( ~w4195 & w7961 ) | ( ~w4195 & w7967 ) | ( w7961 & w7967 ) ;
  assign w7974 = ~w7961 & w7973 ;
  assign w7975 = w7972 | w7974 ;
  assign w7976 = ( w3941 & w7969 ) | ( w3941 & ~w7975 ) | ( w7969 & ~w7975 ) ;
  assign w7977 = w3941 & w7976 ;
  assign w7978 = w7611 | w7616 ;
  assign w7979 = w7867 & ~w7978 ;
  assign w7980 = w7614 ^ w7979 ;
  assign w7981 = ( ~w3941 & w7969 ) | ( ~w3941 & w7975 ) | ( w7969 & w7975 ) ;
  assign w7982 = ~w7969 & w7981 ;
  assign w7983 = w7980 | w7982 ;
  assign w7984 = ( w3695 & w7977 ) | ( w3695 & ~w7983 ) | ( w7977 & ~w7983 ) ;
  assign w7985 = w3695 & w7984 ;
  assign w7986 = w7619 | w7624 ;
  assign w7987 = w7867 & ~w7986 ;
  assign w7988 = w7622 ^ w7987 ;
  assign w7989 = ( ~w3695 & w7977 ) | ( ~w3695 & w7983 ) | ( w7977 & w7983 ) ;
  assign w7990 = ~w7977 & w7989 ;
  assign w7991 = w7988 | w7990 ;
  assign w7992 = ( w3457 & w7985 ) | ( w3457 & ~w7991 ) | ( w7985 & ~w7991 ) ;
  assign w7993 = w3457 & w7992 ;
  assign w7994 = w7627 | w7632 ;
  assign w7995 = w7867 & ~w7994 ;
  assign w7996 = w7630 ^ w7995 ;
  assign w7997 = ( ~w3457 & w7985 ) | ( ~w3457 & w7991 ) | ( w7985 & w7991 ) ;
  assign w7998 = ~w7985 & w7997 ;
  assign w7999 = w7996 | w7998 ;
  assign w8000 = ( w3227 & w7993 ) | ( w3227 & ~w7999 ) | ( w7993 & ~w7999 ) ;
  assign w8001 = w3227 & w8000 ;
  assign w8002 = w7635 | w7640 ;
  assign w8003 = w7867 & ~w8002 ;
  assign w8004 = w7638 ^ w8003 ;
  assign w8005 = ( ~w3227 & w7993 ) | ( ~w3227 & w7999 ) | ( w7993 & w7999 ) ;
  assign w8006 = ~w7993 & w8005 ;
  assign w8007 = w8004 | w8006 ;
  assign w8008 = ( w3005 & w8001 ) | ( w3005 & ~w8007 ) | ( w8001 & ~w8007 ) ;
  assign w8009 = w3005 & w8008 ;
  assign w8010 = w7643 | w7648 ;
  assign w8011 = w7867 & ~w8010 ;
  assign w8012 = w7646 ^ w8011 ;
  assign w8013 = ( ~w3005 & w8001 ) | ( ~w3005 & w8007 ) | ( w8001 & w8007 ) ;
  assign w8014 = ~w8001 & w8013 ;
  assign w8015 = w8012 | w8014 ;
  assign w8016 = ( w2791 & w8009 ) | ( w2791 & ~w8015 ) | ( w8009 & ~w8015 ) ;
  assign w8017 = w2791 & w8016 ;
  assign w8018 = w7651 | w7656 ;
  assign w8019 = w7867 & ~w8018 ;
  assign w8020 = w7654 ^ w8019 ;
  assign w8021 = ( ~w2791 & w8009 ) | ( ~w2791 & w8015 ) | ( w8009 & w8015 ) ;
  assign w8022 = ~w8009 & w8021 ;
  assign w8023 = w8020 | w8022 ;
  assign w8024 = ( w2585 & w8017 ) | ( w2585 & ~w8023 ) | ( w8017 & ~w8023 ) ;
  assign w8025 = w2585 & w8024 ;
  assign w8026 = w7659 | w7664 ;
  assign w8027 = w7867 & ~w8026 ;
  assign w8028 = w7662 ^ w8027 ;
  assign w8029 = ( ~w2585 & w8017 ) | ( ~w2585 & w8023 ) | ( w8017 & w8023 ) ;
  assign w8030 = ~w8017 & w8029 ;
  assign w8031 = w8028 | w8030 ;
  assign w8032 = ( w2387 & w8025 ) | ( w2387 & ~w8031 ) | ( w8025 & ~w8031 ) ;
  assign w8033 = w2387 & w8032 ;
  assign w8034 = w7667 | w7672 ;
  assign w8035 = w7867 & ~w8034 ;
  assign w8036 = w7670 ^ w8035 ;
  assign w8037 = ( ~w2387 & w8025 ) | ( ~w2387 & w8031 ) | ( w8025 & w8031 ) ;
  assign w8038 = ~w8025 & w8037 ;
  assign w8039 = w8036 | w8038 ;
  assign w8040 = ( w2197 & w8033 ) | ( w2197 & ~w8039 ) | ( w8033 & ~w8039 ) ;
  assign w8041 = w2197 & w8040 ;
  assign w8042 = ( ~w2197 & w8033 ) | ( ~w2197 & w8039 ) | ( w8033 & w8039 ) ;
  assign w8043 = ~w8033 & w8042 ;
  assign w8044 = w7675 | w7677 ;
  assign w8045 = w7867 & ~w8044 ;
  assign w8046 = w7680 ^ w8045 ;
  assign w8047 = w8043 | w8046 ;
  assign w8048 = ( w2015 & w8041 ) | ( w2015 & ~w8047 ) | ( w8041 & ~w8047 ) ;
  assign w8049 = w2015 & w8048 ;
  assign w8050 = w7683 | w7688 ;
  assign w8051 = w7867 & ~w8050 ;
  assign w8052 = w7686 ^ w8051 ;
  assign w8053 = ( ~w2015 & w8041 ) | ( ~w2015 & w8047 ) | ( w8041 & w8047 ) ;
  assign w8054 = ~w8041 & w8053 ;
  assign w8055 = w8052 | w8054 ;
  assign w8056 = ( w1841 & w8049 ) | ( w1841 & ~w8055 ) | ( w8049 & ~w8055 ) ;
  assign w8057 = w1841 & w8056 ;
  assign w8058 = w7691 | w7696 ;
  assign w8059 = w7867 & ~w8058 ;
  assign w8060 = w7694 ^ w8059 ;
  assign w8061 = ( ~w1841 & w8049 ) | ( ~w1841 & w8055 ) | ( w8049 & w8055 ) ;
  assign w8062 = ~w8049 & w8061 ;
  assign w8063 = w8060 | w8062 ;
  assign w8064 = ( w1675 & w8057 ) | ( w1675 & ~w8063 ) | ( w8057 & ~w8063 ) ;
  assign w8065 = w1675 & w8064 ;
  assign w8066 = w7699 | w7704 ;
  assign w8067 = w7867 & ~w8066 ;
  assign w8068 = w7702 ^ w8067 ;
  assign w8069 = ( ~w1675 & w8057 ) | ( ~w1675 & w8063 ) | ( w8057 & w8063 ) ;
  assign w8070 = ~w8057 & w8069 ;
  assign w8071 = w8068 | w8070 ;
  assign w8072 = ( w1517 & w8065 ) | ( w1517 & ~w8071 ) | ( w8065 & ~w8071 ) ;
  assign w8073 = w1517 & w8072 ;
  assign w8074 = w7707 | w7712 ;
  assign w8075 = w7867 & ~w8074 ;
  assign w8076 = w7710 ^ w8075 ;
  assign w8077 = ( ~w1517 & w8065 ) | ( ~w1517 & w8071 ) | ( w8065 & w8071 ) ;
  assign w8078 = ~w8065 & w8077 ;
  assign w8079 = w8076 | w8078 ;
  assign w8080 = ( w1367 & w8073 ) | ( w1367 & ~w8079 ) | ( w8073 & ~w8079 ) ;
  assign w8081 = w1367 & w8080 ;
  assign w8082 = w7715 | w7720 ;
  assign w8083 = w7867 & ~w8082 ;
  assign w8084 = w7718 ^ w8083 ;
  assign w8085 = ( ~w1367 & w8073 ) | ( ~w1367 & w8079 ) | ( w8073 & w8079 ) ;
  assign w8086 = ~w8073 & w8085 ;
  assign w8087 = w8084 | w8086 ;
  assign w8088 = ( w1225 & w8081 ) | ( w1225 & ~w8087 ) | ( w8081 & ~w8087 ) ;
  assign w8089 = w1225 & w8088 ;
  assign w8090 = w7723 | w7728 ;
  assign w8091 = w7867 & ~w8090 ;
  assign w8092 = w7726 ^ w8091 ;
  assign w8093 = ( ~w1225 & w8081 ) | ( ~w1225 & w8087 ) | ( w8081 & w8087 ) ;
  assign w8094 = ~w8081 & w8093 ;
  assign w8095 = w8092 | w8094 ;
  assign w8096 = ( w1091 & w8089 ) | ( w1091 & ~w8095 ) | ( w8089 & ~w8095 ) ;
  assign w8097 = w1091 & w8096 ;
  assign w8098 = w7731 | w7736 ;
  assign w8099 = w7867 & ~w8098 ;
  assign w8100 = w7734 ^ w8099 ;
  assign w8101 = ( ~w1091 & w8089 ) | ( ~w1091 & w8095 ) | ( w8089 & w8095 ) ;
  assign w8102 = ~w8089 & w8101 ;
  assign w8103 = w8100 | w8102 ;
  assign w8104 = ( w965 & w8097 ) | ( w965 & ~w8103 ) | ( w8097 & ~w8103 ) ;
  assign w8105 = w965 & w8104 ;
  assign w8106 = w7739 | w7744 ;
  assign w8107 = w7867 & ~w8106 ;
  assign w8108 = w7742 ^ w8107 ;
  assign w8109 = ( ~w965 & w8097 ) | ( ~w965 & w8103 ) | ( w8097 & w8103 ) ;
  assign w8110 = ~w8097 & w8109 ;
  assign w8111 = w8108 | w8110 ;
  assign w8112 = ( w847 & w8105 ) | ( w847 & ~w8111 ) | ( w8105 & ~w8111 ) ;
  assign w8113 = w847 & w8112 ;
  assign w8114 = w7747 | w7752 ;
  assign w8115 = w7867 & ~w8114 ;
  assign w8116 = w7750 ^ w8115 ;
  assign w8117 = ( ~w847 & w8105 ) | ( ~w847 & w8111 ) | ( w8105 & w8111 ) ;
  assign w8118 = ~w8105 & w8117 ;
  assign w8119 = w8116 | w8118 ;
  assign w8120 = ( w737 & w8113 ) | ( w737 & ~w8119 ) | ( w8113 & ~w8119 ) ;
  assign w8121 = w737 & w8120 ;
  assign w8122 = w7755 | w7760 ;
  assign w8123 = w7867 & ~w8122 ;
  assign w8124 = w7758 ^ w8123 ;
  assign w8125 = ( ~w737 & w8113 ) | ( ~w737 & w8119 ) | ( w8113 & w8119 ) ;
  assign w8126 = ~w8113 & w8125 ;
  assign w8127 = w8124 | w8126 ;
  assign w8128 = ( w635 & w8121 ) | ( w635 & ~w8127 ) | ( w8121 & ~w8127 ) ;
  assign w8129 = w635 & w8128 ;
  assign w8130 = w7763 | w7768 ;
  assign w8131 = w7867 & ~w8130 ;
  assign w8132 = w7766 ^ w8131 ;
  assign w8133 = ( ~w635 & w8121 ) | ( ~w635 & w8127 ) | ( w8121 & w8127 ) ;
  assign w8134 = ~w8121 & w8133 ;
  assign w8135 = w8132 | w8134 ;
  assign w8136 = ( w541 & w8129 ) | ( w541 & ~w8135 ) | ( w8129 & ~w8135 ) ;
  assign w8137 = w541 & w8136 ;
  assign w8138 = w7771 | w7776 ;
  assign w8139 = w7867 & ~w8138 ;
  assign w8140 = w7774 ^ w8139 ;
  assign w8141 = ( ~w541 & w8129 ) | ( ~w541 & w8135 ) | ( w8129 & w8135 ) ;
  assign w8142 = ~w8129 & w8141 ;
  assign w8143 = w8140 | w8142 ;
  assign w8144 = ( w455 & w8137 ) | ( w455 & ~w8143 ) | ( w8137 & ~w8143 ) ;
  assign w8145 = w455 & w8144 ;
  assign w8146 = w7779 | w7784 ;
  assign w8147 = w7867 & ~w8146 ;
  assign w8148 = w7782 ^ w8147 ;
  assign w8149 = ( ~w455 & w8137 ) | ( ~w455 & w8143 ) | ( w8137 & w8143 ) ;
  assign w8150 = ~w8137 & w8149 ;
  assign w8151 = w8148 | w8150 ;
  assign w8152 = ( w377 & w8145 ) | ( w377 & ~w8151 ) | ( w8145 & ~w8151 ) ;
  assign w8153 = w377 & w8152 ;
  assign w8154 = w7787 | w7792 ;
  assign w8155 = w7867 & ~w8154 ;
  assign w8156 = w7790 ^ w8155 ;
  assign w8157 = ( ~w377 & w8145 ) | ( ~w377 & w8151 ) | ( w8145 & w8151 ) ;
  assign w8158 = ~w8145 & w8157 ;
  assign w8159 = w8156 | w8158 ;
  assign w8160 = ( w307 & w8153 ) | ( w307 & ~w8159 ) | ( w8153 & ~w8159 ) ;
  assign w8161 = w307 & w8160 ;
  assign w8162 = w7795 | w7800 ;
  assign w8163 = w7867 & ~w8162 ;
  assign w8164 = w7798 ^ w8163 ;
  assign w8165 = ( ~w307 & w8153 ) | ( ~w307 & w8159 ) | ( w8153 & w8159 ) ;
  assign w8166 = ~w8153 & w8165 ;
  assign w8167 = w8164 | w8166 ;
  assign w8168 = ( w246 & w8161 ) | ( w246 & ~w8167 ) | ( w8161 & ~w8167 ) ;
  assign w8169 = w246 & w8168 ;
  assign w8170 = w7803 | w7808 ;
  assign w8171 = w7867 & ~w8170 ;
  assign w8172 = w7806 ^ w8171 ;
  assign w8173 = ( ~w246 & w8161 ) | ( ~w246 & w8167 ) | ( w8161 & w8167 ) ;
  assign w8174 = ~w8161 & w8173 ;
  assign w8175 = w8172 | w8174 ;
  assign w8176 = ( w185 & w8169 ) | ( w185 & ~w8175 ) | ( w8169 & ~w8175 ) ;
  assign w8177 = w185 & w8176 ;
  assign w8178 = w7811 | w7816 ;
  assign w8179 = w7867 & ~w8178 ;
  assign w8180 = w7814 ^ w8179 ;
  assign w8181 = ( ~w185 & w8169 ) | ( ~w185 & w8175 ) | ( w8169 & w8175 ) ;
  assign w8182 = ~w8169 & w8181 ;
  assign w8183 = w8180 | w8182 ;
  assign w8184 = ( w145 & w8177 ) | ( w145 & ~w8183 ) | ( w8177 & ~w8183 ) ;
  assign w8185 = w145 & w8184 ;
  assign w8186 = w7819 | w7824 ;
  assign w8187 = w7867 & ~w8186 ;
  assign w8188 = w7822 ^ w8187 ;
  assign w8189 = ( ~w145 & w8177 ) | ( ~w145 & w8183 ) | ( w8177 & w8183 ) ;
  assign w8190 = ~w8177 & w8189 ;
  assign w8191 = w8188 | w8190 ;
  assign w8192 = ( w132 & w8185 ) | ( w132 & ~w8191 ) | ( w8185 & ~w8191 ) ;
  assign w8193 = w132 & w8192 ;
  assign w8194 = w7827 | w7832 ;
  assign w8195 = w7867 & ~w8194 ;
  assign w8196 = w7830 ^ w8195 ;
  assign w8197 = ( ~w132 & w8185 ) | ( ~w132 & w8191 ) | ( w8185 & w8191 ) ;
  assign w8198 = ~w8185 & w8197 ;
  assign w8199 = w8196 | w8198 ;
  assign w8200 = ~w8193 & w8199 ;
  assign w8201 = w7835 | w7840 ;
  assign w8202 = w7867 & ~w8201 ;
  assign w8203 = w7838 ^ w8202 ;
  assign w8204 = ( ~w7853 & w8200 ) | ( ~w7853 & w8203 ) | ( w8200 & w8203 ) ;
  assign w8205 = w7842 & ~w8204 ;
  assign w8206 = ~w7845 & w7867 ;
  assign w8207 = ( w8204 & ~w8205 ) | ( w8204 & w8206 ) | ( ~w8205 & w8206 ) ;
  assign w8208 = w7853 | w8207 ;
  assign w8209 = ~w129 & w8208 ;
  assign w8210 = ( w8193 & w8199 ) | ( w8193 & w8203 ) | ( w8199 & w8203 ) ;
  assign w8211 = ~w8193 & w8210 ;
  assign w8212 = ( w129 & w7842 ) | ( w129 & w7845 ) | ( w7842 & w7845 ) ;
  assign w8213 = ( w7845 & ~w7867 ) | ( w7845 & w8212 ) | ( ~w7867 & w8212 ) ;
  assign w8214 = w7842 & w8213 ;
  assign w8215 = w8212 ^ w8214 ;
  assign w8216 = ( w7485 & w7490 ) | ( w7485 & w7517 ) | ( w7490 & w7517 ) ;
  assign w8217 = w7517 & ~w8216 ;
  assign w8218 = w7488 ^ w8217 ;
  assign w8219 = ( ~w7857 & w7864 ) | ( ~w7857 & w8218 ) | ( w7864 & w8218 ) ;
  assign w8220 = ~w7864 & w8219 ;
  assign w8221 = ( ~w7851 & w7853 ) | ( ~w7851 & w8220 ) | ( w7853 & w8220 ) ;
  assign w8222 = ~w7853 & w8221 ;
  assign w8223 = w8211 | w8222 ;
  assign w8224 = ( w8209 & ~w8211 ) | ( w8209 & w8215 ) | ( ~w8211 & w8215 ) ;
  assign w8225 = w8223 | w8224 ;
  assign w8226 = ( ~\pi041 & \pi042 ) | ( ~\pi041 & w7867 ) | ( \pi042 & w7867 ) ;
  assign w8227 = ( ~\pi040 & \pi042 ) | ( ~\pi040 & w8226 ) | ( \pi042 & w8226 ) ;
  assign w8228 = ( ~\pi042 & w7867 ) | ( ~\pi042 & w8225 ) | ( w7867 & w8225 ) ;
  assign w8229 = w8227 & w8228 ;
  assign w8230 = ( w7853 & w7857 ) | ( w7853 & ~w7864 ) | ( w7857 & ~w7864 ) ;
  assign w8231 = \pi041 & ~w8230 ;
  assign w8232 = \pi040 | \pi042 ;
  assign w8233 = ( ~w8230 & w8231 ) | ( ~w8230 & w8232 ) | ( w8231 & w8232 ) ;
  assign w8234 = ~w7864 & w8233 ;
  assign w8235 = ~w7851 & w8234 ;
  assign w8236 = ( \pi042 & w8225 ) | ( \pi042 & ~w8234 ) | ( w8225 & ~w8234 ) ;
  assign w8237 = w8235 & ~w8236 ;
  assign w8238 = ~\pi042 & w8225 ;
  assign w8239 = \pi043 ^ w8238 ;
  assign w8240 = w8237 | w8239 ;
  assign w8241 = ( w7517 & w8229 ) | ( w7517 & ~w8240 ) | ( w8229 & ~w8240 ) ;
  assign w8242 = w7517 & w8241 ;
  assign w8243 = ( ~w7517 & w8229 ) | ( ~w7517 & w8240 ) | ( w8229 & w8240 ) ;
  assign w8244 = ~w8229 & w8243 ;
  assign w8245 = w7867 & ~w8222 ;
  assign w8246 = ~w8211 & w8245 ;
  assign w8247 = ~w8224 & w8246 ;
  assign w8248 = \pi043 & w8225 ;
  assign w8249 = ( \pi042 & w8225 ) | ( \pi042 & ~w8248 ) | ( w8225 & ~w8248 ) ;
  assign w8250 = ( ~\pi042 & w8247 ) | ( ~\pi042 & w8249 ) | ( w8247 & w8249 ) ;
  assign w8251 = \pi044 ^ w8250 ;
  assign w8252 = w8244 | w8251 ;
  assign w8253 = ( w7175 & w8242 ) | ( w7175 & ~w8252 ) | ( w8242 & ~w8252 ) ;
  assign w8254 = w7175 & w8253 ;
  assign w8255 = ( w7871 & ~w7879 ) | ( w7871 & w8225 ) | ( ~w7879 & w8225 ) ;
  assign w8256 = ~w7871 & w8255 ;
  assign w8257 = \pi045 ^ w8256 ;
  assign w8258 = w7880 ^ w8257 ;
  assign w8259 = ( ~w7175 & w8242 ) | ( ~w7175 & w8252 ) | ( w8242 & w8252 ) ;
  assign w8260 = ~w8242 & w8259 ;
  assign w8261 = w8258 | w8260 ;
  assign w8262 = ( w6841 & w8254 ) | ( w6841 & ~w8261 ) | ( w8254 & ~w8261 ) ;
  assign w8263 = w6841 & w8262 ;
  assign w8264 = w7884 | w7886 ;
  assign w8265 = w8225 & ~w8264 ;
  assign w8266 = w7893 ^ w8265 ;
  assign w8267 = ( ~w6841 & w8254 ) | ( ~w6841 & w8261 ) | ( w8254 & w8261 ) ;
  assign w8268 = ~w8254 & w8267 ;
  assign w8269 = w8266 | w8268 ;
  assign w8270 = ( w6515 & w8263 ) | ( w6515 & ~w8269 ) | ( w8263 & ~w8269 ) ;
  assign w8271 = w6515 & w8270 ;
  assign w8272 = w7896 | w7902 ;
  assign w8273 = w8225 & ~w8272 ;
  assign w8274 = w7900 ^ w8273 ;
  assign w8275 = ( ~w6515 & w8263 ) | ( ~w6515 & w8269 ) | ( w8263 & w8269 ) ;
  assign w8276 = ~w8263 & w8275 ;
  assign w8277 = w8274 | w8276 ;
  assign w8278 = ( w6197 & w8271 ) | ( w6197 & ~w8277 ) | ( w8271 & ~w8277 ) ;
  assign w8279 = w6197 & w8278 ;
  assign w8280 = w7905 | w7910 ;
  assign w8281 = w8225 & ~w8280 ;
  assign w8282 = w7908 ^ w8281 ;
  assign w8283 = ( ~w6197 & w8271 ) | ( ~w6197 & w8277 ) | ( w8271 & w8277 ) ;
  assign w8284 = ~w8271 & w8283 ;
  assign w8285 = w8282 | w8284 ;
  assign w8286 = ( w5887 & w8279 ) | ( w5887 & ~w8285 ) | ( w8279 & ~w8285 ) ;
  assign w8287 = w5887 & w8286 ;
  assign w8288 = w7913 | w7918 ;
  assign w8289 = w8225 & ~w8288 ;
  assign w8290 = w7916 ^ w8289 ;
  assign w8291 = ( ~w5887 & w8279 ) | ( ~w5887 & w8285 ) | ( w8279 & w8285 ) ;
  assign w8292 = ~w8279 & w8291 ;
  assign w8293 = w8290 | w8292 ;
  assign w8294 = ( w5585 & w8287 ) | ( w5585 & ~w8293 ) | ( w8287 & ~w8293 ) ;
  assign w8295 = w5585 & w8294 ;
  assign w8296 = w7921 | w7926 ;
  assign w8297 = w8225 & ~w8296 ;
  assign w8298 = w7924 ^ w8297 ;
  assign w8299 = ( ~w5585 & w8287 ) | ( ~w5585 & w8293 ) | ( w8287 & w8293 ) ;
  assign w8300 = ~w8287 & w8299 ;
  assign w8301 = w8298 | w8300 ;
  assign w8302 = ( w5291 & w8295 ) | ( w5291 & ~w8301 ) | ( w8295 & ~w8301 ) ;
  assign w8303 = w5291 & w8302 ;
  assign w8304 = w7929 | w7934 ;
  assign w8305 = w8225 & ~w8304 ;
  assign w8306 = w7932 ^ w8305 ;
  assign w8307 = ( ~w5291 & w8295 ) | ( ~w5291 & w8301 ) | ( w8295 & w8301 ) ;
  assign w8308 = ~w8295 & w8307 ;
  assign w8309 = w8306 | w8308 ;
  assign w8310 = ( w5005 & w8303 ) | ( w5005 & ~w8309 ) | ( w8303 & ~w8309 ) ;
  assign w8311 = w5005 & w8310 ;
  assign w8312 = w7937 | w7942 ;
  assign w8313 = w8225 & ~w8312 ;
  assign w8314 = w7940 ^ w8313 ;
  assign w8315 = ( ~w5005 & w8303 ) | ( ~w5005 & w8309 ) | ( w8303 & w8309 ) ;
  assign w8316 = ~w8303 & w8315 ;
  assign w8317 = w8314 | w8316 ;
  assign w8318 = ( w4727 & w8311 ) | ( w4727 & ~w8317 ) | ( w8311 & ~w8317 ) ;
  assign w8319 = w4727 & w8318 ;
  assign w8320 = w7945 | w7950 ;
  assign w8321 = w8225 & ~w8320 ;
  assign w8322 = w7948 ^ w8321 ;
  assign w8323 = ( ~w4727 & w8311 ) | ( ~w4727 & w8317 ) | ( w8311 & w8317 ) ;
  assign w8324 = ~w8311 & w8323 ;
  assign w8325 = w8322 | w8324 ;
  assign w8326 = ( w4457 & w8319 ) | ( w4457 & ~w8325 ) | ( w8319 & ~w8325 ) ;
  assign w8327 = w4457 & w8326 ;
  assign w8328 = w7953 | w7958 ;
  assign w8329 = w8225 & ~w8328 ;
  assign w8330 = w7956 ^ w8329 ;
  assign w8331 = ( ~w4457 & w8319 ) | ( ~w4457 & w8325 ) | ( w8319 & w8325 ) ;
  assign w8332 = ~w8319 & w8331 ;
  assign w8333 = w8330 | w8332 ;
  assign w8334 = ( w4195 & w8327 ) | ( w4195 & ~w8333 ) | ( w8327 & ~w8333 ) ;
  assign w8335 = w4195 & w8334 ;
  assign w8336 = w7961 | w7966 ;
  assign w8337 = w8225 & ~w8336 ;
  assign w8338 = w7964 ^ w8337 ;
  assign w8339 = ( ~w4195 & w8327 ) | ( ~w4195 & w8333 ) | ( w8327 & w8333 ) ;
  assign w8340 = ~w8327 & w8339 ;
  assign w8341 = w8338 | w8340 ;
  assign w8342 = ( w3941 & w8335 ) | ( w3941 & ~w8341 ) | ( w8335 & ~w8341 ) ;
  assign w8343 = w3941 & w8342 ;
  assign w8344 = w7969 | w7974 ;
  assign w8345 = w8225 & ~w8344 ;
  assign w8346 = w7972 ^ w8345 ;
  assign w8347 = ( ~w3941 & w8335 ) | ( ~w3941 & w8341 ) | ( w8335 & w8341 ) ;
  assign w8348 = ~w8335 & w8347 ;
  assign w8349 = w8346 | w8348 ;
  assign w8350 = ( w3695 & w8343 ) | ( w3695 & ~w8349 ) | ( w8343 & ~w8349 ) ;
  assign w8351 = w3695 & w8350 ;
  assign w8352 = w7977 | w7982 ;
  assign w8353 = w8225 & ~w8352 ;
  assign w8354 = w7980 ^ w8353 ;
  assign w8355 = ( ~w3695 & w8343 ) | ( ~w3695 & w8349 ) | ( w8343 & w8349 ) ;
  assign w8356 = ~w8343 & w8355 ;
  assign w8357 = w8354 | w8356 ;
  assign w8358 = ( w3457 & w8351 ) | ( w3457 & ~w8357 ) | ( w8351 & ~w8357 ) ;
  assign w8359 = w3457 & w8358 ;
  assign w8360 = w7985 | w7990 ;
  assign w8361 = w8225 & ~w8360 ;
  assign w8362 = w7988 ^ w8361 ;
  assign w8363 = ( ~w3457 & w8351 ) | ( ~w3457 & w8357 ) | ( w8351 & w8357 ) ;
  assign w8364 = ~w8351 & w8363 ;
  assign w8365 = w8362 | w8364 ;
  assign w8366 = ( w3227 & w8359 ) | ( w3227 & ~w8365 ) | ( w8359 & ~w8365 ) ;
  assign w8367 = w3227 & w8366 ;
  assign w8368 = w7993 | w7998 ;
  assign w8369 = w8225 & ~w8368 ;
  assign w8370 = w7996 ^ w8369 ;
  assign w8371 = ( ~w3227 & w8359 ) | ( ~w3227 & w8365 ) | ( w8359 & w8365 ) ;
  assign w8372 = ~w8359 & w8371 ;
  assign w8373 = w8370 | w8372 ;
  assign w8374 = ( w3005 & w8367 ) | ( w3005 & ~w8373 ) | ( w8367 & ~w8373 ) ;
  assign w8375 = w3005 & w8374 ;
  assign w8376 = w8001 | w8006 ;
  assign w8377 = w8225 & ~w8376 ;
  assign w8378 = w8004 ^ w8377 ;
  assign w8379 = ( ~w3005 & w8367 ) | ( ~w3005 & w8373 ) | ( w8367 & w8373 ) ;
  assign w8380 = ~w8367 & w8379 ;
  assign w8381 = w8378 | w8380 ;
  assign w8382 = ( w2791 & w8375 ) | ( w2791 & ~w8381 ) | ( w8375 & ~w8381 ) ;
  assign w8383 = w2791 & w8382 ;
  assign w8384 = w8009 | w8014 ;
  assign w8385 = w8225 & ~w8384 ;
  assign w8386 = w8012 ^ w8385 ;
  assign w8387 = ( ~w2791 & w8375 ) | ( ~w2791 & w8381 ) | ( w8375 & w8381 ) ;
  assign w8388 = ~w8375 & w8387 ;
  assign w8389 = w8386 | w8388 ;
  assign w8390 = ( w2585 & w8383 ) | ( w2585 & ~w8389 ) | ( w8383 & ~w8389 ) ;
  assign w8391 = w2585 & w8390 ;
  assign w8392 = w8017 | w8022 ;
  assign w8393 = w8225 & ~w8392 ;
  assign w8394 = w8020 ^ w8393 ;
  assign w8395 = ( ~w2585 & w8383 ) | ( ~w2585 & w8389 ) | ( w8383 & w8389 ) ;
  assign w8396 = ~w8383 & w8395 ;
  assign w8397 = w8394 | w8396 ;
  assign w8398 = ( w2387 & w8391 ) | ( w2387 & ~w8397 ) | ( w8391 & ~w8397 ) ;
  assign w8399 = w2387 & w8398 ;
  assign w8400 = w8025 | w8030 ;
  assign w8401 = w8225 & ~w8400 ;
  assign w8402 = w8028 ^ w8401 ;
  assign w8403 = ( ~w2387 & w8391 ) | ( ~w2387 & w8397 ) | ( w8391 & w8397 ) ;
  assign w8404 = ~w8391 & w8403 ;
  assign w8405 = w8402 | w8404 ;
  assign w8406 = ( w2197 & w8399 ) | ( w2197 & ~w8405 ) | ( w8399 & ~w8405 ) ;
  assign w8407 = w2197 & w8406 ;
  assign w8408 = w8033 | w8038 ;
  assign w8409 = w8225 & ~w8408 ;
  assign w8410 = w8036 ^ w8409 ;
  assign w8411 = ( ~w2197 & w8399 ) | ( ~w2197 & w8405 ) | ( w8399 & w8405 ) ;
  assign w8412 = ~w8399 & w8411 ;
  assign w8413 = w8410 | w8412 ;
  assign w8414 = ( w2015 & w8407 ) | ( w2015 & ~w8413 ) | ( w8407 & ~w8413 ) ;
  assign w8415 = w2015 & w8414 ;
  assign w8416 = ( ~w2015 & w8407 ) | ( ~w2015 & w8413 ) | ( w8407 & w8413 ) ;
  assign w8417 = ~w8407 & w8416 ;
  assign w8418 = w8041 | w8043 ;
  assign w8419 = w8225 & ~w8418 ;
  assign w8420 = w8046 ^ w8419 ;
  assign w8421 = w8417 | w8420 ;
  assign w8422 = ( w1841 & w8415 ) | ( w1841 & ~w8421 ) | ( w8415 & ~w8421 ) ;
  assign w8423 = w1841 & w8422 ;
  assign w8424 = w8049 | w8054 ;
  assign w8425 = w8225 & ~w8424 ;
  assign w8426 = w8052 ^ w8425 ;
  assign w8427 = ( ~w1841 & w8415 ) | ( ~w1841 & w8421 ) | ( w8415 & w8421 ) ;
  assign w8428 = ~w8415 & w8427 ;
  assign w8429 = w8426 | w8428 ;
  assign w8430 = ( w1675 & w8423 ) | ( w1675 & ~w8429 ) | ( w8423 & ~w8429 ) ;
  assign w8431 = w1675 & w8430 ;
  assign w8432 = w8057 | w8062 ;
  assign w8433 = w8225 & ~w8432 ;
  assign w8434 = w8060 ^ w8433 ;
  assign w8435 = ( ~w1675 & w8423 ) | ( ~w1675 & w8429 ) | ( w8423 & w8429 ) ;
  assign w8436 = ~w8423 & w8435 ;
  assign w8437 = w8434 | w8436 ;
  assign w8438 = ( w1517 & w8431 ) | ( w1517 & ~w8437 ) | ( w8431 & ~w8437 ) ;
  assign w8439 = w1517 & w8438 ;
  assign w8440 = w8065 | w8070 ;
  assign w8441 = w8225 & ~w8440 ;
  assign w8442 = w8068 ^ w8441 ;
  assign w8443 = ( ~w1517 & w8431 ) | ( ~w1517 & w8437 ) | ( w8431 & w8437 ) ;
  assign w8444 = ~w8431 & w8443 ;
  assign w8445 = w8442 | w8444 ;
  assign w8446 = ( w1367 & w8439 ) | ( w1367 & ~w8445 ) | ( w8439 & ~w8445 ) ;
  assign w8447 = w1367 & w8446 ;
  assign w8448 = w8073 | w8078 ;
  assign w8449 = w8225 & ~w8448 ;
  assign w8450 = w8076 ^ w8449 ;
  assign w8451 = ( ~w1367 & w8439 ) | ( ~w1367 & w8445 ) | ( w8439 & w8445 ) ;
  assign w8452 = ~w8439 & w8451 ;
  assign w8453 = w8450 | w8452 ;
  assign w8454 = ( w1225 & w8447 ) | ( w1225 & ~w8453 ) | ( w8447 & ~w8453 ) ;
  assign w8455 = w1225 & w8454 ;
  assign w8456 = w8081 | w8086 ;
  assign w8457 = w8225 & ~w8456 ;
  assign w8458 = w8084 ^ w8457 ;
  assign w8459 = ( ~w1225 & w8447 ) | ( ~w1225 & w8453 ) | ( w8447 & w8453 ) ;
  assign w8460 = ~w8447 & w8459 ;
  assign w8461 = w8458 | w8460 ;
  assign w8462 = ( w1091 & w8455 ) | ( w1091 & ~w8461 ) | ( w8455 & ~w8461 ) ;
  assign w8463 = w1091 & w8462 ;
  assign w8464 = w8089 | w8094 ;
  assign w8465 = w8225 & ~w8464 ;
  assign w8466 = w8092 ^ w8465 ;
  assign w8467 = ( ~w1091 & w8455 ) | ( ~w1091 & w8461 ) | ( w8455 & w8461 ) ;
  assign w8468 = ~w8455 & w8467 ;
  assign w8469 = w8466 | w8468 ;
  assign w8470 = ( w965 & w8463 ) | ( w965 & ~w8469 ) | ( w8463 & ~w8469 ) ;
  assign w8471 = w965 & w8470 ;
  assign w8472 = w8097 | w8102 ;
  assign w8473 = w8225 & ~w8472 ;
  assign w8474 = w8100 ^ w8473 ;
  assign w8475 = ( ~w965 & w8463 ) | ( ~w965 & w8469 ) | ( w8463 & w8469 ) ;
  assign w8476 = ~w8463 & w8475 ;
  assign w8477 = w8474 | w8476 ;
  assign w8478 = ( w847 & w8471 ) | ( w847 & ~w8477 ) | ( w8471 & ~w8477 ) ;
  assign w8479 = w847 & w8478 ;
  assign w8480 = w8105 | w8110 ;
  assign w8481 = w8225 & ~w8480 ;
  assign w8482 = w8108 ^ w8481 ;
  assign w8483 = ( ~w847 & w8471 ) | ( ~w847 & w8477 ) | ( w8471 & w8477 ) ;
  assign w8484 = ~w8471 & w8483 ;
  assign w8485 = w8482 | w8484 ;
  assign w8486 = ( w737 & w8479 ) | ( w737 & ~w8485 ) | ( w8479 & ~w8485 ) ;
  assign w8487 = w737 & w8486 ;
  assign w8488 = w8113 | w8118 ;
  assign w8489 = w8225 & ~w8488 ;
  assign w8490 = w8116 ^ w8489 ;
  assign w8491 = ( ~w737 & w8479 ) | ( ~w737 & w8485 ) | ( w8479 & w8485 ) ;
  assign w8492 = ~w8479 & w8491 ;
  assign w8493 = w8490 | w8492 ;
  assign w8494 = ( w635 & w8487 ) | ( w635 & ~w8493 ) | ( w8487 & ~w8493 ) ;
  assign w8495 = w635 & w8494 ;
  assign w8496 = w8121 | w8126 ;
  assign w8497 = w8225 & ~w8496 ;
  assign w8498 = w8124 ^ w8497 ;
  assign w8499 = ( ~w635 & w8487 ) | ( ~w635 & w8493 ) | ( w8487 & w8493 ) ;
  assign w8500 = ~w8487 & w8499 ;
  assign w8501 = w8498 | w8500 ;
  assign w8502 = ( w541 & w8495 ) | ( w541 & ~w8501 ) | ( w8495 & ~w8501 ) ;
  assign w8503 = w541 & w8502 ;
  assign w8504 = w8129 | w8134 ;
  assign w8505 = w8225 & ~w8504 ;
  assign w8506 = w8132 ^ w8505 ;
  assign w8507 = ( ~w541 & w8495 ) | ( ~w541 & w8501 ) | ( w8495 & w8501 ) ;
  assign w8508 = ~w8495 & w8507 ;
  assign w8509 = w8506 | w8508 ;
  assign w8510 = ( w455 & w8503 ) | ( w455 & ~w8509 ) | ( w8503 & ~w8509 ) ;
  assign w8511 = w455 & w8510 ;
  assign w8512 = w8137 | w8142 ;
  assign w8513 = w8225 & ~w8512 ;
  assign w8514 = w8140 ^ w8513 ;
  assign w8515 = ( ~w455 & w8503 ) | ( ~w455 & w8509 ) | ( w8503 & w8509 ) ;
  assign w8516 = ~w8503 & w8515 ;
  assign w8517 = w8514 | w8516 ;
  assign w8518 = ( w377 & w8511 ) | ( w377 & ~w8517 ) | ( w8511 & ~w8517 ) ;
  assign w8519 = w377 & w8518 ;
  assign w8520 = w8145 | w8150 ;
  assign w8521 = w8225 & ~w8520 ;
  assign w8522 = w8148 ^ w8521 ;
  assign w8523 = ( ~w377 & w8511 ) | ( ~w377 & w8517 ) | ( w8511 & w8517 ) ;
  assign w8524 = ~w8511 & w8523 ;
  assign w8525 = w8522 | w8524 ;
  assign w8526 = ( w307 & w8519 ) | ( w307 & ~w8525 ) | ( w8519 & ~w8525 ) ;
  assign w8527 = w307 & w8526 ;
  assign w8528 = w8153 | w8158 ;
  assign w8529 = w8225 & ~w8528 ;
  assign w8530 = w8156 ^ w8529 ;
  assign w8531 = ( ~w307 & w8519 ) | ( ~w307 & w8525 ) | ( w8519 & w8525 ) ;
  assign w8532 = ~w8519 & w8531 ;
  assign w8533 = w8530 | w8532 ;
  assign w8534 = ( w246 & w8527 ) | ( w246 & ~w8533 ) | ( w8527 & ~w8533 ) ;
  assign w8535 = w246 & w8534 ;
  assign w8536 = w8161 | w8166 ;
  assign w8537 = w8225 & ~w8536 ;
  assign w8538 = w8164 ^ w8537 ;
  assign w8539 = ( ~w246 & w8527 ) | ( ~w246 & w8533 ) | ( w8527 & w8533 ) ;
  assign w8540 = ~w8527 & w8539 ;
  assign w8541 = w8538 | w8540 ;
  assign w8542 = ( w185 & w8535 ) | ( w185 & ~w8541 ) | ( w8535 & ~w8541 ) ;
  assign w8543 = w185 & w8542 ;
  assign w8544 = w8169 | w8174 ;
  assign w8545 = w8225 & ~w8544 ;
  assign w8546 = w8172 ^ w8545 ;
  assign w8547 = ( ~w185 & w8535 ) | ( ~w185 & w8541 ) | ( w8535 & w8541 ) ;
  assign w8548 = ~w8535 & w8547 ;
  assign w8549 = w8546 | w8548 ;
  assign w8550 = ( w145 & w8543 ) | ( w145 & ~w8549 ) | ( w8543 & ~w8549 ) ;
  assign w8551 = w145 & w8550 ;
  assign w8552 = w8177 | w8182 ;
  assign w8553 = w8225 & ~w8552 ;
  assign w8554 = w8180 ^ w8553 ;
  assign w8555 = ( ~w145 & w8543 ) | ( ~w145 & w8549 ) | ( w8543 & w8549 ) ;
  assign w8556 = ~w8543 & w8555 ;
  assign w8557 = w8554 | w8556 ;
  assign w8558 = ( w132 & w8551 ) | ( w132 & ~w8557 ) | ( w8551 & ~w8557 ) ;
  assign w8559 = w132 & w8558 ;
  assign w8560 = w8185 | w8190 ;
  assign w8561 = w8225 & ~w8560 ;
  assign w8562 = w8188 ^ w8561 ;
  assign w8563 = ( ~w132 & w8551 ) | ( ~w132 & w8557 ) | ( w8551 & w8557 ) ;
  assign w8564 = ~w8551 & w8563 ;
  assign w8565 = w8562 | w8564 ;
  assign w8566 = ~w8559 & w8565 ;
  assign w8567 = w8193 | w8198 ;
  assign w8568 = w8225 & ~w8567 ;
  assign w8569 = w8196 ^ w8568 ;
  assign w8570 = ( ~w8211 & w8566 ) | ( ~w8211 & w8569 ) | ( w8566 & w8569 ) ;
  assign w8571 = w8200 & ~w8570 ;
  assign w8572 = ~w8203 & w8225 ;
  assign w8573 = ( w8570 & ~w8571 ) | ( w8570 & w8572 ) | ( ~w8571 & w8572 ) ;
  assign w8574 = w8211 | w8573 ;
  assign w8575 = ~w129 & w8574 ;
  assign w8576 = ( w8559 & w8565 ) | ( w8559 & w8569 ) | ( w8565 & w8569 ) ;
  assign w8577 = ~w8559 & w8576 ;
  assign w8578 = ( w129 & w8200 ) | ( w129 & w8203 ) | ( w8200 & w8203 ) ;
  assign w8579 = ( w8203 & ~w8225 ) | ( w8203 & w8578 ) | ( ~w8225 & w8578 ) ;
  assign w8580 = w8200 & w8579 ;
  assign w8581 = w8578 ^ w8580 ;
  assign w8582 = ( w7835 & w7840 ) | ( w7835 & w7867 ) | ( w7840 & w7867 ) ;
  assign w8583 = w7867 & ~w8582 ;
  assign w8584 = w7838 ^ w8583 ;
  assign w8585 = ( ~w8215 & w8222 ) | ( ~w8215 & w8584 ) | ( w8222 & w8584 ) ;
  assign w8586 = ~w8222 & w8585 ;
  assign w8587 = ( ~w8209 & w8211 ) | ( ~w8209 & w8586 ) | ( w8211 & w8586 ) ;
  assign w8588 = ~w8211 & w8587 ;
  assign w8589 = w8577 | w8588 ;
  assign w8590 = ( w8575 & ~w8577 ) | ( w8575 & w8581 ) | ( ~w8577 & w8581 ) ;
  assign w8591 = w8589 | w8590 ;
  assign w8592 = ( ~\pi039 & \pi040 ) | ( ~\pi039 & w8225 ) | ( \pi040 & w8225 ) ;
  assign w8593 = ( ~\pi038 & \pi040 ) | ( ~\pi038 & w8592 ) | ( \pi040 & w8592 ) ;
  assign w8594 = ( ~\pi040 & w8225 ) | ( ~\pi040 & w8591 ) | ( w8225 & w8591 ) ;
  assign w8595 = w8593 & w8594 ;
  assign w8596 = ( w8211 & w8215 ) | ( w8211 & ~w8222 ) | ( w8215 & ~w8222 ) ;
  assign w8597 = \pi039 & ~w8596 ;
  assign w8598 = \pi038 | \pi040 ;
  assign w8599 = ( ~w8596 & w8597 ) | ( ~w8596 & w8598 ) | ( w8597 & w8598 ) ;
  assign w8600 = ~w8222 & w8599 ;
  assign w8601 = ~w8209 & w8600 ;
  assign w8602 = ( \pi040 & w8591 ) | ( \pi040 & ~w8600 ) | ( w8591 & ~w8600 ) ;
  assign w8603 = w8601 & ~w8602 ;
  assign w8604 = ~\pi040 & w8591 ;
  assign w8605 = \pi041 ^ w8604 ;
  assign w8606 = w8603 | w8605 ;
  assign w8607 = ( w7867 & w8595 ) | ( w7867 & ~w8606 ) | ( w8595 & ~w8606 ) ;
  assign w8608 = w7867 & w8607 ;
  assign w8609 = ( ~w7867 & w8595 ) | ( ~w7867 & w8606 ) | ( w8595 & w8606 ) ;
  assign w8610 = ~w8595 & w8609 ;
  assign w8611 = w8225 & ~w8588 ;
  assign w8612 = ~w8577 & w8611 ;
  assign w8613 = ~w8590 & w8612 ;
  assign w8614 = \pi041 & w8591 ;
  assign w8615 = ( \pi040 & w8591 ) | ( \pi040 & ~w8614 ) | ( w8591 & ~w8614 ) ;
  assign w8616 = ( ~\pi040 & w8613 ) | ( ~\pi040 & w8615 ) | ( w8613 & w8615 ) ;
  assign w8617 = \pi042 ^ w8616 ;
  assign w8618 = w8610 | w8617 ;
  assign w8619 = ( w7517 & w8608 ) | ( w7517 & ~w8618 ) | ( w8608 & ~w8618 ) ;
  assign w8620 = w7517 & w8619 ;
  assign w8621 = ( w8229 & ~w8237 ) | ( w8229 & w8591 ) | ( ~w8237 & w8591 ) ;
  assign w8622 = ~w8229 & w8621 ;
  assign w8623 = \pi043 ^ w8622 ;
  assign w8624 = w8238 ^ w8623 ;
  assign w8625 = ( ~w7517 & w8608 ) | ( ~w7517 & w8618 ) | ( w8608 & w8618 ) ;
  assign w8626 = ~w8608 & w8625 ;
  assign w8627 = w8624 | w8626 ;
  assign w8628 = ( w7175 & w8620 ) | ( w7175 & ~w8627 ) | ( w8620 & ~w8627 ) ;
  assign w8629 = w7175 & w8628 ;
  assign w8630 = w8242 | w8244 ;
  assign w8631 = w8591 & ~w8630 ;
  assign w8632 = w8251 ^ w8631 ;
  assign w8633 = ( ~w7175 & w8620 ) | ( ~w7175 & w8627 ) | ( w8620 & w8627 ) ;
  assign w8634 = ~w8620 & w8633 ;
  assign w8635 = w8632 | w8634 ;
  assign w8636 = ( w6841 & w8629 ) | ( w6841 & ~w8635 ) | ( w8629 & ~w8635 ) ;
  assign w8637 = w6841 & w8636 ;
  assign w8638 = w8254 | w8260 ;
  assign w8639 = w8591 & ~w8638 ;
  assign w8640 = w8258 ^ w8639 ;
  assign w8641 = ( ~w6841 & w8629 ) | ( ~w6841 & w8635 ) | ( w8629 & w8635 ) ;
  assign w8642 = ~w8629 & w8641 ;
  assign w8643 = w8640 | w8642 ;
  assign w8644 = ( w6515 & w8637 ) | ( w6515 & ~w8643 ) | ( w8637 & ~w8643 ) ;
  assign w8645 = w6515 & w8644 ;
  assign w8646 = w8263 | w8268 ;
  assign w8647 = w8591 & ~w8646 ;
  assign w8648 = w8266 ^ w8647 ;
  assign w8649 = ( ~w6515 & w8637 ) | ( ~w6515 & w8643 ) | ( w8637 & w8643 ) ;
  assign w8650 = ~w8637 & w8649 ;
  assign w8651 = w8648 | w8650 ;
  assign w8652 = ( w6197 & w8645 ) | ( w6197 & ~w8651 ) | ( w8645 & ~w8651 ) ;
  assign w8653 = w6197 & w8652 ;
  assign w8654 = w8271 | w8276 ;
  assign w8655 = w8591 & ~w8654 ;
  assign w8656 = w8274 ^ w8655 ;
  assign w8657 = ( ~w6197 & w8645 ) | ( ~w6197 & w8651 ) | ( w8645 & w8651 ) ;
  assign w8658 = ~w8645 & w8657 ;
  assign w8659 = w8656 | w8658 ;
  assign w8660 = ( w5887 & w8653 ) | ( w5887 & ~w8659 ) | ( w8653 & ~w8659 ) ;
  assign w8661 = w5887 & w8660 ;
  assign w8662 = w8279 | w8284 ;
  assign w8663 = w8591 & ~w8662 ;
  assign w8664 = w8282 ^ w8663 ;
  assign w8665 = ( ~w5887 & w8653 ) | ( ~w5887 & w8659 ) | ( w8653 & w8659 ) ;
  assign w8666 = ~w8653 & w8665 ;
  assign w8667 = w8664 | w8666 ;
  assign w8668 = ( w5585 & w8661 ) | ( w5585 & ~w8667 ) | ( w8661 & ~w8667 ) ;
  assign w8669 = w5585 & w8668 ;
  assign w8670 = w8287 | w8292 ;
  assign w8671 = w8591 & ~w8670 ;
  assign w8672 = w8290 ^ w8671 ;
  assign w8673 = ( ~w5585 & w8661 ) | ( ~w5585 & w8667 ) | ( w8661 & w8667 ) ;
  assign w8674 = ~w8661 & w8673 ;
  assign w8675 = w8672 | w8674 ;
  assign w8676 = ( w5291 & w8669 ) | ( w5291 & ~w8675 ) | ( w8669 & ~w8675 ) ;
  assign w8677 = w5291 & w8676 ;
  assign w8678 = w8295 | w8300 ;
  assign w8679 = w8591 & ~w8678 ;
  assign w8680 = w8298 ^ w8679 ;
  assign w8681 = ( ~w5291 & w8669 ) | ( ~w5291 & w8675 ) | ( w8669 & w8675 ) ;
  assign w8682 = ~w8669 & w8681 ;
  assign w8683 = w8680 | w8682 ;
  assign w8684 = ( w5005 & w8677 ) | ( w5005 & ~w8683 ) | ( w8677 & ~w8683 ) ;
  assign w8685 = w5005 & w8684 ;
  assign w8686 = w8303 | w8308 ;
  assign w8687 = w8591 & ~w8686 ;
  assign w8688 = w8306 ^ w8687 ;
  assign w8689 = ( ~w5005 & w8677 ) | ( ~w5005 & w8683 ) | ( w8677 & w8683 ) ;
  assign w8690 = ~w8677 & w8689 ;
  assign w8691 = w8688 | w8690 ;
  assign w8692 = ( w4727 & w8685 ) | ( w4727 & ~w8691 ) | ( w8685 & ~w8691 ) ;
  assign w8693 = w4727 & w8692 ;
  assign w8694 = w8311 | w8316 ;
  assign w8695 = w8591 & ~w8694 ;
  assign w8696 = w8314 ^ w8695 ;
  assign w8697 = ( ~w4727 & w8685 ) | ( ~w4727 & w8691 ) | ( w8685 & w8691 ) ;
  assign w8698 = ~w8685 & w8697 ;
  assign w8699 = w8696 | w8698 ;
  assign w8700 = ( w4457 & w8693 ) | ( w4457 & ~w8699 ) | ( w8693 & ~w8699 ) ;
  assign w8701 = w4457 & w8700 ;
  assign w8702 = w8319 | w8324 ;
  assign w8703 = w8591 & ~w8702 ;
  assign w8704 = w8322 ^ w8703 ;
  assign w8705 = ( ~w4457 & w8693 ) | ( ~w4457 & w8699 ) | ( w8693 & w8699 ) ;
  assign w8706 = ~w8693 & w8705 ;
  assign w8707 = w8704 | w8706 ;
  assign w8708 = ( w4195 & w8701 ) | ( w4195 & ~w8707 ) | ( w8701 & ~w8707 ) ;
  assign w8709 = w4195 & w8708 ;
  assign w8710 = w8327 | w8332 ;
  assign w8711 = w8591 & ~w8710 ;
  assign w8712 = w8330 ^ w8711 ;
  assign w8713 = ( ~w4195 & w8701 ) | ( ~w4195 & w8707 ) | ( w8701 & w8707 ) ;
  assign w8714 = ~w8701 & w8713 ;
  assign w8715 = w8712 | w8714 ;
  assign w8716 = ( w3941 & w8709 ) | ( w3941 & ~w8715 ) | ( w8709 & ~w8715 ) ;
  assign w8717 = w3941 & w8716 ;
  assign w8718 = w8335 | w8340 ;
  assign w8719 = w8591 & ~w8718 ;
  assign w8720 = w8338 ^ w8719 ;
  assign w8721 = ( ~w3941 & w8709 ) | ( ~w3941 & w8715 ) | ( w8709 & w8715 ) ;
  assign w8722 = ~w8709 & w8721 ;
  assign w8723 = w8720 | w8722 ;
  assign w8724 = ( w3695 & w8717 ) | ( w3695 & ~w8723 ) | ( w8717 & ~w8723 ) ;
  assign w8725 = w3695 & w8724 ;
  assign w8726 = w8343 | w8348 ;
  assign w8727 = w8591 & ~w8726 ;
  assign w8728 = w8346 ^ w8727 ;
  assign w8729 = ( ~w3695 & w8717 ) | ( ~w3695 & w8723 ) | ( w8717 & w8723 ) ;
  assign w8730 = ~w8717 & w8729 ;
  assign w8731 = w8728 | w8730 ;
  assign w8732 = ( w3457 & w8725 ) | ( w3457 & ~w8731 ) | ( w8725 & ~w8731 ) ;
  assign w8733 = w3457 & w8732 ;
  assign w8734 = w8351 | w8356 ;
  assign w8735 = w8591 & ~w8734 ;
  assign w8736 = w8354 ^ w8735 ;
  assign w8737 = ( ~w3457 & w8725 ) | ( ~w3457 & w8731 ) | ( w8725 & w8731 ) ;
  assign w8738 = ~w8725 & w8737 ;
  assign w8739 = w8736 | w8738 ;
  assign w8740 = ( w3227 & w8733 ) | ( w3227 & ~w8739 ) | ( w8733 & ~w8739 ) ;
  assign w8741 = w3227 & w8740 ;
  assign w8742 = w8359 | w8364 ;
  assign w8743 = w8591 & ~w8742 ;
  assign w8744 = w8362 ^ w8743 ;
  assign w8745 = ( ~w3227 & w8733 ) | ( ~w3227 & w8739 ) | ( w8733 & w8739 ) ;
  assign w8746 = ~w8733 & w8745 ;
  assign w8747 = w8744 | w8746 ;
  assign w8748 = ( w3005 & w8741 ) | ( w3005 & ~w8747 ) | ( w8741 & ~w8747 ) ;
  assign w8749 = w3005 & w8748 ;
  assign w8750 = w8367 | w8372 ;
  assign w8751 = w8591 & ~w8750 ;
  assign w8752 = w8370 ^ w8751 ;
  assign w8753 = ( ~w3005 & w8741 ) | ( ~w3005 & w8747 ) | ( w8741 & w8747 ) ;
  assign w8754 = ~w8741 & w8753 ;
  assign w8755 = w8752 | w8754 ;
  assign w8756 = ( w2791 & w8749 ) | ( w2791 & ~w8755 ) | ( w8749 & ~w8755 ) ;
  assign w8757 = w2791 & w8756 ;
  assign w8758 = w8375 | w8380 ;
  assign w8759 = w8591 & ~w8758 ;
  assign w8760 = w8378 ^ w8759 ;
  assign w8761 = ( ~w2791 & w8749 ) | ( ~w2791 & w8755 ) | ( w8749 & w8755 ) ;
  assign w8762 = ~w8749 & w8761 ;
  assign w8763 = w8760 | w8762 ;
  assign w8764 = ( w2585 & w8757 ) | ( w2585 & ~w8763 ) | ( w8757 & ~w8763 ) ;
  assign w8765 = w2585 & w8764 ;
  assign w8766 = w8383 | w8388 ;
  assign w8767 = w8591 & ~w8766 ;
  assign w8768 = w8386 ^ w8767 ;
  assign w8769 = ( ~w2585 & w8757 ) | ( ~w2585 & w8763 ) | ( w8757 & w8763 ) ;
  assign w8770 = ~w8757 & w8769 ;
  assign w8771 = w8768 | w8770 ;
  assign w8772 = ( w2387 & w8765 ) | ( w2387 & ~w8771 ) | ( w8765 & ~w8771 ) ;
  assign w8773 = w2387 & w8772 ;
  assign w8774 = w8391 | w8396 ;
  assign w8775 = w8591 & ~w8774 ;
  assign w8776 = w8394 ^ w8775 ;
  assign w8777 = ( ~w2387 & w8765 ) | ( ~w2387 & w8771 ) | ( w8765 & w8771 ) ;
  assign w8778 = ~w8765 & w8777 ;
  assign w8779 = w8776 | w8778 ;
  assign w8780 = ( w2197 & w8773 ) | ( w2197 & ~w8779 ) | ( w8773 & ~w8779 ) ;
  assign w8781 = w2197 & w8780 ;
  assign w8782 = w8399 | w8404 ;
  assign w8783 = w8591 & ~w8782 ;
  assign w8784 = w8402 ^ w8783 ;
  assign w8785 = ( ~w2197 & w8773 ) | ( ~w2197 & w8779 ) | ( w8773 & w8779 ) ;
  assign w8786 = ~w8773 & w8785 ;
  assign w8787 = w8784 | w8786 ;
  assign w8788 = ( w2015 & w8781 ) | ( w2015 & ~w8787 ) | ( w8781 & ~w8787 ) ;
  assign w8789 = w2015 & w8788 ;
  assign w8790 = w8407 | w8412 ;
  assign w8791 = w8591 & ~w8790 ;
  assign w8792 = w8410 ^ w8791 ;
  assign w8793 = ( ~w2015 & w8781 ) | ( ~w2015 & w8787 ) | ( w8781 & w8787 ) ;
  assign w8794 = ~w8781 & w8793 ;
  assign w8795 = w8792 | w8794 ;
  assign w8796 = ( w1841 & w8789 ) | ( w1841 & ~w8795 ) | ( w8789 & ~w8795 ) ;
  assign w8797 = w1841 & w8796 ;
  assign w8798 = ( ~w1841 & w8789 ) | ( ~w1841 & w8795 ) | ( w8789 & w8795 ) ;
  assign w8799 = ~w8789 & w8798 ;
  assign w8800 = w8415 | w8417 ;
  assign w8801 = w8591 & ~w8800 ;
  assign w8802 = w8420 ^ w8801 ;
  assign w8803 = w8799 | w8802 ;
  assign w8804 = ( w1675 & w8797 ) | ( w1675 & ~w8803 ) | ( w8797 & ~w8803 ) ;
  assign w8805 = w1675 & w8804 ;
  assign w8806 = w8423 | w8428 ;
  assign w8807 = w8591 & ~w8806 ;
  assign w8808 = w8426 ^ w8807 ;
  assign w8809 = ( ~w1675 & w8797 ) | ( ~w1675 & w8803 ) | ( w8797 & w8803 ) ;
  assign w8810 = ~w8797 & w8809 ;
  assign w8811 = w8808 | w8810 ;
  assign w8812 = ( w1517 & w8805 ) | ( w1517 & ~w8811 ) | ( w8805 & ~w8811 ) ;
  assign w8813 = w1517 & w8812 ;
  assign w8814 = w8431 | w8436 ;
  assign w8815 = w8591 & ~w8814 ;
  assign w8816 = w8434 ^ w8815 ;
  assign w8817 = ( ~w1517 & w8805 ) | ( ~w1517 & w8811 ) | ( w8805 & w8811 ) ;
  assign w8818 = ~w8805 & w8817 ;
  assign w8819 = w8816 | w8818 ;
  assign w8820 = ( w1367 & w8813 ) | ( w1367 & ~w8819 ) | ( w8813 & ~w8819 ) ;
  assign w8821 = w1367 & w8820 ;
  assign w8822 = w8439 | w8444 ;
  assign w8823 = w8591 & ~w8822 ;
  assign w8824 = w8442 ^ w8823 ;
  assign w8825 = ( ~w1367 & w8813 ) | ( ~w1367 & w8819 ) | ( w8813 & w8819 ) ;
  assign w8826 = ~w8813 & w8825 ;
  assign w8827 = w8824 | w8826 ;
  assign w8828 = ( w1225 & w8821 ) | ( w1225 & ~w8827 ) | ( w8821 & ~w8827 ) ;
  assign w8829 = w1225 & w8828 ;
  assign w8830 = w8447 | w8452 ;
  assign w8831 = w8591 & ~w8830 ;
  assign w8832 = w8450 ^ w8831 ;
  assign w8833 = ( ~w1225 & w8821 ) | ( ~w1225 & w8827 ) | ( w8821 & w8827 ) ;
  assign w8834 = ~w8821 & w8833 ;
  assign w8835 = w8832 | w8834 ;
  assign w8836 = ( w1091 & w8829 ) | ( w1091 & ~w8835 ) | ( w8829 & ~w8835 ) ;
  assign w8837 = w1091 & w8836 ;
  assign w8838 = w8455 | w8460 ;
  assign w8839 = w8591 & ~w8838 ;
  assign w8840 = w8458 ^ w8839 ;
  assign w8841 = ( ~w1091 & w8829 ) | ( ~w1091 & w8835 ) | ( w8829 & w8835 ) ;
  assign w8842 = ~w8829 & w8841 ;
  assign w8843 = w8840 | w8842 ;
  assign w8844 = ( w965 & w8837 ) | ( w965 & ~w8843 ) | ( w8837 & ~w8843 ) ;
  assign w8845 = w965 & w8844 ;
  assign w8846 = w8463 | w8468 ;
  assign w8847 = w8591 & ~w8846 ;
  assign w8848 = w8466 ^ w8847 ;
  assign w8849 = ( ~w965 & w8837 ) | ( ~w965 & w8843 ) | ( w8837 & w8843 ) ;
  assign w8850 = ~w8837 & w8849 ;
  assign w8851 = w8848 | w8850 ;
  assign w8852 = ( w847 & w8845 ) | ( w847 & ~w8851 ) | ( w8845 & ~w8851 ) ;
  assign w8853 = w847 & w8852 ;
  assign w8854 = w8471 | w8476 ;
  assign w8855 = w8591 & ~w8854 ;
  assign w8856 = w8474 ^ w8855 ;
  assign w8857 = ( ~w847 & w8845 ) | ( ~w847 & w8851 ) | ( w8845 & w8851 ) ;
  assign w8858 = ~w8845 & w8857 ;
  assign w8859 = w8856 | w8858 ;
  assign w8860 = ( w737 & w8853 ) | ( w737 & ~w8859 ) | ( w8853 & ~w8859 ) ;
  assign w8861 = w737 & w8860 ;
  assign w8862 = w8479 | w8484 ;
  assign w8863 = w8591 & ~w8862 ;
  assign w8864 = w8482 ^ w8863 ;
  assign w8865 = ( ~w737 & w8853 ) | ( ~w737 & w8859 ) | ( w8853 & w8859 ) ;
  assign w8866 = ~w8853 & w8865 ;
  assign w8867 = w8864 | w8866 ;
  assign w8868 = ( w635 & w8861 ) | ( w635 & ~w8867 ) | ( w8861 & ~w8867 ) ;
  assign w8869 = w635 & w8868 ;
  assign w8870 = w8487 | w8492 ;
  assign w8871 = w8591 & ~w8870 ;
  assign w8872 = w8490 ^ w8871 ;
  assign w8873 = ( ~w635 & w8861 ) | ( ~w635 & w8867 ) | ( w8861 & w8867 ) ;
  assign w8874 = ~w8861 & w8873 ;
  assign w8875 = w8872 | w8874 ;
  assign w8876 = ( w541 & w8869 ) | ( w541 & ~w8875 ) | ( w8869 & ~w8875 ) ;
  assign w8877 = w541 & w8876 ;
  assign w8878 = w8495 | w8500 ;
  assign w8879 = w8591 & ~w8878 ;
  assign w8880 = w8498 ^ w8879 ;
  assign w8881 = ( ~w541 & w8869 ) | ( ~w541 & w8875 ) | ( w8869 & w8875 ) ;
  assign w8882 = ~w8869 & w8881 ;
  assign w8883 = w8880 | w8882 ;
  assign w8884 = ( w455 & w8877 ) | ( w455 & ~w8883 ) | ( w8877 & ~w8883 ) ;
  assign w8885 = w455 & w8884 ;
  assign w8886 = w8503 | w8508 ;
  assign w8887 = w8591 & ~w8886 ;
  assign w8888 = w8506 ^ w8887 ;
  assign w8889 = ( ~w455 & w8877 ) | ( ~w455 & w8883 ) | ( w8877 & w8883 ) ;
  assign w8890 = ~w8877 & w8889 ;
  assign w8891 = w8888 | w8890 ;
  assign w8892 = ( w377 & w8885 ) | ( w377 & ~w8891 ) | ( w8885 & ~w8891 ) ;
  assign w8893 = w377 & w8892 ;
  assign w8894 = w8511 | w8516 ;
  assign w8895 = w8591 & ~w8894 ;
  assign w8896 = w8514 ^ w8895 ;
  assign w8897 = ( ~w377 & w8885 ) | ( ~w377 & w8891 ) | ( w8885 & w8891 ) ;
  assign w8898 = ~w8885 & w8897 ;
  assign w8899 = w8896 | w8898 ;
  assign w8900 = ( w307 & w8893 ) | ( w307 & ~w8899 ) | ( w8893 & ~w8899 ) ;
  assign w8901 = w307 & w8900 ;
  assign w8902 = w8519 | w8524 ;
  assign w8903 = w8591 & ~w8902 ;
  assign w8904 = w8522 ^ w8903 ;
  assign w8905 = ( ~w307 & w8893 ) | ( ~w307 & w8899 ) | ( w8893 & w8899 ) ;
  assign w8906 = ~w8893 & w8905 ;
  assign w8907 = w8904 | w8906 ;
  assign w8908 = ( w246 & w8901 ) | ( w246 & ~w8907 ) | ( w8901 & ~w8907 ) ;
  assign w8909 = w246 & w8908 ;
  assign w8910 = w8527 | w8532 ;
  assign w8911 = w8591 & ~w8910 ;
  assign w8912 = w8530 ^ w8911 ;
  assign w8913 = ( ~w246 & w8901 ) | ( ~w246 & w8907 ) | ( w8901 & w8907 ) ;
  assign w8914 = ~w8901 & w8913 ;
  assign w8915 = w8912 | w8914 ;
  assign w8916 = ( w185 & w8909 ) | ( w185 & ~w8915 ) | ( w8909 & ~w8915 ) ;
  assign w8917 = w185 & w8916 ;
  assign w8918 = w8535 | w8540 ;
  assign w8919 = w8591 & ~w8918 ;
  assign w8920 = w8538 ^ w8919 ;
  assign w8921 = ( ~w185 & w8909 ) | ( ~w185 & w8915 ) | ( w8909 & w8915 ) ;
  assign w8922 = ~w8909 & w8921 ;
  assign w8923 = w8920 | w8922 ;
  assign w8924 = ( w145 & w8917 ) | ( w145 & ~w8923 ) | ( w8917 & ~w8923 ) ;
  assign w8925 = w145 & w8924 ;
  assign w8926 = w8543 | w8548 ;
  assign w8927 = w8591 & ~w8926 ;
  assign w8928 = w8546 ^ w8927 ;
  assign w8929 = ( ~w145 & w8917 ) | ( ~w145 & w8923 ) | ( w8917 & w8923 ) ;
  assign w8930 = ~w8917 & w8929 ;
  assign w8931 = w8928 | w8930 ;
  assign w8932 = ( w132 & w8925 ) | ( w132 & ~w8931 ) | ( w8925 & ~w8931 ) ;
  assign w8933 = w132 & w8932 ;
  assign w8934 = w8551 | w8556 ;
  assign w8935 = w8591 & ~w8934 ;
  assign w8936 = w8554 ^ w8935 ;
  assign w8937 = ( ~w132 & w8925 ) | ( ~w132 & w8931 ) | ( w8925 & w8931 ) ;
  assign w8938 = ~w8925 & w8937 ;
  assign w8939 = w8936 | w8938 ;
  assign w8940 = ~w8933 & w8939 ;
  assign w8941 = w8559 | w8564 ;
  assign w8942 = w8591 & ~w8941 ;
  assign w8943 = w8562 ^ w8942 ;
  assign w8944 = ( ~w8577 & w8940 ) | ( ~w8577 & w8943 ) | ( w8940 & w8943 ) ;
  assign w8945 = w8566 & ~w8944 ;
  assign w8946 = ~w8569 & w8591 ;
  assign w8947 = ( w8944 & ~w8945 ) | ( w8944 & w8946 ) | ( ~w8945 & w8946 ) ;
  assign w8948 = w8577 | w8947 ;
  assign w8949 = ~w129 & w8948 ;
  assign w8950 = ( w8933 & w8939 ) | ( w8933 & w8943 ) | ( w8939 & w8943 ) ;
  assign w8951 = ~w8933 & w8950 ;
  assign w8952 = ( w129 & w8566 ) | ( w129 & w8569 ) | ( w8566 & w8569 ) ;
  assign w8953 = ( w8569 & ~w8591 ) | ( w8569 & w8952 ) | ( ~w8591 & w8952 ) ;
  assign w8954 = w8566 & w8953 ;
  assign w8955 = w8952 ^ w8954 ;
  assign w8956 = ( w8193 & w8198 ) | ( w8193 & w8225 ) | ( w8198 & w8225 ) ;
  assign w8957 = w8225 & ~w8956 ;
  assign w8958 = w8196 ^ w8957 ;
  assign w8959 = ( ~w8581 & w8588 ) | ( ~w8581 & w8958 ) | ( w8588 & w8958 ) ;
  assign w8960 = ~w8588 & w8959 ;
  assign w8961 = ( ~w8575 & w8577 ) | ( ~w8575 & w8960 ) | ( w8577 & w8960 ) ;
  assign w8962 = ~w8577 & w8961 ;
  assign w8963 = w8951 | w8962 ;
  assign w8964 = ( w8949 & ~w8951 ) | ( w8949 & w8955 ) | ( ~w8951 & w8955 ) ;
  assign w8965 = w8963 | w8964 ;
  assign w8966 = ( ~\pi037 & \pi038 ) | ( ~\pi037 & w8591 ) | ( \pi038 & w8591 ) ;
  assign w8967 = ( ~\pi036 & \pi038 ) | ( ~\pi036 & w8966 ) | ( \pi038 & w8966 ) ;
  assign w8968 = ( ~\pi038 & w8591 ) | ( ~\pi038 & w8965 ) | ( w8591 & w8965 ) ;
  assign w8969 = w8967 & w8968 ;
  assign w8970 = ( w8577 & w8581 ) | ( w8577 & ~w8588 ) | ( w8581 & ~w8588 ) ;
  assign w8971 = \pi037 & ~w8970 ;
  assign w8972 = \pi036 | \pi038 ;
  assign w8973 = ( ~w8970 & w8971 ) | ( ~w8970 & w8972 ) | ( w8971 & w8972 ) ;
  assign w8974 = ~w8588 & w8973 ;
  assign w8975 = ~w8575 & w8974 ;
  assign w8976 = ( \pi038 & w8965 ) | ( \pi038 & ~w8974 ) | ( w8965 & ~w8974 ) ;
  assign w8977 = w8975 & ~w8976 ;
  assign w8978 = ~\pi038 & w8965 ;
  assign w8979 = \pi039 ^ w8978 ;
  assign w8980 = w8977 | w8979 ;
  assign w8981 = ( w8225 & w8969 ) | ( w8225 & ~w8980 ) | ( w8969 & ~w8980 ) ;
  assign w8982 = w8225 & w8981 ;
  assign w8983 = ( ~w8225 & w8969 ) | ( ~w8225 & w8980 ) | ( w8969 & w8980 ) ;
  assign w8984 = ~w8969 & w8983 ;
  assign w8985 = w8591 & ~w8962 ;
  assign w8986 = ~w8951 & w8985 ;
  assign w8987 = ~w8964 & w8986 ;
  assign w8988 = \pi039 & w8965 ;
  assign w8989 = ( \pi038 & w8965 ) | ( \pi038 & ~w8988 ) | ( w8965 & ~w8988 ) ;
  assign w8990 = ( ~\pi038 & w8987 ) | ( ~\pi038 & w8989 ) | ( w8987 & w8989 ) ;
  assign w8991 = \pi040 ^ w8990 ;
  assign w8992 = w8984 | w8991 ;
  assign w8993 = ( w7867 & w8982 ) | ( w7867 & ~w8992 ) | ( w8982 & ~w8992 ) ;
  assign w8994 = w7867 & w8993 ;
  assign w8995 = ( w8595 & ~w8603 ) | ( w8595 & w8965 ) | ( ~w8603 & w8965 ) ;
  assign w8996 = ~w8595 & w8995 ;
  assign w8997 = \pi041 ^ w8996 ;
  assign w8998 = w8604 ^ w8997 ;
  assign w8999 = ( ~w7867 & w8982 ) | ( ~w7867 & w8992 ) | ( w8982 & w8992 ) ;
  assign w9000 = ~w8982 & w8999 ;
  assign w9001 = w8998 | w9000 ;
  assign w9002 = ( w7517 & w8994 ) | ( w7517 & ~w9001 ) | ( w8994 & ~w9001 ) ;
  assign w9003 = w7517 & w9002 ;
  assign w9004 = w8608 | w8610 ;
  assign w9005 = w8965 & ~w9004 ;
  assign w9006 = w8617 ^ w9005 ;
  assign w9007 = ( ~w7517 & w8994 ) | ( ~w7517 & w9001 ) | ( w8994 & w9001 ) ;
  assign w9008 = ~w8994 & w9007 ;
  assign w9009 = w9006 | w9008 ;
  assign w9010 = ( w7175 & w9003 ) | ( w7175 & ~w9009 ) | ( w9003 & ~w9009 ) ;
  assign w9011 = w7175 & w9010 ;
  assign w9012 = w8620 | w8626 ;
  assign w9013 = w8965 & ~w9012 ;
  assign w9014 = w8624 ^ w9013 ;
  assign w9015 = ( ~w7175 & w9003 ) | ( ~w7175 & w9009 ) | ( w9003 & w9009 ) ;
  assign w9016 = ~w9003 & w9015 ;
  assign w9017 = w9014 | w9016 ;
  assign w9018 = ( w6841 & w9011 ) | ( w6841 & ~w9017 ) | ( w9011 & ~w9017 ) ;
  assign w9019 = w6841 & w9018 ;
  assign w9020 = w8629 | w8634 ;
  assign w9021 = w8965 & ~w9020 ;
  assign w9022 = w8632 ^ w9021 ;
  assign w9023 = ( ~w6841 & w9011 ) | ( ~w6841 & w9017 ) | ( w9011 & w9017 ) ;
  assign w9024 = ~w9011 & w9023 ;
  assign w9025 = w9022 | w9024 ;
  assign w9026 = ( w6515 & w9019 ) | ( w6515 & ~w9025 ) | ( w9019 & ~w9025 ) ;
  assign w9027 = w6515 & w9026 ;
  assign w9028 = w8637 | w8642 ;
  assign w9029 = w8965 & ~w9028 ;
  assign w9030 = w8640 ^ w9029 ;
  assign w9031 = ( ~w6515 & w9019 ) | ( ~w6515 & w9025 ) | ( w9019 & w9025 ) ;
  assign w9032 = ~w9019 & w9031 ;
  assign w9033 = w9030 | w9032 ;
  assign w9034 = ( w6197 & w9027 ) | ( w6197 & ~w9033 ) | ( w9027 & ~w9033 ) ;
  assign w9035 = w6197 & w9034 ;
  assign w9036 = w8645 | w8650 ;
  assign w9037 = w8965 & ~w9036 ;
  assign w9038 = w8648 ^ w9037 ;
  assign w9039 = ( ~w6197 & w9027 ) | ( ~w6197 & w9033 ) | ( w9027 & w9033 ) ;
  assign w9040 = ~w9027 & w9039 ;
  assign w9041 = w9038 | w9040 ;
  assign w9042 = ( w5887 & w9035 ) | ( w5887 & ~w9041 ) | ( w9035 & ~w9041 ) ;
  assign w9043 = w5887 & w9042 ;
  assign w9044 = w8653 | w8658 ;
  assign w9045 = w8965 & ~w9044 ;
  assign w9046 = w8656 ^ w9045 ;
  assign w9047 = ( ~w5887 & w9035 ) | ( ~w5887 & w9041 ) | ( w9035 & w9041 ) ;
  assign w9048 = ~w9035 & w9047 ;
  assign w9049 = w9046 | w9048 ;
  assign w9050 = ( w5585 & w9043 ) | ( w5585 & ~w9049 ) | ( w9043 & ~w9049 ) ;
  assign w9051 = w5585 & w9050 ;
  assign w9052 = w8661 | w8666 ;
  assign w9053 = w8965 & ~w9052 ;
  assign w9054 = w8664 ^ w9053 ;
  assign w9055 = ( ~w5585 & w9043 ) | ( ~w5585 & w9049 ) | ( w9043 & w9049 ) ;
  assign w9056 = ~w9043 & w9055 ;
  assign w9057 = w9054 | w9056 ;
  assign w9058 = ( w5291 & w9051 ) | ( w5291 & ~w9057 ) | ( w9051 & ~w9057 ) ;
  assign w9059 = w5291 & w9058 ;
  assign w9060 = w8669 | w8674 ;
  assign w9061 = w8965 & ~w9060 ;
  assign w9062 = w8672 ^ w9061 ;
  assign w9063 = ( ~w5291 & w9051 ) | ( ~w5291 & w9057 ) | ( w9051 & w9057 ) ;
  assign w9064 = ~w9051 & w9063 ;
  assign w9065 = w9062 | w9064 ;
  assign w9066 = ( w5005 & w9059 ) | ( w5005 & ~w9065 ) | ( w9059 & ~w9065 ) ;
  assign w9067 = w5005 & w9066 ;
  assign w9068 = w8677 | w8682 ;
  assign w9069 = w8965 & ~w9068 ;
  assign w9070 = w8680 ^ w9069 ;
  assign w9071 = ( ~w5005 & w9059 ) | ( ~w5005 & w9065 ) | ( w9059 & w9065 ) ;
  assign w9072 = ~w9059 & w9071 ;
  assign w9073 = w9070 | w9072 ;
  assign w9074 = ( w4727 & w9067 ) | ( w4727 & ~w9073 ) | ( w9067 & ~w9073 ) ;
  assign w9075 = w4727 & w9074 ;
  assign w9076 = w8685 | w8690 ;
  assign w9077 = w8965 & ~w9076 ;
  assign w9078 = w8688 ^ w9077 ;
  assign w9079 = ( ~w4727 & w9067 ) | ( ~w4727 & w9073 ) | ( w9067 & w9073 ) ;
  assign w9080 = ~w9067 & w9079 ;
  assign w9081 = w9078 | w9080 ;
  assign w9082 = ( w4457 & w9075 ) | ( w4457 & ~w9081 ) | ( w9075 & ~w9081 ) ;
  assign w9083 = w4457 & w9082 ;
  assign w9084 = w8693 | w8698 ;
  assign w9085 = w8965 & ~w9084 ;
  assign w9086 = w8696 ^ w9085 ;
  assign w9087 = ( ~w4457 & w9075 ) | ( ~w4457 & w9081 ) | ( w9075 & w9081 ) ;
  assign w9088 = ~w9075 & w9087 ;
  assign w9089 = w9086 | w9088 ;
  assign w9090 = ( w4195 & w9083 ) | ( w4195 & ~w9089 ) | ( w9083 & ~w9089 ) ;
  assign w9091 = w4195 & w9090 ;
  assign w9092 = w8701 | w8706 ;
  assign w9093 = w8965 & ~w9092 ;
  assign w9094 = w8704 ^ w9093 ;
  assign w9095 = ( ~w4195 & w9083 ) | ( ~w4195 & w9089 ) | ( w9083 & w9089 ) ;
  assign w9096 = ~w9083 & w9095 ;
  assign w9097 = w9094 | w9096 ;
  assign w9098 = ( w3941 & w9091 ) | ( w3941 & ~w9097 ) | ( w9091 & ~w9097 ) ;
  assign w9099 = w3941 & w9098 ;
  assign w9100 = w8709 | w8714 ;
  assign w9101 = w8965 & ~w9100 ;
  assign w9102 = w8712 ^ w9101 ;
  assign w9103 = ( ~w3941 & w9091 ) | ( ~w3941 & w9097 ) | ( w9091 & w9097 ) ;
  assign w9104 = ~w9091 & w9103 ;
  assign w9105 = w9102 | w9104 ;
  assign w9106 = ( w3695 & w9099 ) | ( w3695 & ~w9105 ) | ( w9099 & ~w9105 ) ;
  assign w9107 = w3695 & w9106 ;
  assign w9108 = w8717 | w8722 ;
  assign w9109 = w8965 & ~w9108 ;
  assign w9110 = w8720 ^ w9109 ;
  assign w9111 = ( ~w3695 & w9099 ) | ( ~w3695 & w9105 ) | ( w9099 & w9105 ) ;
  assign w9112 = ~w9099 & w9111 ;
  assign w9113 = w9110 | w9112 ;
  assign w9114 = ( w3457 & w9107 ) | ( w3457 & ~w9113 ) | ( w9107 & ~w9113 ) ;
  assign w9115 = w3457 & w9114 ;
  assign w9116 = w8725 | w8730 ;
  assign w9117 = w8965 & ~w9116 ;
  assign w9118 = w8728 ^ w9117 ;
  assign w9119 = ( ~w3457 & w9107 ) | ( ~w3457 & w9113 ) | ( w9107 & w9113 ) ;
  assign w9120 = ~w9107 & w9119 ;
  assign w9121 = w9118 | w9120 ;
  assign w9122 = ( w3227 & w9115 ) | ( w3227 & ~w9121 ) | ( w9115 & ~w9121 ) ;
  assign w9123 = w3227 & w9122 ;
  assign w9124 = w8733 | w8738 ;
  assign w9125 = w8965 & ~w9124 ;
  assign w9126 = w8736 ^ w9125 ;
  assign w9127 = ( ~w3227 & w9115 ) | ( ~w3227 & w9121 ) | ( w9115 & w9121 ) ;
  assign w9128 = ~w9115 & w9127 ;
  assign w9129 = w9126 | w9128 ;
  assign w9130 = ( w3005 & w9123 ) | ( w3005 & ~w9129 ) | ( w9123 & ~w9129 ) ;
  assign w9131 = w3005 & w9130 ;
  assign w9132 = w8741 | w8746 ;
  assign w9133 = w8965 & ~w9132 ;
  assign w9134 = w8744 ^ w9133 ;
  assign w9135 = ( ~w3005 & w9123 ) | ( ~w3005 & w9129 ) | ( w9123 & w9129 ) ;
  assign w9136 = ~w9123 & w9135 ;
  assign w9137 = w9134 | w9136 ;
  assign w9138 = ( w2791 & w9131 ) | ( w2791 & ~w9137 ) | ( w9131 & ~w9137 ) ;
  assign w9139 = w2791 & w9138 ;
  assign w9140 = w8749 | w8754 ;
  assign w9141 = w8965 & ~w9140 ;
  assign w9142 = w8752 ^ w9141 ;
  assign w9143 = ( ~w2791 & w9131 ) | ( ~w2791 & w9137 ) | ( w9131 & w9137 ) ;
  assign w9144 = ~w9131 & w9143 ;
  assign w9145 = w9142 | w9144 ;
  assign w9146 = ( w2585 & w9139 ) | ( w2585 & ~w9145 ) | ( w9139 & ~w9145 ) ;
  assign w9147 = w2585 & w9146 ;
  assign w9148 = w8757 | w8762 ;
  assign w9149 = w8965 & ~w9148 ;
  assign w9150 = w8760 ^ w9149 ;
  assign w9151 = ( ~w2585 & w9139 ) | ( ~w2585 & w9145 ) | ( w9139 & w9145 ) ;
  assign w9152 = ~w9139 & w9151 ;
  assign w9153 = w9150 | w9152 ;
  assign w9154 = ( w2387 & w9147 ) | ( w2387 & ~w9153 ) | ( w9147 & ~w9153 ) ;
  assign w9155 = w2387 & w9154 ;
  assign w9156 = w8765 | w8770 ;
  assign w9157 = w8965 & ~w9156 ;
  assign w9158 = w8768 ^ w9157 ;
  assign w9159 = ( ~w2387 & w9147 ) | ( ~w2387 & w9153 ) | ( w9147 & w9153 ) ;
  assign w9160 = ~w9147 & w9159 ;
  assign w9161 = w9158 | w9160 ;
  assign w9162 = ( w2197 & w9155 ) | ( w2197 & ~w9161 ) | ( w9155 & ~w9161 ) ;
  assign w9163 = w2197 & w9162 ;
  assign w9164 = w8773 | w8778 ;
  assign w9165 = w8965 & ~w9164 ;
  assign w9166 = w8776 ^ w9165 ;
  assign w9167 = ( ~w2197 & w9155 ) | ( ~w2197 & w9161 ) | ( w9155 & w9161 ) ;
  assign w9168 = ~w9155 & w9167 ;
  assign w9169 = w9166 | w9168 ;
  assign w9170 = ( w2015 & w9163 ) | ( w2015 & ~w9169 ) | ( w9163 & ~w9169 ) ;
  assign w9171 = w2015 & w9170 ;
  assign w9172 = w8781 | w8786 ;
  assign w9173 = w8965 & ~w9172 ;
  assign w9174 = w8784 ^ w9173 ;
  assign w9175 = ( ~w2015 & w9163 ) | ( ~w2015 & w9169 ) | ( w9163 & w9169 ) ;
  assign w9176 = ~w9163 & w9175 ;
  assign w9177 = w9174 | w9176 ;
  assign w9178 = ( w1841 & w9171 ) | ( w1841 & ~w9177 ) | ( w9171 & ~w9177 ) ;
  assign w9179 = w1841 & w9178 ;
  assign w9180 = w8789 | w8794 ;
  assign w9181 = w8965 & ~w9180 ;
  assign w9182 = w8792 ^ w9181 ;
  assign w9183 = ( ~w1841 & w9171 ) | ( ~w1841 & w9177 ) | ( w9171 & w9177 ) ;
  assign w9184 = ~w9171 & w9183 ;
  assign w9185 = w9182 | w9184 ;
  assign w9186 = ( w1675 & w9179 ) | ( w1675 & ~w9185 ) | ( w9179 & ~w9185 ) ;
  assign w9187 = w1675 & w9186 ;
  assign w9188 = ( ~w1675 & w9179 ) | ( ~w1675 & w9185 ) | ( w9179 & w9185 ) ;
  assign w9189 = ~w9179 & w9188 ;
  assign w9190 = w8797 | w8799 ;
  assign w9191 = w8965 & ~w9190 ;
  assign w9192 = w8802 ^ w9191 ;
  assign w9193 = w9189 | w9192 ;
  assign w9194 = ( w1517 & w9187 ) | ( w1517 & ~w9193 ) | ( w9187 & ~w9193 ) ;
  assign w9195 = w1517 & w9194 ;
  assign w9196 = w8805 | w8810 ;
  assign w9197 = w8965 & ~w9196 ;
  assign w9198 = w8808 ^ w9197 ;
  assign w9199 = ( ~w1517 & w9187 ) | ( ~w1517 & w9193 ) | ( w9187 & w9193 ) ;
  assign w9200 = ~w9187 & w9199 ;
  assign w9201 = w9198 | w9200 ;
  assign w9202 = ( w1367 & w9195 ) | ( w1367 & ~w9201 ) | ( w9195 & ~w9201 ) ;
  assign w9203 = w1367 & w9202 ;
  assign w9204 = w8813 | w8818 ;
  assign w9205 = w8965 & ~w9204 ;
  assign w9206 = w8816 ^ w9205 ;
  assign w9207 = ( ~w1367 & w9195 ) | ( ~w1367 & w9201 ) | ( w9195 & w9201 ) ;
  assign w9208 = ~w9195 & w9207 ;
  assign w9209 = w9206 | w9208 ;
  assign w9210 = ( w1225 & w9203 ) | ( w1225 & ~w9209 ) | ( w9203 & ~w9209 ) ;
  assign w9211 = w1225 & w9210 ;
  assign w9212 = w8821 | w8826 ;
  assign w9213 = w8965 & ~w9212 ;
  assign w9214 = w8824 ^ w9213 ;
  assign w9215 = ( ~w1225 & w9203 ) | ( ~w1225 & w9209 ) | ( w9203 & w9209 ) ;
  assign w9216 = ~w9203 & w9215 ;
  assign w9217 = w9214 | w9216 ;
  assign w9218 = ( w1091 & w9211 ) | ( w1091 & ~w9217 ) | ( w9211 & ~w9217 ) ;
  assign w9219 = w1091 & w9218 ;
  assign w9220 = w8829 | w8834 ;
  assign w9221 = w8965 & ~w9220 ;
  assign w9222 = w8832 ^ w9221 ;
  assign w9223 = ( ~w1091 & w9211 ) | ( ~w1091 & w9217 ) | ( w9211 & w9217 ) ;
  assign w9224 = ~w9211 & w9223 ;
  assign w9225 = w9222 | w9224 ;
  assign w9226 = ( w965 & w9219 ) | ( w965 & ~w9225 ) | ( w9219 & ~w9225 ) ;
  assign w9227 = w965 & w9226 ;
  assign w9228 = w8837 | w8842 ;
  assign w9229 = w8965 & ~w9228 ;
  assign w9230 = w8840 ^ w9229 ;
  assign w9231 = ( ~w965 & w9219 ) | ( ~w965 & w9225 ) | ( w9219 & w9225 ) ;
  assign w9232 = ~w9219 & w9231 ;
  assign w9233 = w9230 | w9232 ;
  assign w9234 = ( w847 & w9227 ) | ( w847 & ~w9233 ) | ( w9227 & ~w9233 ) ;
  assign w9235 = w847 & w9234 ;
  assign w9236 = w8845 | w8850 ;
  assign w9237 = w8965 & ~w9236 ;
  assign w9238 = w8848 ^ w9237 ;
  assign w9239 = ( ~w847 & w9227 ) | ( ~w847 & w9233 ) | ( w9227 & w9233 ) ;
  assign w9240 = ~w9227 & w9239 ;
  assign w9241 = w9238 | w9240 ;
  assign w9242 = ( w737 & w9235 ) | ( w737 & ~w9241 ) | ( w9235 & ~w9241 ) ;
  assign w9243 = w737 & w9242 ;
  assign w9244 = w8853 | w8858 ;
  assign w9245 = w8965 & ~w9244 ;
  assign w9246 = w8856 ^ w9245 ;
  assign w9247 = ( ~w737 & w9235 ) | ( ~w737 & w9241 ) | ( w9235 & w9241 ) ;
  assign w9248 = ~w9235 & w9247 ;
  assign w9249 = w9246 | w9248 ;
  assign w9250 = ( w635 & w9243 ) | ( w635 & ~w9249 ) | ( w9243 & ~w9249 ) ;
  assign w9251 = w635 & w9250 ;
  assign w9252 = w8861 | w8866 ;
  assign w9253 = w8965 & ~w9252 ;
  assign w9254 = w8864 ^ w9253 ;
  assign w9255 = ( ~w635 & w9243 ) | ( ~w635 & w9249 ) | ( w9243 & w9249 ) ;
  assign w9256 = ~w9243 & w9255 ;
  assign w9257 = w9254 | w9256 ;
  assign w9258 = ( w541 & w9251 ) | ( w541 & ~w9257 ) | ( w9251 & ~w9257 ) ;
  assign w9259 = w541 & w9258 ;
  assign w9260 = w8869 | w8874 ;
  assign w9261 = w8965 & ~w9260 ;
  assign w9262 = w8872 ^ w9261 ;
  assign w9263 = ( ~w541 & w9251 ) | ( ~w541 & w9257 ) | ( w9251 & w9257 ) ;
  assign w9264 = ~w9251 & w9263 ;
  assign w9265 = w9262 | w9264 ;
  assign w9266 = ( w455 & w9259 ) | ( w455 & ~w9265 ) | ( w9259 & ~w9265 ) ;
  assign w9267 = w455 & w9266 ;
  assign w9268 = w8877 | w8882 ;
  assign w9269 = w8965 & ~w9268 ;
  assign w9270 = w8880 ^ w9269 ;
  assign w9271 = ( ~w455 & w9259 ) | ( ~w455 & w9265 ) | ( w9259 & w9265 ) ;
  assign w9272 = ~w9259 & w9271 ;
  assign w9273 = w9270 | w9272 ;
  assign w9274 = ( w377 & w9267 ) | ( w377 & ~w9273 ) | ( w9267 & ~w9273 ) ;
  assign w9275 = w377 & w9274 ;
  assign w9276 = w8885 | w8890 ;
  assign w9277 = w8965 & ~w9276 ;
  assign w9278 = w8888 ^ w9277 ;
  assign w9279 = ( ~w377 & w9267 ) | ( ~w377 & w9273 ) | ( w9267 & w9273 ) ;
  assign w9280 = ~w9267 & w9279 ;
  assign w9281 = w9278 | w9280 ;
  assign w9282 = ( w307 & w9275 ) | ( w307 & ~w9281 ) | ( w9275 & ~w9281 ) ;
  assign w9283 = w307 & w9282 ;
  assign w9284 = w8893 | w8898 ;
  assign w9285 = w8965 & ~w9284 ;
  assign w9286 = w8896 ^ w9285 ;
  assign w9287 = ( ~w307 & w9275 ) | ( ~w307 & w9281 ) | ( w9275 & w9281 ) ;
  assign w9288 = ~w9275 & w9287 ;
  assign w9289 = w9286 | w9288 ;
  assign w9290 = ( w246 & w9283 ) | ( w246 & ~w9289 ) | ( w9283 & ~w9289 ) ;
  assign w9291 = w246 & w9290 ;
  assign w9292 = w8901 | w8906 ;
  assign w9293 = w8965 & ~w9292 ;
  assign w9294 = w8904 ^ w9293 ;
  assign w9295 = ( ~w246 & w9283 ) | ( ~w246 & w9289 ) | ( w9283 & w9289 ) ;
  assign w9296 = ~w9283 & w9295 ;
  assign w9297 = w9294 | w9296 ;
  assign w9298 = ( w185 & w9291 ) | ( w185 & ~w9297 ) | ( w9291 & ~w9297 ) ;
  assign w9299 = w185 & w9298 ;
  assign w9300 = w8909 | w8914 ;
  assign w9301 = w8965 & ~w9300 ;
  assign w9302 = w8912 ^ w9301 ;
  assign w9303 = ( ~w185 & w9291 ) | ( ~w185 & w9297 ) | ( w9291 & w9297 ) ;
  assign w9304 = ~w9291 & w9303 ;
  assign w9305 = w9302 | w9304 ;
  assign w9306 = ( w145 & w9299 ) | ( w145 & ~w9305 ) | ( w9299 & ~w9305 ) ;
  assign w9307 = w145 & w9306 ;
  assign w9308 = w8917 | w8922 ;
  assign w9309 = w8965 & ~w9308 ;
  assign w9310 = w8920 ^ w9309 ;
  assign w9311 = ( ~w145 & w9299 ) | ( ~w145 & w9305 ) | ( w9299 & w9305 ) ;
  assign w9312 = ~w9299 & w9311 ;
  assign w9313 = w9310 | w9312 ;
  assign w9314 = ( w132 & w9307 ) | ( w132 & ~w9313 ) | ( w9307 & ~w9313 ) ;
  assign w9315 = w132 & w9314 ;
  assign w9316 = w8925 | w8930 ;
  assign w9317 = w8965 & ~w9316 ;
  assign w9318 = w8928 ^ w9317 ;
  assign w9319 = ( ~w132 & w9307 ) | ( ~w132 & w9313 ) | ( w9307 & w9313 ) ;
  assign w9320 = ~w9307 & w9319 ;
  assign w9321 = w9318 | w9320 ;
  assign w9322 = ~w9315 & w9321 ;
  assign w9323 = w8933 | w8938 ;
  assign w9324 = w8965 & ~w9323 ;
  assign w9325 = w8936 ^ w9324 ;
  assign w9326 = ( ~w8951 & w9322 ) | ( ~w8951 & w9325 ) | ( w9322 & w9325 ) ;
  assign w9327 = w8940 & ~w9326 ;
  assign w9328 = ~w8943 & w8965 ;
  assign w9329 = ( w9326 & ~w9327 ) | ( w9326 & w9328 ) | ( ~w9327 & w9328 ) ;
  assign w9330 = w8951 | w9329 ;
  assign w9331 = ~w129 & w9330 ;
  assign w9332 = ( w9315 & w9321 ) | ( w9315 & w9325 ) | ( w9321 & w9325 ) ;
  assign w9333 = ~w9315 & w9332 ;
  assign w9334 = ( w129 & w8940 ) | ( w129 & w8943 ) | ( w8940 & w8943 ) ;
  assign w9335 = ( w8943 & ~w8965 ) | ( w8943 & w9334 ) | ( ~w8965 & w9334 ) ;
  assign w9336 = w8940 & w9335 ;
  assign w9337 = w9334 ^ w9336 ;
  assign w9338 = ( w8559 & w8564 ) | ( w8559 & w8591 ) | ( w8564 & w8591 ) ;
  assign w9339 = w8591 & ~w9338 ;
  assign w9340 = w8562 ^ w9339 ;
  assign w9341 = ( ~w8955 & w8962 ) | ( ~w8955 & w9340 ) | ( w8962 & w9340 ) ;
  assign w9342 = ~w8962 & w9341 ;
  assign w9343 = ( ~w8949 & w8951 ) | ( ~w8949 & w9342 ) | ( w8951 & w9342 ) ;
  assign w9344 = ~w8951 & w9343 ;
  assign w9345 = w9333 | w9344 ;
  assign w9346 = ( w9331 & ~w9333 ) | ( w9331 & w9337 ) | ( ~w9333 & w9337 ) ;
  assign w9347 = w9345 | w9346 ;
  assign w9348 = ( ~\pi035 & \pi036 ) | ( ~\pi035 & w8965 ) | ( \pi036 & w8965 ) ;
  assign w9349 = ( ~\pi034 & \pi036 ) | ( ~\pi034 & w9348 ) | ( \pi036 & w9348 ) ;
  assign w9350 = ( ~\pi036 & w8965 ) | ( ~\pi036 & w9347 ) | ( w8965 & w9347 ) ;
  assign w9351 = w9349 & w9350 ;
  assign w9352 = ( w8951 & w8955 ) | ( w8951 & ~w8962 ) | ( w8955 & ~w8962 ) ;
  assign w9353 = \pi035 & ~w9352 ;
  assign w9354 = \pi034 | \pi036 ;
  assign w9355 = ( ~w9352 & w9353 ) | ( ~w9352 & w9354 ) | ( w9353 & w9354 ) ;
  assign w9356 = ~w8962 & w9355 ;
  assign w9357 = ~w8949 & w9356 ;
  assign w9358 = ( \pi036 & w9347 ) | ( \pi036 & ~w9356 ) | ( w9347 & ~w9356 ) ;
  assign w9359 = w9357 & ~w9358 ;
  assign w9360 = ~\pi036 & w9347 ;
  assign w9361 = \pi037 ^ w9360 ;
  assign w9362 = w9359 | w9361 ;
  assign w9363 = ( w8591 & w9351 ) | ( w8591 & ~w9362 ) | ( w9351 & ~w9362 ) ;
  assign w9364 = w8591 & w9363 ;
  assign w9365 = ( ~w8591 & w9351 ) | ( ~w8591 & w9362 ) | ( w9351 & w9362 ) ;
  assign w9366 = ~w9351 & w9365 ;
  assign w9367 = w8965 & ~w9344 ;
  assign w9368 = ~w9333 & w9367 ;
  assign w9369 = ~w9346 & w9368 ;
  assign w9370 = \pi037 & w9347 ;
  assign w9371 = ( \pi036 & w9347 ) | ( \pi036 & ~w9370 ) | ( w9347 & ~w9370 ) ;
  assign w9372 = ( ~\pi036 & w9369 ) | ( ~\pi036 & w9371 ) | ( w9369 & w9371 ) ;
  assign w9373 = \pi038 ^ w9372 ;
  assign w9374 = w9366 | w9373 ;
  assign w9375 = ( w8225 & w9364 ) | ( w8225 & ~w9374 ) | ( w9364 & ~w9374 ) ;
  assign w9376 = w8225 & w9375 ;
  assign w9377 = ( w8969 & ~w8977 ) | ( w8969 & w9347 ) | ( ~w8977 & w9347 ) ;
  assign w9378 = ~w8969 & w9377 ;
  assign w9379 = \pi039 ^ w9378 ;
  assign w9380 = w8978 ^ w9379 ;
  assign w9381 = ( ~w8225 & w9364 ) | ( ~w8225 & w9374 ) | ( w9364 & w9374 ) ;
  assign w9382 = ~w9364 & w9381 ;
  assign w9383 = w9380 | w9382 ;
  assign w9384 = ( w7867 & w9376 ) | ( w7867 & ~w9383 ) | ( w9376 & ~w9383 ) ;
  assign w9385 = w7867 & w9384 ;
  assign w9386 = w8982 | w8984 ;
  assign w9387 = w9347 & ~w9386 ;
  assign w9388 = w8991 ^ w9387 ;
  assign w9389 = ( ~w7867 & w9376 ) | ( ~w7867 & w9383 ) | ( w9376 & w9383 ) ;
  assign w9390 = ~w9376 & w9389 ;
  assign w9391 = w9388 | w9390 ;
  assign w9392 = ( w7517 & w9385 ) | ( w7517 & ~w9391 ) | ( w9385 & ~w9391 ) ;
  assign w9393 = w7517 & w9392 ;
  assign w9394 = w8994 | w9000 ;
  assign w9395 = w9347 & ~w9394 ;
  assign w9396 = w8998 ^ w9395 ;
  assign w9397 = ( ~w7517 & w9385 ) | ( ~w7517 & w9391 ) | ( w9385 & w9391 ) ;
  assign w9398 = ~w9385 & w9397 ;
  assign w9399 = w9396 | w9398 ;
  assign w9400 = ( w7175 & w9393 ) | ( w7175 & ~w9399 ) | ( w9393 & ~w9399 ) ;
  assign w9401 = w7175 & w9400 ;
  assign w9402 = w9003 | w9008 ;
  assign w9403 = w9347 & ~w9402 ;
  assign w9404 = w9006 ^ w9403 ;
  assign w9405 = ( ~w7175 & w9393 ) | ( ~w7175 & w9399 ) | ( w9393 & w9399 ) ;
  assign w9406 = ~w9393 & w9405 ;
  assign w9407 = w9404 | w9406 ;
  assign w9408 = ( w6841 & w9401 ) | ( w6841 & ~w9407 ) | ( w9401 & ~w9407 ) ;
  assign w9409 = w6841 & w9408 ;
  assign w9410 = w9011 | w9016 ;
  assign w9411 = w9347 & ~w9410 ;
  assign w9412 = w9014 ^ w9411 ;
  assign w9413 = ( ~w6841 & w9401 ) | ( ~w6841 & w9407 ) | ( w9401 & w9407 ) ;
  assign w9414 = ~w9401 & w9413 ;
  assign w9415 = w9412 | w9414 ;
  assign w9416 = ( w6515 & w9409 ) | ( w6515 & ~w9415 ) | ( w9409 & ~w9415 ) ;
  assign w9417 = w6515 & w9416 ;
  assign w9418 = w9019 | w9024 ;
  assign w9419 = w9347 & ~w9418 ;
  assign w9420 = w9022 ^ w9419 ;
  assign w9421 = ( ~w6515 & w9409 ) | ( ~w6515 & w9415 ) | ( w9409 & w9415 ) ;
  assign w9422 = ~w9409 & w9421 ;
  assign w9423 = w9420 | w9422 ;
  assign w9424 = ( w6197 & w9417 ) | ( w6197 & ~w9423 ) | ( w9417 & ~w9423 ) ;
  assign w9425 = w6197 & w9424 ;
  assign w9426 = w9027 | w9032 ;
  assign w9427 = w9347 & ~w9426 ;
  assign w9428 = w9030 ^ w9427 ;
  assign w9429 = ( ~w6197 & w9417 ) | ( ~w6197 & w9423 ) | ( w9417 & w9423 ) ;
  assign w9430 = ~w9417 & w9429 ;
  assign w9431 = w9428 | w9430 ;
  assign w9432 = ( w5887 & w9425 ) | ( w5887 & ~w9431 ) | ( w9425 & ~w9431 ) ;
  assign w9433 = w5887 & w9432 ;
  assign w9434 = w9035 | w9040 ;
  assign w9435 = w9347 & ~w9434 ;
  assign w9436 = w9038 ^ w9435 ;
  assign w9437 = ( ~w5887 & w9425 ) | ( ~w5887 & w9431 ) | ( w9425 & w9431 ) ;
  assign w9438 = ~w9425 & w9437 ;
  assign w9439 = w9436 | w9438 ;
  assign w9440 = ( w5585 & w9433 ) | ( w5585 & ~w9439 ) | ( w9433 & ~w9439 ) ;
  assign w9441 = w5585 & w9440 ;
  assign w9442 = w9043 | w9048 ;
  assign w9443 = w9347 & ~w9442 ;
  assign w9444 = w9046 ^ w9443 ;
  assign w9445 = ( ~w5585 & w9433 ) | ( ~w5585 & w9439 ) | ( w9433 & w9439 ) ;
  assign w9446 = ~w9433 & w9445 ;
  assign w9447 = w9444 | w9446 ;
  assign w9448 = ( w5291 & w9441 ) | ( w5291 & ~w9447 ) | ( w9441 & ~w9447 ) ;
  assign w9449 = w5291 & w9448 ;
  assign w9450 = w9051 | w9056 ;
  assign w9451 = w9347 & ~w9450 ;
  assign w9452 = w9054 ^ w9451 ;
  assign w9453 = ( ~w5291 & w9441 ) | ( ~w5291 & w9447 ) | ( w9441 & w9447 ) ;
  assign w9454 = ~w9441 & w9453 ;
  assign w9455 = w9452 | w9454 ;
  assign w9456 = ( w5005 & w9449 ) | ( w5005 & ~w9455 ) | ( w9449 & ~w9455 ) ;
  assign w9457 = w5005 & w9456 ;
  assign w9458 = w9059 | w9064 ;
  assign w9459 = w9347 & ~w9458 ;
  assign w9460 = w9062 ^ w9459 ;
  assign w9461 = ( ~w5005 & w9449 ) | ( ~w5005 & w9455 ) | ( w9449 & w9455 ) ;
  assign w9462 = ~w9449 & w9461 ;
  assign w9463 = w9460 | w9462 ;
  assign w9464 = ( w4727 & w9457 ) | ( w4727 & ~w9463 ) | ( w9457 & ~w9463 ) ;
  assign w9465 = w4727 & w9464 ;
  assign w9466 = w9067 | w9072 ;
  assign w9467 = w9347 & ~w9466 ;
  assign w9468 = w9070 ^ w9467 ;
  assign w9469 = ( ~w4727 & w9457 ) | ( ~w4727 & w9463 ) | ( w9457 & w9463 ) ;
  assign w9470 = ~w9457 & w9469 ;
  assign w9471 = w9468 | w9470 ;
  assign w9472 = ( w4457 & w9465 ) | ( w4457 & ~w9471 ) | ( w9465 & ~w9471 ) ;
  assign w9473 = w4457 & w9472 ;
  assign w9474 = w9075 | w9080 ;
  assign w9475 = w9347 & ~w9474 ;
  assign w9476 = w9078 ^ w9475 ;
  assign w9477 = ( ~w4457 & w9465 ) | ( ~w4457 & w9471 ) | ( w9465 & w9471 ) ;
  assign w9478 = ~w9465 & w9477 ;
  assign w9479 = w9476 | w9478 ;
  assign w9480 = ( w4195 & w9473 ) | ( w4195 & ~w9479 ) | ( w9473 & ~w9479 ) ;
  assign w9481 = w4195 & w9480 ;
  assign w9482 = w9083 | w9088 ;
  assign w9483 = w9347 & ~w9482 ;
  assign w9484 = w9086 ^ w9483 ;
  assign w9485 = ( ~w4195 & w9473 ) | ( ~w4195 & w9479 ) | ( w9473 & w9479 ) ;
  assign w9486 = ~w9473 & w9485 ;
  assign w9487 = w9484 | w9486 ;
  assign w9488 = ( w3941 & w9481 ) | ( w3941 & ~w9487 ) | ( w9481 & ~w9487 ) ;
  assign w9489 = w3941 & w9488 ;
  assign w9490 = w9091 | w9096 ;
  assign w9491 = w9347 & ~w9490 ;
  assign w9492 = w9094 ^ w9491 ;
  assign w9493 = ( ~w3941 & w9481 ) | ( ~w3941 & w9487 ) | ( w9481 & w9487 ) ;
  assign w9494 = ~w9481 & w9493 ;
  assign w9495 = w9492 | w9494 ;
  assign w9496 = ( w3695 & w9489 ) | ( w3695 & ~w9495 ) | ( w9489 & ~w9495 ) ;
  assign w9497 = w3695 & w9496 ;
  assign w9498 = w9099 | w9104 ;
  assign w9499 = w9347 & ~w9498 ;
  assign w9500 = w9102 ^ w9499 ;
  assign w9501 = ( ~w3695 & w9489 ) | ( ~w3695 & w9495 ) | ( w9489 & w9495 ) ;
  assign w9502 = ~w9489 & w9501 ;
  assign w9503 = w9500 | w9502 ;
  assign w9504 = ( w3457 & w9497 ) | ( w3457 & ~w9503 ) | ( w9497 & ~w9503 ) ;
  assign w9505 = w3457 & w9504 ;
  assign w9506 = w9107 | w9112 ;
  assign w9507 = w9347 & ~w9506 ;
  assign w9508 = w9110 ^ w9507 ;
  assign w9509 = ( ~w3457 & w9497 ) | ( ~w3457 & w9503 ) | ( w9497 & w9503 ) ;
  assign w9510 = ~w9497 & w9509 ;
  assign w9511 = w9508 | w9510 ;
  assign w9512 = ( w3227 & w9505 ) | ( w3227 & ~w9511 ) | ( w9505 & ~w9511 ) ;
  assign w9513 = w3227 & w9512 ;
  assign w9514 = w9115 | w9120 ;
  assign w9515 = w9347 & ~w9514 ;
  assign w9516 = w9118 ^ w9515 ;
  assign w9517 = ( ~w3227 & w9505 ) | ( ~w3227 & w9511 ) | ( w9505 & w9511 ) ;
  assign w9518 = ~w9505 & w9517 ;
  assign w9519 = w9516 | w9518 ;
  assign w9520 = ( w3005 & w9513 ) | ( w3005 & ~w9519 ) | ( w9513 & ~w9519 ) ;
  assign w9521 = w3005 & w9520 ;
  assign w9522 = w9123 | w9128 ;
  assign w9523 = w9347 & ~w9522 ;
  assign w9524 = w9126 ^ w9523 ;
  assign w9525 = ( ~w3005 & w9513 ) | ( ~w3005 & w9519 ) | ( w9513 & w9519 ) ;
  assign w9526 = ~w9513 & w9525 ;
  assign w9527 = w9524 | w9526 ;
  assign w9528 = ( w2791 & w9521 ) | ( w2791 & ~w9527 ) | ( w9521 & ~w9527 ) ;
  assign w9529 = w2791 & w9528 ;
  assign w9530 = w9131 | w9136 ;
  assign w9531 = w9347 & ~w9530 ;
  assign w9532 = w9134 ^ w9531 ;
  assign w9533 = ( ~w2791 & w9521 ) | ( ~w2791 & w9527 ) | ( w9521 & w9527 ) ;
  assign w9534 = ~w9521 & w9533 ;
  assign w9535 = w9532 | w9534 ;
  assign w9536 = ( w2585 & w9529 ) | ( w2585 & ~w9535 ) | ( w9529 & ~w9535 ) ;
  assign w9537 = w2585 & w9536 ;
  assign w9538 = w9139 | w9144 ;
  assign w9539 = w9347 & ~w9538 ;
  assign w9540 = w9142 ^ w9539 ;
  assign w9541 = ( ~w2585 & w9529 ) | ( ~w2585 & w9535 ) | ( w9529 & w9535 ) ;
  assign w9542 = ~w9529 & w9541 ;
  assign w9543 = w9540 | w9542 ;
  assign w9544 = ( w2387 & w9537 ) | ( w2387 & ~w9543 ) | ( w9537 & ~w9543 ) ;
  assign w9545 = w2387 & w9544 ;
  assign w9546 = w9147 | w9152 ;
  assign w9547 = w9347 & ~w9546 ;
  assign w9548 = w9150 ^ w9547 ;
  assign w9549 = ( ~w2387 & w9537 ) | ( ~w2387 & w9543 ) | ( w9537 & w9543 ) ;
  assign w9550 = ~w9537 & w9549 ;
  assign w9551 = w9548 | w9550 ;
  assign w9552 = ( w2197 & w9545 ) | ( w2197 & ~w9551 ) | ( w9545 & ~w9551 ) ;
  assign w9553 = w2197 & w9552 ;
  assign w9554 = w9155 | w9160 ;
  assign w9555 = w9347 & ~w9554 ;
  assign w9556 = w9158 ^ w9555 ;
  assign w9557 = ( ~w2197 & w9545 ) | ( ~w2197 & w9551 ) | ( w9545 & w9551 ) ;
  assign w9558 = ~w9545 & w9557 ;
  assign w9559 = w9556 | w9558 ;
  assign w9560 = ( w2015 & w9553 ) | ( w2015 & ~w9559 ) | ( w9553 & ~w9559 ) ;
  assign w9561 = w2015 & w9560 ;
  assign w9562 = w9163 | w9168 ;
  assign w9563 = w9347 & ~w9562 ;
  assign w9564 = w9166 ^ w9563 ;
  assign w9565 = ( ~w2015 & w9553 ) | ( ~w2015 & w9559 ) | ( w9553 & w9559 ) ;
  assign w9566 = ~w9553 & w9565 ;
  assign w9567 = w9564 | w9566 ;
  assign w9568 = ( w1841 & w9561 ) | ( w1841 & ~w9567 ) | ( w9561 & ~w9567 ) ;
  assign w9569 = w1841 & w9568 ;
  assign w9570 = w9171 | w9176 ;
  assign w9571 = w9347 & ~w9570 ;
  assign w9572 = w9174 ^ w9571 ;
  assign w9573 = ( ~w1841 & w9561 ) | ( ~w1841 & w9567 ) | ( w9561 & w9567 ) ;
  assign w9574 = ~w9561 & w9573 ;
  assign w9575 = w9572 | w9574 ;
  assign w9576 = ( w1675 & w9569 ) | ( w1675 & ~w9575 ) | ( w9569 & ~w9575 ) ;
  assign w9577 = w1675 & w9576 ;
  assign w9578 = w9179 | w9184 ;
  assign w9579 = w9347 & ~w9578 ;
  assign w9580 = w9182 ^ w9579 ;
  assign w9581 = ( ~w1675 & w9569 ) | ( ~w1675 & w9575 ) | ( w9569 & w9575 ) ;
  assign w9582 = ~w9569 & w9581 ;
  assign w9583 = w9580 | w9582 ;
  assign w9584 = ( w1517 & w9577 ) | ( w1517 & ~w9583 ) | ( w9577 & ~w9583 ) ;
  assign w9585 = w1517 & w9584 ;
  assign w9586 = ( ~w1517 & w9577 ) | ( ~w1517 & w9583 ) | ( w9577 & w9583 ) ;
  assign w9587 = ~w9577 & w9586 ;
  assign w9588 = w9187 | w9189 ;
  assign w9589 = w9347 & ~w9588 ;
  assign w9590 = w9192 ^ w9589 ;
  assign w9591 = w9587 | w9590 ;
  assign w9592 = ( w1367 & w9585 ) | ( w1367 & ~w9591 ) | ( w9585 & ~w9591 ) ;
  assign w9593 = w1367 & w9592 ;
  assign w9594 = w9195 | w9200 ;
  assign w9595 = w9347 & ~w9594 ;
  assign w9596 = w9198 ^ w9595 ;
  assign w9597 = ( ~w1367 & w9585 ) | ( ~w1367 & w9591 ) | ( w9585 & w9591 ) ;
  assign w9598 = ~w9585 & w9597 ;
  assign w9599 = w9596 | w9598 ;
  assign w9600 = ( w1225 & w9593 ) | ( w1225 & ~w9599 ) | ( w9593 & ~w9599 ) ;
  assign w9601 = w1225 & w9600 ;
  assign w9602 = w9203 | w9208 ;
  assign w9603 = w9347 & ~w9602 ;
  assign w9604 = w9206 ^ w9603 ;
  assign w9605 = ( ~w1225 & w9593 ) | ( ~w1225 & w9599 ) | ( w9593 & w9599 ) ;
  assign w9606 = ~w9593 & w9605 ;
  assign w9607 = w9604 | w9606 ;
  assign w9608 = ( w1091 & w9601 ) | ( w1091 & ~w9607 ) | ( w9601 & ~w9607 ) ;
  assign w9609 = w1091 & w9608 ;
  assign w9610 = w9211 | w9216 ;
  assign w9611 = w9347 & ~w9610 ;
  assign w9612 = w9214 ^ w9611 ;
  assign w9613 = ( ~w1091 & w9601 ) | ( ~w1091 & w9607 ) | ( w9601 & w9607 ) ;
  assign w9614 = ~w9601 & w9613 ;
  assign w9615 = w9612 | w9614 ;
  assign w9616 = ( w965 & w9609 ) | ( w965 & ~w9615 ) | ( w9609 & ~w9615 ) ;
  assign w9617 = w965 & w9616 ;
  assign w9618 = w9219 | w9224 ;
  assign w9619 = w9347 & ~w9618 ;
  assign w9620 = w9222 ^ w9619 ;
  assign w9621 = ( ~w965 & w9609 ) | ( ~w965 & w9615 ) | ( w9609 & w9615 ) ;
  assign w9622 = ~w9609 & w9621 ;
  assign w9623 = w9620 | w9622 ;
  assign w9624 = ( w847 & w9617 ) | ( w847 & ~w9623 ) | ( w9617 & ~w9623 ) ;
  assign w9625 = w847 & w9624 ;
  assign w9626 = w9227 | w9232 ;
  assign w9627 = w9347 & ~w9626 ;
  assign w9628 = w9230 ^ w9627 ;
  assign w9629 = ( ~w847 & w9617 ) | ( ~w847 & w9623 ) | ( w9617 & w9623 ) ;
  assign w9630 = ~w9617 & w9629 ;
  assign w9631 = w9628 | w9630 ;
  assign w9632 = ( w737 & w9625 ) | ( w737 & ~w9631 ) | ( w9625 & ~w9631 ) ;
  assign w9633 = w737 & w9632 ;
  assign w9634 = w9235 | w9240 ;
  assign w9635 = w9347 & ~w9634 ;
  assign w9636 = w9238 ^ w9635 ;
  assign w9637 = ( ~w737 & w9625 ) | ( ~w737 & w9631 ) | ( w9625 & w9631 ) ;
  assign w9638 = ~w9625 & w9637 ;
  assign w9639 = w9636 | w9638 ;
  assign w9640 = ( w635 & w9633 ) | ( w635 & ~w9639 ) | ( w9633 & ~w9639 ) ;
  assign w9641 = w635 & w9640 ;
  assign w9642 = w9243 | w9248 ;
  assign w9643 = w9347 & ~w9642 ;
  assign w9644 = w9246 ^ w9643 ;
  assign w9645 = ( ~w635 & w9633 ) | ( ~w635 & w9639 ) | ( w9633 & w9639 ) ;
  assign w9646 = ~w9633 & w9645 ;
  assign w9647 = w9644 | w9646 ;
  assign w9648 = ( w541 & w9641 ) | ( w541 & ~w9647 ) | ( w9641 & ~w9647 ) ;
  assign w9649 = w541 & w9648 ;
  assign w9650 = w9251 | w9256 ;
  assign w9651 = w9347 & ~w9650 ;
  assign w9652 = w9254 ^ w9651 ;
  assign w9653 = ( ~w541 & w9641 ) | ( ~w541 & w9647 ) | ( w9641 & w9647 ) ;
  assign w9654 = ~w9641 & w9653 ;
  assign w9655 = w9652 | w9654 ;
  assign w9656 = ( w455 & w9649 ) | ( w455 & ~w9655 ) | ( w9649 & ~w9655 ) ;
  assign w9657 = w455 & w9656 ;
  assign w9658 = w9259 | w9264 ;
  assign w9659 = w9347 & ~w9658 ;
  assign w9660 = w9262 ^ w9659 ;
  assign w9661 = ( ~w455 & w9649 ) | ( ~w455 & w9655 ) | ( w9649 & w9655 ) ;
  assign w9662 = ~w9649 & w9661 ;
  assign w9663 = w9660 | w9662 ;
  assign w9664 = ( w377 & w9657 ) | ( w377 & ~w9663 ) | ( w9657 & ~w9663 ) ;
  assign w9665 = w377 & w9664 ;
  assign w9666 = w9267 | w9272 ;
  assign w9667 = w9347 & ~w9666 ;
  assign w9668 = w9270 ^ w9667 ;
  assign w9669 = ( ~w377 & w9657 ) | ( ~w377 & w9663 ) | ( w9657 & w9663 ) ;
  assign w9670 = ~w9657 & w9669 ;
  assign w9671 = w9668 | w9670 ;
  assign w9672 = ( w307 & w9665 ) | ( w307 & ~w9671 ) | ( w9665 & ~w9671 ) ;
  assign w9673 = w307 & w9672 ;
  assign w9674 = w9275 | w9280 ;
  assign w9675 = w9347 & ~w9674 ;
  assign w9676 = w9278 ^ w9675 ;
  assign w9677 = ( ~w307 & w9665 ) | ( ~w307 & w9671 ) | ( w9665 & w9671 ) ;
  assign w9678 = ~w9665 & w9677 ;
  assign w9679 = w9676 | w9678 ;
  assign w9680 = ( w246 & w9673 ) | ( w246 & ~w9679 ) | ( w9673 & ~w9679 ) ;
  assign w9681 = w246 & w9680 ;
  assign w9682 = w9283 | w9288 ;
  assign w9683 = w9347 & ~w9682 ;
  assign w9684 = w9286 ^ w9683 ;
  assign w9685 = ( ~w246 & w9673 ) | ( ~w246 & w9679 ) | ( w9673 & w9679 ) ;
  assign w9686 = ~w9673 & w9685 ;
  assign w9687 = w9684 | w9686 ;
  assign w9688 = ( w185 & w9681 ) | ( w185 & ~w9687 ) | ( w9681 & ~w9687 ) ;
  assign w9689 = w185 & w9688 ;
  assign w9690 = w9291 | w9296 ;
  assign w9691 = w9347 & ~w9690 ;
  assign w9692 = w9294 ^ w9691 ;
  assign w9693 = ( ~w185 & w9681 ) | ( ~w185 & w9687 ) | ( w9681 & w9687 ) ;
  assign w9694 = ~w9681 & w9693 ;
  assign w9695 = w9692 | w9694 ;
  assign w9696 = ( w145 & w9689 ) | ( w145 & ~w9695 ) | ( w9689 & ~w9695 ) ;
  assign w9697 = w145 & w9696 ;
  assign w9698 = w9299 | w9304 ;
  assign w9699 = w9347 & ~w9698 ;
  assign w9700 = w9302 ^ w9699 ;
  assign w9701 = ( ~w145 & w9689 ) | ( ~w145 & w9695 ) | ( w9689 & w9695 ) ;
  assign w9702 = ~w9689 & w9701 ;
  assign w9703 = w9700 | w9702 ;
  assign w9704 = ( w132 & w9697 ) | ( w132 & ~w9703 ) | ( w9697 & ~w9703 ) ;
  assign w9705 = w132 & w9704 ;
  assign w9706 = w9307 | w9312 ;
  assign w9707 = w9347 & ~w9706 ;
  assign w9708 = w9310 ^ w9707 ;
  assign w9709 = ( ~w132 & w9697 ) | ( ~w132 & w9703 ) | ( w9697 & w9703 ) ;
  assign w9710 = ~w9697 & w9709 ;
  assign w9711 = w9708 | w9710 ;
  assign w9712 = ~w9705 & w9711 ;
  assign w9713 = w9315 | w9320 ;
  assign w9714 = w9347 & ~w9713 ;
  assign w9715 = w9318 ^ w9714 ;
  assign w9716 = ( ~w9333 & w9712 ) | ( ~w9333 & w9715 ) | ( w9712 & w9715 ) ;
  assign w9717 = w9322 & ~w9716 ;
  assign w9718 = ~w9325 & w9347 ;
  assign w9719 = ( w9716 & ~w9717 ) | ( w9716 & w9718 ) | ( ~w9717 & w9718 ) ;
  assign w9720 = w9333 | w9719 ;
  assign w9721 = ~w129 & w9720 ;
  assign w9722 = ( w9705 & w9711 ) | ( w9705 & w9715 ) | ( w9711 & w9715 ) ;
  assign w9723 = ~w9705 & w9722 ;
  assign w9724 = ( w129 & w9322 ) | ( w129 & w9325 ) | ( w9322 & w9325 ) ;
  assign w9725 = ( w9325 & ~w9347 ) | ( w9325 & w9724 ) | ( ~w9347 & w9724 ) ;
  assign w9726 = w9322 & w9725 ;
  assign w9727 = w9724 ^ w9726 ;
  assign w9728 = ( w8933 & w8938 ) | ( w8933 & w8965 ) | ( w8938 & w8965 ) ;
  assign w9729 = w8965 & ~w9728 ;
  assign w9730 = w8936 ^ w9729 ;
  assign w9731 = ( ~w9337 & w9344 ) | ( ~w9337 & w9730 ) | ( w9344 & w9730 ) ;
  assign w9732 = ~w9344 & w9731 ;
  assign w9733 = ( ~w9331 & w9333 ) | ( ~w9331 & w9732 ) | ( w9333 & w9732 ) ;
  assign w9734 = ~w9333 & w9733 ;
  assign w9735 = w9723 | w9734 ;
  assign w9736 = ( w9721 & ~w9723 ) | ( w9721 & w9727 ) | ( ~w9723 & w9727 ) ;
  assign w9737 = w9735 | w9736 ;
  assign w9738 = ( ~\pi033 & \pi034 ) | ( ~\pi033 & w9347 ) | ( \pi034 & w9347 ) ;
  assign w9739 = ( ~\pi032 & \pi034 ) | ( ~\pi032 & w9738 ) | ( \pi034 & w9738 ) ;
  assign w9740 = ( ~\pi034 & w9347 ) | ( ~\pi034 & w9737 ) | ( w9347 & w9737 ) ;
  assign w9741 = w9739 & w9740 ;
  assign w9742 = ( w9333 & w9337 ) | ( w9333 & ~w9344 ) | ( w9337 & ~w9344 ) ;
  assign w9743 = \pi033 & ~w9742 ;
  assign w9744 = \pi032 | \pi034 ;
  assign w9745 = ( ~w9742 & w9743 ) | ( ~w9742 & w9744 ) | ( w9743 & w9744 ) ;
  assign w9746 = ~w9344 & w9745 ;
  assign w9747 = ~w9331 & w9746 ;
  assign w9748 = ( \pi034 & w9737 ) | ( \pi034 & ~w9746 ) | ( w9737 & ~w9746 ) ;
  assign w9749 = w9747 & ~w9748 ;
  assign w9750 = ~\pi034 & w9737 ;
  assign w9751 = \pi035 ^ w9750 ;
  assign w9752 = w9749 | w9751 ;
  assign w9753 = ( w8965 & w9741 ) | ( w8965 & ~w9752 ) | ( w9741 & ~w9752 ) ;
  assign w9754 = w8965 & w9753 ;
  assign w9755 = ( ~w8965 & w9741 ) | ( ~w8965 & w9752 ) | ( w9741 & w9752 ) ;
  assign w9756 = ~w9741 & w9755 ;
  assign w9757 = w9347 & ~w9734 ;
  assign w9758 = ~w9723 & w9757 ;
  assign w9759 = ~w9736 & w9758 ;
  assign w9760 = \pi035 & w9737 ;
  assign w9761 = ( \pi034 & w9737 ) | ( \pi034 & ~w9760 ) | ( w9737 & ~w9760 ) ;
  assign w9762 = ( ~\pi034 & w9759 ) | ( ~\pi034 & w9761 ) | ( w9759 & w9761 ) ;
  assign w9763 = \pi036 ^ w9762 ;
  assign w9764 = w9756 | w9763 ;
  assign w9765 = ( w8591 & w9754 ) | ( w8591 & ~w9764 ) | ( w9754 & ~w9764 ) ;
  assign w9766 = w8591 & w9765 ;
  assign w9767 = ( w9351 & ~w9359 ) | ( w9351 & w9737 ) | ( ~w9359 & w9737 ) ;
  assign w9768 = ~w9351 & w9767 ;
  assign w9769 = \pi037 ^ w9768 ;
  assign w9770 = w9360 ^ w9769 ;
  assign w9771 = ( ~w8591 & w9754 ) | ( ~w8591 & w9764 ) | ( w9754 & w9764 ) ;
  assign w9772 = ~w9754 & w9771 ;
  assign w9773 = w9770 | w9772 ;
  assign w9774 = ( w8225 & w9766 ) | ( w8225 & ~w9773 ) | ( w9766 & ~w9773 ) ;
  assign w9775 = w8225 & w9774 ;
  assign w9776 = w9364 | w9366 ;
  assign w9777 = w9737 & ~w9776 ;
  assign w9778 = w9373 ^ w9777 ;
  assign w9779 = ( ~w8225 & w9766 ) | ( ~w8225 & w9773 ) | ( w9766 & w9773 ) ;
  assign w9780 = ~w9766 & w9779 ;
  assign w9781 = w9778 | w9780 ;
  assign w9782 = ( w7867 & w9775 ) | ( w7867 & ~w9781 ) | ( w9775 & ~w9781 ) ;
  assign w9783 = w7867 & w9782 ;
  assign w9784 = w9376 | w9382 ;
  assign w9785 = w9737 & ~w9784 ;
  assign w9786 = w9380 ^ w9785 ;
  assign w9787 = ( ~w7867 & w9775 ) | ( ~w7867 & w9781 ) | ( w9775 & w9781 ) ;
  assign w9788 = ~w9775 & w9787 ;
  assign w9789 = w9786 | w9788 ;
  assign w9790 = ( w7517 & w9783 ) | ( w7517 & ~w9789 ) | ( w9783 & ~w9789 ) ;
  assign w9791 = w7517 & w9790 ;
  assign w9792 = w9385 | w9390 ;
  assign w9793 = w9737 & ~w9792 ;
  assign w9794 = w9388 ^ w9793 ;
  assign w9795 = ( ~w7517 & w9783 ) | ( ~w7517 & w9789 ) | ( w9783 & w9789 ) ;
  assign w9796 = ~w9783 & w9795 ;
  assign w9797 = w9794 | w9796 ;
  assign w9798 = ( w7175 & w9791 ) | ( w7175 & ~w9797 ) | ( w9791 & ~w9797 ) ;
  assign w9799 = w7175 & w9798 ;
  assign w9800 = w9393 | w9398 ;
  assign w9801 = w9737 & ~w9800 ;
  assign w9802 = w9396 ^ w9801 ;
  assign w9803 = ( ~w7175 & w9791 ) | ( ~w7175 & w9797 ) | ( w9791 & w9797 ) ;
  assign w9804 = ~w9791 & w9803 ;
  assign w9805 = w9802 | w9804 ;
  assign w9806 = ( w6841 & w9799 ) | ( w6841 & ~w9805 ) | ( w9799 & ~w9805 ) ;
  assign w9807 = w6841 & w9806 ;
  assign w9808 = w9401 | w9406 ;
  assign w9809 = w9737 & ~w9808 ;
  assign w9810 = w9404 ^ w9809 ;
  assign w9811 = ( ~w6841 & w9799 ) | ( ~w6841 & w9805 ) | ( w9799 & w9805 ) ;
  assign w9812 = ~w9799 & w9811 ;
  assign w9813 = w9810 | w9812 ;
  assign w9814 = ( w6515 & w9807 ) | ( w6515 & ~w9813 ) | ( w9807 & ~w9813 ) ;
  assign w9815 = w6515 & w9814 ;
  assign w9816 = w9409 | w9414 ;
  assign w9817 = w9737 & ~w9816 ;
  assign w9818 = w9412 ^ w9817 ;
  assign w9819 = ( ~w6515 & w9807 ) | ( ~w6515 & w9813 ) | ( w9807 & w9813 ) ;
  assign w9820 = ~w9807 & w9819 ;
  assign w9821 = w9818 | w9820 ;
  assign w9822 = ( w6197 & w9815 ) | ( w6197 & ~w9821 ) | ( w9815 & ~w9821 ) ;
  assign w9823 = w6197 & w9822 ;
  assign w9824 = w9417 | w9422 ;
  assign w9825 = w9737 & ~w9824 ;
  assign w9826 = w9420 ^ w9825 ;
  assign w9827 = ( ~w6197 & w9815 ) | ( ~w6197 & w9821 ) | ( w9815 & w9821 ) ;
  assign w9828 = ~w9815 & w9827 ;
  assign w9829 = w9826 | w9828 ;
  assign w9830 = ( w5887 & w9823 ) | ( w5887 & ~w9829 ) | ( w9823 & ~w9829 ) ;
  assign w9831 = w5887 & w9830 ;
  assign w9832 = w9425 | w9430 ;
  assign w9833 = w9737 & ~w9832 ;
  assign w9834 = w9428 ^ w9833 ;
  assign w9835 = ( ~w5887 & w9823 ) | ( ~w5887 & w9829 ) | ( w9823 & w9829 ) ;
  assign w9836 = ~w9823 & w9835 ;
  assign w9837 = w9834 | w9836 ;
  assign w9838 = ( w5585 & w9831 ) | ( w5585 & ~w9837 ) | ( w9831 & ~w9837 ) ;
  assign w9839 = w5585 & w9838 ;
  assign w9840 = w9433 | w9438 ;
  assign w9841 = w9737 & ~w9840 ;
  assign w9842 = w9436 ^ w9841 ;
  assign w9843 = ( ~w5585 & w9831 ) | ( ~w5585 & w9837 ) | ( w9831 & w9837 ) ;
  assign w9844 = ~w9831 & w9843 ;
  assign w9845 = w9842 | w9844 ;
  assign w9846 = ( w5291 & w9839 ) | ( w5291 & ~w9845 ) | ( w9839 & ~w9845 ) ;
  assign w9847 = w5291 & w9846 ;
  assign w9848 = w9441 | w9446 ;
  assign w9849 = w9737 & ~w9848 ;
  assign w9850 = w9444 ^ w9849 ;
  assign w9851 = ( ~w5291 & w9839 ) | ( ~w5291 & w9845 ) | ( w9839 & w9845 ) ;
  assign w9852 = ~w9839 & w9851 ;
  assign w9853 = w9850 | w9852 ;
  assign w9854 = ( w5005 & w9847 ) | ( w5005 & ~w9853 ) | ( w9847 & ~w9853 ) ;
  assign w9855 = w5005 & w9854 ;
  assign w9856 = w9449 | w9454 ;
  assign w9857 = w9737 & ~w9856 ;
  assign w9858 = w9452 ^ w9857 ;
  assign w9859 = ( ~w5005 & w9847 ) | ( ~w5005 & w9853 ) | ( w9847 & w9853 ) ;
  assign w9860 = ~w9847 & w9859 ;
  assign w9861 = w9858 | w9860 ;
  assign w9862 = ( w4727 & w9855 ) | ( w4727 & ~w9861 ) | ( w9855 & ~w9861 ) ;
  assign w9863 = w4727 & w9862 ;
  assign w9864 = w9457 | w9462 ;
  assign w9865 = w9737 & ~w9864 ;
  assign w9866 = w9460 ^ w9865 ;
  assign w9867 = ( ~w4727 & w9855 ) | ( ~w4727 & w9861 ) | ( w9855 & w9861 ) ;
  assign w9868 = ~w9855 & w9867 ;
  assign w9869 = w9866 | w9868 ;
  assign w9870 = ( w4457 & w9863 ) | ( w4457 & ~w9869 ) | ( w9863 & ~w9869 ) ;
  assign w9871 = w4457 & w9870 ;
  assign w9872 = w9465 | w9470 ;
  assign w9873 = w9737 & ~w9872 ;
  assign w9874 = w9468 ^ w9873 ;
  assign w9875 = ( ~w4457 & w9863 ) | ( ~w4457 & w9869 ) | ( w9863 & w9869 ) ;
  assign w9876 = ~w9863 & w9875 ;
  assign w9877 = w9874 | w9876 ;
  assign w9878 = ( w4195 & w9871 ) | ( w4195 & ~w9877 ) | ( w9871 & ~w9877 ) ;
  assign w9879 = w4195 & w9878 ;
  assign w9880 = w9473 | w9478 ;
  assign w9881 = w9737 & ~w9880 ;
  assign w9882 = w9476 ^ w9881 ;
  assign w9883 = ( ~w4195 & w9871 ) | ( ~w4195 & w9877 ) | ( w9871 & w9877 ) ;
  assign w9884 = ~w9871 & w9883 ;
  assign w9885 = w9882 | w9884 ;
  assign w9886 = ( w3941 & w9879 ) | ( w3941 & ~w9885 ) | ( w9879 & ~w9885 ) ;
  assign w9887 = w3941 & w9886 ;
  assign w9888 = w9481 | w9486 ;
  assign w9889 = w9737 & ~w9888 ;
  assign w9890 = w9484 ^ w9889 ;
  assign w9891 = ( ~w3941 & w9879 ) | ( ~w3941 & w9885 ) | ( w9879 & w9885 ) ;
  assign w9892 = ~w9879 & w9891 ;
  assign w9893 = w9890 | w9892 ;
  assign w9894 = ( w3695 & w9887 ) | ( w3695 & ~w9893 ) | ( w9887 & ~w9893 ) ;
  assign w9895 = w3695 & w9894 ;
  assign w9896 = w9489 | w9494 ;
  assign w9897 = w9737 & ~w9896 ;
  assign w9898 = w9492 ^ w9897 ;
  assign w9899 = ( ~w3695 & w9887 ) | ( ~w3695 & w9893 ) | ( w9887 & w9893 ) ;
  assign w9900 = ~w9887 & w9899 ;
  assign w9901 = w9898 | w9900 ;
  assign w9902 = ( w3457 & w9895 ) | ( w3457 & ~w9901 ) | ( w9895 & ~w9901 ) ;
  assign w9903 = w3457 & w9902 ;
  assign w9904 = w9497 | w9502 ;
  assign w9905 = w9737 & ~w9904 ;
  assign w9906 = w9500 ^ w9905 ;
  assign w9907 = ( ~w3457 & w9895 ) | ( ~w3457 & w9901 ) | ( w9895 & w9901 ) ;
  assign w9908 = ~w9895 & w9907 ;
  assign w9909 = w9906 | w9908 ;
  assign w9910 = ( w3227 & w9903 ) | ( w3227 & ~w9909 ) | ( w9903 & ~w9909 ) ;
  assign w9911 = w3227 & w9910 ;
  assign w9912 = w9505 | w9510 ;
  assign w9913 = w9737 & ~w9912 ;
  assign w9914 = w9508 ^ w9913 ;
  assign w9915 = ( ~w3227 & w9903 ) | ( ~w3227 & w9909 ) | ( w9903 & w9909 ) ;
  assign w9916 = ~w9903 & w9915 ;
  assign w9917 = w9914 | w9916 ;
  assign w9918 = ( w3005 & w9911 ) | ( w3005 & ~w9917 ) | ( w9911 & ~w9917 ) ;
  assign w9919 = w3005 & w9918 ;
  assign w9920 = w9513 | w9518 ;
  assign w9921 = w9737 & ~w9920 ;
  assign w9922 = w9516 ^ w9921 ;
  assign w9923 = ( ~w3005 & w9911 ) | ( ~w3005 & w9917 ) | ( w9911 & w9917 ) ;
  assign w9924 = ~w9911 & w9923 ;
  assign w9925 = w9922 | w9924 ;
  assign w9926 = ( w2791 & w9919 ) | ( w2791 & ~w9925 ) | ( w9919 & ~w9925 ) ;
  assign w9927 = w2791 & w9926 ;
  assign w9928 = w9521 | w9526 ;
  assign w9929 = w9737 & ~w9928 ;
  assign w9930 = w9524 ^ w9929 ;
  assign w9931 = ( ~w2791 & w9919 ) | ( ~w2791 & w9925 ) | ( w9919 & w9925 ) ;
  assign w9932 = ~w9919 & w9931 ;
  assign w9933 = w9930 | w9932 ;
  assign w9934 = ( w2585 & w9927 ) | ( w2585 & ~w9933 ) | ( w9927 & ~w9933 ) ;
  assign w9935 = w2585 & w9934 ;
  assign w9936 = w9529 | w9534 ;
  assign w9937 = w9737 & ~w9936 ;
  assign w9938 = w9532 ^ w9937 ;
  assign w9939 = ( ~w2585 & w9927 ) | ( ~w2585 & w9933 ) | ( w9927 & w9933 ) ;
  assign w9940 = ~w9927 & w9939 ;
  assign w9941 = w9938 | w9940 ;
  assign w9942 = ( w2387 & w9935 ) | ( w2387 & ~w9941 ) | ( w9935 & ~w9941 ) ;
  assign w9943 = w2387 & w9942 ;
  assign w9944 = w9537 | w9542 ;
  assign w9945 = w9737 & ~w9944 ;
  assign w9946 = w9540 ^ w9945 ;
  assign w9947 = ( ~w2387 & w9935 ) | ( ~w2387 & w9941 ) | ( w9935 & w9941 ) ;
  assign w9948 = ~w9935 & w9947 ;
  assign w9949 = w9946 | w9948 ;
  assign w9950 = ( w2197 & w9943 ) | ( w2197 & ~w9949 ) | ( w9943 & ~w9949 ) ;
  assign w9951 = w2197 & w9950 ;
  assign w9952 = w9545 | w9550 ;
  assign w9953 = w9737 & ~w9952 ;
  assign w9954 = w9548 ^ w9953 ;
  assign w9955 = ( ~w2197 & w9943 ) | ( ~w2197 & w9949 ) | ( w9943 & w9949 ) ;
  assign w9956 = ~w9943 & w9955 ;
  assign w9957 = w9954 | w9956 ;
  assign w9958 = ( w2015 & w9951 ) | ( w2015 & ~w9957 ) | ( w9951 & ~w9957 ) ;
  assign w9959 = w2015 & w9958 ;
  assign w9960 = w9553 | w9558 ;
  assign w9961 = w9737 & ~w9960 ;
  assign w9962 = w9556 ^ w9961 ;
  assign w9963 = ( ~w2015 & w9951 ) | ( ~w2015 & w9957 ) | ( w9951 & w9957 ) ;
  assign w9964 = ~w9951 & w9963 ;
  assign w9965 = w9962 | w9964 ;
  assign w9966 = ( w1841 & w9959 ) | ( w1841 & ~w9965 ) | ( w9959 & ~w9965 ) ;
  assign w9967 = w1841 & w9966 ;
  assign w9968 = w9561 | w9566 ;
  assign w9969 = w9737 & ~w9968 ;
  assign w9970 = w9564 ^ w9969 ;
  assign w9971 = ( ~w1841 & w9959 ) | ( ~w1841 & w9965 ) | ( w9959 & w9965 ) ;
  assign w9972 = ~w9959 & w9971 ;
  assign w9973 = w9970 | w9972 ;
  assign w9974 = ( w1675 & w9967 ) | ( w1675 & ~w9973 ) | ( w9967 & ~w9973 ) ;
  assign w9975 = w1675 & w9974 ;
  assign w9976 = w9569 | w9574 ;
  assign w9977 = w9737 & ~w9976 ;
  assign w9978 = w9572 ^ w9977 ;
  assign w9979 = ( ~w1675 & w9967 ) | ( ~w1675 & w9973 ) | ( w9967 & w9973 ) ;
  assign w9980 = ~w9967 & w9979 ;
  assign w9981 = w9978 | w9980 ;
  assign w9982 = ( w1517 & w9975 ) | ( w1517 & ~w9981 ) | ( w9975 & ~w9981 ) ;
  assign w9983 = w1517 & w9982 ;
  assign w9984 = w9577 | w9582 ;
  assign w9985 = w9737 & ~w9984 ;
  assign w9986 = w9580 ^ w9985 ;
  assign w9987 = ( ~w1517 & w9975 ) | ( ~w1517 & w9981 ) | ( w9975 & w9981 ) ;
  assign w9988 = ~w9975 & w9987 ;
  assign w9989 = w9986 | w9988 ;
  assign w9990 = ( w1367 & w9983 ) | ( w1367 & ~w9989 ) | ( w9983 & ~w9989 ) ;
  assign w9991 = w1367 & w9990 ;
  assign w9992 = ( ~w1367 & w9983 ) | ( ~w1367 & w9989 ) | ( w9983 & w9989 ) ;
  assign w9993 = ~w9983 & w9992 ;
  assign w9994 = w9585 | w9587 ;
  assign w9995 = w9737 & ~w9994 ;
  assign w9996 = w9590 ^ w9995 ;
  assign w9997 = w9993 | w9996 ;
  assign w9998 = ( w1225 & w9991 ) | ( w1225 & ~w9997 ) | ( w9991 & ~w9997 ) ;
  assign w9999 = w1225 & w9998 ;
  assign w10000 = w9593 | w9598 ;
  assign w10001 = w9737 & ~w10000 ;
  assign w10002 = w9596 ^ w10001 ;
  assign w10003 = ( ~w1225 & w9991 ) | ( ~w1225 & w9997 ) | ( w9991 & w9997 ) ;
  assign w10004 = ~w9991 & w10003 ;
  assign w10005 = w10002 | w10004 ;
  assign w10006 = ( w1091 & w9999 ) | ( w1091 & ~w10005 ) | ( w9999 & ~w10005 ) ;
  assign w10007 = w1091 & w10006 ;
  assign w10008 = w9601 | w9606 ;
  assign w10009 = w9737 & ~w10008 ;
  assign w10010 = w9604 ^ w10009 ;
  assign w10011 = ( ~w1091 & w9999 ) | ( ~w1091 & w10005 ) | ( w9999 & w10005 ) ;
  assign w10012 = ~w9999 & w10011 ;
  assign w10013 = w10010 | w10012 ;
  assign w10014 = ( w965 & w10007 ) | ( w965 & ~w10013 ) | ( w10007 & ~w10013 ) ;
  assign w10015 = w965 & w10014 ;
  assign w10016 = w9609 | w9614 ;
  assign w10017 = w9737 & ~w10016 ;
  assign w10018 = w9612 ^ w10017 ;
  assign w10019 = ( ~w965 & w10007 ) | ( ~w965 & w10013 ) | ( w10007 & w10013 ) ;
  assign w10020 = ~w10007 & w10019 ;
  assign w10021 = w10018 | w10020 ;
  assign w10022 = ( w847 & w10015 ) | ( w847 & ~w10021 ) | ( w10015 & ~w10021 ) ;
  assign w10023 = w847 & w10022 ;
  assign w10024 = w9617 | w9622 ;
  assign w10025 = w9737 & ~w10024 ;
  assign w10026 = w9620 ^ w10025 ;
  assign w10027 = ( ~w847 & w10015 ) | ( ~w847 & w10021 ) | ( w10015 & w10021 ) ;
  assign w10028 = ~w10015 & w10027 ;
  assign w10029 = w10026 | w10028 ;
  assign w10030 = ( w737 & w10023 ) | ( w737 & ~w10029 ) | ( w10023 & ~w10029 ) ;
  assign w10031 = w737 & w10030 ;
  assign w10032 = w9625 | w9630 ;
  assign w10033 = w9737 & ~w10032 ;
  assign w10034 = w9628 ^ w10033 ;
  assign w10035 = ( ~w737 & w10023 ) | ( ~w737 & w10029 ) | ( w10023 & w10029 ) ;
  assign w10036 = ~w10023 & w10035 ;
  assign w10037 = w10034 | w10036 ;
  assign w10038 = ( w635 & w10031 ) | ( w635 & ~w10037 ) | ( w10031 & ~w10037 ) ;
  assign w10039 = w635 & w10038 ;
  assign w10040 = w9633 | w9638 ;
  assign w10041 = w9737 & ~w10040 ;
  assign w10042 = w9636 ^ w10041 ;
  assign w10043 = ( ~w635 & w10031 ) | ( ~w635 & w10037 ) | ( w10031 & w10037 ) ;
  assign w10044 = ~w10031 & w10043 ;
  assign w10045 = w10042 | w10044 ;
  assign w10046 = ( w541 & w10039 ) | ( w541 & ~w10045 ) | ( w10039 & ~w10045 ) ;
  assign w10047 = w541 & w10046 ;
  assign w10048 = w9641 | w9646 ;
  assign w10049 = w9737 & ~w10048 ;
  assign w10050 = w9644 ^ w10049 ;
  assign w10051 = ( ~w541 & w10039 ) | ( ~w541 & w10045 ) | ( w10039 & w10045 ) ;
  assign w10052 = ~w10039 & w10051 ;
  assign w10053 = w10050 | w10052 ;
  assign w10054 = ( w455 & w10047 ) | ( w455 & ~w10053 ) | ( w10047 & ~w10053 ) ;
  assign w10055 = w455 & w10054 ;
  assign w10056 = w9649 | w9654 ;
  assign w10057 = w9737 & ~w10056 ;
  assign w10058 = w9652 ^ w10057 ;
  assign w10059 = ( ~w455 & w10047 ) | ( ~w455 & w10053 ) | ( w10047 & w10053 ) ;
  assign w10060 = ~w10047 & w10059 ;
  assign w10061 = w10058 | w10060 ;
  assign w10062 = ( w377 & w10055 ) | ( w377 & ~w10061 ) | ( w10055 & ~w10061 ) ;
  assign w10063 = w377 & w10062 ;
  assign w10064 = w9657 | w9662 ;
  assign w10065 = w9737 & ~w10064 ;
  assign w10066 = w9660 ^ w10065 ;
  assign w10067 = ( ~w377 & w10055 ) | ( ~w377 & w10061 ) | ( w10055 & w10061 ) ;
  assign w10068 = ~w10055 & w10067 ;
  assign w10069 = w10066 | w10068 ;
  assign w10070 = ( w307 & w10063 ) | ( w307 & ~w10069 ) | ( w10063 & ~w10069 ) ;
  assign w10071 = w307 & w10070 ;
  assign w10072 = w9665 | w9670 ;
  assign w10073 = w9737 & ~w10072 ;
  assign w10074 = w9668 ^ w10073 ;
  assign w10075 = ( ~w307 & w10063 ) | ( ~w307 & w10069 ) | ( w10063 & w10069 ) ;
  assign w10076 = ~w10063 & w10075 ;
  assign w10077 = w10074 | w10076 ;
  assign w10078 = ( w246 & w10071 ) | ( w246 & ~w10077 ) | ( w10071 & ~w10077 ) ;
  assign w10079 = w246 & w10078 ;
  assign w10080 = w9673 | w9678 ;
  assign w10081 = w9737 & ~w10080 ;
  assign w10082 = w9676 ^ w10081 ;
  assign w10083 = ( ~w246 & w10071 ) | ( ~w246 & w10077 ) | ( w10071 & w10077 ) ;
  assign w10084 = ~w10071 & w10083 ;
  assign w10085 = w10082 | w10084 ;
  assign w10086 = ( w185 & w10079 ) | ( w185 & ~w10085 ) | ( w10079 & ~w10085 ) ;
  assign w10087 = w185 & w10086 ;
  assign w10088 = w9681 | w9686 ;
  assign w10089 = w9737 & ~w10088 ;
  assign w10090 = w9684 ^ w10089 ;
  assign w10091 = ( ~w185 & w10079 ) | ( ~w185 & w10085 ) | ( w10079 & w10085 ) ;
  assign w10092 = ~w10079 & w10091 ;
  assign w10093 = w10090 | w10092 ;
  assign w10094 = ( w145 & w10087 ) | ( w145 & ~w10093 ) | ( w10087 & ~w10093 ) ;
  assign w10095 = w145 & w10094 ;
  assign w10096 = w9689 | w9694 ;
  assign w10097 = w9737 & ~w10096 ;
  assign w10098 = w9692 ^ w10097 ;
  assign w10099 = ( ~w145 & w10087 ) | ( ~w145 & w10093 ) | ( w10087 & w10093 ) ;
  assign w10100 = ~w10087 & w10099 ;
  assign w10101 = w10098 | w10100 ;
  assign w10102 = ( w132 & w10095 ) | ( w132 & ~w10101 ) | ( w10095 & ~w10101 ) ;
  assign w10103 = w132 & w10102 ;
  assign w10104 = w9697 | w9702 ;
  assign w10105 = w9737 & ~w10104 ;
  assign w10106 = w9700 ^ w10105 ;
  assign w10107 = ( ~w132 & w10095 ) | ( ~w132 & w10101 ) | ( w10095 & w10101 ) ;
  assign w10108 = ~w10095 & w10107 ;
  assign w10109 = w10106 | w10108 ;
  assign w10110 = ~w10103 & w10109 ;
  assign w10111 = w9705 | w9710 ;
  assign w10112 = w9737 & ~w10111 ;
  assign w10113 = w9708 ^ w10112 ;
  assign w10114 = ( ~w9723 & w10110 ) | ( ~w9723 & w10113 ) | ( w10110 & w10113 ) ;
  assign w10115 = w9712 & ~w10114 ;
  assign w10116 = ~w9715 & w9737 ;
  assign w10117 = ( w10114 & ~w10115 ) | ( w10114 & w10116 ) | ( ~w10115 & w10116 ) ;
  assign w10118 = w9723 | w10117 ;
  assign w10119 = ~w129 & w10118 ;
  assign w10120 = ( w10103 & w10109 ) | ( w10103 & w10113 ) | ( w10109 & w10113 ) ;
  assign w10121 = ~w10103 & w10120 ;
  assign w10122 = ( w129 & w9712 ) | ( w129 & w9715 ) | ( w9712 & w9715 ) ;
  assign w10123 = ( w9715 & ~w9737 ) | ( w9715 & w10122 ) | ( ~w9737 & w10122 ) ;
  assign w10124 = w9712 & w10123 ;
  assign w10125 = w10122 ^ w10124 ;
  assign w10126 = ( w9315 & w9320 ) | ( w9315 & w9347 ) | ( w9320 & w9347 ) ;
  assign w10127 = w9347 & ~w10126 ;
  assign w10128 = w9318 ^ w10127 ;
  assign w10129 = ( ~w9727 & w9734 ) | ( ~w9727 & w10128 ) | ( w9734 & w10128 ) ;
  assign w10130 = ~w9734 & w10129 ;
  assign w10131 = ( ~w9721 & w9723 ) | ( ~w9721 & w10130 ) | ( w9723 & w10130 ) ;
  assign w10132 = ~w9723 & w10131 ;
  assign w10133 = w10121 | w10132 ;
  assign w10134 = ( w10119 & ~w10121 ) | ( w10119 & w10125 ) | ( ~w10121 & w10125 ) ;
  assign w10135 = w10133 | w10134 ;
  assign w10136 = ( ~\pi031 & \pi032 ) | ( ~\pi031 & w9737 ) | ( \pi032 & w9737 ) ;
  assign w10137 = ( ~\pi030 & \pi032 ) | ( ~\pi030 & w10136 ) | ( \pi032 & w10136 ) ;
  assign w10138 = ( ~\pi032 & w9737 ) | ( ~\pi032 & w10135 ) | ( w9737 & w10135 ) ;
  assign w10139 = w10137 & w10138 ;
  assign w10140 = ( w9723 & w9727 ) | ( w9723 & ~w9734 ) | ( w9727 & ~w9734 ) ;
  assign w10141 = \pi031 & ~w10140 ;
  assign w10142 = \pi030 | \pi032 ;
  assign w10143 = ( ~w10140 & w10141 ) | ( ~w10140 & w10142 ) | ( w10141 & w10142 ) ;
  assign w10144 = ~w9734 & w10143 ;
  assign w10145 = ~w9721 & w10144 ;
  assign w10146 = ( \pi032 & w10135 ) | ( \pi032 & ~w10144 ) | ( w10135 & ~w10144 ) ;
  assign w10147 = w10145 & ~w10146 ;
  assign w10148 = ~\pi032 & w10135 ;
  assign w10149 = \pi033 ^ w10148 ;
  assign w10150 = w10147 | w10149 ;
  assign w10151 = ( w9347 & w10139 ) | ( w9347 & ~w10150 ) | ( w10139 & ~w10150 ) ;
  assign w10152 = w9347 & w10151 ;
  assign w10153 = ( ~w9347 & w10139 ) | ( ~w9347 & w10150 ) | ( w10139 & w10150 ) ;
  assign w10154 = ~w10139 & w10153 ;
  assign w10155 = w9737 & ~w10132 ;
  assign w10156 = ~w10121 & w10155 ;
  assign w10157 = ~w10134 & w10156 ;
  assign w10158 = \pi033 & w10135 ;
  assign w10159 = ( \pi032 & w10135 ) | ( \pi032 & ~w10158 ) | ( w10135 & ~w10158 ) ;
  assign w10160 = ( ~\pi032 & w10157 ) | ( ~\pi032 & w10159 ) | ( w10157 & w10159 ) ;
  assign w10161 = \pi034 ^ w10160 ;
  assign w10162 = w10154 | w10161 ;
  assign w10163 = ( w8965 & w10152 ) | ( w8965 & ~w10162 ) | ( w10152 & ~w10162 ) ;
  assign w10164 = w8965 & w10163 ;
  assign w10165 = ( w9741 & ~w9749 ) | ( w9741 & w10135 ) | ( ~w9749 & w10135 ) ;
  assign w10166 = ~w9741 & w10165 ;
  assign w10167 = \pi035 ^ w10166 ;
  assign w10168 = w9750 ^ w10167 ;
  assign w10169 = ( ~w8965 & w10152 ) | ( ~w8965 & w10162 ) | ( w10152 & w10162 ) ;
  assign w10170 = ~w10152 & w10169 ;
  assign w10171 = w10168 | w10170 ;
  assign w10172 = ( w8591 & w10164 ) | ( w8591 & ~w10171 ) | ( w10164 & ~w10171 ) ;
  assign w10173 = w8591 & w10172 ;
  assign w10174 = w9754 | w9756 ;
  assign w10175 = w10135 & ~w10174 ;
  assign w10176 = w9763 ^ w10175 ;
  assign w10177 = ( ~w8591 & w10164 ) | ( ~w8591 & w10171 ) | ( w10164 & w10171 ) ;
  assign w10178 = ~w10164 & w10177 ;
  assign w10179 = w10176 | w10178 ;
  assign w10180 = ( w8225 & w10173 ) | ( w8225 & ~w10179 ) | ( w10173 & ~w10179 ) ;
  assign w10181 = w8225 & w10180 ;
  assign w10182 = w9766 | w9772 ;
  assign w10183 = w10135 & ~w10182 ;
  assign w10184 = w9770 ^ w10183 ;
  assign w10185 = ( ~w8225 & w10173 ) | ( ~w8225 & w10179 ) | ( w10173 & w10179 ) ;
  assign w10186 = ~w10173 & w10185 ;
  assign w10187 = w10184 | w10186 ;
  assign w10188 = ( w7867 & w10181 ) | ( w7867 & ~w10187 ) | ( w10181 & ~w10187 ) ;
  assign w10189 = w7867 & w10188 ;
  assign w10190 = w9775 | w9780 ;
  assign w10191 = w10135 & ~w10190 ;
  assign w10192 = w9778 ^ w10191 ;
  assign w10193 = ( ~w7867 & w10181 ) | ( ~w7867 & w10187 ) | ( w10181 & w10187 ) ;
  assign w10194 = ~w10181 & w10193 ;
  assign w10195 = w10192 | w10194 ;
  assign w10196 = ( w7517 & w10189 ) | ( w7517 & ~w10195 ) | ( w10189 & ~w10195 ) ;
  assign w10197 = w7517 & w10196 ;
  assign w10198 = w9783 | w9788 ;
  assign w10199 = w10135 & ~w10198 ;
  assign w10200 = w9786 ^ w10199 ;
  assign w10201 = ( ~w7517 & w10189 ) | ( ~w7517 & w10195 ) | ( w10189 & w10195 ) ;
  assign w10202 = ~w10189 & w10201 ;
  assign w10203 = w10200 | w10202 ;
  assign w10204 = ( w7175 & w10197 ) | ( w7175 & ~w10203 ) | ( w10197 & ~w10203 ) ;
  assign w10205 = w7175 & w10204 ;
  assign w10206 = w9791 | w9796 ;
  assign w10207 = w10135 & ~w10206 ;
  assign w10208 = w9794 ^ w10207 ;
  assign w10209 = ( ~w7175 & w10197 ) | ( ~w7175 & w10203 ) | ( w10197 & w10203 ) ;
  assign w10210 = ~w10197 & w10209 ;
  assign w10211 = w10208 | w10210 ;
  assign w10212 = ( w6841 & w10205 ) | ( w6841 & ~w10211 ) | ( w10205 & ~w10211 ) ;
  assign w10213 = w6841 & w10212 ;
  assign w10214 = w9799 | w9804 ;
  assign w10215 = w10135 & ~w10214 ;
  assign w10216 = w9802 ^ w10215 ;
  assign w10217 = ( ~w6841 & w10205 ) | ( ~w6841 & w10211 ) | ( w10205 & w10211 ) ;
  assign w10218 = ~w10205 & w10217 ;
  assign w10219 = w10216 | w10218 ;
  assign w10220 = ( w6515 & w10213 ) | ( w6515 & ~w10219 ) | ( w10213 & ~w10219 ) ;
  assign w10221 = w6515 & w10220 ;
  assign w10222 = w9807 | w9812 ;
  assign w10223 = w10135 & ~w10222 ;
  assign w10224 = w9810 ^ w10223 ;
  assign w10225 = ( ~w6515 & w10213 ) | ( ~w6515 & w10219 ) | ( w10213 & w10219 ) ;
  assign w10226 = ~w10213 & w10225 ;
  assign w10227 = w10224 | w10226 ;
  assign w10228 = ( w6197 & w10221 ) | ( w6197 & ~w10227 ) | ( w10221 & ~w10227 ) ;
  assign w10229 = w6197 & w10228 ;
  assign w10230 = w9815 | w9820 ;
  assign w10231 = w10135 & ~w10230 ;
  assign w10232 = w9818 ^ w10231 ;
  assign w10233 = ( ~w6197 & w10221 ) | ( ~w6197 & w10227 ) | ( w10221 & w10227 ) ;
  assign w10234 = ~w10221 & w10233 ;
  assign w10235 = w10232 | w10234 ;
  assign w10236 = ( w5887 & w10229 ) | ( w5887 & ~w10235 ) | ( w10229 & ~w10235 ) ;
  assign w10237 = w5887 & w10236 ;
  assign w10238 = w9823 | w9828 ;
  assign w10239 = w10135 & ~w10238 ;
  assign w10240 = w9826 ^ w10239 ;
  assign w10241 = ( ~w5887 & w10229 ) | ( ~w5887 & w10235 ) | ( w10229 & w10235 ) ;
  assign w10242 = ~w10229 & w10241 ;
  assign w10243 = w10240 | w10242 ;
  assign w10244 = ( w5585 & w10237 ) | ( w5585 & ~w10243 ) | ( w10237 & ~w10243 ) ;
  assign w10245 = w5585 & w10244 ;
  assign w10246 = w9831 | w9836 ;
  assign w10247 = w10135 & ~w10246 ;
  assign w10248 = w9834 ^ w10247 ;
  assign w10249 = ( ~w5585 & w10237 ) | ( ~w5585 & w10243 ) | ( w10237 & w10243 ) ;
  assign w10250 = ~w10237 & w10249 ;
  assign w10251 = w10248 | w10250 ;
  assign w10252 = ( w5291 & w10245 ) | ( w5291 & ~w10251 ) | ( w10245 & ~w10251 ) ;
  assign w10253 = w5291 & w10252 ;
  assign w10254 = w9839 | w9844 ;
  assign w10255 = w10135 & ~w10254 ;
  assign w10256 = w9842 ^ w10255 ;
  assign w10257 = ( ~w5291 & w10245 ) | ( ~w5291 & w10251 ) | ( w10245 & w10251 ) ;
  assign w10258 = ~w10245 & w10257 ;
  assign w10259 = w10256 | w10258 ;
  assign w10260 = ( w5005 & w10253 ) | ( w5005 & ~w10259 ) | ( w10253 & ~w10259 ) ;
  assign w10261 = w5005 & w10260 ;
  assign w10262 = w9847 | w9852 ;
  assign w10263 = w10135 & ~w10262 ;
  assign w10264 = w9850 ^ w10263 ;
  assign w10265 = ( ~w5005 & w10253 ) | ( ~w5005 & w10259 ) | ( w10253 & w10259 ) ;
  assign w10266 = ~w10253 & w10265 ;
  assign w10267 = w10264 | w10266 ;
  assign w10268 = ( w4727 & w10261 ) | ( w4727 & ~w10267 ) | ( w10261 & ~w10267 ) ;
  assign w10269 = w4727 & w10268 ;
  assign w10270 = w9855 | w9860 ;
  assign w10271 = w10135 & ~w10270 ;
  assign w10272 = w9858 ^ w10271 ;
  assign w10273 = ( ~w4727 & w10261 ) | ( ~w4727 & w10267 ) | ( w10261 & w10267 ) ;
  assign w10274 = ~w10261 & w10273 ;
  assign w10275 = w10272 | w10274 ;
  assign w10276 = ( w4457 & w10269 ) | ( w4457 & ~w10275 ) | ( w10269 & ~w10275 ) ;
  assign w10277 = w4457 & w10276 ;
  assign w10278 = w9863 | w9868 ;
  assign w10279 = w10135 & ~w10278 ;
  assign w10280 = w9866 ^ w10279 ;
  assign w10281 = ( ~w4457 & w10269 ) | ( ~w4457 & w10275 ) | ( w10269 & w10275 ) ;
  assign w10282 = ~w10269 & w10281 ;
  assign w10283 = w10280 | w10282 ;
  assign w10284 = ( w4195 & w10277 ) | ( w4195 & ~w10283 ) | ( w10277 & ~w10283 ) ;
  assign w10285 = w4195 & w10284 ;
  assign w10286 = w9871 | w9876 ;
  assign w10287 = w10135 & ~w10286 ;
  assign w10288 = w9874 ^ w10287 ;
  assign w10289 = ( ~w4195 & w10277 ) | ( ~w4195 & w10283 ) | ( w10277 & w10283 ) ;
  assign w10290 = ~w10277 & w10289 ;
  assign w10291 = w10288 | w10290 ;
  assign w10292 = ( w3941 & w10285 ) | ( w3941 & ~w10291 ) | ( w10285 & ~w10291 ) ;
  assign w10293 = w3941 & w10292 ;
  assign w10294 = w9879 | w9884 ;
  assign w10295 = w10135 & ~w10294 ;
  assign w10296 = w9882 ^ w10295 ;
  assign w10297 = ( ~w3941 & w10285 ) | ( ~w3941 & w10291 ) | ( w10285 & w10291 ) ;
  assign w10298 = ~w10285 & w10297 ;
  assign w10299 = w10296 | w10298 ;
  assign w10300 = ( w3695 & w10293 ) | ( w3695 & ~w10299 ) | ( w10293 & ~w10299 ) ;
  assign w10301 = w3695 & w10300 ;
  assign w10302 = w9887 | w9892 ;
  assign w10303 = w10135 & ~w10302 ;
  assign w10304 = w9890 ^ w10303 ;
  assign w10305 = ( ~w3695 & w10293 ) | ( ~w3695 & w10299 ) | ( w10293 & w10299 ) ;
  assign w10306 = ~w10293 & w10305 ;
  assign w10307 = w10304 | w10306 ;
  assign w10308 = ( w3457 & w10301 ) | ( w3457 & ~w10307 ) | ( w10301 & ~w10307 ) ;
  assign w10309 = w3457 & w10308 ;
  assign w10310 = w9895 | w9900 ;
  assign w10311 = w10135 & ~w10310 ;
  assign w10312 = w9898 ^ w10311 ;
  assign w10313 = ( ~w3457 & w10301 ) | ( ~w3457 & w10307 ) | ( w10301 & w10307 ) ;
  assign w10314 = ~w10301 & w10313 ;
  assign w10315 = w10312 | w10314 ;
  assign w10316 = ( w3227 & w10309 ) | ( w3227 & ~w10315 ) | ( w10309 & ~w10315 ) ;
  assign w10317 = w3227 & w10316 ;
  assign w10318 = w9903 | w9908 ;
  assign w10319 = w10135 & ~w10318 ;
  assign w10320 = w9906 ^ w10319 ;
  assign w10321 = ( ~w3227 & w10309 ) | ( ~w3227 & w10315 ) | ( w10309 & w10315 ) ;
  assign w10322 = ~w10309 & w10321 ;
  assign w10323 = w10320 | w10322 ;
  assign w10324 = ( w3005 & w10317 ) | ( w3005 & ~w10323 ) | ( w10317 & ~w10323 ) ;
  assign w10325 = w3005 & w10324 ;
  assign w10326 = w9911 | w9916 ;
  assign w10327 = w10135 & ~w10326 ;
  assign w10328 = w9914 ^ w10327 ;
  assign w10329 = ( ~w3005 & w10317 ) | ( ~w3005 & w10323 ) | ( w10317 & w10323 ) ;
  assign w10330 = ~w10317 & w10329 ;
  assign w10331 = w10328 | w10330 ;
  assign w10332 = ( w2791 & w10325 ) | ( w2791 & ~w10331 ) | ( w10325 & ~w10331 ) ;
  assign w10333 = w2791 & w10332 ;
  assign w10334 = w9919 | w9924 ;
  assign w10335 = w10135 & ~w10334 ;
  assign w10336 = w9922 ^ w10335 ;
  assign w10337 = ( ~w2791 & w10325 ) | ( ~w2791 & w10331 ) | ( w10325 & w10331 ) ;
  assign w10338 = ~w10325 & w10337 ;
  assign w10339 = w10336 | w10338 ;
  assign w10340 = ( w2585 & w10333 ) | ( w2585 & ~w10339 ) | ( w10333 & ~w10339 ) ;
  assign w10341 = w2585 & w10340 ;
  assign w10342 = w9927 | w9932 ;
  assign w10343 = w10135 & ~w10342 ;
  assign w10344 = w9930 ^ w10343 ;
  assign w10345 = ( ~w2585 & w10333 ) | ( ~w2585 & w10339 ) | ( w10333 & w10339 ) ;
  assign w10346 = ~w10333 & w10345 ;
  assign w10347 = w10344 | w10346 ;
  assign w10348 = ( w2387 & w10341 ) | ( w2387 & ~w10347 ) | ( w10341 & ~w10347 ) ;
  assign w10349 = w2387 & w10348 ;
  assign w10350 = w9935 | w9940 ;
  assign w10351 = w10135 & ~w10350 ;
  assign w10352 = w9938 ^ w10351 ;
  assign w10353 = ( ~w2387 & w10341 ) | ( ~w2387 & w10347 ) | ( w10341 & w10347 ) ;
  assign w10354 = ~w10341 & w10353 ;
  assign w10355 = w10352 | w10354 ;
  assign w10356 = ( w2197 & w10349 ) | ( w2197 & ~w10355 ) | ( w10349 & ~w10355 ) ;
  assign w10357 = w2197 & w10356 ;
  assign w10358 = w9943 | w9948 ;
  assign w10359 = w10135 & ~w10358 ;
  assign w10360 = w9946 ^ w10359 ;
  assign w10361 = ( ~w2197 & w10349 ) | ( ~w2197 & w10355 ) | ( w10349 & w10355 ) ;
  assign w10362 = ~w10349 & w10361 ;
  assign w10363 = w10360 | w10362 ;
  assign w10364 = ( w2015 & w10357 ) | ( w2015 & ~w10363 ) | ( w10357 & ~w10363 ) ;
  assign w10365 = w2015 & w10364 ;
  assign w10366 = w9951 | w9956 ;
  assign w10367 = w10135 & ~w10366 ;
  assign w10368 = w9954 ^ w10367 ;
  assign w10369 = ( ~w2015 & w10357 ) | ( ~w2015 & w10363 ) | ( w10357 & w10363 ) ;
  assign w10370 = ~w10357 & w10369 ;
  assign w10371 = w10368 | w10370 ;
  assign w10372 = ( w1841 & w10365 ) | ( w1841 & ~w10371 ) | ( w10365 & ~w10371 ) ;
  assign w10373 = w1841 & w10372 ;
  assign w10374 = w9959 | w9964 ;
  assign w10375 = w10135 & ~w10374 ;
  assign w10376 = w9962 ^ w10375 ;
  assign w10377 = ( ~w1841 & w10365 ) | ( ~w1841 & w10371 ) | ( w10365 & w10371 ) ;
  assign w10378 = ~w10365 & w10377 ;
  assign w10379 = w10376 | w10378 ;
  assign w10380 = ( w1675 & w10373 ) | ( w1675 & ~w10379 ) | ( w10373 & ~w10379 ) ;
  assign w10381 = w1675 & w10380 ;
  assign w10382 = w9967 | w9972 ;
  assign w10383 = w10135 & ~w10382 ;
  assign w10384 = w9970 ^ w10383 ;
  assign w10385 = ( ~w1675 & w10373 ) | ( ~w1675 & w10379 ) | ( w10373 & w10379 ) ;
  assign w10386 = ~w10373 & w10385 ;
  assign w10387 = w10384 | w10386 ;
  assign w10388 = ( w1517 & w10381 ) | ( w1517 & ~w10387 ) | ( w10381 & ~w10387 ) ;
  assign w10389 = w1517 & w10388 ;
  assign w10390 = w9975 | w9980 ;
  assign w10391 = w10135 & ~w10390 ;
  assign w10392 = w9978 ^ w10391 ;
  assign w10393 = ( ~w1517 & w10381 ) | ( ~w1517 & w10387 ) | ( w10381 & w10387 ) ;
  assign w10394 = ~w10381 & w10393 ;
  assign w10395 = w10392 | w10394 ;
  assign w10396 = ( w1367 & w10389 ) | ( w1367 & ~w10395 ) | ( w10389 & ~w10395 ) ;
  assign w10397 = w1367 & w10396 ;
  assign w10398 = w9983 | w9988 ;
  assign w10399 = w10135 & ~w10398 ;
  assign w10400 = w9986 ^ w10399 ;
  assign w10401 = ( ~w1367 & w10389 ) | ( ~w1367 & w10395 ) | ( w10389 & w10395 ) ;
  assign w10402 = ~w10389 & w10401 ;
  assign w10403 = w10400 | w10402 ;
  assign w10404 = ( w1225 & w10397 ) | ( w1225 & ~w10403 ) | ( w10397 & ~w10403 ) ;
  assign w10405 = w1225 & w10404 ;
  assign w10406 = ( ~w1225 & w10397 ) | ( ~w1225 & w10403 ) | ( w10397 & w10403 ) ;
  assign w10407 = ~w10397 & w10406 ;
  assign w10408 = w9991 | w9993 ;
  assign w10409 = w10135 & ~w10408 ;
  assign w10410 = w9996 ^ w10409 ;
  assign w10411 = w10407 | w10410 ;
  assign w10412 = ( w1091 & w10405 ) | ( w1091 & ~w10411 ) | ( w10405 & ~w10411 ) ;
  assign w10413 = w1091 & w10412 ;
  assign w10414 = w9999 | w10004 ;
  assign w10415 = w10135 & ~w10414 ;
  assign w10416 = w10002 ^ w10415 ;
  assign w10417 = ( ~w1091 & w10405 ) | ( ~w1091 & w10411 ) | ( w10405 & w10411 ) ;
  assign w10418 = ~w10405 & w10417 ;
  assign w10419 = w10416 | w10418 ;
  assign w10420 = ( w965 & w10413 ) | ( w965 & ~w10419 ) | ( w10413 & ~w10419 ) ;
  assign w10421 = w965 & w10420 ;
  assign w10422 = w10007 | w10012 ;
  assign w10423 = w10135 & ~w10422 ;
  assign w10424 = w10010 ^ w10423 ;
  assign w10425 = ( ~w965 & w10413 ) | ( ~w965 & w10419 ) | ( w10413 & w10419 ) ;
  assign w10426 = ~w10413 & w10425 ;
  assign w10427 = w10424 | w10426 ;
  assign w10428 = ( w847 & w10421 ) | ( w847 & ~w10427 ) | ( w10421 & ~w10427 ) ;
  assign w10429 = w847 & w10428 ;
  assign w10430 = w10015 | w10020 ;
  assign w10431 = w10135 & ~w10430 ;
  assign w10432 = w10018 ^ w10431 ;
  assign w10433 = ( ~w847 & w10421 ) | ( ~w847 & w10427 ) | ( w10421 & w10427 ) ;
  assign w10434 = ~w10421 & w10433 ;
  assign w10435 = w10432 | w10434 ;
  assign w10436 = ( w737 & w10429 ) | ( w737 & ~w10435 ) | ( w10429 & ~w10435 ) ;
  assign w10437 = w737 & w10436 ;
  assign w10438 = w10023 | w10028 ;
  assign w10439 = w10135 & ~w10438 ;
  assign w10440 = w10026 ^ w10439 ;
  assign w10441 = ( ~w737 & w10429 ) | ( ~w737 & w10435 ) | ( w10429 & w10435 ) ;
  assign w10442 = ~w10429 & w10441 ;
  assign w10443 = w10440 | w10442 ;
  assign w10444 = ( w635 & w10437 ) | ( w635 & ~w10443 ) | ( w10437 & ~w10443 ) ;
  assign w10445 = w635 & w10444 ;
  assign w10446 = w10031 | w10036 ;
  assign w10447 = w10135 & ~w10446 ;
  assign w10448 = w10034 ^ w10447 ;
  assign w10449 = ( ~w635 & w10437 ) | ( ~w635 & w10443 ) | ( w10437 & w10443 ) ;
  assign w10450 = ~w10437 & w10449 ;
  assign w10451 = w10448 | w10450 ;
  assign w10452 = ( w541 & w10445 ) | ( w541 & ~w10451 ) | ( w10445 & ~w10451 ) ;
  assign w10453 = w541 & w10452 ;
  assign w10454 = w10039 | w10044 ;
  assign w10455 = w10135 & ~w10454 ;
  assign w10456 = w10042 ^ w10455 ;
  assign w10457 = ( ~w541 & w10445 ) | ( ~w541 & w10451 ) | ( w10445 & w10451 ) ;
  assign w10458 = ~w10445 & w10457 ;
  assign w10459 = w10456 | w10458 ;
  assign w10460 = ( w455 & w10453 ) | ( w455 & ~w10459 ) | ( w10453 & ~w10459 ) ;
  assign w10461 = w455 & w10460 ;
  assign w10462 = w10047 | w10052 ;
  assign w10463 = w10135 & ~w10462 ;
  assign w10464 = w10050 ^ w10463 ;
  assign w10465 = ( ~w455 & w10453 ) | ( ~w455 & w10459 ) | ( w10453 & w10459 ) ;
  assign w10466 = ~w10453 & w10465 ;
  assign w10467 = w10464 | w10466 ;
  assign w10468 = ( w377 & w10461 ) | ( w377 & ~w10467 ) | ( w10461 & ~w10467 ) ;
  assign w10469 = w377 & w10468 ;
  assign w10470 = w10055 | w10060 ;
  assign w10471 = w10135 & ~w10470 ;
  assign w10472 = w10058 ^ w10471 ;
  assign w10473 = ( ~w377 & w10461 ) | ( ~w377 & w10467 ) | ( w10461 & w10467 ) ;
  assign w10474 = ~w10461 & w10473 ;
  assign w10475 = w10472 | w10474 ;
  assign w10476 = ( w307 & w10469 ) | ( w307 & ~w10475 ) | ( w10469 & ~w10475 ) ;
  assign w10477 = w307 & w10476 ;
  assign w10478 = w10063 | w10068 ;
  assign w10479 = w10135 & ~w10478 ;
  assign w10480 = w10066 ^ w10479 ;
  assign w10481 = ( ~w307 & w10469 ) | ( ~w307 & w10475 ) | ( w10469 & w10475 ) ;
  assign w10482 = ~w10469 & w10481 ;
  assign w10483 = w10480 | w10482 ;
  assign w10484 = ( w246 & w10477 ) | ( w246 & ~w10483 ) | ( w10477 & ~w10483 ) ;
  assign w10485 = w246 & w10484 ;
  assign w10486 = w10071 | w10076 ;
  assign w10487 = w10135 & ~w10486 ;
  assign w10488 = w10074 ^ w10487 ;
  assign w10489 = ( ~w246 & w10477 ) | ( ~w246 & w10483 ) | ( w10477 & w10483 ) ;
  assign w10490 = ~w10477 & w10489 ;
  assign w10491 = w10488 | w10490 ;
  assign w10492 = ( w185 & w10485 ) | ( w185 & ~w10491 ) | ( w10485 & ~w10491 ) ;
  assign w10493 = w185 & w10492 ;
  assign w10494 = w10079 | w10084 ;
  assign w10495 = w10135 & ~w10494 ;
  assign w10496 = w10082 ^ w10495 ;
  assign w10497 = ( ~w185 & w10485 ) | ( ~w185 & w10491 ) | ( w10485 & w10491 ) ;
  assign w10498 = ~w10485 & w10497 ;
  assign w10499 = w10496 | w10498 ;
  assign w10500 = ( w145 & w10493 ) | ( w145 & ~w10499 ) | ( w10493 & ~w10499 ) ;
  assign w10501 = w145 & w10500 ;
  assign w10502 = w10087 | w10092 ;
  assign w10503 = w10135 & ~w10502 ;
  assign w10504 = w10090 ^ w10503 ;
  assign w10505 = ( ~w145 & w10493 ) | ( ~w145 & w10499 ) | ( w10493 & w10499 ) ;
  assign w10506 = ~w10493 & w10505 ;
  assign w10507 = w10504 | w10506 ;
  assign w10508 = ( w132 & w10501 ) | ( w132 & ~w10507 ) | ( w10501 & ~w10507 ) ;
  assign w10509 = w132 & w10508 ;
  assign w10510 = w10095 | w10100 ;
  assign w10511 = w10135 & ~w10510 ;
  assign w10512 = w10098 ^ w10511 ;
  assign w10513 = ( ~w132 & w10501 ) | ( ~w132 & w10507 ) | ( w10501 & w10507 ) ;
  assign w10514 = ~w10501 & w10513 ;
  assign w10515 = w10512 | w10514 ;
  assign w10516 = ~w10509 & w10515 ;
  assign w10517 = w10103 | w10108 ;
  assign w10518 = w10135 & ~w10517 ;
  assign w10519 = w10106 ^ w10518 ;
  assign w10520 = ( ~w10121 & w10516 ) | ( ~w10121 & w10519 ) | ( w10516 & w10519 ) ;
  assign w10521 = w10110 & ~w10520 ;
  assign w10522 = ~w10113 & w10135 ;
  assign w10523 = ( w10520 & ~w10521 ) | ( w10520 & w10522 ) | ( ~w10521 & w10522 ) ;
  assign w10524 = w10121 | w10523 ;
  assign w10525 = ~w129 & w10524 ;
  assign w10526 = ( w10509 & w10515 ) | ( w10509 & w10519 ) | ( w10515 & w10519 ) ;
  assign w10527 = ~w10509 & w10526 ;
  assign w10528 = ( w129 & w10110 ) | ( w129 & w10113 ) | ( w10110 & w10113 ) ;
  assign w10529 = ( w10113 & ~w10135 ) | ( w10113 & w10528 ) | ( ~w10135 & w10528 ) ;
  assign w10530 = w10110 & w10529 ;
  assign w10531 = w10528 ^ w10530 ;
  assign w10532 = ( w9705 & w9710 ) | ( w9705 & w9737 ) | ( w9710 & w9737 ) ;
  assign w10533 = w9737 & ~w10532 ;
  assign w10534 = w9708 ^ w10533 ;
  assign w10535 = ( ~w10125 & w10132 ) | ( ~w10125 & w10534 ) | ( w10132 & w10534 ) ;
  assign w10536 = ~w10132 & w10535 ;
  assign w10537 = ( ~w10119 & w10121 ) | ( ~w10119 & w10536 ) | ( w10121 & w10536 ) ;
  assign w10538 = ~w10121 & w10537 ;
  assign w10539 = w10527 | w10538 ;
  assign w10540 = ( w10525 & ~w10527 ) | ( w10525 & w10531 ) | ( ~w10527 & w10531 ) ;
  assign w10541 = w10539 | w10540 ;
  assign w10542 = ( ~\pi029 & \pi030 ) | ( ~\pi029 & w10135 ) | ( \pi030 & w10135 ) ;
  assign w10543 = ( ~\pi028 & \pi030 ) | ( ~\pi028 & w10542 ) | ( \pi030 & w10542 ) ;
  assign w10544 = ( ~\pi030 & w10135 ) | ( ~\pi030 & w10541 ) | ( w10135 & w10541 ) ;
  assign w10545 = w10543 & w10544 ;
  assign w10546 = ( w10121 & w10125 ) | ( w10121 & ~w10132 ) | ( w10125 & ~w10132 ) ;
  assign w10547 = \pi029 & ~w10546 ;
  assign w10548 = \pi028 | \pi030 ;
  assign w10549 = ( ~w10546 & w10547 ) | ( ~w10546 & w10548 ) | ( w10547 & w10548 ) ;
  assign w10550 = ~w10132 & w10549 ;
  assign w10551 = ~w10119 & w10550 ;
  assign w10552 = ( \pi030 & w10541 ) | ( \pi030 & ~w10550 ) | ( w10541 & ~w10550 ) ;
  assign w10553 = w10551 & ~w10552 ;
  assign w10554 = ~\pi030 & w10541 ;
  assign w10555 = \pi031 ^ w10554 ;
  assign w10556 = w10553 | w10555 ;
  assign w10557 = ( w9737 & w10545 ) | ( w9737 & ~w10556 ) | ( w10545 & ~w10556 ) ;
  assign w10558 = w9737 & w10557 ;
  assign w10559 = ( ~w9737 & w10545 ) | ( ~w9737 & w10556 ) | ( w10545 & w10556 ) ;
  assign w10560 = ~w10545 & w10559 ;
  assign w10561 = w10135 & ~w10538 ;
  assign w10562 = ~w10527 & w10561 ;
  assign w10563 = ~w10540 & w10562 ;
  assign w10564 = \pi031 & w10541 ;
  assign w10565 = ( \pi030 & w10541 ) | ( \pi030 & ~w10564 ) | ( w10541 & ~w10564 ) ;
  assign w10566 = ( ~\pi030 & w10563 ) | ( ~\pi030 & w10565 ) | ( w10563 & w10565 ) ;
  assign w10567 = \pi032 ^ w10566 ;
  assign w10568 = w10560 | w10567 ;
  assign w10569 = ( w9347 & w10558 ) | ( w9347 & ~w10568 ) | ( w10558 & ~w10568 ) ;
  assign w10570 = w9347 & w10569 ;
  assign w10571 = ( w10139 & ~w10147 ) | ( w10139 & w10541 ) | ( ~w10147 & w10541 ) ;
  assign w10572 = ~w10139 & w10571 ;
  assign w10573 = \pi033 ^ w10572 ;
  assign w10574 = w10148 ^ w10573 ;
  assign w10575 = ( ~w9347 & w10558 ) | ( ~w9347 & w10568 ) | ( w10558 & w10568 ) ;
  assign w10576 = ~w10558 & w10575 ;
  assign w10577 = w10574 | w10576 ;
  assign w10578 = ( w8965 & w10570 ) | ( w8965 & ~w10577 ) | ( w10570 & ~w10577 ) ;
  assign w10579 = w8965 & w10578 ;
  assign w10580 = w10152 | w10154 ;
  assign w10581 = w10541 & ~w10580 ;
  assign w10582 = w10161 ^ w10581 ;
  assign w10583 = ( ~w8965 & w10570 ) | ( ~w8965 & w10577 ) | ( w10570 & w10577 ) ;
  assign w10584 = ~w10570 & w10583 ;
  assign w10585 = w10582 | w10584 ;
  assign w10586 = ( w8591 & w10579 ) | ( w8591 & ~w10585 ) | ( w10579 & ~w10585 ) ;
  assign w10587 = w8591 & w10586 ;
  assign w10588 = w10164 | w10170 ;
  assign w10589 = w10541 & ~w10588 ;
  assign w10590 = w10168 ^ w10589 ;
  assign w10591 = ( ~w8591 & w10579 ) | ( ~w8591 & w10585 ) | ( w10579 & w10585 ) ;
  assign w10592 = ~w10579 & w10591 ;
  assign w10593 = w10590 | w10592 ;
  assign w10594 = ( w8225 & w10587 ) | ( w8225 & ~w10593 ) | ( w10587 & ~w10593 ) ;
  assign w10595 = w8225 & w10594 ;
  assign w10596 = w10173 | w10178 ;
  assign w10597 = w10541 & ~w10596 ;
  assign w10598 = w10176 ^ w10597 ;
  assign w10599 = ( ~w8225 & w10587 ) | ( ~w8225 & w10593 ) | ( w10587 & w10593 ) ;
  assign w10600 = ~w10587 & w10599 ;
  assign w10601 = w10598 | w10600 ;
  assign w10602 = ( w7867 & w10595 ) | ( w7867 & ~w10601 ) | ( w10595 & ~w10601 ) ;
  assign w10603 = w7867 & w10602 ;
  assign w10604 = w10181 | w10186 ;
  assign w10605 = w10541 & ~w10604 ;
  assign w10606 = w10184 ^ w10605 ;
  assign w10607 = ( ~w7867 & w10595 ) | ( ~w7867 & w10601 ) | ( w10595 & w10601 ) ;
  assign w10608 = ~w10595 & w10607 ;
  assign w10609 = w10606 | w10608 ;
  assign w10610 = ( w7517 & w10603 ) | ( w7517 & ~w10609 ) | ( w10603 & ~w10609 ) ;
  assign w10611 = w7517 & w10610 ;
  assign w10612 = w10189 | w10194 ;
  assign w10613 = w10541 & ~w10612 ;
  assign w10614 = w10192 ^ w10613 ;
  assign w10615 = ( ~w7517 & w10603 ) | ( ~w7517 & w10609 ) | ( w10603 & w10609 ) ;
  assign w10616 = ~w10603 & w10615 ;
  assign w10617 = w10614 | w10616 ;
  assign w10618 = ( w7175 & w10611 ) | ( w7175 & ~w10617 ) | ( w10611 & ~w10617 ) ;
  assign w10619 = w7175 & w10618 ;
  assign w10620 = w10197 | w10202 ;
  assign w10621 = w10541 & ~w10620 ;
  assign w10622 = w10200 ^ w10621 ;
  assign w10623 = ( ~w7175 & w10611 ) | ( ~w7175 & w10617 ) | ( w10611 & w10617 ) ;
  assign w10624 = ~w10611 & w10623 ;
  assign w10625 = w10622 | w10624 ;
  assign w10626 = ( w6841 & w10619 ) | ( w6841 & ~w10625 ) | ( w10619 & ~w10625 ) ;
  assign w10627 = w6841 & w10626 ;
  assign w10628 = w10205 | w10210 ;
  assign w10629 = w10541 & ~w10628 ;
  assign w10630 = w10208 ^ w10629 ;
  assign w10631 = ( ~w6841 & w10619 ) | ( ~w6841 & w10625 ) | ( w10619 & w10625 ) ;
  assign w10632 = ~w10619 & w10631 ;
  assign w10633 = w10630 | w10632 ;
  assign w10634 = ( w6515 & w10627 ) | ( w6515 & ~w10633 ) | ( w10627 & ~w10633 ) ;
  assign w10635 = w6515 & w10634 ;
  assign w10636 = w10213 | w10218 ;
  assign w10637 = w10541 & ~w10636 ;
  assign w10638 = w10216 ^ w10637 ;
  assign w10639 = ( ~w6515 & w10627 ) | ( ~w6515 & w10633 ) | ( w10627 & w10633 ) ;
  assign w10640 = ~w10627 & w10639 ;
  assign w10641 = w10638 | w10640 ;
  assign w10642 = ( w6197 & w10635 ) | ( w6197 & ~w10641 ) | ( w10635 & ~w10641 ) ;
  assign w10643 = w6197 & w10642 ;
  assign w10644 = w10221 | w10226 ;
  assign w10645 = w10541 & ~w10644 ;
  assign w10646 = w10224 ^ w10645 ;
  assign w10647 = ( ~w6197 & w10635 ) | ( ~w6197 & w10641 ) | ( w10635 & w10641 ) ;
  assign w10648 = ~w10635 & w10647 ;
  assign w10649 = w10646 | w10648 ;
  assign w10650 = ( w5887 & w10643 ) | ( w5887 & ~w10649 ) | ( w10643 & ~w10649 ) ;
  assign w10651 = w5887 & w10650 ;
  assign w10652 = w10229 | w10234 ;
  assign w10653 = w10541 & ~w10652 ;
  assign w10654 = w10232 ^ w10653 ;
  assign w10655 = ( ~w5887 & w10643 ) | ( ~w5887 & w10649 ) | ( w10643 & w10649 ) ;
  assign w10656 = ~w10643 & w10655 ;
  assign w10657 = w10654 | w10656 ;
  assign w10658 = ( w5585 & w10651 ) | ( w5585 & ~w10657 ) | ( w10651 & ~w10657 ) ;
  assign w10659 = w5585 & w10658 ;
  assign w10660 = w10237 | w10242 ;
  assign w10661 = w10541 & ~w10660 ;
  assign w10662 = w10240 ^ w10661 ;
  assign w10663 = ( ~w5585 & w10651 ) | ( ~w5585 & w10657 ) | ( w10651 & w10657 ) ;
  assign w10664 = ~w10651 & w10663 ;
  assign w10665 = w10662 | w10664 ;
  assign w10666 = ( w5291 & w10659 ) | ( w5291 & ~w10665 ) | ( w10659 & ~w10665 ) ;
  assign w10667 = w5291 & w10666 ;
  assign w10668 = w10245 | w10250 ;
  assign w10669 = w10541 & ~w10668 ;
  assign w10670 = w10248 ^ w10669 ;
  assign w10671 = ( ~w5291 & w10659 ) | ( ~w5291 & w10665 ) | ( w10659 & w10665 ) ;
  assign w10672 = ~w10659 & w10671 ;
  assign w10673 = w10670 | w10672 ;
  assign w10674 = ( w5005 & w10667 ) | ( w5005 & ~w10673 ) | ( w10667 & ~w10673 ) ;
  assign w10675 = w5005 & w10674 ;
  assign w10676 = w10253 | w10258 ;
  assign w10677 = w10541 & ~w10676 ;
  assign w10678 = w10256 ^ w10677 ;
  assign w10679 = ( ~w5005 & w10667 ) | ( ~w5005 & w10673 ) | ( w10667 & w10673 ) ;
  assign w10680 = ~w10667 & w10679 ;
  assign w10681 = w10678 | w10680 ;
  assign w10682 = ( w4727 & w10675 ) | ( w4727 & ~w10681 ) | ( w10675 & ~w10681 ) ;
  assign w10683 = w4727 & w10682 ;
  assign w10684 = w10261 | w10266 ;
  assign w10685 = w10541 & ~w10684 ;
  assign w10686 = w10264 ^ w10685 ;
  assign w10687 = ( ~w4727 & w10675 ) | ( ~w4727 & w10681 ) | ( w10675 & w10681 ) ;
  assign w10688 = ~w10675 & w10687 ;
  assign w10689 = w10686 | w10688 ;
  assign w10690 = ( w4457 & w10683 ) | ( w4457 & ~w10689 ) | ( w10683 & ~w10689 ) ;
  assign w10691 = w4457 & w10690 ;
  assign w10692 = w10269 | w10274 ;
  assign w10693 = w10541 & ~w10692 ;
  assign w10694 = w10272 ^ w10693 ;
  assign w10695 = ( ~w4457 & w10683 ) | ( ~w4457 & w10689 ) | ( w10683 & w10689 ) ;
  assign w10696 = ~w10683 & w10695 ;
  assign w10697 = w10694 | w10696 ;
  assign w10698 = ( w4195 & w10691 ) | ( w4195 & ~w10697 ) | ( w10691 & ~w10697 ) ;
  assign w10699 = w4195 & w10698 ;
  assign w10700 = w10277 | w10282 ;
  assign w10701 = w10541 & ~w10700 ;
  assign w10702 = w10280 ^ w10701 ;
  assign w10703 = ( ~w4195 & w10691 ) | ( ~w4195 & w10697 ) | ( w10691 & w10697 ) ;
  assign w10704 = ~w10691 & w10703 ;
  assign w10705 = w10702 | w10704 ;
  assign w10706 = ( w3941 & w10699 ) | ( w3941 & ~w10705 ) | ( w10699 & ~w10705 ) ;
  assign w10707 = w3941 & w10706 ;
  assign w10708 = w10285 | w10290 ;
  assign w10709 = w10541 & ~w10708 ;
  assign w10710 = w10288 ^ w10709 ;
  assign w10711 = ( ~w3941 & w10699 ) | ( ~w3941 & w10705 ) | ( w10699 & w10705 ) ;
  assign w10712 = ~w10699 & w10711 ;
  assign w10713 = w10710 | w10712 ;
  assign w10714 = ( w3695 & w10707 ) | ( w3695 & ~w10713 ) | ( w10707 & ~w10713 ) ;
  assign w10715 = w3695 & w10714 ;
  assign w10716 = w10293 | w10298 ;
  assign w10717 = w10541 & ~w10716 ;
  assign w10718 = w10296 ^ w10717 ;
  assign w10719 = ( ~w3695 & w10707 ) | ( ~w3695 & w10713 ) | ( w10707 & w10713 ) ;
  assign w10720 = ~w10707 & w10719 ;
  assign w10721 = w10718 | w10720 ;
  assign w10722 = ( w3457 & w10715 ) | ( w3457 & ~w10721 ) | ( w10715 & ~w10721 ) ;
  assign w10723 = w3457 & w10722 ;
  assign w10724 = w10301 | w10306 ;
  assign w10725 = w10541 & ~w10724 ;
  assign w10726 = w10304 ^ w10725 ;
  assign w10727 = ( ~w3457 & w10715 ) | ( ~w3457 & w10721 ) | ( w10715 & w10721 ) ;
  assign w10728 = ~w10715 & w10727 ;
  assign w10729 = w10726 | w10728 ;
  assign w10730 = ( w3227 & w10723 ) | ( w3227 & ~w10729 ) | ( w10723 & ~w10729 ) ;
  assign w10731 = w3227 & w10730 ;
  assign w10732 = w10309 | w10314 ;
  assign w10733 = w10541 & ~w10732 ;
  assign w10734 = w10312 ^ w10733 ;
  assign w10735 = ( ~w3227 & w10723 ) | ( ~w3227 & w10729 ) | ( w10723 & w10729 ) ;
  assign w10736 = ~w10723 & w10735 ;
  assign w10737 = w10734 | w10736 ;
  assign w10738 = ( w3005 & w10731 ) | ( w3005 & ~w10737 ) | ( w10731 & ~w10737 ) ;
  assign w10739 = w3005 & w10738 ;
  assign w10740 = w10317 | w10322 ;
  assign w10741 = w10541 & ~w10740 ;
  assign w10742 = w10320 ^ w10741 ;
  assign w10743 = ( ~w3005 & w10731 ) | ( ~w3005 & w10737 ) | ( w10731 & w10737 ) ;
  assign w10744 = ~w10731 & w10743 ;
  assign w10745 = w10742 | w10744 ;
  assign w10746 = ( w2791 & w10739 ) | ( w2791 & ~w10745 ) | ( w10739 & ~w10745 ) ;
  assign w10747 = w2791 & w10746 ;
  assign w10748 = w10325 | w10330 ;
  assign w10749 = w10541 & ~w10748 ;
  assign w10750 = w10328 ^ w10749 ;
  assign w10751 = ( ~w2791 & w10739 ) | ( ~w2791 & w10745 ) | ( w10739 & w10745 ) ;
  assign w10752 = ~w10739 & w10751 ;
  assign w10753 = w10750 | w10752 ;
  assign w10754 = ( w2585 & w10747 ) | ( w2585 & ~w10753 ) | ( w10747 & ~w10753 ) ;
  assign w10755 = w2585 & w10754 ;
  assign w10756 = w10333 | w10338 ;
  assign w10757 = w10541 & ~w10756 ;
  assign w10758 = w10336 ^ w10757 ;
  assign w10759 = ( ~w2585 & w10747 ) | ( ~w2585 & w10753 ) | ( w10747 & w10753 ) ;
  assign w10760 = ~w10747 & w10759 ;
  assign w10761 = w10758 | w10760 ;
  assign w10762 = ( w2387 & w10755 ) | ( w2387 & ~w10761 ) | ( w10755 & ~w10761 ) ;
  assign w10763 = w2387 & w10762 ;
  assign w10764 = w10341 | w10346 ;
  assign w10765 = w10541 & ~w10764 ;
  assign w10766 = w10344 ^ w10765 ;
  assign w10767 = ( ~w2387 & w10755 ) | ( ~w2387 & w10761 ) | ( w10755 & w10761 ) ;
  assign w10768 = ~w10755 & w10767 ;
  assign w10769 = w10766 | w10768 ;
  assign w10770 = ( w2197 & w10763 ) | ( w2197 & ~w10769 ) | ( w10763 & ~w10769 ) ;
  assign w10771 = w2197 & w10770 ;
  assign w10772 = w10349 | w10354 ;
  assign w10773 = w10541 & ~w10772 ;
  assign w10774 = w10352 ^ w10773 ;
  assign w10775 = ( ~w2197 & w10763 ) | ( ~w2197 & w10769 ) | ( w10763 & w10769 ) ;
  assign w10776 = ~w10763 & w10775 ;
  assign w10777 = w10774 | w10776 ;
  assign w10778 = ( w2015 & w10771 ) | ( w2015 & ~w10777 ) | ( w10771 & ~w10777 ) ;
  assign w10779 = w2015 & w10778 ;
  assign w10780 = w10357 | w10362 ;
  assign w10781 = w10541 & ~w10780 ;
  assign w10782 = w10360 ^ w10781 ;
  assign w10783 = ( ~w2015 & w10771 ) | ( ~w2015 & w10777 ) | ( w10771 & w10777 ) ;
  assign w10784 = ~w10771 & w10783 ;
  assign w10785 = w10782 | w10784 ;
  assign w10786 = ( w1841 & w10779 ) | ( w1841 & ~w10785 ) | ( w10779 & ~w10785 ) ;
  assign w10787 = w1841 & w10786 ;
  assign w10788 = w10365 | w10370 ;
  assign w10789 = w10541 & ~w10788 ;
  assign w10790 = w10368 ^ w10789 ;
  assign w10791 = ( ~w1841 & w10779 ) | ( ~w1841 & w10785 ) | ( w10779 & w10785 ) ;
  assign w10792 = ~w10779 & w10791 ;
  assign w10793 = w10790 | w10792 ;
  assign w10794 = ( w1675 & w10787 ) | ( w1675 & ~w10793 ) | ( w10787 & ~w10793 ) ;
  assign w10795 = w1675 & w10794 ;
  assign w10796 = w10373 | w10378 ;
  assign w10797 = w10541 & ~w10796 ;
  assign w10798 = w10376 ^ w10797 ;
  assign w10799 = ( ~w1675 & w10787 ) | ( ~w1675 & w10793 ) | ( w10787 & w10793 ) ;
  assign w10800 = ~w10787 & w10799 ;
  assign w10801 = w10798 | w10800 ;
  assign w10802 = ( w1517 & w10795 ) | ( w1517 & ~w10801 ) | ( w10795 & ~w10801 ) ;
  assign w10803 = w1517 & w10802 ;
  assign w10804 = w10381 | w10386 ;
  assign w10805 = w10541 & ~w10804 ;
  assign w10806 = w10384 ^ w10805 ;
  assign w10807 = ( ~w1517 & w10795 ) | ( ~w1517 & w10801 ) | ( w10795 & w10801 ) ;
  assign w10808 = ~w10795 & w10807 ;
  assign w10809 = w10806 | w10808 ;
  assign w10810 = ( w1367 & w10803 ) | ( w1367 & ~w10809 ) | ( w10803 & ~w10809 ) ;
  assign w10811 = w1367 & w10810 ;
  assign w10812 = w10389 | w10394 ;
  assign w10813 = w10541 & ~w10812 ;
  assign w10814 = w10392 ^ w10813 ;
  assign w10815 = ( ~w1367 & w10803 ) | ( ~w1367 & w10809 ) | ( w10803 & w10809 ) ;
  assign w10816 = ~w10803 & w10815 ;
  assign w10817 = w10814 | w10816 ;
  assign w10818 = ( w1225 & w10811 ) | ( w1225 & ~w10817 ) | ( w10811 & ~w10817 ) ;
  assign w10819 = w1225 & w10818 ;
  assign w10820 = w10397 | w10402 ;
  assign w10821 = w10541 & ~w10820 ;
  assign w10822 = w10400 ^ w10821 ;
  assign w10823 = ( ~w1225 & w10811 ) | ( ~w1225 & w10817 ) | ( w10811 & w10817 ) ;
  assign w10824 = ~w10811 & w10823 ;
  assign w10825 = w10822 | w10824 ;
  assign w10826 = ( w1091 & w10819 ) | ( w1091 & ~w10825 ) | ( w10819 & ~w10825 ) ;
  assign w10827 = w1091 & w10826 ;
  assign w10828 = ( ~w1091 & w10819 ) | ( ~w1091 & w10825 ) | ( w10819 & w10825 ) ;
  assign w10829 = ~w10819 & w10828 ;
  assign w10830 = w10405 | w10407 ;
  assign w10831 = w10541 & ~w10830 ;
  assign w10832 = w10410 ^ w10831 ;
  assign w10833 = w10829 | w10832 ;
  assign w10834 = ( w965 & w10827 ) | ( w965 & ~w10833 ) | ( w10827 & ~w10833 ) ;
  assign w10835 = w965 & w10834 ;
  assign w10836 = w10413 | w10418 ;
  assign w10837 = w10541 & ~w10836 ;
  assign w10838 = w10416 ^ w10837 ;
  assign w10839 = ( ~w965 & w10827 ) | ( ~w965 & w10833 ) | ( w10827 & w10833 ) ;
  assign w10840 = ~w10827 & w10839 ;
  assign w10841 = w10838 | w10840 ;
  assign w10842 = ( w847 & w10835 ) | ( w847 & ~w10841 ) | ( w10835 & ~w10841 ) ;
  assign w10843 = w847 & w10842 ;
  assign w10844 = w10421 | w10426 ;
  assign w10845 = w10541 & ~w10844 ;
  assign w10846 = w10424 ^ w10845 ;
  assign w10847 = ( ~w847 & w10835 ) | ( ~w847 & w10841 ) | ( w10835 & w10841 ) ;
  assign w10848 = ~w10835 & w10847 ;
  assign w10849 = w10846 | w10848 ;
  assign w10850 = ( w737 & w10843 ) | ( w737 & ~w10849 ) | ( w10843 & ~w10849 ) ;
  assign w10851 = w737 & w10850 ;
  assign w10852 = w10429 | w10434 ;
  assign w10853 = w10541 & ~w10852 ;
  assign w10854 = w10432 ^ w10853 ;
  assign w10855 = ( ~w737 & w10843 ) | ( ~w737 & w10849 ) | ( w10843 & w10849 ) ;
  assign w10856 = ~w10843 & w10855 ;
  assign w10857 = w10854 | w10856 ;
  assign w10858 = ( w635 & w10851 ) | ( w635 & ~w10857 ) | ( w10851 & ~w10857 ) ;
  assign w10859 = w635 & w10858 ;
  assign w10860 = w10437 | w10442 ;
  assign w10861 = w10541 & ~w10860 ;
  assign w10862 = w10440 ^ w10861 ;
  assign w10863 = ( ~w635 & w10851 ) | ( ~w635 & w10857 ) | ( w10851 & w10857 ) ;
  assign w10864 = ~w10851 & w10863 ;
  assign w10865 = w10862 | w10864 ;
  assign w10866 = ( w541 & w10859 ) | ( w541 & ~w10865 ) | ( w10859 & ~w10865 ) ;
  assign w10867 = w541 & w10866 ;
  assign w10868 = w10445 | w10450 ;
  assign w10869 = w10541 & ~w10868 ;
  assign w10870 = w10448 ^ w10869 ;
  assign w10871 = ( ~w541 & w10859 ) | ( ~w541 & w10865 ) | ( w10859 & w10865 ) ;
  assign w10872 = ~w10859 & w10871 ;
  assign w10873 = w10870 | w10872 ;
  assign w10874 = ( w455 & w10867 ) | ( w455 & ~w10873 ) | ( w10867 & ~w10873 ) ;
  assign w10875 = w455 & w10874 ;
  assign w10876 = w10453 | w10458 ;
  assign w10877 = w10541 & ~w10876 ;
  assign w10878 = w10456 ^ w10877 ;
  assign w10879 = ( ~w455 & w10867 ) | ( ~w455 & w10873 ) | ( w10867 & w10873 ) ;
  assign w10880 = ~w10867 & w10879 ;
  assign w10881 = w10878 | w10880 ;
  assign w10882 = ( w377 & w10875 ) | ( w377 & ~w10881 ) | ( w10875 & ~w10881 ) ;
  assign w10883 = w377 & w10882 ;
  assign w10884 = w10461 | w10466 ;
  assign w10885 = w10541 & ~w10884 ;
  assign w10886 = w10464 ^ w10885 ;
  assign w10887 = ( ~w377 & w10875 ) | ( ~w377 & w10881 ) | ( w10875 & w10881 ) ;
  assign w10888 = ~w10875 & w10887 ;
  assign w10889 = w10886 | w10888 ;
  assign w10890 = ( w307 & w10883 ) | ( w307 & ~w10889 ) | ( w10883 & ~w10889 ) ;
  assign w10891 = w307 & w10890 ;
  assign w10892 = w10469 | w10474 ;
  assign w10893 = w10541 & ~w10892 ;
  assign w10894 = w10472 ^ w10893 ;
  assign w10895 = ( ~w307 & w10883 ) | ( ~w307 & w10889 ) | ( w10883 & w10889 ) ;
  assign w10896 = ~w10883 & w10895 ;
  assign w10897 = w10894 | w10896 ;
  assign w10898 = ( w246 & w10891 ) | ( w246 & ~w10897 ) | ( w10891 & ~w10897 ) ;
  assign w10899 = w246 & w10898 ;
  assign w10900 = w10477 | w10482 ;
  assign w10901 = w10541 & ~w10900 ;
  assign w10902 = w10480 ^ w10901 ;
  assign w10903 = ( ~w246 & w10891 ) | ( ~w246 & w10897 ) | ( w10891 & w10897 ) ;
  assign w10904 = ~w10891 & w10903 ;
  assign w10905 = w10902 | w10904 ;
  assign w10906 = ( w185 & w10899 ) | ( w185 & ~w10905 ) | ( w10899 & ~w10905 ) ;
  assign w10907 = w185 & w10906 ;
  assign w10908 = w10485 | w10490 ;
  assign w10909 = w10541 & ~w10908 ;
  assign w10910 = w10488 ^ w10909 ;
  assign w10911 = ( ~w185 & w10899 ) | ( ~w185 & w10905 ) | ( w10899 & w10905 ) ;
  assign w10912 = ~w10899 & w10911 ;
  assign w10913 = w10910 | w10912 ;
  assign w10914 = ( w145 & w10907 ) | ( w145 & ~w10913 ) | ( w10907 & ~w10913 ) ;
  assign w10915 = w145 & w10914 ;
  assign w10916 = w10493 | w10498 ;
  assign w10917 = w10541 & ~w10916 ;
  assign w10918 = w10496 ^ w10917 ;
  assign w10919 = ( ~w145 & w10907 ) | ( ~w145 & w10913 ) | ( w10907 & w10913 ) ;
  assign w10920 = ~w10907 & w10919 ;
  assign w10921 = w10918 | w10920 ;
  assign w10922 = ( w132 & w10915 ) | ( w132 & ~w10921 ) | ( w10915 & ~w10921 ) ;
  assign w10923 = w132 & w10922 ;
  assign w10924 = w10501 | w10506 ;
  assign w10925 = w10541 & ~w10924 ;
  assign w10926 = w10504 ^ w10925 ;
  assign w10927 = ( ~w132 & w10915 ) | ( ~w132 & w10921 ) | ( w10915 & w10921 ) ;
  assign w10928 = ~w10915 & w10927 ;
  assign w10929 = w10926 | w10928 ;
  assign w10930 = ~w10923 & w10929 ;
  assign w10931 = w10509 | w10514 ;
  assign w10932 = w10541 & ~w10931 ;
  assign w10933 = w10512 ^ w10932 ;
  assign w10934 = ( ~w10527 & w10930 ) | ( ~w10527 & w10933 ) | ( w10930 & w10933 ) ;
  assign w10935 = w10516 & ~w10934 ;
  assign w10936 = ~w10519 & w10541 ;
  assign w10937 = ( w10934 & ~w10935 ) | ( w10934 & w10936 ) | ( ~w10935 & w10936 ) ;
  assign w10938 = w10527 | w10937 ;
  assign w10939 = ~w129 & w10938 ;
  assign w10940 = ( w10923 & w10929 ) | ( w10923 & w10933 ) | ( w10929 & w10933 ) ;
  assign w10941 = ~w10923 & w10940 ;
  assign w10942 = ( w129 & w10516 ) | ( w129 & w10519 ) | ( w10516 & w10519 ) ;
  assign w10943 = ( w10519 & ~w10541 ) | ( w10519 & w10942 ) | ( ~w10541 & w10942 ) ;
  assign w10944 = w10516 & w10943 ;
  assign w10945 = w10942 ^ w10944 ;
  assign w10946 = ( w10103 & w10108 ) | ( w10103 & w10135 ) | ( w10108 & w10135 ) ;
  assign w10947 = w10135 & ~w10946 ;
  assign w10948 = w10106 ^ w10947 ;
  assign w10949 = ( ~w10531 & w10538 ) | ( ~w10531 & w10948 ) | ( w10538 & w10948 ) ;
  assign w10950 = ~w10538 & w10949 ;
  assign w10951 = ( ~w10525 & w10527 ) | ( ~w10525 & w10950 ) | ( w10527 & w10950 ) ;
  assign w10952 = ~w10527 & w10951 ;
  assign w10953 = w10941 | w10952 ;
  assign w10954 = ( w10939 & ~w10941 ) | ( w10939 & w10945 ) | ( ~w10941 & w10945 ) ;
  assign w10955 = w10953 | w10954 ;
  assign w10956 = ( ~\pi027 & \pi028 ) | ( ~\pi027 & w10541 ) | ( \pi028 & w10541 ) ;
  assign w10957 = ( ~\pi026 & \pi028 ) | ( ~\pi026 & w10956 ) | ( \pi028 & w10956 ) ;
  assign w10958 = ( ~\pi028 & w10541 ) | ( ~\pi028 & w10955 ) | ( w10541 & w10955 ) ;
  assign w10959 = w10957 & w10958 ;
  assign w10960 = ( w10527 & w10531 ) | ( w10527 & ~w10538 ) | ( w10531 & ~w10538 ) ;
  assign w10961 = \pi027 & ~w10960 ;
  assign w10962 = \pi026 | \pi028 ;
  assign w10963 = ( ~w10960 & w10961 ) | ( ~w10960 & w10962 ) | ( w10961 & w10962 ) ;
  assign w10964 = ~w10538 & w10963 ;
  assign w10965 = ~w10525 & w10964 ;
  assign w10966 = ( \pi028 & w10955 ) | ( \pi028 & ~w10964 ) | ( w10955 & ~w10964 ) ;
  assign w10967 = w10965 & ~w10966 ;
  assign w10968 = ~\pi028 & w10955 ;
  assign w10969 = \pi029 ^ w10968 ;
  assign w10970 = w10967 | w10969 ;
  assign w10971 = ( w10135 & w10959 ) | ( w10135 & ~w10970 ) | ( w10959 & ~w10970 ) ;
  assign w10972 = w10135 & w10971 ;
  assign w10973 = ( ~w10135 & w10959 ) | ( ~w10135 & w10970 ) | ( w10959 & w10970 ) ;
  assign w10974 = ~w10959 & w10973 ;
  assign w10975 = w10541 & ~w10952 ;
  assign w10976 = ~w10941 & w10975 ;
  assign w10977 = ~w10954 & w10976 ;
  assign w10978 = \pi029 & w10955 ;
  assign w10979 = ( \pi028 & w10955 ) | ( \pi028 & ~w10978 ) | ( w10955 & ~w10978 ) ;
  assign w10980 = ( ~\pi028 & w10977 ) | ( ~\pi028 & w10979 ) | ( w10977 & w10979 ) ;
  assign w10981 = \pi030 ^ w10980 ;
  assign w10982 = w10974 | w10981 ;
  assign w10983 = ( w9737 & w10972 ) | ( w9737 & ~w10982 ) | ( w10972 & ~w10982 ) ;
  assign w10984 = w9737 & w10983 ;
  assign w10985 = ( w10545 & ~w10553 ) | ( w10545 & w10955 ) | ( ~w10553 & w10955 ) ;
  assign w10986 = ~w10545 & w10985 ;
  assign w10987 = \pi031 ^ w10986 ;
  assign w10988 = w10554 ^ w10987 ;
  assign w10989 = ( ~w9737 & w10972 ) | ( ~w9737 & w10982 ) | ( w10972 & w10982 ) ;
  assign w10990 = ~w10972 & w10989 ;
  assign w10991 = w10988 | w10990 ;
  assign w10992 = ( w9347 & w10984 ) | ( w9347 & ~w10991 ) | ( w10984 & ~w10991 ) ;
  assign w10993 = w9347 & w10992 ;
  assign w10994 = w10558 | w10560 ;
  assign w10995 = w10955 & ~w10994 ;
  assign w10996 = w10567 ^ w10995 ;
  assign w10997 = ( ~w9347 & w10984 ) | ( ~w9347 & w10991 ) | ( w10984 & w10991 ) ;
  assign w10998 = ~w10984 & w10997 ;
  assign w10999 = w10996 | w10998 ;
  assign w11000 = ( w8965 & w10993 ) | ( w8965 & ~w10999 ) | ( w10993 & ~w10999 ) ;
  assign w11001 = w8965 & w11000 ;
  assign w11002 = w10570 | w10576 ;
  assign w11003 = w10955 & ~w11002 ;
  assign w11004 = w10574 ^ w11003 ;
  assign w11005 = ( ~w8965 & w10993 ) | ( ~w8965 & w10999 ) | ( w10993 & w10999 ) ;
  assign w11006 = ~w10993 & w11005 ;
  assign w11007 = w11004 | w11006 ;
  assign w11008 = ( w8591 & w11001 ) | ( w8591 & ~w11007 ) | ( w11001 & ~w11007 ) ;
  assign w11009 = w8591 & w11008 ;
  assign w11010 = w10579 | w10584 ;
  assign w11011 = w10955 & ~w11010 ;
  assign w11012 = w10582 ^ w11011 ;
  assign w11013 = ( ~w8591 & w11001 ) | ( ~w8591 & w11007 ) | ( w11001 & w11007 ) ;
  assign w11014 = ~w11001 & w11013 ;
  assign w11015 = w11012 | w11014 ;
  assign w11016 = ( w8225 & w11009 ) | ( w8225 & ~w11015 ) | ( w11009 & ~w11015 ) ;
  assign w11017 = w8225 & w11016 ;
  assign w11018 = w10587 | w10592 ;
  assign w11019 = w10955 & ~w11018 ;
  assign w11020 = w10590 ^ w11019 ;
  assign w11021 = ( ~w8225 & w11009 ) | ( ~w8225 & w11015 ) | ( w11009 & w11015 ) ;
  assign w11022 = ~w11009 & w11021 ;
  assign w11023 = w11020 | w11022 ;
  assign w11024 = ( w7867 & w11017 ) | ( w7867 & ~w11023 ) | ( w11017 & ~w11023 ) ;
  assign w11025 = w7867 & w11024 ;
  assign w11026 = w10595 | w10600 ;
  assign w11027 = w10955 & ~w11026 ;
  assign w11028 = w10598 ^ w11027 ;
  assign w11029 = ( ~w7867 & w11017 ) | ( ~w7867 & w11023 ) | ( w11017 & w11023 ) ;
  assign w11030 = ~w11017 & w11029 ;
  assign w11031 = w11028 | w11030 ;
  assign w11032 = ( w7517 & w11025 ) | ( w7517 & ~w11031 ) | ( w11025 & ~w11031 ) ;
  assign w11033 = w7517 & w11032 ;
  assign w11034 = w10603 | w10608 ;
  assign w11035 = w10955 & ~w11034 ;
  assign w11036 = w10606 ^ w11035 ;
  assign w11037 = ( ~w7517 & w11025 ) | ( ~w7517 & w11031 ) | ( w11025 & w11031 ) ;
  assign w11038 = ~w11025 & w11037 ;
  assign w11039 = w11036 | w11038 ;
  assign w11040 = ( w7175 & w11033 ) | ( w7175 & ~w11039 ) | ( w11033 & ~w11039 ) ;
  assign w11041 = w7175 & w11040 ;
  assign w11042 = w10611 | w10616 ;
  assign w11043 = w10955 & ~w11042 ;
  assign w11044 = w10614 ^ w11043 ;
  assign w11045 = ( ~w7175 & w11033 ) | ( ~w7175 & w11039 ) | ( w11033 & w11039 ) ;
  assign w11046 = ~w11033 & w11045 ;
  assign w11047 = w11044 | w11046 ;
  assign w11048 = ( w6841 & w11041 ) | ( w6841 & ~w11047 ) | ( w11041 & ~w11047 ) ;
  assign w11049 = w6841 & w11048 ;
  assign w11050 = w10619 | w10624 ;
  assign w11051 = w10955 & ~w11050 ;
  assign w11052 = w10622 ^ w11051 ;
  assign w11053 = ( ~w6841 & w11041 ) | ( ~w6841 & w11047 ) | ( w11041 & w11047 ) ;
  assign w11054 = ~w11041 & w11053 ;
  assign w11055 = w11052 | w11054 ;
  assign w11056 = ( w6515 & w11049 ) | ( w6515 & ~w11055 ) | ( w11049 & ~w11055 ) ;
  assign w11057 = w6515 & w11056 ;
  assign w11058 = w10627 | w10632 ;
  assign w11059 = w10955 & ~w11058 ;
  assign w11060 = w10630 ^ w11059 ;
  assign w11061 = ( ~w6515 & w11049 ) | ( ~w6515 & w11055 ) | ( w11049 & w11055 ) ;
  assign w11062 = ~w11049 & w11061 ;
  assign w11063 = w11060 | w11062 ;
  assign w11064 = ( w6197 & w11057 ) | ( w6197 & ~w11063 ) | ( w11057 & ~w11063 ) ;
  assign w11065 = w6197 & w11064 ;
  assign w11066 = w10635 | w10640 ;
  assign w11067 = w10955 & ~w11066 ;
  assign w11068 = w10638 ^ w11067 ;
  assign w11069 = ( ~w6197 & w11057 ) | ( ~w6197 & w11063 ) | ( w11057 & w11063 ) ;
  assign w11070 = ~w11057 & w11069 ;
  assign w11071 = w11068 | w11070 ;
  assign w11072 = ( w5887 & w11065 ) | ( w5887 & ~w11071 ) | ( w11065 & ~w11071 ) ;
  assign w11073 = w5887 & w11072 ;
  assign w11074 = w10643 | w10648 ;
  assign w11075 = w10955 & ~w11074 ;
  assign w11076 = w10646 ^ w11075 ;
  assign w11077 = ( ~w5887 & w11065 ) | ( ~w5887 & w11071 ) | ( w11065 & w11071 ) ;
  assign w11078 = ~w11065 & w11077 ;
  assign w11079 = w11076 | w11078 ;
  assign w11080 = ( w5585 & w11073 ) | ( w5585 & ~w11079 ) | ( w11073 & ~w11079 ) ;
  assign w11081 = w5585 & w11080 ;
  assign w11082 = w10651 | w10656 ;
  assign w11083 = w10955 & ~w11082 ;
  assign w11084 = w10654 ^ w11083 ;
  assign w11085 = ( ~w5585 & w11073 ) | ( ~w5585 & w11079 ) | ( w11073 & w11079 ) ;
  assign w11086 = ~w11073 & w11085 ;
  assign w11087 = w11084 | w11086 ;
  assign w11088 = ( w5291 & w11081 ) | ( w5291 & ~w11087 ) | ( w11081 & ~w11087 ) ;
  assign w11089 = w5291 & w11088 ;
  assign w11090 = w10659 | w10664 ;
  assign w11091 = w10955 & ~w11090 ;
  assign w11092 = w10662 ^ w11091 ;
  assign w11093 = ( ~w5291 & w11081 ) | ( ~w5291 & w11087 ) | ( w11081 & w11087 ) ;
  assign w11094 = ~w11081 & w11093 ;
  assign w11095 = w11092 | w11094 ;
  assign w11096 = ( w5005 & w11089 ) | ( w5005 & ~w11095 ) | ( w11089 & ~w11095 ) ;
  assign w11097 = w5005 & w11096 ;
  assign w11098 = w10667 | w10672 ;
  assign w11099 = w10955 & ~w11098 ;
  assign w11100 = w10670 ^ w11099 ;
  assign w11101 = ( ~w5005 & w11089 ) | ( ~w5005 & w11095 ) | ( w11089 & w11095 ) ;
  assign w11102 = ~w11089 & w11101 ;
  assign w11103 = w11100 | w11102 ;
  assign w11104 = ( w4727 & w11097 ) | ( w4727 & ~w11103 ) | ( w11097 & ~w11103 ) ;
  assign w11105 = w4727 & w11104 ;
  assign w11106 = w10675 | w10680 ;
  assign w11107 = w10955 & ~w11106 ;
  assign w11108 = w10678 ^ w11107 ;
  assign w11109 = ( ~w4727 & w11097 ) | ( ~w4727 & w11103 ) | ( w11097 & w11103 ) ;
  assign w11110 = ~w11097 & w11109 ;
  assign w11111 = w11108 | w11110 ;
  assign w11112 = ( w4457 & w11105 ) | ( w4457 & ~w11111 ) | ( w11105 & ~w11111 ) ;
  assign w11113 = w4457 & w11112 ;
  assign w11114 = w10683 | w10688 ;
  assign w11115 = w10955 & ~w11114 ;
  assign w11116 = w10686 ^ w11115 ;
  assign w11117 = ( ~w4457 & w11105 ) | ( ~w4457 & w11111 ) | ( w11105 & w11111 ) ;
  assign w11118 = ~w11105 & w11117 ;
  assign w11119 = w11116 | w11118 ;
  assign w11120 = ( w4195 & w11113 ) | ( w4195 & ~w11119 ) | ( w11113 & ~w11119 ) ;
  assign w11121 = w4195 & w11120 ;
  assign w11122 = w10691 | w10696 ;
  assign w11123 = w10955 & ~w11122 ;
  assign w11124 = w10694 ^ w11123 ;
  assign w11125 = ( ~w4195 & w11113 ) | ( ~w4195 & w11119 ) | ( w11113 & w11119 ) ;
  assign w11126 = ~w11113 & w11125 ;
  assign w11127 = w11124 | w11126 ;
  assign w11128 = ( w3941 & w11121 ) | ( w3941 & ~w11127 ) | ( w11121 & ~w11127 ) ;
  assign w11129 = w3941 & w11128 ;
  assign w11130 = w10699 | w10704 ;
  assign w11131 = w10955 & ~w11130 ;
  assign w11132 = w10702 ^ w11131 ;
  assign w11133 = ( ~w3941 & w11121 ) | ( ~w3941 & w11127 ) | ( w11121 & w11127 ) ;
  assign w11134 = ~w11121 & w11133 ;
  assign w11135 = w11132 | w11134 ;
  assign w11136 = ( w3695 & w11129 ) | ( w3695 & ~w11135 ) | ( w11129 & ~w11135 ) ;
  assign w11137 = w3695 & w11136 ;
  assign w11138 = w10707 | w10712 ;
  assign w11139 = w10955 & ~w11138 ;
  assign w11140 = w10710 ^ w11139 ;
  assign w11141 = ( ~w3695 & w11129 ) | ( ~w3695 & w11135 ) | ( w11129 & w11135 ) ;
  assign w11142 = ~w11129 & w11141 ;
  assign w11143 = w11140 | w11142 ;
  assign w11144 = ( w3457 & w11137 ) | ( w3457 & ~w11143 ) | ( w11137 & ~w11143 ) ;
  assign w11145 = w3457 & w11144 ;
  assign w11146 = w10715 | w10720 ;
  assign w11147 = w10955 & ~w11146 ;
  assign w11148 = w10718 ^ w11147 ;
  assign w11149 = ( ~w3457 & w11137 ) | ( ~w3457 & w11143 ) | ( w11137 & w11143 ) ;
  assign w11150 = ~w11137 & w11149 ;
  assign w11151 = w11148 | w11150 ;
  assign w11152 = ( w3227 & w11145 ) | ( w3227 & ~w11151 ) | ( w11145 & ~w11151 ) ;
  assign w11153 = w3227 & w11152 ;
  assign w11154 = w10723 | w10728 ;
  assign w11155 = w10955 & ~w11154 ;
  assign w11156 = w10726 ^ w11155 ;
  assign w11157 = ( ~w3227 & w11145 ) | ( ~w3227 & w11151 ) | ( w11145 & w11151 ) ;
  assign w11158 = ~w11145 & w11157 ;
  assign w11159 = w11156 | w11158 ;
  assign w11160 = ( w3005 & w11153 ) | ( w3005 & ~w11159 ) | ( w11153 & ~w11159 ) ;
  assign w11161 = w3005 & w11160 ;
  assign w11162 = w10731 | w10736 ;
  assign w11163 = w10955 & ~w11162 ;
  assign w11164 = w10734 ^ w11163 ;
  assign w11165 = ( ~w3005 & w11153 ) | ( ~w3005 & w11159 ) | ( w11153 & w11159 ) ;
  assign w11166 = ~w11153 & w11165 ;
  assign w11167 = w11164 | w11166 ;
  assign w11168 = ( w2791 & w11161 ) | ( w2791 & ~w11167 ) | ( w11161 & ~w11167 ) ;
  assign w11169 = w2791 & w11168 ;
  assign w11170 = w10739 | w10744 ;
  assign w11171 = w10955 & ~w11170 ;
  assign w11172 = w10742 ^ w11171 ;
  assign w11173 = ( ~w2791 & w11161 ) | ( ~w2791 & w11167 ) | ( w11161 & w11167 ) ;
  assign w11174 = ~w11161 & w11173 ;
  assign w11175 = w11172 | w11174 ;
  assign w11176 = ( w2585 & w11169 ) | ( w2585 & ~w11175 ) | ( w11169 & ~w11175 ) ;
  assign w11177 = w2585 & w11176 ;
  assign w11178 = w10747 | w10752 ;
  assign w11179 = w10955 & ~w11178 ;
  assign w11180 = w10750 ^ w11179 ;
  assign w11181 = ( ~w2585 & w11169 ) | ( ~w2585 & w11175 ) | ( w11169 & w11175 ) ;
  assign w11182 = ~w11169 & w11181 ;
  assign w11183 = w11180 | w11182 ;
  assign w11184 = ( w2387 & w11177 ) | ( w2387 & ~w11183 ) | ( w11177 & ~w11183 ) ;
  assign w11185 = w2387 & w11184 ;
  assign w11186 = w10755 | w10760 ;
  assign w11187 = w10955 & ~w11186 ;
  assign w11188 = w10758 ^ w11187 ;
  assign w11189 = ( ~w2387 & w11177 ) | ( ~w2387 & w11183 ) | ( w11177 & w11183 ) ;
  assign w11190 = ~w11177 & w11189 ;
  assign w11191 = w11188 | w11190 ;
  assign w11192 = ( w2197 & w11185 ) | ( w2197 & ~w11191 ) | ( w11185 & ~w11191 ) ;
  assign w11193 = w2197 & w11192 ;
  assign w11194 = w10763 | w10768 ;
  assign w11195 = w10955 & ~w11194 ;
  assign w11196 = w10766 ^ w11195 ;
  assign w11197 = ( ~w2197 & w11185 ) | ( ~w2197 & w11191 ) | ( w11185 & w11191 ) ;
  assign w11198 = ~w11185 & w11197 ;
  assign w11199 = w11196 | w11198 ;
  assign w11200 = ( w2015 & w11193 ) | ( w2015 & ~w11199 ) | ( w11193 & ~w11199 ) ;
  assign w11201 = w2015 & w11200 ;
  assign w11202 = w10771 | w10776 ;
  assign w11203 = w10955 & ~w11202 ;
  assign w11204 = w10774 ^ w11203 ;
  assign w11205 = ( ~w2015 & w11193 ) | ( ~w2015 & w11199 ) | ( w11193 & w11199 ) ;
  assign w11206 = ~w11193 & w11205 ;
  assign w11207 = w11204 | w11206 ;
  assign w11208 = ( w1841 & w11201 ) | ( w1841 & ~w11207 ) | ( w11201 & ~w11207 ) ;
  assign w11209 = w1841 & w11208 ;
  assign w11210 = w10779 | w10784 ;
  assign w11211 = w10955 & ~w11210 ;
  assign w11212 = w10782 ^ w11211 ;
  assign w11213 = ( ~w1841 & w11201 ) | ( ~w1841 & w11207 ) | ( w11201 & w11207 ) ;
  assign w11214 = ~w11201 & w11213 ;
  assign w11215 = w11212 | w11214 ;
  assign w11216 = ( w1675 & w11209 ) | ( w1675 & ~w11215 ) | ( w11209 & ~w11215 ) ;
  assign w11217 = w1675 & w11216 ;
  assign w11218 = w10787 | w10792 ;
  assign w11219 = w10955 & ~w11218 ;
  assign w11220 = w10790 ^ w11219 ;
  assign w11221 = ( ~w1675 & w11209 ) | ( ~w1675 & w11215 ) | ( w11209 & w11215 ) ;
  assign w11222 = ~w11209 & w11221 ;
  assign w11223 = w11220 | w11222 ;
  assign w11224 = ( w1517 & w11217 ) | ( w1517 & ~w11223 ) | ( w11217 & ~w11223 ) ;
  assign w11225 = w1517 & w11224 ;
  assign w11226 = w10795 | w10800 ;
  assign w11227 = w10955 & ~w11226 ;
  assign w11228 = w10798 ^ w11227 ;
  assign w11229 = ( ~w1517 & w11217 ) | ( ~w1517 & w11223 ) | ( w11217 & w11223 ) ;
  assign w11230 = ~w11217 & w11229 ;
  assign w11231 = w11228 | w11230 ;
  assign w11232 = ( w1367 & w11225 ) | ( w1367 & ~w11231 ) | ( w11225 & ~w11231 ) ;
  assign w11233 = w1367 & w11232 ;
  assign w11234 = w10803 | w10808 ;
  assign w11235 = w10955 & ~w11234 ;
  assign w11236 = w10806 ^ w11235 ;
  assign w11237 = ( ~w1367 & w11225 ) | ( ~w1367 & w11231 ) | ( w11225 & w11231 ) ;
  assign w11238 = ~w11225 & w11237 ;
  assign w11239 = w11236 | w11238 ;
  assign w11240 = ( w1225 & w11233 ) | ( w1225 & ~w11239 ) | ( w11233 & ~w11239 ) ;
  assign w11241 = w1225 & w11240 ;
  assign w11242 = w10811 | w10816 ;
  assign w11243 = w10955 & ~w11242 ;
  assign w11244 = w10814 ^ w11243 ;
  assign w11245 = ( ~w1225 & w11233 ) | ( ~w1225 & w11239 ) | ( w11233 & w11239 ) ;
  assign w11246 = ~w11233 & w11245 ;
  assign w11247 = w11244 | w11246 ;
  assign w11248 = ( w1091 & w11241 ) | ( w1091 & ~w11247 ) | ( w11241 & ~w11247 ) ;
  assign w11249 = w1091 & w11248 ;
  assign w11250 = w10819 | w10824 ;
  assign w11251 = w10955 & ~w11250 ;
  assign w11252 = w10822 ^ w11251 ;
  assign w11253 = ( ~w1091 & w11241 ) | ( ~w1091 & w11247 ) | ( w11241 & w11247 ) ;
  assign w11254 = ~w11241 & w11253 ;
  assign w11255 = w11252 | w11254 ;
  assign w11256 = ( w965 & w11249 ) | ( w965 & ~w11255 ) | ( w11249 & ~w11255 ) ;
  assign w11257 = w965 & w11256 ;
  assign w11258 = ( ~w965 & w11249 ) | ( ~w965 & w11255 ) | ( w11249 & w11255 ) ;
  assign w11259 = ~w11249 & w11258 ;
  assign w11260 = w10827 | w10829 ;
  assign w11261 = w10955 & ~w11260 ;
  assign w11262 = w10832 ^ w11261 ;
  assign w11263 = w11259 | w11262 ;
  assign w11264 = ( w847 & w11257 ) | ( w847 & ~w11263 ) | ( w11257 & ~w11263 ) ;
  assign w11265 = w847 & w11264 ;
  assign w11266 = w10835 | w10840 ;
  assign w11267 = w10955 & ~w11266 ;
  assign w11268 = w10838 ^ w11267 ;
  assign w11269 = ( ~w847 & w11257 ) | ( ~w847 & w11263 ) | ( w11257 & w11263 ) ;
  assign w11270 = ~w11257 & w11269 ;
  assign w11271 = w11268 | w11270 ;
  assign w11272 = ( w737 & w11265 ) | ( w737 & ~w11271 ) | ( w11265 & ~w11271 ) ;
  assign w11273 = w737 & w11272 ;
  assign w11274 = w10843 | w10848 ;
  assign w11275 = w10955 & ~w11274 ;
  assign w11276 = w10846 ^ w11275 ;
  assign w11277 = ( ~w737 & w11265 ) | ( ~w737 & w11271 ) | ( w11265 & w11271 ) ;
  assign w11278 = ~w11265 & w11277 ;
  assign w11279 = w11276 | w11278 ;
  assign w11280 = ( w635 & w11273 ) | ( w635 & ~w11279 ) | ( w11273 & ~w11279 ) ;
  assign w11281 = w635 & w11280 ;
  assign w11282 = w10851 | w10856 ;
  assign w11283 = w10955 & ~w11282 ;
  assign w11284 = w10854 ^ w11283 ;
  assign w11285 = ( ~w635 & w11273 ) | ( ~w635 & w11279 ) | ( w11273 & w11279 ) ;
  assign w11286 = ~w11273 & w11285 ;
  assign w11287 = w11284 | w11286 ;
  assign w11288 = ( w541 & w11281 ) | ( w541 & ~w11287 ) | ( w11281 & ~w11287 ) ;
  assign w11289 = w541 & w11288 ;
  assign w11290 = w10859 | w10864 ;
  assign w11291 = w10955 & ~w11290 ;
  assign w11292 = w10862 ^ w11291 ;
  assign w11293 = ( ~w541 & w11281 ) | ( ~w541 & w11287 ) | ( w11281 & w11287 ) ;
  assign w11294 = ~w11281 & w11293 ;
  assign w11295 = w11292 | w11294 ;
  assign w11296 = ( w455 & w11289 ) | ( w455 & ~w11295 ) | ( w11289 & ~w11295 ) ;
  assign w11297 = w455 & w11296 ;
  assign w11298 = w10867 | w10872 ;
  assign w11299 = w10955 & ~w11298 ;
  assign w11300 = w10870 ^ w11299 ;
  assign w11301 = ( ~w455 & w11289 ) | ( ~w455 & w11295 ) | ( w11289 & w11295 ) ;
  assign w11302 = ~w11289 & w11301 ;
  assign w11303 = w11300 | w11302 ;
  assign w11304 = ( w377 & w11297 ) | ( w377 & ~w11303 ) | ( w11297 & ~w11303 ) ;
  assign w11305 = w377 & w11304 ;
  assign w11306 = w10875 | w10880 ;
  assign w11307 = w10955 & ~w11306 ;
  assign w11308 = w10878 ^ w11307 ;
  assign w11309 = ( ~w377 & w11297 ) | ( ~w377 & w11303 ) | ( w11297 & w11303 ) ;
  assign w11310 = ~w11297 & w11309 ;
  assign w11311 = w11308 | w11310 ;
  assign w11312 = ( w307 & w11305 ) | ( w307 & ~w11311 ) | ( w11305 & ~w11311 ) ;
  assign w11313 = w307 & w11312 ;
  assign w11314 = w10883 | w10888 ;
  assign w11315 = w10955 & ~w11314 ;
  assign w11316 = w10886 ^ w11315 ;
  assign w11317 = ( ~w307 & w11305 ) | ( ~w307 & w11311 ) | ( w11305 & w11311 ) ;
  assign w11318 = ~w11305 & w11317 ;
  assign w11319 = w11316 | w11318 ;
  assign w11320 = ( w246 & w11313 ) | ( w246 & ~w11319 ) | ( w11313 & ~w11319 ) ;
  assign w11321 = w246 & w11320 ;
  assign w11322 = w10891 | w10896 ;
  assign w11323 = w10955 & ~w11322 ;
  assign w11324 = w10894 ^ w11323 ;
  assign w11325 = ( ~w246 & w11313 ) | ( ~w246 & w11319 ) | ( w11313 & w11319 ) ;
  assign w11326 = ~w11313 & w11325 ;
  assign w11327 = w11324 | w11326 ;
  assign w11328 = ( w185 & w11321 ) | ( w185 & ~w11327 ) | ( w11321 & ~w11327 ) ;
  assign w11329 = w185 & w11328 ;
  assign w11330 = w10899 | w10904 ;
  assign w11331 = w10955 & ~w11330 ;
  assign w11332 = w10902 ^ w11331 ;
  assign w11333 = ( ~w185 & w11321 ) | ( ~w185 & w11327 ) | ( w11321 & w11327 ) ;
  assign w11334 = ~w11321 & w11333 ;
  assign w11335 = w11332 | w11334 ;
  assign w11336 = ( w145 & w11329 ) | ( w145 & ~w11335 ) | ( w11329 & ~w11335 ) ;
  assign w11337 = w145 & w11336 ;
  assign w11338 = w10907 | w10912 ;
  assign w11339 = w10955 & ~w11338 ;
  assign w11340 = w10910 ^ w11339 ;
  assign w11341 = ( ~w145 & w11329 ) | ( ~w145 & w11335 ) | ( w11329 & w11335 ) ;
  assign w11342 = ~w11329 & w11341 ;
  assign w11343 = w11340 | w11342 ;
  assign w11344 = ( w132 & w11337 ) | ( w132 & ~w11343 ) | ( w11337 & ~w11343 ) ;
  assign w11345 = w132 & w11344 ;
  assign w11346 = w10915 | w10920 ;
  assign w11347 = w10955 & ~w11346 ;
  assign w11348 = w10918 ^ w11347 ;
  assign w11349 = ( ~w132 & w11337 ) | ( ~w132 & w11343 ) | ( w11337 & w11343 ) ;
  assign w11350 = ~w11337 & w11349 ;
  assign w11351 = w11348 | w11350 ;
  assign w11352 = ~w11345 & w11351 ;
  assign w11353 = w10923 | w10928 ;
  assign w11354 = w10955 & ~w11353 ;
  assign w11355 = w10926 ^ w11354 ;
  assign w11356 = ( ~w10941 & w11352 ) | ( ~w10941 & w11355 ) | ( w11352 & w11355 ) ;
  assign w11357 = w10930 & ~w11356 ;
  assign w11358 = ~w10933 & w10955 ;
  assign w11359 = ( w11356 & ~w11357 ) | ( w11356 & w11358 ) | ( ~w11357 & w11358 ) ;
  assign w11360 = w10941 | w11359 ;
  assign w11361 = ~w129 & w11360 ;
  assign w11362 = ( w11345 & w11351 ) | ( w11345 & w11355 ) | ( w11351 & w11355 ) ;
  assign w11363 = ~w11345 & w11362 ;
  assign w11364 = ( w129 & w10930 ) | ( w129 & w10933 ) | ( w10930 & w10933 ) ;
  assign w11365 = ( w10933 & ~w10955 ) | ( w10933 & w11364 ) | ( ~w10955 & w11364 ) ;
  assign w11366 = w10930 & w11365 ;
  assign w11367 = w11364 ^ w11366 ;
  assign w11368 = ( w10509 & w10514 ) | ( w10509 & w10541 ) | ( w10514 & w10541 ) ;
  assign w11369 = w10541 & ~w11368 ;
  assign w11370 = w10512 ^ w11369 ;
  assign w11371 = ( ~w10945 & w10952 ) | ( ~w10945 & w11370 ) | ( w10952 & w11370 ) ;
  assign w11372 = ~w10952 & w11371 ;
  assign w11373 = ( ~w10939 & w10941 ) | ( ~w10939 & w11372 ) | ( w10941 & w11372 ) ;
  assign w11374 = ~w10941 & w11373 ;
  assign w11375 = w11363 | w11374 ;
  assign w11376 = ( w11361 & ~w11363 ) | ( w11361 & w11367 ) | ( ~w11363 & w11367 ) ;
  assign w11377 = w11375 | w11376 ;
  assign w11378 = ( ~\pi025 & \pi026 ) | ( ~\pi025 & w10955 ) | ( \pi026 & w10955 ) ;
  assign w11379 = ( ~\pi024 & \pi026 ) | ( ~\pi024 & w11378 ) | ( \pi026 & w11378 ) ;
  assign w11380 = ( ~\pi026 & w10955 ) | ( ~\pi026 & w11377 ) | ( w10955 & w11377 ) ;
  assign w11381 = w11379 & w11380 ;
  assign w11382 = ( w10941 & w10945 ) | ( w10941 & ~w10952 ) | ( w10945 & ~w10952 ) ;
  assign w11383 = \pi025 & ~w11382 ;
  assign w11384 = \pi024 | \pi026 ;
  assign w11385 = ( ~w11382 & w11383 ) | ( ~w11382 & w11384 ) | ( w11383 & w11384 ) ;
  assign w11386 = ~w10952 & w11385 ;
  assign w11387 = ~w10939 & w11386 ;
  assign w11388 = ( \pi026 & w11377 ) | ( \pi026 & ~w11386 ) | ( w11377 & ~w11386 ) ;
  assign w11389 = w11387 & ~w11388 ;
  assign w11390 = ~\pi026 & w11377 ;
  assign w11391 = \pi027 ^ w11390 ;
  assign w11392 = w11389 | w11391 ;
  assign w11393 = ( w10541 & w11381 ) | ( w10541 & ~w11392 ) | ( w11381 & ~w11392 ) ;
  assign w11394 = w10541 & w11393 ;
  assign w11395 = ( ~w10541 & w11381 ) | ( ~w10541 & w11392 ) | ( w11381 & w11392 ) ;
  assign w11396 = ~w11381 & w11395 ;
  assign w11397 = w10955 & ~w11374 ;
  assign w11398 = ~w11363 & w11397 ;
  assign w11399 = ~w11376 & w11398 ;
  assign w11400 = \pi027 & w11377 ;
  assign w11401 = ( \pi026 & w11377 ) | ( \pi026 & ~w11400 ) | ( w11377 & ~w11400 ) ;
  assign w11402 = ( ~\pi026 & w11399 ) | ( ~\pi026 & w11401 ) | ( w11399 & w11401 ) ;
  assign w11403 = \pi028 ^ w11402 ;
  assign w11404 = w11396 | w11403 ;
  assign w11405 = ( w10135 & w11394 ) | ( w10135 & ~w11404 ) | ( w11394 & ~w11404 ) ;
  assign w11406 = w10135 & w11405 ;
  assign w11407 = ( w10959 & ~w10967 ) | ( w10959 & w11377 ) | ( ~w10967 & w11377 ) ;
  assign w11408 = ~w10959 & w11407 ;
  assign w11409 = \pi029 ^ w11408 ;
  assign w11410 = w10968 ^ w11409 ;
  assign w11411 = ( ~w10135 & w11394 ) | ( ~w10135 & w11404 ) | ( w11394 & w11404 ) ;
  assign w11412 = ~w11394 & w11411 ;
  assign w11413 = w11410 | w11412 ;
  assign w11414 = ( w9737 & w11406 ) | ( w9737 & ~w11413 ) | ( w11406 & ~w11413 ) ;
  assign w11415 = w9737 & w11414 ;
  assign w11416 = w10972 | w10974 ;
  assign w11417 = w11377 & ~w11416 ;
  assign w11418 = w10981 ^ w11417 ;
  assign w11419 = ( ~w9737 & w11406 ) | ( ~w9737 & w11413 ) | ( w11406 & w11413 ) ;
  assign w11420 = ~w11406 & w11419 ;
  assign w11421 = w11418 | w11420 ;
  assign w11422 = ( w9347 & w11415 ) | ( w9347 & ~w11421 ) | ( w11415 & ~w11421 ) ;
  assign w11423 = w9347 & w11422 ;
  assign w11424 = w10984 | w10990 ;
  assign w11425 = w11377 & ~w11424 ;
  assign w11426 = w10988 ^ w11425 ;
  assign w11427 = ( ~w9347 & w11415 ) | ( ~w9347 & w11421 ) | ( w11415 & w11421 ) ;
  assign w11428 = ~w11415 & w11427 ;
  assign w11429 = w11426 | w11428 ;
  assign w11430 = ( w8965 & w11423 ) | ( w8965 & ~w11429 ) | ( w11423 & ~w11429 ) ;
  assign w11431 = w8965 & w11430 ;
  assign w11432 = w10993 | w10998 ;
  assign w11433 = w11377 & ~w11432 ;
  assign w11434 = w10996 ^ w11433 ;
  assign w11435 = ( ~w8965 & w11423 ) | ( ~w8965 & w11429 ) | ( w11423 & w11429 ) ;
  assign w11436 = ~w11423 & w11435 ;
  assign w11437 = w11434 | w11436 ;
  assign w11438 = ( w8591 & w11431 ) | ( w8591 & ~w11437 ) | ( w11431 & ~w11437 ) ;
  assign w11439 = w8591 & w11438 ;
  assign w11440 = w11001 | w11006 ;
  assign w11441 = w11377 & ~w11440 ;
  assign w11442 = w11004 ^ w11441 ;
  assign w11443 = ( ~w8591 & w11431 ) | ( ~w8591 & w11437 ) | ( w11431 & w11437 ) ;
  assign w11444 = ~w11431 & w11443 ;
  assign w11445 = w11442 | w11444 ;
  assign w11446 = ( w8225 & w11439 ) | ( w8225 & ~w11445 ) | ( w11439 & ~w11445 ) ;
  assign w11447 = w8225 & w11446 ;
  assign w11448 = w11009 | w11014 ;
  assign w11449 = w11377 & ~w11448 ;
  assign w11450 = w11012 ^ w11449 ;
  assign w11451 = ( ~w8225 & w11439 ) | ( ~w8225 & w11445 ) | ( w11439 & w11445 ) ;
  assign w11452 = ~w11439 & w11451 ;
  assign w11453 = w11450 | w11452 ;
  assign w11454 = ( w7867 & w11447 ) | ( w7867 & ~w11453 ) | ( w11447 & ~w11453 ) ;
  assign w11455 = w7867 & w11454 ;
  assign w11456 = w11017 | w11022 ;
  assign w11457 = w11377 & ~w11456 ;
  assign w11458 = w11020 ^ w11457 ;
  assign w11459 = ( ~w7867 & w11447 ) | ( ~w7867 & w11453 ) | ( w11447 & w11453 ) ;
  assign w11460 = ~w11447 & w11459 ;
  assign w11461 = w11458 | w11460 ;
  assign w11462 = ( w7517 & w11455 ) | ( w7517 & ~w11461 ) | ( w11455 & ~w11461 ) ;
  assign w11463 = w7517 & w11462 ;
  assign w11464 = w11025 | w11030 ;
  assign w11465 = w11377 & ~w11464 ;
  assign w11466 = w11028 ^ w11465 ;
  assign w11467 = ( ~w7517 & w11455 ) | ( ~w7517 & w11461 ) | ( w11455 & w11461 ) ;
  assign w11468 = ~w11455 & w11467 ;
  assign w11469 = w11466 | w11468 ;
  assign w11470 = ( w7175 & w11463 ) | ( w7175 & ~w11469 ) | ( w11463 & ~w11469 ) ;
  assign w11471 = w7175 & w11470 ;
  assign w11472 = w11033 | w11038 ;
  assign w11473 = w11377 & ~w11472 ;
  assign w11474 = w11036 ^ w11473 ;
  assign w11475 = ( ~w7175 & w11463 ) | ( ~w7175 & w11469 ) | ( w11463 & w11469 ) ;
  assign w11476 = ~w11463 & w11475 ;
  assign w11477 = w11474 | w11476 ;
  assign w11478 = ( w6841 & w11471 ) | ( w6841 & ~w11477 ) | ( w11471 & ~w11477 ) ;
  assign w11479 = w6841 & w11478 ;
  assign w11480 = w11041 | w11046 ;
  assign w11481 = w11377 & ~w11480 ;
  assign w11482 = w11044 ^ w11481 ;
  assign w11483 = ( ~w6841 & w11471 ) | ( ~w6841 & w11477 ) | ( w11471 & w11477 ) ;
  assign w11484 = ~w11471 & w11483 ;
  assign w11485 = w11482 | w11484 ;
  assign w11486 = ( w6515 & w11479 ) | ( w6515 & ~w11485 ) | ( w11479 & ~w11485 ) ;
  assign w11487 = w6515 & w11486 ;
  assign w11488 = w11049 | w11054 ;
  assign w11489 = w11377 & ~w11488 ;
  assign w11490 = w11052 ^ w11489 ;
  assign w11491 = ( ~w6515 & w11479 ) | ( ~w6515 & w11485 ) | ( w11479 & w11485 ) ;
  assign w11492 = ~w11479 & w11491 ;
  assign w11493 = w11490 | w11492 ;
  assign w11494 = ( w6197 & w11487 ) | ( w6197 & ~w11493 ) | ( w11487 & ~w11493 ) ;
  assign w11495 = w6197 & w11494 ;
  assign w11496 = w11057 | w11062 ;
  assign w11497 = w11377 & ~w11496 ;
  assign w11498 = w11060 ^ w11497 ;
  assign w11499 = ( ~w6197 & w11487 ) | ( ~w6197 & w11493 ) | ( w11487 & w11493 ) ;
  assign w11500 = ~w11487 & w11499 ;
  assign w11501 = w11498 | w11500 ;
  assign w11502 = ( w5887 & w11495 ) | ( w5887 & ~w11501 ) | ( w11495 & ~w11501 ) ;
  assign w11503 = w5887 & w11502 ;
  assign w11504 = w11065 | w11070 ;
  assign w11505 = w11377 & ~w11504 ;
  assign w11506 = w11068 ^ w11505 ;
  assign w11507 = ( ~w5887 & w11495 ) | ( ~w5887 & w11501 ) | ( w11495 & w11501 ) ;
  assign w11508 = ~w11495 & w11507 ;
  assign w11509 = w11506 | w11508 ;
  assign w11510 = ( w5585 & w11503 ) | ( w5585 & ~w11509 ) | ( w11503 & ~w11509 ) ;
  assign w11511 = w5585 & w11510 ;
  assign w11512 = w11073 | w11078 ;
  assign w11513 = w11377 & ~w11512 ;
  assign w11514 = w11076 ^ w11513 ;
  assign w11515 = ( ~w5585 & w11503 ) | ( ~w5585 & w11509 ) | ( w11503 & w11509 ) ;
  assign w11516 = ~w11503 & w11515 ;
  assign w11517 = w11514 | w11516 ;
  assign w11518 = ( w5291 & w11511 ) | ( w5291 & ~w11517 ) | ( w11511 & ~w11517 ) ;
  assign w11519 = w5291 & w11518 ;
  assign w11520 = w11081 | w11086 ;
  assign w11521 = w11377 & ~w11520 ;
  assign w11522 = w11084 ^ w11521 ;
  assign w11523 = ( ~w5291 & w11511 ) | ( ~w5291 & w11517 ) | ( w11511 & w11517 ) ;
  assign w11524 = ~w11511 & w11523 ;
  assign w11525 = w11522 | w11524 ;
  assign w11526 = ( w5005 & w11519 ) | ( w5005 & ~w11525 ) | ( w11519 & ~w11525 ) ;
  assign w11527 = w5005 & w11526 ;
  assign w11528 = w11089 | w11094 ;
  assign w11529 = w11377 & ~w11528 ;
  assign w11530 = w11092 ^ w11529 ;
  assign w11531 = ( ~w5005 & w11519 ) | ( ~w5005 & w11525 ) | ( w11519 & w11525 ) ;
  assign w11532 = ~w11519 & w11531 ;
  assign w11533 = w11530 | w11532 ;
  assign w11534 = ( w4727 & w11527 ) | ( w4727 & ~w11533 ) | ( w11527 & ~w11533 ) ;
  assign w11535 = w4727 & w11534 ;
  assign w11536 = w11097 | w11102 ;
  assign w11537 = w11377 & ~w11536 ;
  assign w11538 = w11100 ^ w11537 ;
  assign w11539 = ( ~w4727 & w11527 ) | ( ~w4727 & w11533 ) | ( w11527 & w11533 ) ;
  assign w11540 = ~w11527 & w11539 ;
  assign w11541 = w11538 | w11540 ;
  assign w11542 = ( w4457 & w11535 ) | ( w4457 & ~w11541 ) | ( w11535 & ~w11541 ) ;
  assign w11543 = w4457 & w11542 ;
  assign w11544 = w11105 | w11110 ;
  assign w11545 = w11377 & ~w11544 ;
  assign w11546 = w11108 ^ w11545 ;
  assign w11547 = ( ~w4457 & w11535 ) | ( ~w4457 & w11541 ) | ( w11535 & w11541 ) ;
  assign w11548 = ~w11535 & w11547 ;
  assign w11549 = w11546 | w11548 ;
  assign w11550 = ( w4195 & w11543 ) | ( w4195 & ~w11549 ) | ( w11543 & ~w11549 ) ;
  assign w11551 = w4195 & w11550 ;
  assign w11552 = w11113 | w11118 ;
  assign w11553 = w11377 & ~w11552 ;
  assign w11554 = w11116 ^ w11553 ;
  assign w11555 = ( ~w4195 & w11543 ) | ( ~w4195 & w11549 ) | ( w11543 & w11549 ) ;
  assign w11556 = ~w11543 & w11555 ;
  assign w11557 = w11554 | w11556 ;
  assign w11558 = ( w3941 & w11551 ) | ( w3941 & ~w11557 ) | ( w11551 & ~w11557 ) ;
  assign w11559 = w3941 & w11558 ;
  assign w11560 = w11121 | w11126 ;
  assign w11561 = w11377 & ~w11560 ;
  assign w11562 = w11124 ^ w11561 ;
  assign w11563 = ( ~w3941 & w11551 ) | ( ~w3941 & w11557 ) | ( w11551 & w11557 ) ;
  assign w11564 = ~w11551 & w11563 ;
  assign w11565 = w11562 | w11564 ;
  assign w11566 = ( w3695 & w11559 ) | ( w3695 & ~w11565 ) | ( w11559 & ~w11565 ) ;
  assign w11567 = w3695 & w11566 ;
  assign w11568 = w11129 | w11134 ;
  assign w11569 = w11377 & ~w11568 ;
  assign w11570 = w11132 ^ w11569 ;
  assign w11571 = ( ~w3695 & w11559 ) | ( ~w3695 & w11565 ) | ( w11559 & w11565 ) ;
  assign w11572 = ~w11559 & w11571 ;
  assign w11573 = w11570 | w11572 ;
  assign w11574 = ( w3457 & w11567 ) | ( w3457 & ~w11573 ) | ( w11567 & ~w11573 ) ;
  assign w11575 = w3457 & w11574 ;
  assign w11576 = w11137 | w11142 ;
  assign w11577 = w11377 & ~w11576 ;
  assign w11578 = w11140 ^ w11577 ;
  assign w11579 = ( ~w3457 & w11567 ) | ( ~w3457 & w11573 ) | ( w11567 & w11573 ) ;
  assign w11580 = ~w11567 & w11579 ;
  assign w11581 = w11578 | w11580 ;
  assign w11582 = ( w3227 & w11575 ) | ( w3227 & ~w11581 ) | ( w11575 & ~w11581 ) ;
  assign w11583 = w3227 & w11582 ;
  assign w11584 = w11145 | w11150 ;
  assign w11585 = w11377 & ~w11584 ;
  assign w11586 = w11148 ^ w11585 ;
  assign w11587 = ( ~w3227 & w11575 ) | ( ~w3227 & w11581 ) | ( w11575 & w11581 ) ;
  assign w11588 = ~w11575 & w11587 ;
  assign w11589 = w11586 | w11588 ;
  assign w11590 = ( w3005 & w11583 ) | ( w3005 & ~w11589 ) | ( w11583 & ~w11589 ) ;
  assign w11591 = w3005 & w11590 ;
  assign w11592 = w11153 | w11158 ;
  assign w11593 = w11377 & ~w11592 ;
  assign w11594 = w11156 ^ w11593 ;
  assign w11595 = ( ~w3005 & w11583 ) | ( ~w3005 & w11589 ) | ( w11583 & w11589 ) ;
  assign w11596 = ~w11583 & w11595 ;
  assign w11597 = w11594 | w11596 ;
  assign w11598 = ( w2791 & w11591 ) | ( w2791 & ~w11597 ) | ( w11591 & ~w11597 ) ;
  assign w11599 = w2791 & w11598 ;
  assign w11600 = w11161 | w11166 ;
  assign w11601 = w11377 & ~w11600 ;
  assign w11602 = w11164 ^ w11601 ;
  assign w11603 = ( ~w2791 & w11591 ) | ( ~w2791 & w11597 ) | ( w11591 & w11597 ) ;
  assign w11604 = ~w11591 & w11603 ;
  assign w11605 = w11602 | w11604 ;
  assign w11606 = ( w2585 & w11599 ) | ( w2585 & ~w11605 ) | ( w11599 & ~w11605 ) ;
  assign w11607 = w2585 & w11606 ;
  assign w11608 = w11169 | w11174 ;
  assign w11609 = w11377 & ~w11608 ;
  assign w11610 = w11172 ^ w11609 ;
  assign w11611 = ( ~w2585 & w11599 ) | ( ~w2585 & w11605 ) | ( w11599 & w11605 ) ;
  assign w11612 = ~w11599 & w11611 ;
  assign w11613 = w11610 | w11612 ;
  assign w11614 = ( w2387 & w11607 ) | ( w2387 & ~w11613 ) | ( w11607 & ~w11613 ) ;
  assign w11615 = w2387 & w11614 ;
  assign w11616 = w11177 | w11182 ;
  assign w11617 = w11377 & ~w11616 ;
  assign w11618 = w11180 ^ w11617 ;
  assign w11619 = ( ~w2387 & w11607 ) | ( ~w2387 & w11613 ) | ( w11607 & w11613 ) ;
  assign w11620 = ~w11607 & w11619 ;
  assign w11621 = w11618 | w11620 ;
  assign w11622 = ( w2197 & w11615 ) | ( w2197 & ~w11621 ) | ( w11615 & ~w11621 ) ;
  assign w11623 = w2197 & w11622 ;
  assign w11624 = w11185 | w11190 ;
  assign w11625 = w11377 & ~w11624 ;
  assign w11626 = w11188 ^ w11625 ;
  assign w11627 = ( ~w2197 & w11615 ) | ( ~w2197 & w11621 ) | ( w11615 & w11621 ) ;
  assign w11628 = ~w11615 & w11627 ;
  assign w11629 = w11626 | w11628 ;
  assign w11630 = ( w2015 & w11623 ) | ( w2015 & ~w11629 ) | ( w11623 & ~w11629 ) ;
  assign w11631 = w2015 & w11630 ;
  assign w11632 = w11193 | w11198 ;
  assign w11633 = w11377 & ~w11632 ;
  assign w11634 = w11196 ^ w11633 ;
  assign w11635 = ( ~w2015 & w11623 ) | ( ~w2015 & w11629 ) | ( w11623 & w11629 ) ;
  assign w11636 = ~w11623 & w11635 ;
  assign w11637 = w11634 | w11636 ;
  assign w11638 = ( w1841 & w11631 ) | ( w1841 & ~w11637 ) | ( w11631 & ~w11637 ) ;
  assign w11639 = w1841 & w11638 ;
  assign w11640 = w11201 | w11206 ;
  assign w11641 = w11377 & ~w11640 ;
  assign w11642 = w11204 ^ w11641 ;
  assign w11643 = ( ~w1841 & w11631 ) | ( ~w1841 & w11637 ) | ( w11631 & w11637 ) ;
  assign w11644 = ~w11631 & w11643 ;
  assign w11645 = w11642 | w11644 ;
  assign w11646 = ( w1675 & w11639 ) | ( w1675 & ~w11645 ) | ( w11639 & ~w11645 ) ;
  assign w11647 = w1675 & w11646 ;
  assign w11648 = w11209 | w11214 ;
  assign w11649 = w11377 & ~w11648 ;
  assign w11650 = w11212 ^ w11649 ;
  assign w11651 = ( ~w1675 & w11639 ) | ( ~w1675 & w11645 ) | ( w11639 & w11645 ) ;
  assign w11652 = ~w11639 & w11651 ;
  assign w11653 = w11650 | w11652 ;
  assign w11654 = ( w1517 & w11647 ) | ( w1517 & ~w11653 ) | ( w11647 & ~w11653 ) ;
  assign w11655 = w1517 & w11654 ;
  assign w11656 = w11217 | w11222 ;
  assign w11657 = w11377 & ~w11656 ;
  assign w11658 = w11220 ^ w11657 ;
  assign w11659 = ( ~w1517 & w11647 ) | ( ~w1517 & w11653 ) | ( w11647 & w11653 ) ;
  assign w11660 = ~w11647 & w11659 ;
  assign w11661 = w11658 | w11660 ;
  assign w11662 = ( w1367 & w11655 ) | ( w1367 & ~w11661 ) | ( w11655 & ~w11661 ) ;
  assign w11663 = w1367 & w11662 ;
  assign w11664 = w11225 | w11230 ;
  assign w11665 = w11377 & ~w11664 ;
  assign w11666 = w11228 ^ w11665 ;
  assign w11667 = ( ~w1367 & w11655 ) | ( ~w1367 & w11661 ) | ( w11655 & w11661 ) ;
  assign w11668 = ~w11655 & w11667 ;
  assign w11669 = w11666 | w11668 ;
  assign w11670 = ( w1225 & w11663 ) | ( w1225 & ~w11669 ) | ( w11663 & ~w11669 ) ;
  assign w11671 = w1225 & w11670 ;
  assign w11672 = w11233 | w11238 ;
  assign w11673 = w11377 & ~w11672 ;
  assign w11674 = w11236 ^ w11673 ;
  assign w11675 = ( ~w1225 & w11663 ) | ( ~w1225 & w11669 ) | ( w11663 & w11669 ) ;
  assign w11676 = ~w11663 & w11675 ;
  assign w11677 = w11674 | w11676 ;
  assign w11678 = ( w1091 & w11671 ) | ( w1091 & ~w11677 ) | ( w11671 & ~w11677 ) ;
  assign w11679 = w1091 & w11678 ;
  assign w11680 = w11241 | w11246 ;
  assign w11681 = w11377 & ~w11680 ;
  assign w11682 = w11244 ^ w11681 ;
  assign w11683 = ( ~w1091 & w11671 ) | ( ~w1091 & w11677 ) | ( w11671 & w11677 ) ;
  assign w11684 = ~w11671 & w11683 ;
  assign w11685 = w11682 | w11684 ;
  assign w11686 = ( w965 & w11679 ) | ( w965 & ~w11685 ) | ( w11679 & ~w11685 ) ;
  assign w11687 = w965 & w11686 ;
  assign w11688 = w11249 | w11254 ;
  assign w11689 = w11377 & ~w11688 ;
  assign w11690 = w11252 ^ w11689 ;
  assign w11691 = ( ~w965 & w11679 ) | ( ~w965 & w11685 ) | ( w11679 & w11685 ) ;
  assign w11692 = ~w11679 & w11691 ;
  assign w11693 = w11690 | w11692 ;
  assign w11694 = ( w847 & w11687 ) | ( w847 & ~w11693 ) | ( w11687 & ~w11693 ) ;
  assign w11695 = w847 & w11694 ;
  assign w11696 = ( ~w847 & w11687 ) | ( ~w847 & w11693 ) | ( w11687 & w11693 ) ;
  assign w11697 = ~w11687 & w11696 ;
  assign w11698 = w11257 | w11259 ;
  assign w11699 = w11377 & ~w11698 ;
  assign w11700 = w11262 ^ w11699 ;
  assign w11701 = w11697 | w11700 ;
  assign w11702 = ( w737 & w11695 ) | ( w737 & ~w11701 ) | ( w11695 & ~w11701 ) ;
  assign w11703 = w737 & w11702 ;
  assign w11704 = w11265 | w11270 ;
  assign w11705 = w11377 & ~w11704 ;
  assign w11706 = w11268 ^ w11705 ;
  assign w11707 = ( ~w737 & w11695 ) | ( ~w737 & w11701 ) | ( w11695 & w11701 ) ;
  assign w11708 = ~w11695 & w11707 ;
  assign w11709 = w11706 | w11708 ;
  assign w11710 = ( w635 & w11703 ) | ( w635 & ~w11709 ) | ( w11703 & ~w11709 ) ;
  assign w11711 = w635 & w11710 ;
  assign w11712 = w11273 | w11278 ;
  assign w11713 = w11377 & ~w11712 ;
  assign w11714 = w11276 ^ w11713 ;
  assign w11715 = ( ~w635 & w11703 ) | ( ~w635 & w11709 ) | ( w11703 & w11709 ) ;
  assign w11716 = ~w11703 & w11715 ;
  assign w11717 = w11714 | w11716 ;
  assign w11718 = ( w541 & w11711 ) | ( w541 & ~w11717 ) | ( w11711 & ~w11717 ) ;
  assign w11719 = w541 & w11718 ;
  assign w11720 = w11281 | w11286 ;
  assign w11721 = w11377 & ~w11720 ;
  assign w11722 = w11284 ^ w11721 ;
  assign w11723 = ( ~w541 & w11711 ) | ( ~w541 & w11717 ) | ( w11711 & w11717 ) ;
  assign w11724 = ~w11711 & w11723 ;
  assign w11725 = w11722 | w11724 ;
  assign w11726 = ( w455 & w11719 ) | ( w455 & ~w11725 ) | ( w11719 & ~w11725 ) ;
  assign w11727 = w455 & w11726 ;
  assign w11728 = w11289 | w11294 ;
  assign w11729 = w11377 & ~w11728 ;
  assign w11730 = w11292 ^ w11729 ;
  assign w11731 = ( ~w455 & w11719 ) | ( ~w455 & w11725 ) | ( w11719 & w11725 ) ;
  assign w11732 = ~w11719 & w11731 ;
  assign w11733 = w11730 | w11732 ;
  assign w11734 = ( w377 & w11727 ) | ( w377 & ~w11733 ) | ( w11727 & ~w11733 ) ;
  assign w11735 = w377 & w11734 ;
  assign w11736 = w11297 | w11302 ;
  assign w11737 = w11377 & ~w11736 ;
  assign w11738 = w11300 ^ w11737 ;
  assign w11739 = ( ~w377 & w11727 ) | ( ~w377 & w11733 ) | ( w11727 & w11733 ) ;
  assign w11740 = ~w11727 & w11739 ;
  assign w11741 = w11738 | w11740 ;
  assign w11742 = ( w307 & w11735 ) | ( w307 & ~w11741 ) | ( w11735 & ~w11741 ) ;
  assign w11743 = w307 & w11742 ;
  assign w11744 = w11305 | w11310 ;
  assign w11745 = w11377 & ~w11744 ;
  assign w11746 = w11308 ^ w11745 ;
  assign w11747 = ( ~w307 & w11735 ) | ( ~w307 & w11741 ) | ( w11735 & w11741 ) ;
  assign w11748 = ~w11735 & w11747 ;
  assign w11749 = w11746 | w11748 ;
  assign w11750 = ( w246 & w11743 ) | ( w246 & ~w11749 ) | ( w11743 & ~w11749 ) ;
  assign w11751 = w246 & w11750 ;
  assign w11752 = w11313 | w11318 ;
  assign w11753 = w11377 & ~w11752 ;
  assign w11754 = w11316 ^ w11753 ;
  assign w11755 = ( ~w246 & w11743 ) | ( ~w246 & w11749 ) | ( w11743 & w11749 ) ;
  assign w11756 = ~w11743 & w11755 ;
  assign w11757 = w11754 | w11756 ;
  assign w11758 = ( w185 & w11751 ) | ( w185 & ~w11757 ) | ( w11751 & ~w11757 ) ;
  assign w11759 = w185 & w11758 ;
  assign w11760 = w11321 | w11326 ;
  assign w11761 = w11377 & ~w11760 ;
  assign w11762 = w11324 ^ w11761 ;
  assign w11763 = ( ~w185 & w11751 ) | ( ~w185 & w11757 ) | ( w11751 & w11757 ) ;
  assign w11764 = ~w11751 & w11763 ;
  assign w11765 = w11762 | w11764 ;
  assign w11766 = ( w145 & w11759 ) | ( w145 & ~w11765 ) | ( w11759 & ~w11765 ) ;
  assign w11767 = w145 & w11766 ;
  assign w11768 = w11329 | w11334 ;
  assign w11769 = w11377 & ~w11768 ;
  assign w11770 = w11332 ^ w11769 ;
  assign w11771 = ( ~w145 & w11759 ) | ( ~w145 & w11765 ) | ( w11759 & w11765 ) ;
  assign w11772 = ~w11759 & w11771 ;
  assign w11773 = w11770 | w11772 ;
  assign w11774 = ( w132 & w11767 ) | ( w132 & ~w11773 ) | ( w11767 & ~w11773 ) ;
  assign w11775 = w132 & w11774 ;
  assign w11776 = w11337 | w11342 ;
  assign w11777 = w11377 & ~w11776 ;
  assign w11778 = w11340 ^ w11777 ;
  assign w11779 = ( ~w132 & w11767 ) | ( ~w132 & w11773 ) | ( w11767 & w11773 ) ;
  assign w11780 = ~w11767 & w11779 ;
  assign w11781 = w11778 | w11780 ;
  assign w11782 = ~w11775 & w11781 ;
  assign w11783 = w11345 | w11350 ;
  assign w11784 = w11377 & ~w11783 ;
  assign w11785 = w11348 ^ w11784 ;
  assign w11786 = ( ~w11363 & w11782 ) | ( ~w11363 & w11785 ) | ( w11782 & w11785 ) ;
  assign w11787 = w11352 & ~w11786 ;
  assign w11788 = ~w11355 & w11377 ;
  assign w11789 = ( w11786 & ~w11787 ) | ( w11786 & w11788 ) | ( ~w11787 & w11788 ) ;
  assign w11790 = w11363 | w11789 ;
  assign w11791 = ~w129 & w11790 ;
  assign w11792 = ( w11775 & w11781 ) | ( w11775 & w11785 ) | ( w11781 & w11785 ) ;
  assign w11793 = ~w11775 & w11792 ;
  assign w11794 = ( w129 & w11352 ) | ( w129 & w11355 ) | ( w11352 & w11355 ) ;
  assign w11795 = ( w11355 & ~w11377 ) | ( w11355 & w11794 ) | ( ~w11377 & w11794 ) ;
  assign w11796 = w11352 & w11795 ;
  assign w11797 = w11794 ^ w11796 ;
  assign w11798 = ( w10923 & w10928 ) | ( w10923 & w10955 ) | ( w10928 & w10955 ) ;
  assign w11799 = w10955 & ~w11798 ;
  assign w11800 = w10926 ^ w11799 ;
  assign w11801 = ( ~w11367 & w11374 ) | ( ~w11367 & w11800 ) | ( w11374 & w11800 ) ;
  assign w11802 = ~w11374 & w11801 ;
  assign w11803 = ( ~w11361 & w11363 ) | ( ~w11361 & w11802 ) | ( w11363 & w11802 ) ;
  assign w11804 = ~w11363 & w11803 ;
  assign w11805 = w11793 | w11804 ;
  assign w11806 = ( w11791 & ~w11793 ) | ( w11791 & w11797 ) | ( ~w11793 & w11797 ) ;
  assign w11807 = w11805 | w11806 ;
  assign w11808 = ( ~\pi023 & \pi024 ) | ( ~\pi023 & w11377 ) | ( \pi024 & w11377 ) ;
  assign w11809 = ( ~\pi022 & \pi024 ) | ( ~\pi022 & w11808 ) | ( \pi024 & w11808 ) ;
  assign w11810 = ( ~\pi024 & w11377 ) | ( ~\pi024 & w11807 ) | ( w11377 & w11807 ) ;
  assign w11811 = w11809 & w11810 ;
  assign w11812 = ( w11363 & w11367 ) | ( w11363 & ~w11374 ) | ( w11367 & ~w11374 ) ;
  assign w11813 = \pi023 & ~w11812 ;
  assign w11814 = \pi022 | \pi024 ;
  assign w11815 = ( ~w11812 & w11813 ) | ( ~w11812 & w11814 ) | ( w11813 & w11814 ) ;
  assign w11816 = ~w11374 & w11815 ;
  assign w11817 = ~w11361 & w11816 ;
  assign w11818 = ( \pi024 & w11807 ) | ( \pi024 & ~w11816 ) | ( w11807 & ~w11816 ) ;
  assign w11819 = w11817 & ~w11818 ;
  assign w11820 = ~\pi024 & w11807 ;
  assign w11821 = \pi025 ^ w11820 ;
  assign w11822 = w11819 | w11821 ;
  assign w11823 = ( w10955 & w11811 ) | ( w10955 & ~w11822 ) | ( w11811 & ~w11822 ) ;
  assign w11824 = w10955 & w11823 ;
  assign w11825 = ( ~w10955 & w11811 ) | ( ~w10955 & w11822 ) | ( w11811 & w11822 ) ;
  assign w11826 = ~w11811 & w11825 ;
  assign w11827 = w11377 & ~w11804 ;
  assign w11828 = ~w11793 & w11827 ;
  assign w11829 = ~w11806 & w11828 ;
  assign w11830 = \pi025 & w11807 ;
  assign w11831 = ( \pi024 & w11807 ) | ( \pi024 & ~w11830 ) | ( w11807 & ~w11830 ) ;
  assign w11832 = ( ~\pi024 & w11829 ) | ( ~\pi024 & w11831 ) | ( w11829 & w11831 ) ;
  assign w11833 = \pi026 ^ w11832 ;
  assign w11834 = w11826 | w11833 ;
  assign w11835 = ( w10541 & w11824 ) | ( w10541 & ~w11834 ) | ( w11824 & ~w11834 ) ;
  assign w11836 = w10541 & w11835 ;
  assign w11837 = ( w11381 & ~w11389 ) | ( w11381 & w11807 ) | ( ~w11389 & w11807 ) ;
  assign w11838 = ~w11381 & w11837 ;
  assign w11839 = \pi027 ^ w11838 ;
  assign w11840 = w11390 ^ w11839 ;
  assign w11841 = ( ~w10541 & w11824 ) | ( ~w10541 & w11834 ) | ( w11824 & w11834 ) ;
  assign w11842 = ~w11824 & w11841 ;
  assign w11843 = w11840 | w11842 ;
  assign w11844 = ( w10135 & w11836 ) | ( w10135 & ~w11843 ) | ( w11836 & ~w11843 ) ;
  assign w11845 = w10135 & w11844 ;
  assign w11846 = w11394 | w11396 ;
  assign w11847 = w11807 & ~w11846 ;
  assign w11848 = w11403 ^ w11847 ;
  assign w11849 = ( ~w10135 & w11836 ) | ( ~w10135 & w11843 ) | ( w11836 & w11843 ) ;
  assign w11850 = ~w11836 & w11849 ;
  assign w11851 = w11848 | w11850 ;
  assign w11852 = ( w9737 & w11845 ) | ( w9737 & ~w11851 ) | ( w11845 & ~w11851 ) ;
  assign w11853 = w9737 & w11852 ;
  assign w11854 = w11406 | w11412 ;
  assign w11855 = w11807 & ~w11854 ;
  assign w11856 = w11410 ^ w11855 ;
  assign w11857 = ( ~w9737 & w11845 ) | ( ~w9737 & w11851 ) | ( w11845 & w11851 ) ;
  assign w11858 = ~w11845 & w11857 ;
  assign w11859 = w11856 | w11858 ;
  assign w11860 = ( w9347 & w11853 ) | ( w9347 & ~w11859 ) | ( w11853 & ~w11859 ) ;
  assign w11861 = w9347 & w11860 ;
  assign w11862 = w11415 | w11420 ;
  assign w11863 = w11807 & ~w11862 ;
  assign w11864 = w11418 ^ w11863 ;
  assign w11865 = ( ~w9347 & w11853 ) | ( ~w9347 & w11859 ) | ( w11853 & w11859 ) ;
  assign w11866 = ~w11853 & w11865 ;
  assign w11867 = w11864 | w11866 ;
  assign w11868 = ( w8965 & w11861 ) | ( w8965 & ~w11867 ) | ( w11861 & ~w11867 ) ;
  assign w11869 = w8965 & w11868 ;
  assign w11870 = w11423 | w11428 ;
  assign w11871 = w11807 & ~w11870 ;
  assign w11872 = w11426 ^ w11871 ;
  assign w11873 = ( ~w8965 & w11861 ) | ( ~w8965 & w11867 ) | ( w11861 & w11867 ) ;
  assign w11874 = ~w11861 & w11873 ;
  assign w11875 = w11872 | w11874 ;
  assign w11876 = ( w8591 & w11869 ) | ( w8591 & ~w11875 ) | ( w11869 & ~w11875 ) ;
  assign w11877 = w8591 & w11876 ;
  assign w11878 = w11431 | w11436 ;
  assign w11879 = w11807 & ~w11878 ;
  assign w11880 = w11434 ^ w11879 ;
  assign w11881 = ( ~w8591 & w11869 ) | ( ~w8591 & w11875 ) | ( w11869 & w11875 ) ;
  assign w11882 = ~w11869 & w11881 ;
  assign w11883 = w11880 | w11882 ;
  assign w11884 = ( w8225 & w11877 ) | ( w8225 & ~w11883 ) | ( w11877 & ~w11883 ) ;
  assign w11885 = w8225 & w11884 ;
  assign w11886 = w11439 | w11444 ;
  assign w11887 = w11807 & ~w11886 ;
  assign w11888 = w11442 ^ w11887 ;
  assign w11889 = ( ~w8225 & w11877 ) | ( ~w8225 & w11883 ) | ( w11877 & w11883 ) ;
  assign w11890 = ~w11877 & w11889 ;
  assign w11891 = w11888 | w11890 ;
  assign w11892 = ( w7867 & w11885 ) | ( w7867 & ~w11891 ) | ( w11885 & ~w11891 ) ;
  assign w11893 = w7867 & w11892 ;
  assign w11894 = w11447 | w11452 ;
  assign w11895 = w11807 & ~w11894 ;
  assign w11896 = w11450 ^ w11895 ;
  assign w11897 = ( ~w7867 & w11885 ) | ( ~w7867 & w11891 ) | ( w11885 & w11891 ) ;
  assign w11898 = ~w11885 & w11897 ;
  assign w11899 = w11896 | w11898 ;
  assign w11900 = ( w7517 & w11893 ) | ( w7517 & ~w11899 ) | ( w11893 & ~w11899 ) ;
  assign w11901 = w7517 & w11900 ;
  assign w11902 = w11455 | w11460 ;
  assign w11903 = w11807 & ~w11902 ;
  assign w11904 = w11458 ^ w11903 ;
  assign w11905 = ( ~w7517 & w11893 ) | ( ~w7517 & w11899 ) | ( w11893 & w11899 ) ;
  assign w11906 = ~w11893 & w11905 ;
  assign w11907 = w11904 | w11906 ;
  assign w11908 = ( w7175 & w11901 ) | ( w7175 & ~w11907 ) | ( w11901 & ~w11907 ) ;
  assign w11909 = w7175 & w11908 ;
  assign w11910 = w11463 | w11468 ;
  assign w11911 = w11807 & ~w11910 ;
  assign w11912 = w11466 ^ w11911 ;
  assign w11913 = ( ~w7175 & w11901 ) | ( ~w7175 & w11907 ) | ( w11901 & w11907 ) ;
  assign w11914 = ~w11901 & w11913 ;
  assign w11915 = w11912 | w11914 ;
  assign w11916 = ( w6841 & w11909 ) | ( w6841 & ~w11915 ) | ( w11909 & ~w11915 ) ;
  assign w11917 = w6841 & w11916 ;
  assign w11918 = w11471 | w11476 ;
  assign w11919 = w11807 & ~w11918 ;
  assign w11920 = w11474 ^ w11919 ;
  assign w11921 = ( ~w6841 & w11909 ) | ( ~w6841 & w11915 ) | ( w11909 & w11915 ) ;
  assign w11922 = ~w11909 & w11921 ;
  assign w11923 = w11920 | w11922 ;
  assign w11924 = ( w6515 & w11917 ) | ( w6515 & ~w11923 ) | ( w11917 & ~w11923 ) ;
  assign w11925 = w6515 & w11924 ;
  assign w11926 = w11479 | w11484 ;
  assign w11927 = w11807 & ~w11926 ;
  assign w11928 = w11482 ^ w11927 ;
  assign w11929 = ( ~w6515 & w11917 ) | ( ~w6515 & w11923 ) | ( w11917 & w11923 ) ;
  assign w11930 = ~w11917 & w11929 ;
  assign w11931 = w11928 | w11930 ;
  assign w11932 = ( w6197 & w11925 ) | ( w6197 & ~w11931 ) | ( w11925 & ~w11931 ) ;
  assign w11933 = w6197 & w11932 ;
  assign w11934 = w11487 | w11492 ;
  assign w11935 = w11807 & ~w11934 ;
  assign w11936 = w11490 ^ w11935 ;
  assign w11937 = ( ~w6197 & w11925 ) | ( ~w6197 & w11931 ) | ( w11925 & w11931 ) ;
  assign w11938 = ~w11925 & w11937 ;
  assign w11939 = w11936 | w11938 ;
  assign w11940 = ( w5887 & w11933 ) | ( w5887 & ~w11939 ) | ( w11933 & ~w11939 ) ;
  assign w11941 = w5887 & w11940 ;
  assign w11942 = w11495 | w11500 ;
  assign w11943 = w11807 & ~w11942 ;
  assign w11944 = w11498 ^ w11943 ;
  assign w11945 = ( ~w5887 & w11933 ) | ( ~w5887 & w11939 ) | ( w11933 & w11939 ) ;
  assign w11946 = ~w11933 & w11945 ;
  assign w11947 = w11944 | w11946 ;
  assign w11948 = ( w5585 & w11941 ) | ( w5585 & ~w11947 ) | ( w11941 & ~w11947 ) ;
  assign w11949 = w5585 & w11948 ;
  assign w11950 = w11503 | w11508 ;
  assign w11951 = w11807 & ~w11950 ;
  assign w11952 = w11506 ^ w11951 ;
  assign w11953 = ( ~w5585 & w11941 ) | ( ~w5585 & w11947 ) | ( w11941 & w11947 ) ;
  assign w11954 = ~w11941 & w11953 ;
  assign w11955 = w11952 | w11954 ;
  assign w11956 = ( w5291 & w11949 ) | ( w5291 & ~w11955 ) | ( w11949 & ~w11955 ) ;
  assign w11957 = w5291 & w11956 ;
  assign w11958 = w11511 | w11516 ;
  assign w11959 = w11807 & ~w11958 ;
  assign w11960 = w11514 ^ w11959 ;
  assign w11961 = ( ~w5291 & w11949 ) | ( ~w5291 & w11955 ) | ( w11949 & w11955 ) ;
  assign w11962 = ~w11949 & w11961 ;
  assign w11963 = w11960 | w11962 ;
  assign w11964 = ( w5005 & w11957 ) | ( w5005 & ~w11963 ) | ( w11957 & ~w11963 ) ;
  assign w11965 = w5005 & w11964 ;
  assign w11966 = w11519 | w11524 ;
  assign w11967 = w11807 & ~w11966 ;
  assign w11968 = w11522 ^ w11967 ;
  assign w11969 = ( ~w5005 & w11957 ) | ( ~w5005 & w11963 ) | ( w11957 & w11963 ) ;
  assign w11970 = ~w11957 & w11969 ;
  assign w11971 = w11968 | w11970 ;
  assign w11972 = ( w4727 & w11965 ) | ( w4727 & ~w11971 ) | ( w11965 & ~w11971 ) ;
  assign w11973 = w4727 & w11972 ;
  assign w11974 = w11527 | w11532 ;
  assign w11975 = w11807 & ~w11974 ;
  assign w11976 = w11530 ^ w11975 ;
  assign w11977 = ( ~w4727 & w11965 ) | ( ~w4727 & w11971 ) | ( w11965 & w11971 ) ;
  assign w11978 = ~w11965 & w11977 ;
  assign w11979 = w11976 | w11978 ;
  assign w11980 = ( w4457 & w11973 ) | ( w4457 & ~w11979 ) | ( w11973 & ~w11979 ) ;
  assign w11981 = w4457 & w11980 ;
  assign w11982 = w11535 | w11540 ;
  assign w11983 = w11807 & ~w11982 ;
  assign w11984 = w11538 ^ w11983 ;
  assign w11985 = ( ~w4457 & w11973 ) | ( ~w4457 & w11979 ) | ( w11973 & w11979 ) ;
  assign w11986 = ~w11973 & w11985 ;
  assign w11987 = w11984 | w11986 ;
  assign w11988 = ( w4195 & w11981 ) | ( w4195 & ~w11987 ) | ( w11981 & ~w11987 ) ;
  assign w11989 = w4195 & w11988 ;
  assign w11990 = w11543 | w11548 ;
  assign w11991 = w11807 & ~w11990 ;
  assign w11992 = w11546 ^ w11991 ;
  assign w11993 = ( ~w4195 & w11981 ) | ( ~w4195 & w11987 ) | ( w11981 & w11987 ) ;
  assign w11994 = ~w11981 & w11993 ;
  assign w11995 = w11992 | w11994 ;
  assign w11996 = ( w3941 & w11989 ) | ( w3941 & ~w11995 ) | ( w11989 & ~w11995 ) ;
  assign w11997 = w3941 & w11996 ;
  assign w11998 = w11551 | w11556 ;
  assign w11999 = w11807 & ~w11998 ;
  assign w12000 = w11554 ^ w11999 ;
  assign w12001 = ( ~w3941 & w11989 ) | ( ~w3941 & w11995 ) | ( w11989 & w11995 ) ;
  assign w12002 = ~w11989 & w12001 ;
  assign w12003 = w12000 | w12002 ;
  assign w12004 = ( w3695 & w11997 ) | ( w3695 & ~w12003 ) | ( w11997 & ~w12003 ) ;
  assign w12005 = w3695 & w12004 ;
  assign w12006 = w11559 | w11564 ;
  assign w12007 = w11807 & ~w12006 ;
  assign w12008 = w11562 ^ w12007 ;
  assign w12009 = ( ~w3695 & w11997 ) | ( ~w3695 & w12003 ) | ( w11997 & w12003 ) ;
  assign w12010 = ~w11997 & w12009 ;
  assign w12011 = w12008 | w12010 ;
  assign w12012 = ( w3457 & w12005 ) | ( w3457 & ~w12011 ) | ( w12005 & ~w12011 ) ;
  assign w12013 = w3457 & w12012 ;
  assign w12014 = w11567 | w11572 ;
  assign w12015 = w11807 & ~w12014 ;
  assign w12016 = w11570 ^ w12015 ;
  assign w12017 = ( ~w3457 & w12005 ) | ( ~w3457 & w12011 ) | ( w12005 & w12011 ) ;
  assign w12018 = ~w12005 & w12017 ;
  assign w12019 = w12016 | w12018 ;
  assign w12020 = ( w3227 & w12013 ) | ( w3227 & ~w12019 ) | ( w12013 & ~w12019 ) ;
  assign w12021 = w3227 & w12020 ;
  assign w12022 = w11575 | w11580 ;
  assign w12023 = w11807 & ~w12022 ;
  assign w12024 = w11578 ^ w12023 ;
  assign w12025 = ( ~w3227 & w12013 ) | ( ~w3227 & w12019 ) | ( w12013 & w12019 ) ;
  assign w12026 = ~w12013 & w12025 ;
  assign w12027 = w12024 | w12026 ;
  assign w12028 = ( w3005 & w12021 ) | ( w3005 & ~w12027 ) | ( w12021 & ~w12027 ) ;
  assign w12029 = w3005 & w12028 ;
  assign w12030 = w11583 | w11588 ;
  assign w12031 = w11807 & ~w12030 ;
  assign w12032 = w11586 ^ w12031 ;
  assign w12033 = ( ~w3005 & w12021 ) | ( ~w3005 & w12027 ) | ( w12021 & w12027 ) ;
  assign w12034 = ~w12021 & w12033 ;
  assign w12035 = w12032 | w12034 ;
  assign w12036 = ( w2791 & w12029 ) | ( w2791 & ~w12035 ) | ( w12029 & ~w12035 ) ;
  assign w12037 = w2791 & w12036 ;
  assign w12038 = w11591 | w11596 ;
  assign w12039 = w11807 & ~w12038 ;
  assign w12040 = w11594 ^ w12039 ;
  assign w12041 = ( ~w2791 & w12029 ) | ( ~w2791 & w12035 ) | ( w12029 & w12035 ) ;
  assign w12042 = ~w12029 & w12041 ;
  assign w12043 = w12040 | w12042 ;
  assign w12044 = ( w2585 & w12037 ) | ( w2585 & ~w12043 ) | ( w12037 & ~w12043 ) ;
  assign w12045 = w2585 & w12044 ;
  assign w12046 = w11599 | w11604 ;
  assign w12047 = w11807 & ~w12046 ;
  assign w12048 = w11602 ^ w12047 ;
  assign w12049 = ( ~w2585 & w12037 ) | ( ~w2585 & w12043 ) | ( w12037 & w12043 ) ;
  assign w12050 = ~w12037 & w12049 ;
  assign w12051 = w12048 | w12050 ;
  assign w12052 = ( w2387 & w12045 ) | ( w2387 & ~w12051 ) | ( w12045 & ~w12051 ) ;
  assign w12053 = w2387 & w12052 ;
  assign w12054 = w11607 | w11612 ;
  assign w12055 = w11807 & ~w12054 ;
  assign w12056 = w11610 ^ w12055 ;
  assign w12057 = ( ~w2387 & w12045 ) | ( ~w2387 & w12051 ) | ( w12045 & w12051 ) ;
  assign w12058 = ~w12045 & w12057 ;
  assign w12059 = w12056 | w12058 ;
  assign w12060 = ( w2197 & w12053 ) | ( w2197 & ~w12059 ) | ( w12053 & ~w12059 ) ;
  assign w12061 = w2197 & w12060 ;
  assign w12062 = w11615 | w11620 ;
  assign w12063 = w11807 & ~w12062 ;
  assign w12064 = w11618 ^ w12063 ;
  assign w12065 = ( ~w2197 & w12053 ) | ( ~w2197 & w12059 ) | ( w12053 & w12059 ) ;
  assign w12066 = ~w12053 & w12065 ;
  assign w12067 = w12064 | w12066 ;
  assign w12068 = ( w2015 & w12061 ) | ( w2015 & ~w12067 ) | ( w12061 & ~w12067 ) ;
  assign w12069 = w2015 & w12068 ;
  assign w12070 = w11623 | w11628 ;
  assign w12071 = w11807 & ~w12070 ;
  assign w12072 = w11626 ^ w12071 ;
  assign w12073 = ( ~w2015 & w12061 ) | ( ~w2015 & w12067 ) | ( w12061 & w12067 ) ;
  assign w12074 = ~w12061 & w12073 ;
  assign w12075 = w12072 | w12074 ;
  assign w12076 = ( w1841 & w12069 ) | ( w1841 & ~w12075 ) | ( w12069 & ~w12075 ) ;
  assign w12077 = w1841 & w12076 ;
  assign w12078 = w11631 | w11636 ;
  assign w12079 = w11807 & ~w12078 ;
  assign w12080 = w11634 ^ w12079 ;
  assign w12081 = ( ~w1841 & w12069 ) | ( ~w1841 & w12075 ) | ( w12069 & w12075 ) ;
  assign w12082 = ~w12069 & w12081 ;
  assign w12083 = w12080 | w12082 ;
  assign w12084 = ( w1675 & w12077 ) | ( w1675 & ~w12083 ) | ( w12077 & ~w12083 ) ;
  assign w12085 = w1675 & w12084 ;
  assign w12086 = w11639 | w11644 ;
  assign w12087 = w11807 & ~w12086 ;
  assign w12088 = w11642 ^ w12087 ;
  assign w12089 = ( ~w1675 & w12077 ) | ( ~w1675 & w12083 ) | ( w12077 & w12083 ) ;
  assign w12090 = ~w12077 & w12089 ;
  assign w12091 = w12088 | w12090 ;
  assign w12092 = ( w1517 & w12085 ) | ( w1517 & ~w12091 ) | ( w12085 & ~w12091 ) ;
  assign w12093 = w1517 & w12092 ;
  assign w12094 = w11647 | w11652 ;
  assign w12095 = w11807 & ~w12094 ;
  assign w12096 = w11650 ^ w12095 ;
  assign w12097 = ( ~w1517 & w12085 ) | ( ~w1517 & w12091 ) | ( w12085 & w12091 ) ;
  assign w12098 = ~w12085 & w12097 ;
  assign w12099 = w12096 | w12098 ;
  assign w12100 = ( w1367 & w12093 ) | ( w1367 & ~w12099 ) | ( w12093 & ~w12099 ) ;
  assign w12101 = w1367 & w12100 ;
  assign w12102 = w11655 | w11660 ;
  assign w12103 = w11807 & ~w12102 ;
  assign w12104 = w11658 ^ w12103 ;
  assign w12105 = ( ~w1367 & w12093 ) | ( ~w1367 & w12099 ) | ( w12093 & w12099 ) ;
  assign w12106 = ~w12093 & w12105 ;
  assign w12107 = w12104 | w12106 ;
  assign w12108 = ( w1225 & w12101 ) | ( w1225 & ~w12107 ) | ( w12101 & ~w12107 ) ;
  assign w12109 = w1225 & w12108 ;
  assign w12110 = w11663 | w11668 ;
  assign w12111 = w11807 & ~w12110 ;
  assign w12112 = w11666 ^ w12111 ;
  assign w12113 = ( ~w1225 & w12101 ) | ( ~w1225 & w12107 ) | ( w12101 & w12107 ) ;
  assign w12114 = ~w12101 & w12113 ;
  assign w12115 = w12112 | w12114 ;
  assign w12116 = ( w1091 & w12109 ) | ( w1091 & ~w12115 ) | ( w12109 & ~w12115 ) ;
  assign w12117 = w1091 & w12116 ;
  assign w12118 = w11671 | w11676 ;
  assign w12119 = w11807 & ~w12118 ;
  assign w12120 = w11674 ^ w12119 ;
  assign w12121 = ( ~w1091 & w12109 ) | ( ~w1091 & w12115 ) | ( w12109 & w12115 ) ;
  assign w12122 = ~w12109 & w12121 ;
  assign w12123 = w12120 | w12122 ;
  assign w12124 = ( w965 & w12117 ) | ( w965 & ~w12123 ) | ( w12117 & ~w12123 ) ;
  assign w12125 = w965 & w12124 ;
  assign w12126 = w11679 | w11684 ;
  assign w12127 = w11807 & ~w12126 ;
  assign w12128 = w11682 ^ w12127 ;
  assign w12129 = ( ~w965 & w12117 ) | ( ~w965 & w12123 ) | ( w12117 & w12123 ) ;
  assign w12130 = ~w12117 & w12129 ;
  assign w12131 = w12128 | w12130 ;
  assign w12132 = ( w847 & w12125 ) | ( w847 & ~w12131 ) | ( w12125 & ~w12131 ) ;
  assign w12133 = w847 & w12132 ;
  assign w12134 = w11687 | w11692 ;
  assign w12135 = w11807 & ~w12134 ;
  assign w12136 = w11690 ^ w12135 ;
  assign w12137 = ( ~w847 & w12125 ) | ( ~w847 & w12131 ) | ( w12125 & w12131 ) ;
  assign w12138 = ~w12125 & w12137 ;
  assign w12139 = w12136 | w12138 ;
  assign w12140 = ( w737 & w12133 ) | ( w737 & ~w12139 ) | ( w12133 & ~w12139 ) ;
  assign w12141 = w737 & w12140 ;
  assign w12142 = ( ~w737 & w12133 ) | ( ~w737 & w12139 ) | ( w12133 & w12139 ) ;
  assign w12143 = ~w12133 & w12142 ;
  assign w12144 = w11695 | w11697 ;
  assign w12145 = w11807 & ~w12144 ;
  assign w12146 = w11700 ^ w12145 ;
  assign w12147 = w12143 | w12146 ;
  assign w12148 = ( w635 & w12141 ) | ( w635 & ~w12147 ) | ( w12141 & ~w12147 ) ;
  assign w12149 = w635 & w12148 ;
  assign w12150 = w11703 | w11708 ;
  assign w12151 = w11807 & ~w12150 ;
  assign w12152 = w11706 ^ w12151 ;
  assign w12153 = ( ~w635 & w12141 ) | ( ~w635 & w12147 ) | ( w12141 & w12147 ) ;
  assign w12154 = ~w12141 & w12153 ;
  assign w12155 = w12152 | w12154 ;
  assign w12156 = ( w541 & w12149 ) | ( w541 & ~w12155 ) | ( w12149 & ~w12155 ) ;
  assign w12157 = w541 & w12156 ;
  assign w12158 = w11711 | w11716 ;
  assign w12159 = w11807 & ~w12158 ;
  assign w12160 = w11714 ^ w12159 ;
  assign w12161 = ( ~w541 & w12149 ) | ( ~w541 & w12155 ) | ( w12149 & w12155 ) ;
  assign w12162 = ~w12149 & w12161 ;
  assign w12163 = w12160 | w12162 ;
  assign w12164 = ( w455 & w12157 ) | ( w455 & ~w12163 ) | ( w12157 & ~w12163 ) ;
  assign w12165 = w455 & w12164 ;
  assign w12166 = w11719 | w11724 ;
  assign w12167 = w11807 & ~w12166 ;
  assign w12168 = w11722 ^ w12167 ;
  assign w12169 = ( ~w455 & w12157 ) | ( ~w455 & w12163 ) | ( w12157 & w12163 ) ;
  assign w12170 = ~w12157 & w12169 ;
  assign w12171 = w12168 | w12170 ;
  assign w12172 = ( w377 & w12165 ) | ( w377 & ~w12171 ) | ( w12165 & ~w12171 ) ;
  assign w12173 = w377 & w12172 ;
  assign w12174 = w11727 | w11732 ;
  assign w12175 = w11807 & ~w12174 ;
  assign w12176 = w11730 ^ w12175 ;
  assign w12177 = ( ~w377 & w12165 ) | ( ~w377 & w12171 ) | ( w12165 & w12171 ) ;
  assign w12178 = ~w12165 & w12177 ;
  assign w12179 = w12176 | w12178 ;
  assign w12180 = ( w307 & w12173 ) | ( w307 & ~w12179 ) | ( w12173 & ~w12179 ) ;
  assign w12181 = w307 & w12180 ;
  assign w12182 = w11735 | w11740 ;
  assign w12183 = w11807 & ~w12182 ;
  assign w12184 = w11738 ^ w12183 ;
  assign w12185 = ( ~w307 & w12173 ) | ( ~w307 & w12179 ) | ( w12173 & w12179 ) ;
  assign w12186 = ~w12173 & w12185 ;
  assign w12187 = w12184 | w12186 ;
  assign w12188 = ( w246 & w12181 ) | ( w246 & ~w12187 ) | ( w12181 & ~w12187 ) ;
  assign w12189 = w246 & w12188 ;
  assign w12190 = w11743 | w11748 ;
  assign w12191 = w11807 & ~w12190 ;
  assign w12192 = w11746 ^ w12191 ;
  assign w12193 = ( ~w246 & w12181 ) | ( ~w246 & w12187 ) | ( w12181 & w12187 ) ;
  assign w12194 = ~w12181 & w12193 ;
  assign w12195 = w12192 | w12194 ;
  assign w12196 = ( w185 & w12189 ) | ( w185 & ~w12195 ) | ( w12189 & ~w12195 ) ;
  assign w12197 = w185 & w12196 ;
  assign w12198 = w11751 | w11756 ;
  assign w12199 = w11807 & ~w12198 ;
  assign w12200 = w11754 ^ w12199 ;
  assign w12201 = ( ~w185 & w12189 ) | ( ~w185 & w12195 ) | ( w12189 & w12195 ) ;
  assign w12202 = ~w12189 & w12201 ;
  assign w12203 = w12200 | w12202 ;
  assign w12204 = ( w145 & w12197 ) | ( w145 & ~w12203 ) | ( w12197 & ~w12203 ) ;
  assign w12205 = w145 & w12204 ;
  assign w12206 = w11759 | w11764 ;
  assign w12207 = w11807 & ~w12206 ;
  assign w12208 = w11762 ^ w12207 ;
  assign w12209 = ( ~w145 & w12197 ) | ( ~w145 & w12203 ) | ( w12197 & w12203 ) ;
  assign w12210 = ~w12197 & w12209 ;
  assign w12211 = w12208 | w12210 ;
  assign w12212 = ( w132 & w12205 ) | ( w132 & ~w12211 ) | ( w12205 & ~w12211 ) ;
  assign w12213 = w132 & w12212 ;
  assign w12214 = w11767 | w11772 ;
  assign w12215 = w11807 & ~w12214 ;
  assign w12216 = w11770 ^ w12215 ;
  assign w12217 = ( ~w132 & w12205 ) | ( ~w132 & w12211 ) | ( w12205 & w12211 ) ;
  assign w12218 = ~w12205 & w12217 ;
  assign w12219 = w12216 | w12218 ;
  assign w12220 = ~w12213 & w12219 ;
  assign w12221 = w11775 | w11780 ;
  assign w12222 = w11807 & ~w12221 ;
  assign w12223 = w11778 ^ w12222 ;
  assign w12224 = ( ~w11793 & w12220 ) | ( ~w11793 & w12223 ) | ( w12220 & w12223 ) ;
  assign w12225 = w11782 & ~w12224 ;
  assign w12226 = ~w11785 & w11807 ;
  assign w12227 = ( w12224 & ~w12225 ) | ( w12224 & w12226 ) | ( ~w12225 & w12226 ) ;
  assign w12228 = w11793 | w12227 ;
  assign w12229 = ~w129 & w12228 ;
  assign w12230 = ( w12213 & w12219 ) | ( w12213 & w12223 ) | ( w12219 & w12223 ) ;
  assign w12231 = ~w12213 & w12230 ;
  assign w12232 = ( w129 & w11782 ) | ( w129 & w11785 ) | ( w11782 & w11785 ) ;
  assign w12233 = ( w11785 & ~w11807 ) | ( w11785 & w12232 ) | ( ~w11807 & w12232 ) ;
  assign w12234 = w11782 & w12233 ;
  assign w12235 = w12232 ^ w12234 ;
  assign w12236 = ( w11345 & w11350 ) | ( w11345 & w11377 ) | ( w11350 & w11377 ) ;
  assign w12237 = w11377 & ~w12236 ;
  assign w12238 = w11348 ^ w12237 ;
  assign w12239 = ( ~w11797 & w11804 ) | ( ~w11797 & w12238 ) | ( w11804 & w12238 ) ;
  assign w12240 = ~w11804 & w12239 ;
  assign w12241 = ( ~w11791 & w11793 ) | ( ~w11791 & w12240 ) | ( w11793 & w12240 ) ;
  assign w12242 = ~w11793 & w12241 ;
  assign w12243 = w12231 | w12242 ;
  assign w12244 = ( w12229 & ~w12231 ) | ( w12229 & w12235 ) | ( ~w12231 & w12235 ) ;
  assign w12245 = w12243 | w12244 ;
  assign w12246 = ( ~\pi021 & \pi022 ) | ( ~\pi021 & w11807 ) | ( \pi022 & w11807 ) ;
  assign w12247 = ( ~\pi020 & \pi022 ) | ( ~\pi020 & w12246 ) | ( \pi022 & w12246 ) ;
  assign w12248 = ( ~\pi022 & w11807 ) | ( ~\pi022 & w12245 ) | ( w11807 & w12245 ) ;
  assign w12249 = w12247 & w12248 ;
  assign w12250 = ( w11793 & w11797 ) | ( w11793 & ~w11804 ) | ( w11797 & ~w11804 ) ;
  assign w12251 = \pi021 & ~w12250 ;
  assign w12252 = \pi020 | \pi022 ;
  assign w12253 = ( ~w12250 & w12251 ) | ( ~w12250 & w12252 ) | ( w12251 & w12252 ) ;
  assign w12254 = ~w11804 & w12253 ;
  assign w12255 = ~w11791 & w12254 ;
  assign w12256 = ( \pi022 & w12245 ) | ( \pi022 & ~w12254 ) | ( w12245 & ~w12254 ) ;
  assign w12257 = w12255 & ~w12256 ;
  assign w12258 = ~\pi022 & w12245 ;
  assign w12259 = \pi023 ^ w12258 ;
  assign w12260 = w12257 | w12259 ;
  assign w12261 = ( w11377 & w12249 ) | ( w11377 & ~w12260 ) | ( w12249 & ~w12260 ) ;
  assign w12262 = w11377 & w12261 ;
  assign w12263 = ( ~w11377 & w12249 ) | ( ~w11377 & w12260 ) | ( w12249 & w12260 ) ;
  assign w12264 = ~w12249 & w12263 ;
  assign w12265 = w11807 & ~w12242 ;
  assign w12266 = ~w12231 & w12265 ;
  assign w12267 = ~w12244 & w12266 ;
  assign w12268 = \pi023 & w12245 ;
  assign w12269 = ( \pi022 & w12245 ) | ( \pi022 & ~w12268 ) | ( w12245 & ~w12268 ) ;
  assign w12270 = ( ~\pi022 & w12267 ) | ( ~\pi022 & w12269 ) | ( w12267 & w12269 ) ;
  assign w12271 = \pi024 ^ w12270 ;
  assign w12272 = w12264 | w12271 ;
  assign w12273 = ( w10955 & w12262 ) | ( w10955 & ~w12272 ) | ( w12262 & ~w12272 ) ;
  assign w12274 = w10955 & w12273 ;
  assign w12275 = ( w11811 & ~w11819 ) | ( w11811 & w12245 ) | ( ~w11819 & w12245 ) ;
  assign w12276 = ~w11811 & w12275 ;
  assign w12277 = \pi025 ^ w12276 ;
  assign w12278 = w11820 ^ w12277 ;
  assign w12279 = ( ~w10955 & w12262 ) | ( ~w10955 & w12272 ) | ( w12262 & w12272 ) ;
  assign w12280 = ~w12262 & w12279 ;
  assign w12281 = w12278 | w12280 ;
  assign w12282 = ( w10541 & w12274 ) | ( w10541 & ~w12281 ) | ( w12274 & ~w12281 ) ;
  assign w12283 = w10541 & w12282 ;
  assign w12284 = w11824 | w11826 ;
  assign w12285 = w12245 & ~w12284 ;
  assign w12286 = w11833 ^ w12285 ;
  assign w12287 = ( ~w10541 & w12274 ) | ( ~w10541 & w12281 ) | ( w12274 & w12281 ) ;
  assign w12288 = ~w12274 & w12287 ;
  assign w12289 = w12286 | w12288 ;
  assign w12290 = ( w10135 & w12283 ) | ( w10135 & ~w12289 ) | ( w12283 & ~w12289 ) ;
  assign w12291 = w10135 & w12290 ;
  assign w12292 = w11836 | w11842 ;
  assign w12293 = w12245 & ~w12292 ;
  assign w12294 = w11840 ^ w12293 ;
  assign w12295 = ( ~w10135 & w12283 ) | ( ~w10135 & w12289 ) | ( w12283 & w12289 ) ;
  assign w12296 = ~w12283 & w12295 ;
  assign w12297 = w12294 | w12296 ;
  assign w12298 = ( w9737 & w12291 ) | ( w9737 & ~w12297 ) | ( w12291 & ~w12297 ) ;
  assign w12299 = w9737 & w12298 ;
  assign w12300 = w11845 | w11850 ;
  assign w12301 = w12245 & ~w12300 ;
  assign w12302 = w11848 ^ w12301 ;
  assign w12303 = ( ~w9737 & w12291 ) | ( ~w9737 & w12297 ) | ( w12291 & w12297 ) ;
  assign w12304 = ~w12291 & w12303 ;
  assign w12305 = w12302 | w12304 ;
  assign w12306 = ( w9347 & w12299 ) | ( w9347 & ~w12305 ) | ( w12299 & ~w12305 ) ;
  assign w12307 = w9347 & w12306 ;
  assign w12308 = w11853 | w11858 ;
  assign w12309 = w12245 & ~w12308 ;
  assign w12310 = w11856 ^ w12309 ;
  assign w12311 = ( ~w9347 & w12299 ) | ( ~w9347 & w12305 ) | ( w12299 & w12305 ) ;
  assign w12312 = ~w12299 & w12311 ;
  assign w12313 = w12310 | w12312 ;
  assign w12314 = ( w8965 & w12307 ) | ( w8965 & ~w12313 ) | ( w12307 & ~w12313 ) ;
  assign w12315 = w8965 & w12314 ;
  assign w12316 = w11861 | w11866 ;
  assign w12317 = w12245 & ~w12316 ;
  assign w12318 = w11864 ^ w12317 ;
  assign w12319 = ( ~w8965 & w12307 ) | ( ~w8965 & w12313 ) | ( w12307 & w12313 ) ;
  assign w12320 = ~w12307 & w12319 ;
  assign w12321 = w12318 | w12320 ;
  assign w12322 = ( w8591 & w12315 ) | ( w8591 & ~w12321 ) | ( w12315 & ~w12321 ) ;
  assign w12323 = w8591 & w12322 ;
  assign w12324 = w11869 | w11874 ;
  assign w12325 = w12245 & ~w12324 ;
  assign w12326 = w11872 ^ w12325 ;
  assign w12327 = ( ~w8591 & w12315 ) | ( ~w8591 & w12321 ) | ( w12315 & w12321 ) ;
  assign w12328 = ~w12315 & w12327 ;
  assign w12329 = w12326 | w12328 ;
  assign w12330 = ( w8225 & w12323 ) | ( w8225 & ~w12329 ) | ( w12323 & ~w12329 ) ;
  assign w12331 = w8225 & w12330 ;
  assign w12332 = w11877 | w11882 ;
  assign w12333 = w12245 & ~w12332 ;
  assign w12334 = w11880 ^ w12333 ;
  assign w12335 = ( ~w8225 & w12323 ) | ( ~w8225 & w12329 ) | ( w12323 & w12329 ) ;
  assign w12336 = ~w12323 & w12335 ;
  assign w12337 = w12334 | w12336 ;
  assign w12338 = ( w7867 & w12331 ) | ( w7867 & ~w12337 ) | ( w12331 & ~w12337 ) ;
  assign w12339 = w7867 & w12338 ;
  assign w12340 = w11885 | w11890 ;
  assign w12341 = w12245 & ~w12340 ;
  assign w12342 = w11888 ^ w12341 ;
  assign w12343 = ( ~w7867 & w12331 ) | ( ~w7867 & w12337 ) | ( w12331 & w12337 ) ;
  assign w12344 = ~w12331 & w12343 ;
  assign w12345 = w12342 | w12344 ;
  assign w12346 = ( w7517 & w12339 ) | ( w7517 & ~w12345 ) | ( w12339 & ~w12345 ) ;
  assign w12347 = w7517 & w12346 ;
  assign w12348 = w11893 | w11898 ;
  assign w12349 = w12245 & ~w12348 ;
  assign w12350 = w11896 ^ w12349 ;
  assign w12351 = ( ~w7517 & w12339 ) | ( ~w7517 & w12345 ) | ( w12339 & w12345 ) ;
  assign w12352 = ~w12339 & w12351 ;
  assign w12353 = w12350 | w12352 ;
  assign w12354 = ( w7175 & w12347 ) | ( w7175 & ~w12353 ) | ( w12347 & ~w12353 ) ;
  assign w12355 = w7175 & w12354 ;
  assign w12356 = w11901 | w11906 ;
  assign w12357 = w12245 & ~w12356 ;
  assign w12358 = w11904 ^ w12357 ;
  assign w12359 = ( ~w7175 & w12347 ) | ( ~w7175 & w12353 ) | ( w12347 & w12353 ) ;
  assign w12360 = ~w12347 & w12359 ;
  assign w12361 = w12358 | w12360 ;
  assign w12362 = ( w6841 & w12355 ) | ( w6841 & ~w12361 ) | ( w12355 & ~w12361 ) ;
  assign w12363 = w6841 & w12362 ;
  assign w12364 = w11909 | w11914 ;
  assign w12365 = w12245 & ~w12364 ;
  assign w12366 = w11912 ^ w12365 ;
  assign w12367 = ( ~w6841 & w12355 ) | ( ~w6841 & w12361 ) | ( w12355 & w12361 ) ;
  assign w12368 = ~w12355 & w12367 ;
  assign w12369 = w12366 | w12368 ;
  assign w12370 = ( w6515 & w12363 ) | ( w6515 & ~w12369 ) | ( w12363 & ~w12369 ) ;
  assign w12371 = w6515 & w12370 ;
  assign w12372 = w11917 | w11922 ;
  assign w12373 = w12245 & ~w12372 ;
  assign w12374 = w11920 ^ w12373 ;
  assign w12375 = ( ~w6515 & w12363 ) | ( ~w6515 & w12369 ) | ( w12363 & w12369 ) ;
  assign w12376 = ~w12363 & w12375 ;
  assign w12377 = w12374 | w12376 ;
  assign w12378 = ( w6197 & w12371 ) | ( w6197 & ~w12377 ) | ( w12371 & ~w12377 ) ;
  assign w12379 = w6197 & w12378 ;
  assign w12380 = w11925 | w11930 ;
  assign w12381 = w12245 & ~w12380 ;
  assign w12382 = w11928 ^ w12381 ;
  assign w12383 = ( ~w6197 & w12371 ) | ( ~w6197 & w12377 ) | ( w12371 & w12377 ) ;
  assign w12384 = ~w12371 & w12383 ;
  assign w12385 = w12382 | w12384 ;
  assign w12386 = ( w5887 & w12379 ) | ( w5887 & ~w12385 ) | ( w12379 & ~w12385 ) ;
  assign w12387 = w5887 & w12386 ;
  assign w12388 = w11933 | w11938 ;
  assign w12389 = w12245 & ~w12388 ;
  assign w12390 = w11936 ^ w12389 ;
  assign w12391 = ( ~w5887 & w12379 ) | ( ~w5887 & w12385 ) | ( w12379 & w12385 ) ;
  assign w12392 = ~w12379 & w12391 ;
  assign w12393 = w12390 | w12392 ;
  assign w12394 = ( w5585 & w12387 ) | ( w5585 & ~w12393 ) | ( w12387 & ~w12393 ) ;
  assign w12395 = w5585 & w12394 ;
  assign w12396 = w11941 | w11946 ;
  assign w12397 = w12245 & ~w12396 ;
  assign w12398 = w11944 ^ w12397 ;
  assign w12399 = ( ~w5585 & w12387 ) | ( ~w5585 & w12393 ) | ( w12387 & w12393 ) ;
  assign w12400 = ~w12387 & w12399 ;
  assign w12401 = w12398 | w12400 ;
  assign w12402 = ( w5291 & w12395 ) | ( w5291 & ~w12401 ) | ( w12395 & ~w12401 ) ;
  assign w12403 = w5291 & w12402 ;
  assign w12404 = w11949 | w11954 ;
  assign w12405 = w12245 & ~w12404 ;
  assign w12406 = w11952 ^ w12405 ;
  assign w12407 = ( ~w5291 & w12395 ) | ( ~w5291 & w12401 ) | ( w12395 & w12401 ) ;
  assign w12408 = ~w12395 & w12407 ;
  assign w12409 = w12406 | w12408 ;
  assign w12410 = ( w5005 & w12403 ) | ( w5005 & ~w12409 ) | ( w12403 & ~w12409 ) ;
  assign w12411 = w5005 & w12410 ;
  assign w12412 = w11957 | w11962 ;
  assign w12413 = w12245 & ~w12412 ;
  assign w12414 = w11960 ^ w12413 ;
  assign w12415 = ( ~w5005 & w12403 ) | ( ~w5005 & w12409 ) | ( w12403 & w12409 ) ;
  assign w12416 = ~w12403 & w12415 ;
  assign w12417 = w12414 | w12416 ;
  assign w12418 = ( w4727 & w12411 ) | ( w4727 & ~w12417 ) | ( w12411 & ~w12417 ) ;
  assign w12419 = w4727 & w12418 ;
  assign w12420 = w11965 | w11970 ;
  assign w12421 = w12245 & ~w12420 ;
  assign w12422 = w11968 ^ w12421 ;
  assign w12423 = ( ~w4727 & w12411 ) | ( ~w4727 & w12417 ) | ( w12411 & w12417 ) ;
  assign w12424 = ~w12411 & w12423 ;
  assign w12425 = w12422 | w12424 ;
  assign w12426 = ( w4457 & w12419 ) | ( w4457 & ~w12425 ) | ( w12419 & ~w12425 ) ;
  assign w12427 = w4457 & w12426 ;
  assign w12428 = w11973 | w11978 ;
  assign w12429 = w12245 & ~w12428 ;
  assign w12430 = w11976 ^ w12429 ;
  assign w12431 = ( ~w4457 & w12419 ) | ( ~w4457 & w12425 ) | ( w12419 & w12425 ) ;
  assign w12432 = ~w12419 & w12431 ;
  assign w12433 = w12430 | w12432 ;
  assign w12434 = ( w4195 & w12427 ) | ( w4195 & ~w12433 ) | ( w12427 & ~w12433 ) ;
  assign w12435 = w4195 & w12434 ;
  assign w12436 = w11981 | w11986 ;
  assign w12437 = w12245 & ~w12436 ;
  assign w12438 = w11984 ^ w12437 ;
  assign w12439 = ( ~w4195 & w12427 ) | ( ~w4195 & w12433 ) | ( w12427 & w12433 ) ;
  assign w12440 = ~w12427 & w12439 ;
  assign w12441 = w12438 | w12440 ;
  assign w12442 = ( w3941 & w12435 ) | ( w3941 & ~w12441 ) | ( w12435 & ~w12441 ) ;
  assign w12443 = w3941 & w12442 ;
  assign w12444 = w11989 | w11994 ;
  assign w12445 = w12245 & ~w12444 ;
  assign w12446 = w11992 ^ w12445 ;
  assign w12447 = ( ~w3941 & w12435 ) | ( ~w3941 & w12441 ) | ( w12435 & w12441 ) ;
  assign w12448 = ~w12435 & w12447 ;
  assign w12449 = w12446 | w12448 ;
  assign w12450 = ( w3695 & w12443 ) | ( w3695 & ~w12449 ) | ( w12443 & ~w12449 ) ;
  assign w12451 = w3695 & w12450 ;
  assign w12452 = w11997 | w12002 ;
  assign w12453 = w12245 & ~w12452 ;
  assign w12454 = w12000 ^ w12453 ;
  assign w12455 = ( ~w3695 & w12443 ) | ( ~w3695 & w12449 ) | ( w12443 & w12449 ) ;
  assign w12456 = ~w12443 & w12455 ;
  assign w12457 = w12454 | w12456 ;
  assign w12458 = ( w3457 & w12451 ) | ( w3457 & ~w12457 ) | ( w12451 & ~w12457 ) ;
  assign w12459 = w3457 & w12458 ;
  assign w12460 = w12005 | w12010 ;
  assign w12461 = w12245 & ~w12460 ;
  assign w12462 = w12008 ^ w12461 ;
  assign w12463 = ( ~w3457 & w12451 ) | ( ~w3457 & w12457 ) | ( w12451 & w12457 ) ;
  assign w12464 = ~w12451 & w12463 ;
  assign w12465 = w12462 | w12464 ;
  assign w12466 = ( w3227 & w12459 ) | ( w3227 & ~w12465 ) | ( w12459 & ~w12465 ) ;
  assign w12467 = w3227 & w12466 ;
  assign w12468 = w12013 | w12018 ;
  assign w12469 = w12245 & ~w12468 ;
  assign w12470 = w12016 ^ w12469 ;
  assign w12471 = ( ~w3227 & w12459 ) | ( ~w3227 & w12465 ) | ( w12459 & w12465 ) ;
  assign w12472 = ~w12459 & w12471 ;
  assign w12473 = w12470 | w12472 ;
  assign w12474 = ( w3005 & w12467 ) | ( w3005 & ~w12473 ) | ( w12467 & ~w12473 ) ;
  assign w12475 = w3005 & w12474 ;
  assign w12476 = w12021 | w12026 ;
  assign w12477 = w12245 & ~w12476 ;
  assign w12478 = w12024 ^ w12477 ;
  assign w12479 = ( ~w3005 & w12467 ) | ( ~w3005 & w12473 ) | ( w12467 & w12473 ) ;
  assign w12480 = ~w12467 & w12479 ;
  assign w12481 = w12478 | w12480 ;
  assign w12482 = ( w2791 & w12475 ) | ( w2791 & ~w12481 ) | ( w12475 & ~w12481 ) ;
  assign w12483 = w2791 & w12482 ;
  assign w12484 = w12029 | w12034 ;
  assign w12485 = w12245 & ~w12484 ;
  assign w12486 = w12032 ^ w12485 ;
  assign w12487 = ( ~w2791 & w12475 ) | ( ~w2791 & w12481 ) | ( w12475 & w12481 ) ;
  assign w12488 = ~w12475 & w12487 ;
  assign w12489 = w12486 | w12488 ;
  assign w12490 = ( w2585 & w12483 ) | ( w2585 & ~w12489 ) | ( w12483 & ~w12489 ) ;
  assign w12491 = w2585 & w12490 ;
  assign w12492 = w12037 | w12042 ;
  assign w12493 = w12245 & ~w12492 ;
  assign w12494 = w12040 ^ w12493 ;
  assign w12495 = ( ~w2585 & w12483 ) | ( ~w2585 & w12489 ) | ( w12483 & w12489 ) ;
  assign w12496 = ~w12483 & w12495 ;
  assign w12497 = w12494 | w12496 ;
  assign w12498 = ( w2387 & w12491 ) | ( w2387 & ~w12497 ) | ( w12491 & ~w12497 ) ;
  assign w12499 = w2387 & w12498 ;
  assign w12500 = w12045 | w12050 ;
  assign w12501 = w12245 & ~w12500 ;
  assign w12502 = w12048 ^ w12501 ;
  assign w12503 = ( ~w2387 & w12491 ) | ( ~w2387 & w12497 ) | ( w12491 & w12497 ) ;
  assign w12504 = ~w12491 & w12503 ;
  assign w12505 = w12502 | w12504 ;
  assign w12506 = ( w2197 & w12499 ) | ( w2197 & ~w12505 ) | ( w12499 & ~w12505 ) ;
  assign w12507 = w2197 & w12506 ;
  assign w12508 = w12053 | w12058 ;
  assign w12509 = w12245 & ~w12508 ;
  assign w12510 = w12056 ^ w12509 ;
  assign w12511 = ( ~w2197 & w12499 ) | ( ~w2197 & w12505 ) | ( w12499 & w12505 ) ;
  assign w12512 = ~w12499 & w12511 ;
  assign w12513 = w12510 | w12512 ;
  assign w12514 = ( w2015 & w12507 ) | ( w2015 & ~w12513 ) | ( w12507 & ~w12513 ) ;
  assign w12515 = w2015 & w12514 ;
  assign w12516 = w12061 | w12066 ;
  assign w12517 = w12245 & ~w12516 ;
  assign w12518 = w12064 ^ w12517 ;
  assign w12519 = ( ~w2015 & w12507 ) | ( ~w2015 & w12513 ) | ( w12507 & w12513 ) ;
  assign w12520 = ~w12507 & w12519 ;
  assign w12521 = w12518 | w12520 ;
  assign w12522 = ( w1841 & w12515 ) | ( w1841 & ~w12521 ) | ( w12515 & ~w12521 ) ;
  assign w12523 = w1841 & w12522 ;
  assign w12524 = w12069 | w12074 ;
  assign w12525 = w12245 & ~w12524 ;
  assign w12526 = w12072 ^ w12525 ;
  assign w12527 = ( ~w1841 & w12515 ) | ( ~w1841 & w12521 ) | ( w12515 & w12521 ) ;
  assign w12528 = ~w12515 & w12527 ;
  assign w12529 = w12526 | w12528 ;
  assign w12530 = ( w1675 & w12523 ) | ( w1675 & ~w12529 ) | ( w12523 & ~w12529 ) ;
  assign w12531 = w1675 & w12530 ;
  assign w12532 = w12077 | w12082 ;
  assign w12533 = w12245 & ~w12532 ;
  assign w12534 = w12080 ^ w12533 ;
  assign w12535 = ( ~w1675 & w12523 ) | ( ~w1675 & w12529 ) | ( w12523 & w12529 ) ;
  assign w12536 = ~w12523 & w12535 ;
  assign w12537 = w12534 | w12536 ;
  assign w12538 = ( w1517 & w12531 ) | ( w1517 & ~w12537 ) | ( w12531 & ~w12537 ) ;
  assign w12539 = w1517 & w12538 ;
  assign w12540 = w12085 | w12090 ;
  assign w12541 = w12245 & ~w12540 ;
  assign w12542 = w12088 ^ w12541 ;
  assign w12543 = ( ~w1517 & w12531 ) | ( ~w1517 & w12537 ) | ( w12531 & w12537 ) ;
  assign w12544 = ~w12531 & w12543 ;
  assign w12545 = w12542 | w12544 ;
  assign w12546 = ( w1367 & w12539 ) | ( w1367 & ~w12545 ) | ( w12539 & ~w12545 ) ;
  assign w12547 = w1367 & w12546 ;
  assign w12548 = w12093 | w12098 ;
  assign w12549 = w12245 & ~w12548 ;
  assign w12550 = w12096 ^ w12549 ;
  assign w12551 = ( ~w1367 & w12539 ) | ( ~w1367 & w12545 ) | ( w12539 & w12545 ) ;
  assign w12552 = ~w12539 & w12551 ;
  assign w12553 = w12550 | w12552 ;
  assign w12554 = ( w1225 & w12547 ) | ( w1225 & ~w12553 ) | ( w12547 & ~w12553 ) ;
  assign w12555 = w1225 & w12554 ;
  assign w12556 = w12101 | w12106 ;
  assign w12557 = w12245 & ~w12556 ;
  assign w12558 = w12104 ^ w12557 ;
  assign w12559 = ( ~w1225 & w12547 ) | ( ~w1225 & w12553 ) | ( w12547 & w12553 ) ;
  assign w12560 = ~w12547 & w12559 ;
  assign w12561 = w12558 | w12560 ;
  assign w12562 = ( w1091 & w12555 ) | ( w1091 & ~w12561 ) | ( w12555 & ~w12561 ) ;
  assign w12563 = w1091 & w12562 ;
  assign w12564 = w12109 | w12114 ;
  assign w12565 = w12245 & ~w12564 ;
  assign w12566 = w12112 ^ w12565 ;
  assign w12567 = ( ~w1091 & w12555 ) | ( ~w1091 & w12561 ) | ( w12555 & w12561 ) ;
  assign w12568 = ~w12555 & w12567 ;
  assign w12569 = w12566 | w12568 ;
  assign w12570 = ( w965 & w12563 ) | ( w965 & ~w12569 ) | ( w12563 & ~w12569 ) ;
  assign w12571 = w965 & w12570 ;
  assign w12572 = w12117 | w12122 ;
  assign w12573 = w12245 & ~w12572 ;
  assign w12574 = w12120 ^ w12573 ;
  assign w12575 = ( ~w965 & w12563 ) | ( ~w965 & w12569 ) | ( w12563 & w12569 ) ;
  assign w12576 = ~w12563 & w12575 ;
  assign w12577 = w12574 | w12576 ;
  assign w12578 = ( w847 & w12571 ) | ( w847 & ~w12577 ) | ( w12571 & ~w12577 ) ;
  assign w12579 = w847 & w12578 ;
  assign w12580 = w12125 | w12130 ;
  assign w12581 = w12245 & ~w12580 ;
  assign w12582 = w12128 ^ w12581 ;
  assign w12583 = ( ~w847 & w12571 ) | ( ~w847 & w12577 ) | ( w12571 & w12577 ) ;
  assign w12584 = ~w12571 & w12583 ;
  assign w12585 = w12582 | w12584 ;
  assign w12586 = ( w737 & w12579 ) | ( w737 & ~w12585 ) | ( w12579 & ~w12585 ) ;
  assign w12587 = w737 & w12586 ;
  assign w12588 = w12133 | w12138 ;
  assign w12589 = w12245 & ~w12588 ;
  assign w12590 = w12136 ^ w12589 ;
  assign w12591 = ( ~w737 & w12579 ) | ( ~w737 & w12585 ) | ( w12579 & w12585 ) ;
  assign w12592 = ~w12579 & w12591 ;
  assign w12593 = w12590 | w12592 ;
  assign w12594 = ( w635 & w12587 ) | ( w635 & ~w12593 ) | ( w12587 & ~w12593 ) ;
  assign w12595 = w635 & w12594 ;
  assign w12596 = ( ~w635 & w12587 ) | ( ~w635 & w12593 ) | ( w12587 & w12593 ) ;
  assign w12597 = ~w12587 & w12596 ;
  assign w12598 = w12141 | w12143 ;
  assign w12599 = w12245 & ~w12598 ;
  assign w12600 = w12146 ^ w12599 ;
  assign w12601 = w12597 | w12600 ;
  assign w12602 = ( w541 & w12595 ) | ( w541 & ~w12601 ) | ( w12595 & ~w12601 ) ;
  assign w12603 = w541 & w12602 ;
  assign w12604 = w12149 | w12154 ;
  assign w12605 = w12245 & ~w12604 ;
  assign w12606 = w12152 ^ w12605 ;
  assign w12607 = ( ~w541 & w12595 ) | ( ~w541 & w12601 ) | ( w12595 & w12601 ) ;
  assign w12608 = ~w12595 & w12607 ;
  assign w12609 = w12606 | w12608 ;
  assign w12610 = ( w455 & w12603 ) | ( w455 & ~w12609 ) | ( w12603 & ~w12609 ) ;
  assign w12611 = w455 & w12610 ;
  assign w12612 = w12157 | w12162 ;
  assign w12613 = w12245 & ~w12612 ;
  assign w12614 = w12160 ^ w12613 ;
  assign w12615 = ( ~w455 & w12603 ) | ( ~w455 & w12609 ) | ( w12603 & w12609 ) ;
  assign w12616 = ~w12603 & w12615 ;
  assign w12617 = w12614 | w12616 ;
  assign w12618 = ( w377 & w12611 ) | ( w377 & ~w12617 ) | ( w12611 & ~w12617 ) ;
  assign w12619 = w377 & w12618 ;
  assign w12620 = w12165 | w12170 ;
  assign w12621 = w12245 & ~w12620 ;
  assign w12622 = w12168 ^ w12621 ;
  assign w12623 = ( ~w377 & w12611 ) | ( ~w377 & w12617 ) | ( w12611 & w12617 ) ;
  assign w12624 = ~w12611 & w12623 ;
  assign w12625 = w12622 | w12624 ;
  assign w12626 = ( w307 & w12619 ) | ( w307 & ~w12625 ) | ( w12619 & ~w12625 ) ;
  assign w12627 = w307 & w12626 ;
  assign w12628 = w12173 | w12178 ;
  assign w12629 = w12245 & ~w12628 ;
  assign w12630 = w12176 ^ w12629 ;
  assign w12631 = ( ~w307 & w12619 ) | ( ~w307 & w12625 ) | ( w12619 & w12625 ) ;
  assign w12632 = ~w12619 & w12631 ;
  assign w12633 = w12630 | w12632 ;
  assign w12634 = ( w246 & w12627 ) | ( w246 & ~w12633 ) | ( w12627 & ~w12633 ) ;
  assign w12635 = w246 & w12634 ;
  assign w12636 = w12181 | w12186 ;
  assign w12637 = w12245 & ~w12636 ;
  assign w12638 = w12184 ^ w12637 ;
  assign w12639 = ( ~w246 & w12627 ) | ( ~w246 & w12633 ) | ( w12627 & w12633 ) ;
  assign w12640 = ~w12627 & w12639 ;
  assign w12641 = w12638 | w12640 ;
  assign w12642 = ( w185 & w12635 ) | ( w185 & ~w12641 ) | ( w12635 & ~w12641 ) ;
  assign w12643 = w185 & w12642 ;
  assign w12644 = w12189 | w12194 ;
  assign w12645 = w12245 & ~w12644 ;
  assign w12646 = w12192 ^ w12645 ;
  assign w12647 = ( ~w185 & w12635 ) | ( ~w185 & w12641 ) | ( w12635 & w12641 ) ;
  assign w12648 = ~w12635 & w12647 ;
  assign w12649 = w12646 | w12648 ;
  assign w12650 = ( w145 & w12643 ) | ( w145 & ~w12649 ) | ( w12643 & ~w12649 ) ;
  assign w12651 = w145 & w12650 ;
  assign w12652 = w12197 | w12202 ;
  assign w12653 = w12245 & ~w12652 ;
  assign w12654 = w12200 ^ w12653 ;
  assign w12655 = ( ~w145 & w12643 ) | ( ~w145 & w12649 ) | ( w12643 & w12649 ) ;
  assign w12656 = ~w12643 & w12655 ;
  assign w12657 = w12654 | w12656 ;
  assign w12658 = ( w132 & w12651 ) | ( w132 & ~w12657 ) | ( w12651 & ~w12657 ) ;
  assign w12659 = w132 & w12658 ;
  assign w12660 = w12205 | w12210 ;
  assign w12661 = w12245 & ~w12660 ;
  assign w12662 = w12208 ^ w12661 ;
  assign w12663 = ( ~w132 & w12651 ) | ( ~w132 & w12657 ) | ( w12651 & w12657 ) ;
  assign w12664 = ~w12651 & w12663 ;
  assign w12665 = w12662 | w12664 ;
  assign w12666 = ~w12659 & w12665 ;
  assign w12667 = w12213 | w12218 ;
  assign w12668 = w12245 & ~w12667 ;
  assign w12669 = w12216 ^ w12668 ;
  assign w12670 = ( ~w12231 & w12666 ) | ( ~w12231 & w12669 ) | ( w12666 & w12669 ) ;
  assign w12671 = w12220 & ~w12670 ;
  assign w12672 = ~w12223 & w12245 ;
  assign w12673 = ( w12670 & ~w12671 ) | ( w12670 & w12672 ) | ( ~w12671 & w12672 ) ;
  assign w12674 = w12231 | w12673 ;
  assign w12675 = ~w129 & w12674 ;
  assign w12676 = ( w12659 & w12665 ) | ( w12659 & w12669 ) | ( w12665 & w12669 ) ;
  assign w12677 = ~w12659 & w12676 ;
  assign w12678 = ( w129 & w12220 ) | ( w129 & w12223 ) | ( w12220 & w12223 ) ;
  assign w12679 = ( w12223 & ~w12245 ) | ( w12223 & w12678 ) | ( ~w12245 & w12678 ) ;
  assign w12680 = w12220 & w12679 ;
  assign w12681 = w12678 ^ w12680 ;
  assign w12682 = ( w11775 & w11780 ) | ( w11775 & w11807 ) | ( w11780 & w11807 ) ;
  assign w12683 = w11807 & ~w12682 ;
  assign w12684 = w11778 ^ w12683 ;
  assign w12685 = ( ~w12235 & w12242 ) | ( ~w12235 & w12684 ) | ( w12242 & w12684 ) ;
  assign w12686 = ~w12242 & w12685 ;
  assign w12687 = ( ~w12229 & w12231 ) | ( ~w12229 & w12686 ) | ( w12231 & w12686 ) ;
  assign w12688 = ~w12231 & w12687 ;
  assign w12689 = w12677 | w12688 ;
  assign w12690 = ( w12675 & ~w12677 ) | ( w12675 & w12681 ) | ( ~w12677 & w12681 ) ;
  assign w12691 = w12689 | w12690 ;
  assign w12692 = ( ~\pi019 & \pi020 ) | ( ~\pi019 & w12245 ) | ( \pi020 & w12245 ) ;
  assign w12693 = ( ~\pi018 & \pi020 ) | ( ~\pi018 & w12692 ) | ( \pi020 & w12692 ) ;
  assign w12694 = ( ~\pi020 & w12245 ) | ( ~\pi020 & w12691 ) | ( w12245 & w12691 ) ;
  assign w12695 = w12693 & w12694 ;
  assign w12696 = ( w12231 & w12235 ) | ( w12231 & ~w12242 ) | ( w12235 & ~w12242 ) ;
  assign w12697 = \pi019 & ~w12696 ;
  assign w12698 = \pi018 | \pi020 ;
  assign w12699 = ( ~w12696 & w12697 ) | ( ~w12696 & w12698 ) | ( w12697 & w12698 ) ;
  assign w12700 = ~w12242 & w12699 ;
  assign w12701 = ~w12229 & w12700 ;
  assign w12702 = ( \pi020 & w12691 ) | ( \pi020 & ~w12700 ) | ( w12691 & ~w12700 ) ;
  assign w12703 = w12701 & ~w12702 ;
  assign w12704 = ~\pi020 & w12691 ;
  assign w12705 = \pi021 ^ w12704 ;
  assign w12706 = w12703 | w12705 ;
  assign w12707 = ( w11807 & w12695 ) | ( w11807 & ~w12706 ) | ( w12695 & ~w12706 ) ;
  assign w12708 = w11807 & w12707 ;
  assign w12709 = ( ~w11807 & w12695 ) | ( ~w11807 & w12706 ) | ( w12695 & w12706 ) ;
  assign w12710 = ~w12695 & w12709 ;
  assign w12711 = w12245 & ~w12688 ;
  assign w12712 = ~w12677 & w12711 ;
  assign w12713 = ~w12690 & w12712 ;
  assign w12714 = \pi021 & w12691 ;
  assign w12715 = ( \pi020 & w12691 ) | ( \pi020 & ~w12714 ) | ( w12691 & ~w12714 ) ;
  assign w12716 = ( ~\pi020 & w12713 ) | ( ~\pi020 & w12715 ) | ( w12713 & w12715 ) ;
  assign w12717 = \pi022 ^ w12716 ;
  assign w12718 = w12710 | w12717 ;
  assign w12719 = ( w11377 & w12708 ) | ( w11377 & ~w12718 ) | ( w12708 & ~w12718 ) ;
  assign w12720 = w11377 & w12719 ;
  assign w12721 = ( w12249 & ~w12257 ) | ( w12249 & w12691 ) | ( ~w12257 & w12691 ) ;
  assign w12722 = ~w12249 & w12721 ;
  assign w12723 = \pi023 ^ w12722 ;
  assign w12724 = w12258 ^ w12723 ;
  assign w12725 = ( ~w11377 & w12708 ) | ( ~w11377 & w12718 ) | ( w12708 & w12718 ) ;
  assign w12726 = ~w12708 & w12725 ;
  assign w12727 = w12724 | w12726 ;
  assign w12728 = ( w10955 & w12720 ) | ( w10955 & ~w12727 ) | ( w12720 & ~w12727 ) ;
  assign w12729 = w10955 & w12728 ;
  assign w12730 = w12262 | w12264 ;
  assign w12731 = w12691 & ~w12730 ;
  assign w12732 = w12271 ^ w12731 ;
  assign w12733 = ( ~w10955 & w12720 ) | ( ~w10955 & w12727 ) | ( w12720 & w12727 ) ;
  assign w12734 = ~w12720 & w12733 ;
  assign w12735 = w12732 | w12734 ;
  assign w12736 = ( w10541 & w12729 ) | ( w10541 & ~w12735 ) | ( w12729 & ~w12735 ) ;
  assign w12737 = w10541 & w12736 ;
  assign w12738 = w12274 | w12280 ;
  assign w12739 = w12691 & ~w12738 ;
  assign w12740 = w12278 ^ w12739 ;
  assign w12741 = ( ~w10541 & w12729 ) | ( ~w10541 & w12735 ) | ( w12729 & w12735 ) ;
  assign w12742 = ~w12729 & w12741 ;
  assign w12743 = w12740 | w12742 ;
  assign w12744 = ( w10135 & w12737 ) | ( w10135 & ~w12743 ) | ( w12737 & ~w12743 ) ;
  assign w12745 = w10135 & w12744 ;
  assign w12746 = w12283 | w12288 ;
  assign w12747 = w12691 & ~w12746 ;
  assign w12748 = w12286 ^ w12747 ;
  assign w12749 = ( ~w10135 & w12737 ) | ( ~w10135 & w12743 ) | ( w12737 & w12743 ) ;
  assign w12750 = ~w12737 & w12749 ;
  assign w12751 = w12748 | w12750 ;
  assign w12752 = ( w9737 & w12745 ) | ( w9737 & ~w12751 ) | ( w12745 & ~w12751 ) ;
  assign w12753 = w9737 & w12752 ;
  assign w12754 = w12291 | w12296 ;
  assign w12755 = w12691 & ~w12754 ;
  assign w12756 = w12294 ^ w12755 ;
  assign w12757 = ( ~w9737 & w12745 ) | ( ~w9737 & w12751 ) | ( w12745 & w12751 ) ;
  assign w12758 = ~w12745 & w12757 ;
  assign w12759 = w12756 | w12758 ;
  assign w12760 = ( w9347 & w12753 ) | ( w9347 & ~w12759 ) | ( w12753 & ~w12759 ) ;
  assign w12761 = w9347 & w12760 ;
  assign w12762 = w12299 | w12304 ;
  assign w12763 = w12691 & ~w12762 ;
  assign w12764 = w12302 ^ w12763 ;
  assign w12765 = ( ~w9347 & w12753 ) | ( ~w9347 & w12759 ) | ( w12753 & w12759 ) ;
  assign w12766 = ~w12753 & w12765 ;
  assign w12767 = w12764 | w12766 ;
  assign w12768 = ( w8965 & w12761 ) | ( w8965 & ~w12767 ) | ( w12761 & ~w12767 ) ;
  assign w12769 = w8965 & w12768 ;
  assign w12770 = w12307 | w12312 ;
  assign w12771 = w12691 & ~w12770 ;
  assign w12772 = w12310 ^ w12771 ;
  assign w12773 = ( ~w8965 & w12761 ) | ( ~w8965 & w12767 ) | ( w12761 & w12767 ) ;
  assign w12774 = ~w12761 & w12773 ;
  assign w12775 = w12772 | w12774 ;
  assign w12776 = ( w8591 & w12769 ) | ( w8591 & ~w12775 ) | ( w12769 & ~w12775 ) ;
  assign w12777 = w8591 & w12776 ;
  assign w12778 = w12315 | w12320 ;
  assign w12779 = w12691 & ~w12778 ;
  assign w12780 = w12318 ^ w12779 ;
  assign w12781 = ( ~w8591 & w12769 ) | ( ~w8591 & w12775 ) | ( w12769 & w12775 ) ;
  assign w12782 = ~w12769 & w12781 ;
  assign w12783 = w12780 | w12782 ;
  assign w12784 = ( w8225 & w12777 ) | ( w8225 & ~w12783 ) | ( w12777 & ~w12783 ) ;
  assign w12785 = w8225 & w12784 ;
  assign w12786 = w12323 | w12328 ;
  assign w12787 = w12691 & ~w12786 ;
  assign w12788 = w12326 ^ w12787 ;
  assign w12789 = ( ~w8225 & w12777 ) | ( ~w8225 & w12783 ) | ( w12777 & w12783 ) ;
  assign w12790 = ~w12777 & w12789 ;
  assign w12791 = w12788 | w12790 ;
  assign w12792 = ( w7867 & w12785 ) | ( w7867 & ~w12791 ) | ( w12785 & ~w12791 ) ;
  assign w12793 = w7867 & w12792 ;
  assign w12794 = w12331 | w12336 ;
  assign w12795 = w12691 & ~w12794 ;
  assign w12796 = w12334 ^ w12795 ;
  assign w12797 = ( ~w7867 & w12785 ) | ( ~w7867 & w12791 ) | ( w12785 & w12791 ) ;
  assign w12798 = ~w12785 & w12797 ;
  assign w12799 = w12796 | w12798 ;
  assign w12800 = ( w7517 & w12793 ) | ( w7517 & ~w12799 ) | ( w12793 & ~w12799 ) ;
  assign w12801 = w7517 & w12800 ;
  assign w12802 = w12339 | w12344 ;
  assign w12803 = w12691 & ~w12802 ;
  assign w12804 = w12342 ^ w12803 ;
  assign w12805 = ( ~w7517 & w12793 ) | ( ~w7517 & w12799 ) | ( w12793 & w12799 ) ;
  assign w12806 = ~w12793 & w12805 ;
  assign w12807 = w12804 | w12806 ;
  assign w12808 = ( w7175 & w12801 ) | ( w7175 & ~w12807 ) | ( w12801 & ~w12807 ) ;
  assign w12809 = w7175 & w12808 ;
  assign w12810 = w12347 | w12352 ;
  assign w12811 = w12691 & ~w12810 ;
  assign w12812 = w12350 ^ w12811 ;
  assign w12813 = ( ~w7175 & w12801 ) | ( ~w7175 & w12807 ) | ( w12801 & w12807 ) ;
  assign w12814 = ~w12801 & w12813 ;
  assign w12815 = w12812 | w12814 ;
  assign w12816 = ( w6841 & w12809 ) | ( w6841 & ~w12815 ) | ( w12809 & ~w12815 ) ;
  assign w12817 = w6841 & w12816 ;
  assign w12818 = w12355 | w12360 ;
  assign w12819 = w12691 & ~w12818 ;
  assign w12820 = w12358 ^ w12819 ;
  assign w12821 = ( ~w6841 & w12809 ) | ( ~w6841 & w12815 ) | ( w12809 & w12815 ) ;
  assign w12822 = ~w12809 & w12821 ;
  assign w12823 = w12820 | w12822 ;
  assign w12824 = ( w6515 & w12817 ) | ( w6515 & ~w12823 ) | ( w12817 & ~w12823 ) ;
  assign w12825 = w6515 & w12824 ;
  assign w12826 = w12363 | w12368 ;
  assign w12827 = w12691 & ~w12826 ;
  assign w12828 = w12366 ^ w12827 ;
  assign w12829 = ( ~w6515 & w12817 ) | ( ~w6515 & w12823 ) | ( w12817 & w12823 ) ;
  assign w12830 = ~w12817 & w12829 ;
  assign w12831 = w12828 | w12830 ;
  assign w12832 = ( w6197 & w12825 ) | ( w6197 & ~w12831 ) | ( w12825 & ~w12831 ) ;
  assign w12833 = w6197 & w12832 ;
  assign w12834 = w12371 | w12376 ;
  assign w12835 = w12691 & ~w12834 ;
  assign w12836 = w12374 ^ w12835 ;
  assign w12837 = ( ~w6197 & w12825 ) | ( ~w6197 & w12831 ) | ( w12825 & w12831 ) ;
  assign w12838 = ~w12825 & w12837 ;
  assign w12839 = w12836 | w12838 ;
  assign w12840 = ( w5887 & w12833 ) | ( w5887 & ~w12839 ) | ( w12833 & ~w12839 ) ;
  assign w12841 = w5887 & w12840 ;
  assign w12842 = w12379 | w12384 ;
  assign w12843 = w12691 & ~w12842 ;
  assign w12844 = w12382 ^ w12843 ;
  assign w12845 = ( ~w5887 & w12833 ) | ( ~w5887 & w12839 ) | ( w12833 & w12839 ) ;
  assign w12846 = ~w12833 & w12845 ;
  assign w12847 = w12844 | w12846 ;
  assign w12848 = ( w5585 & w12841 ) | ( w5585 & ~w12847 ) | ( w12841 & ~w12847 ) ;
  assign w12849 = w5585 & w12848 ;
  assign w12850 = w12387 | w12392 ;
  assign w12851 = w12691 & ~w12850 ;
  assign w12852 = w12390 ^ w12851 ;
  assign w12853 = ( ~w5585 & w12841 ) | ( ~w5585 & w12847 ) | ( w12841 & w12847 ) ;
  assign w12854 = ~w12841 & w12853 ;
  assign w12855 = w12852 | w12854 ;
  assign w12856 = ( w5291 & w12849 ) | ( w5291 & ~w12855 ) | ( w12849 & ~w12855 ) ;
  assign w12857 = w5291 & w12856 ;
  assign w12858 = w12395 | w12400 ;
  assign w12859 = w12691 & ~w12858 ;
  assign w12860 = w12398 ^ w12859 ;
  assign w12861 = ( ~w5291 & w12849 ) | ( ~w5291 & w12855 ) | ( w12849 & w12855 ) ;
  assign w12862 = ~w12849 & w12861 ;
  assign w12863 = w12860 | w12862 ;
  assign w12864 = ( w5005 & w12857 ) | ( w5005 & ~w12863 ) | ( w12857 & ~w12863 ) ;
  assign w12865 = w5005 & w12864 ;
  assign w12866 = w12403 | w12408 ;
  assign w12867 = w12691 & ~w12866 ;
  assign w12868 = w12406 ^ w12867 ;
  assign w12869 = ( ~w5005 & w12857 ) | ( ~w5005 & w12863 ) | ( w12857 & w12863 ) ;
  assign w12870 = ~w12857 & w12869 ;
  assign w12871 = w12868 | w12870 ;
  assign w12872 = ( w4727 & w12865 ) | ( w4727 & ~w12871 ) | ( w12865 & ~w12871 ) ;
  assign w12873 = w4727 & w12872 ;
  assign w12874 = w12411 | w12416 ;
  assign w12875 = w12691 & ~w12874 ;
  assign w12876 = w12414 ^ w12875 ;
  assign w12877 = ( ~w4727 & w12865 ) | ( ~w4727 & w12871 ) | ( w12865 & w12871 ) ;
  assign w12878 = ~w12865 & w12877 ;
  assign w12879 = w12876 | w12878 ;
  assign w12880 = ( w4457 & w12873 ) | ( w4457 & ~w12879 ) | ( w12873 & ~w12879 ) ;
  assign w12881 = w4457 & w12880 ;
  assign w12882 = w12419 | w12424 ;
  assign w12883 = w12691 & ~w12882 ;
  assign w12884 = w12422 ^ w12883 ;
  assign w12885 = ( ~w4457 & w12873 ) | ( ~w4457 & w12879 ) | ( w12873 & w12879 ) ;
  assign w12886 = ~w12873 & w12885 ;
  assign w12887 = w12884 | w12886 ;
  assign w12888 = ( w4195 & w12881 ) | ( w4195 & ~w12887 ) | ( w12881 & ~w12887 ) ;
  assign w12889 = w4195 & w12888 ;
  assign w12890 = w12427 | w12432 ;
  assign w12891 = w12691 & ~w12890 ;
  assign w12892 = w12430 ^ w12891 ;
  assign w12893 = ( ~w4195 & w12881 ) | ( ~w4195 & w12887 ) | ( w12881 & w12887 ) ;
  assign w12894 = ~w12881 & w12893 ;
  assign w12895 = w12892 | w12894 ;
  assign w12896 = ( w3941 & w12889 ) | ( w3941 & ~w12895 ) | ( w12889 & ~w12895 ) ;
  assign w12897 = w3941 & w12896 ;
  assign w12898 = w12435 | w12440 ;
  assign w12899 = w12691 & ~w12898 ;
  assign w12900 = w12438 ^ w12899 ;
  assign w12901 = ( ~w3941 & w12889 ) | ( ~w3941 & w12895 ) | ( w12889 & w12895 ) ;
  assign w12902 = ~w12889 & w12901 ;
  assign w12903 = w12900 | w12902 ;
  assign w12904 = ( w3695 & w12897 ) | ( w3695 & ~w12903 ) | ( w12897 & ~w12903 ) ;
  assign w12905 = w3695 & w12904 ;
  assign w12906 = w12443 | w12448 ;
  assign w12907 = w12691 & ~w12906 ;
  assign w12908 = w12446 ^ w12907 ;
  assign w12909 = ( ~w3695 & w12897 ) | ( ~w3695 & w12903 ) | ( w12897 & w12903 ) ;
  assign w12910 = ~w12897 & w12909 ;
  assign w12911 = w12908 | w12910 ;
  assign w12912 = ( w3457 & w12905 ) | ( w3457 & ~w12911 ) | ( w12905 & ~w12911 ) ;
  assign w12913 = w3457 & w12912 ;
  assign w12914 = w12451 | w12456 ;
  assign w12915 = w12691 & ~w12914 ;
  assign w12916 = w12454 ^ w12915 ;
  assign w12917 = ( ~w3457 & w12905 ) | ( ~w3457 & w12911 ) | ( w12905 & w12911 ) ;
  assign w12918 = ~w12905 & w12917 ;
  assign w12919 = w12916 | w12918 ;
  assign w12920 = ( w3227 & w12913 ) | ( w3227 & ~w12919 ) | ( w12913 & ~w12919 ) ;
  assign w12921 = w3227 & w12920 ;
  assign w12922 = w12459 | w12464 ;
  assign w12923 = w12691 & ~w12922 ;
  assign w12924 = w12462 ^ w12923 ;
  assign w12925 = ( ~w3227 & w12913 ) | ( ~w3227 & w12919 ) | ( w12913 & w12919 ) ;
  assign w12926 = ~w12913 & w12925 ;
  assign w12927 = w12924 | w12926 ;
  assign w12928 = ( w3005 & w12921 ) | ( w3005 & ~w12927 ) | ( w12921 & ~w12927 ) ;
  assign w12929 = w3005 & w12928 ;
  assign w12930 = w12467 | w12472 ;
  assign w12931 = w12691 & ~w12930 ;
  assign w12932 = w12470 ^ w12931 ;
  assign w12933 = ( ~w3005 & w12921 ) | ( ~w3005 & w12927 ) | ( w12921 & w12927 ) ;
  assign w12934 = ~w12921 & w12933 ;
  assign w12935 = w12932 | w12934 ;
  assign w12936 = ( w2791 & w12929 ) | ( w2791 & ~w12935 ) | ( w12929 & ~w12935 ) ;
  assign w12937 = w2791 & w12936 ;
  assign w12938 = w12475 | w12480 ;
  assign w12939 = w12691 & ~w12938 ;
  assign w12940 = w12478 ^ w12939 ;
  assign w12941 = ( ~w2791 & w12929 ) | ( ~w2791 & w12935 ) | ( w12929 & w12935 ) ;
  assign w12942 = ~w12929 & w12941 ;
  assign w12943 = w12940 | w12942 ;
  assign w12944 = ( w2585 & w12937 ) | ( w2585 & ~w12943 ) | ( w12937 & ~w12943 ) ;
  assign w12945 = w2585 & w12944 ;
  assign w12946 = w12483 | w12488 ;
  assign w12947 = w12691 & ~w12946 ;
  assign w12948 = w12486 ^ w12947 ;
  assign w12949 = ( ~w2585 & w12937 ) | ( ~w2585 & w12943 ) | ( w12937 & w12943 ) ;
  assign w12950 = ~w12937 & w12949 ;
  assign w12951 = w12948 | w12950 ;
  assign w12952 = ( w2387 & w12945 ) | ( w2387 & ~w12951 ) | ( w12945 & ~w12951 ) ;
  assign w12953 = w2387 & w12952 ;
  assign w12954 = w12491 | w12496 ;
  assign w12955 = w12691 & ~w12954 ;
  assign w12956 = w12494 ^ w12955 ;
  assign w12957 = ( ~w2387 & w12945 ) | ( ~w2387 & w12951 ) | ( w12945 & w12951 ) ;
  assign w12958 = ~w12945 & w12957 ;
  assign w12959 = w12956 | w12958 ;
  assign w12960 = ( w2197 & w12953 ) | ( w2197 & ~w12959 ) | ( w12953 & ~w12959 ) ;
  assign w12961 = w2197 & w12960 ;
  assign w12962 = w12499 | w12504 ;
  assign w12963 = w12691 & ~w12962 ;
  assign w12964 = w12502 ^ w12963 ;
  assign w12965 = ( ~w2197 & w12953 ) | ( ~w2197 & w12959 ) | ( w12953 & w12959 ) ;
  assign w12966 = ~w12953 & w12965 ;
  assign w12967 = w12964 | w12966 ;
  assign w12968 = ( w2015 & w12961 ) | ( w2015 & ~w12967 ) | ( w12961 & ~w12967 ) ;
  assign w12969 = w2015 & w12968 ;
  assign w12970 = w12507 | w12512 ;
  assign w12971 = w12691 & ~w12970 ;
  assign w12972 = w12510 ^ w12971 ;
  assign w12973 = ( ~w2015 & w12961 ) | ( ~w2015 & w12967 ) | ( w12961 & w12967 ) ;
  assign w12974 = ~w12961 & w12973 ;
  assign w12975 = w12972 | w12974 ;
  assign w12976 = ( w1841 & w12969 ) | ( w1841 & ~w12975 ) | ( w12969 & ~w12975 ) ;
  assign w12977 = w1841 & w12976 ;
  assign w12978 = w12515 | w12520 ;
  assign w12979 = w12691 & ~w12978 ;
  assign w12980 = w12518 ^ w12979 ;
  assign w12981 = ( ~w1841 & w12969 ) | ( ~w1841 & w12975 ) | ( w12969 & w12975 ) ;
  assign w12982 = ~w12969 & w12981 ;
  assign w12983 = w12980 | w12982 ;
  assign w12984 = ( w1675 & w12977 ) | ( w1675 & ~w12983 ) | ( w12977 & ~w12983 ) ;
  assign w12985 = w1675 & w12984 ;
  assign w12986 = w12523 | w12528 ;
  assign w12987 = w12691 & ~w12986 ;
  assign w12988 = w12526 ^ w12987 ;
  assign w12989 = ( ~w1675 & w12977 ) | ( ~w1675 & w12983 ) | ( w12977 & w12983 ) ;
  assign w12990 = ~w12977 & w12989 ;
  assign w12991 = w12988 | w12990 ;
  assign w12992 = ( w1517 & w12985 ) | ( w1517 & ~w12991 ) | ( w12985 & ~w12991 ) ;
  assign w12993 = w1517 & w12992 ;
  assign w12994 = w12531 | w12536 ;
  assign w12995 = w12691 & ~w12994 ;
  assign w12996 = w12534 ^ w12995 ;
  assign w12997 = ( ~w1517 & w12985 ) | ( ~w1517 & w12991 ) | ( w12985 & w12991 ) ;
  assign w12998 = ~w12985 & w12997 ;
  assign w12999 = w12996 | w12998 ;
  assign w13000 = ( w1367 & w12993 ) | ( w1367 & ~w12999 ) | ( w12993 & ~w12999 ) ;
  assign w13001 = w1367 & w13000 ;
  assign w13002 = w12539 | w12544 ;
  assign w13003 = w12691 & ~w13002 ;
  assign w13004 = w12542 ^ w13003 ;
  assign w13005 = ( ~w1367 & w12993 ) | ( ~w1367 & w12999 ) | ( w12993 & w12999 ) ;
  assign w13006 = ~w12993 & w13005 ;
  assign w13007 = w13004 | w13006 ;
  assign w13008 = ( w1225 & w13001 ) | ( w1225 & ~w13007 ) | ( w13001 & ~w13007 ) ;
  assign w13009 = w1225 & w13008 ;
  assign w13010 = w12547 | w12552 ;
  assign w13011 = w12691 & ~w13010 ;
  assign w13012 = w12550 ^ w13011 ;
  assign w13013 = ( ~w1225 & w13001 ) | ( ~w1225 & w13007 ) | ( w13001 & w13007 ) ;
  assign w13014 = ~w13001 & w13013 ;
  assign w13015 = w13012 | w13014 ;
  assign w13016 = ( w1091 & w13009 ) | ( w1091 & ~w13015 ) | ( w13009 & ~w13015 ) ;
  assign w13017 = w1091 & w13016 ;
  assign w13018 = w12555 | w12560 ;
  assign w13019 = w12691 & ~w13018 ;
  assign w13020 = w12558 ^ w13019 ;
  assign w13021 = ( ~w1091 & w13009 ) | ( ~w1091 & w13015 ) | ( w13009 & w13015 ) ;
  assign w13022 = ~w13009 & w13021 ;
  assign w13023 = w13020 | w13022 ;
  assign w13024 = ( w965 & w13017 ) | ( w965 & ~w13023 ) | ( w13017 & ~w13023 ) ;
  assign w13025 = w965 & w13024 ;
  assign w13026 = w12563 | w12568 ;
  assign w13027 = w12691 & ~w13026 ;
  assign w13028 = w12566 ^ w13027 ;
  assign w13029 = ( ~w965 & w13017 ) | ( ~w965 & w13023 ) | ( w13017 & w13023 ) ;
  assign w13030 = ~w13017 & w13029 ;
  assign w13031 = w13028 | w13030 ;
  assign w13032 = ( w847 & w13025 ) | ( w847 & ~w13031 ) | ( w13025 & ~w13031 ) ;
  assign w13033 = w847 & w13032 ;
  assign w13034 = w12571 | w12576 ;
  assign w13035 = w12691 & ~w13034 ;
  assign w13036 = w12574 ^ w13035 ;
  assign w13037 = ( ~w847 & w13025 ) | ( ~w847 & w13031 ) | ( w13025 & w13031 ) ;
  assign w13038 = ~w13025 & w13037 ;
  assign w13039 = w13036 | w13038 ;
  assign w13040 = ( w737 & w13033 ) | ( w737 & ~w13039 ) | ( w13033 & ~w13039 ) ;
  assign w13041 = w737 & w13040 ;
  assign w13042 = w12579 | w12584 ;
  assign w13043 = w12691 & ~w13042 ;
  assign w13044 = w12582 ^ w13043 ;
  assign w13045 = ( ~w737 & w13033 ) | ( ~w737 & w13039 ) | ( w13033 & w13039 ) ;
  assign w13046 = ~w13033 & w13045 ;
  assign w13047 = w13044 | w13046 ;
  assign w13048 = ( w635 & w13041 ) | ( w635 & ~w13047 ) | ( w13041 & ~w13047 ) ;
  assign w13049 = w635 & w13048 ;
  assign w13050 = w12587 | w12592 ;
  assign w13051 = w12691 & ~w13050 ;
  assign w13052 = w12590 ^ w13051 ;
  assign w13053 = ( ~w635 & w13041 ) | ( ~w635 & w13047 ) | ( w13041 & w13047 ) ;
  assign w13054 = ~w13041 & w13053 ;
  assign w13055 = w13052 | w13054 ;
  assign w13056 = ( w541 & w13049 ) | ( w541 & ~w13055 ) | ( w13049 & ~w13055 ) ;
  assign w13057 = w541 & w13056 ;
  assign w13058 = ( ~w541 & w13049 ) | ( ~w541 & w13055 ) | ( w13049 & w13055 ) ;
  assign w13059 = ~w13049 & w13058 ;
  assign w13060 = w12595 | w12597 ;
  assign w13061 = w12691 & ~w13060 ;
  assign w13062 = w12600 ^ w13061 ;
  assign w13063 = w13059 | w13062 ;
  assign w13064 = ( w455 & w13057 ) | ( w455 & ~w13063 ) | ( w13057 & ~w13063 ) ;
  assign w13065 = w455 & w13064 ;
  assign w13066 = w12603 | w12608 ;
  assign w13067 = w12691 & ~w13066 ;
  assign w13068 = w12606 ^ w13067 ;
  assign w13069 = ( ~w455 & w13057 ) | ( ~w455 & w13063 ) | ( w13057 & w13063 ) ;
  assign w13070 = ~w13057 & w13069 ;
  assign w13071 = w13068 | w13070 ;
  assign w13072 = ( w377 & w13065 ) | ( w377 & ~w13071 ) | ( w13065 & ~w13071 ) ;
  assign w13073 = w377 & w13072 ;
  assign w13074 = w12611 | w12616 ;
  assign w13075 = w12691 & ~w13074 ;
  assign w13076 = w12614 ^ w13075 ;
  assign w13077 = ( ~w377 & w13065 ) | ( ~w377 & w13071 ) | ( w13065 & w13071 ) ;
  assign w13078 = ~w13065 & w13077 ;
  assign w13079 = w13076 | w13078 ;
  assign w13080 = ( w307 & w13073 ) | ( w307 & ~w13079 ) | ( w13073 & ~w13079 ) ;
  assign w13081 = w307 & w13080 ;
  assign w13082 = w12619 | w12624 ;
  assign w13083 = w12691 & ~w13082 ;
  assign w13084 = w12622 ^ w13083 ;
  assign w13085 = ( ~w307 & w13073 ) | ( ~w307 & w13079 ) | ( w13073 & w13079 ) ;
  assign w13086 = ~w13073 & w13085 ;
  assign w13087 = w13084 | w13086 ;
  assign w13088 = ( w246 & w13081 ) | ( w246 & ~w13087 ) | ( w13081 & ~w13087 ) ;
  assign w13089 = w246 & w13088 ;
  assign w13090 = w12627 | w12632 ;
  assign w13091 = w12691 & ~w13090 ;
  assign w13092 = w12630 ^ w13091 ;
  assign w13093 = ( ~w246 & w13081 ) | ( ~w246 & w13087 ) | ( w13081 & w13087 ) ;
  assign w13094 = ~w13081 & w13093 ;
  assign w13095 = w13092 | w13094 ;
  assign w13096 = ( w185 & w13089 ) | ( w185 & ~w13095 ) | ( w13089 & ~w13095 ) ;
  assign w13097 = w185 & w13096 ;
  assign w13098 = w12635 | w12640 ;
  assign w13099 = w12691 & ~w13098 ;
  assign w13100 = w12638 ^ w13099 ;
  assign w13101 = ( ~w185 & w13089 ) | ( ~w185 & w13095 ) | ( w13089 & w13095 ) ;
  assign w13102 = ~w13089 & w13101 ;
  assign w13103 = w13100 | w13102 ;
  assign w13104 = ( w145 & w13097 ) | ( w145 & ~w13103 ) | ( w13097 & ~w13103 ) ;
  assign w13105 = w145 & w13104 ;
  assign w13106 = w12643 | w12648 ;
  assign w13107 = w12691 & ~w13106 ;
  assign w13108 = w12646 ^ w13107 ;
  assign w13109 = ( ~w145 & w13097 ) | ( ~w145 & w13103 ) | ( w13097 & w13103 ) ;
  assign w13110 = ~w13097 & w13109 ;
  assign w13111 = w13108 | w13110 ;
  assign w13112 = ( w132 & w13105 ) | ( w132 & ~w13111 ) | ( w13105 & ~w13111 ) ;
  assign w13113 = w132 & w13112 ;
  assign w13114 = w12651 | w12656 ;
  assign w13115 = w12691 & ~w13114 ;
  assign w13116 = w12654 ^ w13115 ;
  assign w13117 = ( ~w132 & w13105 ) | ( ~w132 & w13111 ) | ( w13105 & w13111 ) ;
  assign w13118 = ~w13105 & w13117 ;
  assign w13119 = w13116 | w13118 ;
  assign w13120 = ~w13113 & w13119 ;
  assign w13121 = w12659 | w12664 ;
  assign w13122 = w12691 & ~w13121 ;
  assign w13123 = w12662 ^ w13122 ;
  assign w13124 = ( ~w12677 & w13120 ) | ( ~w12677 & w13123 ) | ( w13120 & w13123 ) ;
  assign w13125 = w12666 & ~w13124 ;
  assign w13126 = ~w12669 & w12691 ;
  assign w13127 = ( w13124 & ~w13125 ) | ( w13124 & w13126 ) | ( ~w13125 & w13126 ) ;
  assign w13128 = w12677 | w13127 ;
  assign w13129 = ~w129 & w13128 ;
  assign w13130 = ( w13113 & w13119 ) | ( w13113 & w13123 ) | ( w13119 & w13123 ) ;
  assign w13131 = ~w13113 & w13130 ;
  assign w13132 = ( w129 & w12666 ) | ( w129 & w12669 ) | ( w12666 & w12669 ) ;
  assign w13133 = ( w12669 & ~w12691 ) | ( w12669 & w13132 ) | ( ~w12691 & w13132 ) ;
  assign w13134 = w12666 & w13133 ;
  assign w13135 = w13132 ^ w13134 ;
  assign w13136 = ( w12213 & w12218 ) | ( w12213 & w12245 ) | ( w12218 & w12245 ) ;
  assign w13137 = w12245 & ~w13136 ;
  assign w13138 = w12216 ^ w13137 ;
  assign w13139 = ( ~w12681 & w12688 ) | ( ~w12681 & w13138 ) | ( w12688 & w13138 ) ;
  assign w13140 = ~w12688 & w13139 ;
  assign w13141 = ( ~w12675 & w12677 ) | ( ~w12675 & w13140 ) | ( w12677 & w13140 ) ;
  assign w13142 = ~w12677 & w13141 ;
  assign w13143 = w13131 | w13142 ;
  assign w13144 = ( w13129 & ~w13131 ) | ( w13129 & w13135 ) | ( ~w13131 & w13135 ) ;
  assign w13145 = w13143 | w13144 ;
  assign w13146 = ( ~\pi017 & \pi018 ) | ( ~\pi017 & w12691 ) | ( \pi018 & w12691 ) ;
  assign w13147 = ( ~\pi016 & \pi018 ) | ( ~\pi016 & w13146 ) | ( \pi018 & w13146 ) ;
  assign w13148 = ( ~\pi018 & w12691 ) | ( ~\pi018 & w13145 ) | ( w12691 & w13145 ) ;
  assign w13149 = w13147 & w13148 ;
  assign w13150 = ( w12677 & w12681 ) | ( w12677 & ~w12688 ) | ( w12681 & ~w12688 ) ;
  assign w13151 = \pi017 & ~w13150 ;
  assign w13152 = \pi016 | \pi018 ;
  assign w13153 = ( ~w13150 & w13151 ) | ( ~w13150 & w13152 ) | ( w13151 & w13152 ) ;
  assign w13154 = ~w12688 & w13153 ;
  assign w13155 = ~w12675 & w13154 ;
  assign w13156 = ( \pi018 & w13145 ) | ( \pi018 & ~w13154 ) | ( w13145 & ~w13154 ) ;
  assign w13157 = w13155 & ~w13156 ;
  assign w13158 = ~\pi018 & w13145 ;
  assign w13159 = \pi019 ^ w13158 ;
  assign w13160 = w13157 | w13159 ;
  assign w13161 = ( w12245 & w13149 ) | ( w12245 & ~w13160 ) | ( w13149 & ~w13160 ) ;
  assign w13162 = w12245 & w13161 ;
  assign w13163 = ( ~w12245 & w13149 ) | ( ~w12245 & w13160 ) | ( w13149 & w13160 ) ;
  assign w13164 = ~w13149 & w13163 ;
  assign w13165 = w12691 & ~w13142 ;
  assign w13166 = ~w13131 & w13165 ;
  assign w13167 = ~w13144 & w13166 ;
  assign w13168 = \pi019 & w13145 ;
  assign w13169 = ( \pi018 & w13145 ) | ( \pi018 & ~w13168 ) | ( w13145 & ~w13168 ) ;
  assign w13170 = ( ~\pi018 & w13167 ) | ( ~\pi018 & w13169 ) | ( w13167 & w13169 ) ;
  assign w13171 = \pi020 ^ w13170 ;
  assign w13172 = w13164 | w13171 ;
  assign w13173 = ( w11807 & w13162 ) | ( w11807 & ~w13172 ) | ( w13162 & ~w13172 ) ;
  assign w13174 = w11807 & w13173 ;
  assign w13175 = ( w12695 & ~w12703 ) | ( w12695 & w13145 ) | ( ~w12703 & w13145 ) ;
  assign w13176 = ~w12695 & w13175 ;
  assign w13177 = \pi021 ^ w13176 ;
  assign w13178 = w12704 ^ w13177 ;
  assign w13179 = ( ~w11807 & w13162 ) | ( ~w11807 & w13172 ) | ( w13162 & w13172 ) ;
  assign w13180 = ~w13162 & w13179 ;
  assign w13181 = w13178 | w13180 ;
  assign w13182 = ( w11377 & w13174 ) | ( w11377 & ~w13181 ) | ( w13174 & ~w13181 ) ;
  assign w13183 = w11377 & w13182 ;
  assign w13184 = w12708 | w12710 ;
  assign w13185 = w13145 & ~w13184 ;
  assign w13186 = w12717 ^ w13185 ;
  assign w13187 = ( ~w11377 & w13174 ) | ( ~w11377 & w13181 ) | ( w13174 & w13181 ) ;
  assign w13188 = ~w13174 & w13187 ;
  assign w13189 = w13186 | w13188 ;
  assign w13190 = ( w10955 & w13183 ) | ( w10955 & ~w13189 ) | ( w13183 & ~w13189 ) ;
  assign w13191 = w10955 & w13190 ;
  assign w13192 = w12720 | w12726 ;
  assign w13193 = w13145 & ~w13192 ;
  assign w13194 = w12724 ^ w13193 ;
  assign w13195 = ( ~w10955 & w13183 ) | ( ~w10955 & w13189 ) | ( w13183 & w13189 ) ;
  assign w13196 = ~w13183 & w13195 ;
  assign w13197 = w13194 | w13196 ;
  assign w13198 = ( w10541 & w13191 ) | ( w10541 & ~w13197 ) | ( w13191 & ~w13197 ) ;
  assign w13199 = w10541 & w13198 ;
  assign w13200 = w12729 | w12734 ;
  assign w13201 = w13145 & ~w13200 ;
  assign w13202 = w12732 ^ w13201 ;
  assign w13203 = ( ~w10541 & w13191 ) | ( ~w10541 & w13197 ) | ( w13191 & w13197 ) ;
  assign w13204 = ~w13191 & w13203 ;
  assign w13205 = w13202 | w13204 ;
  assign w13206 = ( w10135 & w13199 ) | ( w10135 & ~w13205 ) | ( w13199 & ~w13205 ) ;
  assign w13207 = w10135 & w13206 ;
  assign w13208 = w12737 | w12742 ;
  assign w13209 = w13145 & ~w13208 ;
  assign w13210 = w12740 ^ w13209 ;
  assign w13211 = ( ~w10135 & w13199 ) | ( ~w10135 & w13205 ) | ( w13199 & w13205 ) ;
  assign w13212 = ~w13199 & w13211 ;
  assign w13213 = w13210 | w13212 ;
  assign w13214 = ( w9737 & w13207 ) | ( w9737 & ~w13213 ) | ( w13207 & ~w13213 ) ;
  assign w13215 = w9737 & w13214 ;
  assign w13216 = w12745 | w12750 ;
  assign w13217 = w13145 & ~w13216 ;
  assign w13218 = w12748 ^ w13217 ;
  assign w13219 = ( ~w9737 & w13207 ) | ( ~w9737 & w13213 ) | ( w13207 & w13213 ) ;
  assign w13220 = ~w13207 & w13219 ;
  assign w13221 = w13218 | w13220 ;
  assign w13222 = ( w9347 & w13215 ) | ( w9347 & ~w13221 ) | ( w13215 & ~w13221 ) ;
  assign w13223 = w9347 & w13222 ;
  assign w13224 = w12753 | w12758 ;
  assign w13225 = w13145 & ~w13224 ;
  assign w13226 = w12756 ^ w13225 ;
  assign w13227 = ( ~w9347 & w13215 ) | ( ~w9347 & w13221 ) | ( w13215 & w13221 ) ;
  assign w13228 = ~w13215 & w13227 ;
  assign w13229 = w13226 | w13228 ;
  assign w13230 = ( w8965 & w13223 ) | ( w8965 & ~w13229 ) | ( w13223 & ~w13229 ) ;
  assign w13231 = w8965 & w13230 ;
  assign w13232 = w12761 | w12766 ;
  assign w13233 = w13145 & ~w13232 ;
  assign w13234 = w12764 ^ w13233 ;
  assign w13235 = ( ~w8965 & w13223 ) | ( ~w8965 & w13229 ) | ( w13223 & w13229 ) ;
  assign w13236 = ~w13223 & w13235 ;
  assign w13237 = w13234 | w13236 ;
  assign w13238 = ( w8591 & w13231 ) | ( w8591 & ~w13237 ) | ( w13231 & ~w13237 ) ;
  assign w13239 = w8591 & w13238 ;
  assign w13240 = w12769 | w12774 ;
  assign w13241 = w13145 & ~w13240 ;
  assign w13242 = w12772 ^ w13241 ;
  assign w13243 = ( ~w8591 & w13231 ) | ( ~w8591 & w13237 ) | ( w13231 & w13237 ) ;
  assign w13244 = ~w13231 & w13243 ;
  assign w13245 = w13242 | w13244 ;
  assign w13246 = ( w8225 & w13239 ) | ( w8225 & ~w13245 ) | ( w13239 & ~w13245 ) ;
  assign w13247 = w8225 & w13246 ;
  assign w13248 = w12777 | w12782 ;
  assign w13249 = w13145 & ~w13248 ;
  assign w13250 = w12780 ^ w13249 ;
  assign w13251 = ( ~w8225 & w13239 ) | ( ~w8225 & w13245 ) | ( w13239 & w13245 ) ;
  assign w13252 = ~w13239 & w13251 ;
  assign w13253 = w13250 | w13252 ;
  assign w13254 = ( w7867 & w13247 ) | ( w7867 & ~w13253 ) | ( w13247 & ~w13253 ) ;
  assign w13255 = w7867 & w13254 ;
  assign w13256 = w12785 | w12790 ;
  assign w13257 = w13145 & ~w13256 ;
  assign w13258 = w12788 ^ w13257 ;
  assign w13259 = ( ~w7867 & w13247 ) | ( ~w7867 & w13253 ) | ( w13247 & w13253 ) ;
  assign w13260 = ~w13247 & w13259 ;
  assign w13261 = w13258 | w13260 ;
  assign w13262 = ( w7517 & w13255 ) | ( w7517 & ~w13261 ) | ( w13255 & ~w13261 ) ;
  assign w13263 = w7517 & w13262 ;
  assign w13264 = w12793 | w12798 ;
  assign w13265 = w13145 & ~w13264 ;
  assign w13266 = w12796 ^ w13265 ;
  assign w13267 = ( ~w7517 & w13255 ) | ( ~w7517 & w13261 ) | ( w13255 & w13261 ) ;
  assign w13268 = ~w13255 & w13267 ;
  assign w13269 = w13266 | w13268 ;
  assign w13270 = ( w7175 & w13263 ) | ( w7175 & ~w13269 ) | ( w13263 & ~w13269 ) ;
  assign w13271 = w7175 & w13270 ;
  assign w13272 = w12801 | w12806 ;
  assign w13273 = w13145 & ~w13272 ;
  assign w13274 = w12804 ^ w13273 ;
  assign w13275 = ( ~w7175 & w13263 ) | ( ~w7175 & w13269 ) | ( w13263 & w13269 ) ;
  assign w13276 = ~w13263 & w13275 ;
  assign w13277 = w13274 | w13276 ;
  assign w13278 = ( w6841 & w13271 ) | ( w6841 & ~w13277 ) | ( w13271 & ~w13277 ) ;
  assign w13279 = w6841 & w13278 ;
  assign w13280 = w12809 | w12814 ;
  assign w13281 = w13145 & ~w13280 ;
  assign w13282 = w12812 ^ w13281 ;
  assign w13283 = ( ~w6841 & w13271 ) | ( ~w6841 & w13277 ) | ( w13271 & w13277 ) ;
  assign w13284 = ~w13271 & w13283 ;
  assign w13285 = w13282 | w13284 ;
  assign w13286 = ( w6515 & w13279 ) | ( w6515 & ~w13285 ) | ( w13279 & ~w13285 ) ;
  assign w13287 = w6515 & w13286 ;
  assign w13288 = w12817 | w12822 ;
  assign w13289 = w13145 & ~w13288 ;
  assign w13290 = w12820 ^ w13289 ;
  assign w13291 = ( ~w6515 & w13279 ) | ( ~w6515 & w13285 ) | ( w13279 & w13285 ) ;
  assign w13292 = ~w13279 & w13291 ;
  assign w13293 = w13290 | w13292 ;
  assign w13294 = ( w6197 & w13287 ) | ( w6197 & ~w13293 ) | ( w13287 & ~w13293 ) ;
  assign w13295 = w6197 & w13294 ;
  assign w13296 = w12825 | w12830 ;
  assign w13297 = w13145 & ~w13296 ;
  assign w13298 = w12828 ^ w13297 ;
  assign w13299 = ( ~w6197 & w13287 ) | ( ~w6197 & w13293 ) | ( w13287 & w13293 ) ;
  assign w13300 = ~w13287 & w13299 ;
  assign w13301 = w13298 | w13300 ;
  assign w13302 = ( w5887 & w13295 ) | ( w5887 & ~w13301 ) | ( w13295 & ~w13301 ) ;
  assign w13303 = w5887 & w13302 ;
  assign w13304 = w12833 | w12838 ;
  assign w13305 = w13145 & ~w13304 ;
  assign w13306 = w12836 ^ w13305 ;
  assign w13307 = ( ~w5887 & w13295 ) | ( ~w5887 & w13301 ) | ( w13295 & w13301 ) ;
  assign w13308 = ~w13295 & w13307 ;
  assign w13309 = w13306 | w13308 ;
  assign w13310 = ( w5585 & w13303 ) | ( w5585 & ~w13309 ) | ( w13303 & ~w13309 ) ;
  assign w13311 = w5585 & w13310 ;
  assign w13312 = w12841 | w12846 ;
  assign w13313 = w13145 & ~w13312 ;
  assign w13314 = w12844 ^ w13313 ;
  assign w13315 = ( ~w5585 & w13303 ) | ( ~w5585 & w13309 ) | ( w13303 & w13309 ) ;
  assign w13316 = ~w13303 & w13315 ;
  assign w13317 = w13314 | w13316 ;
  assign w13318 = ( w5291 & w13311 ) | ( w5291 & ~w13317 ) | ( w13311 & ~w13317 ) ;
  assign w13319 = w5291 & w13318 ;
  assign w13320 = w12849 | w12854 ;
  assign w13321 = w13145 & ~w13320 ;
  assign w13322 = w12852 ^ w13321 ;
  assign w13323 = ( ~w5291 & w13311 ) | ( ~w5291 & w13317 ) | ( w13311 & w13317 ) ;
  assign w13324 = ~w13311 & w13323 ;
  assign w13325 = w13322 | w13324 ;
  assign w13326 = ( w5005 & w13319 ) | ( w5005 & ~w13325 ) | ( w13319 & ~w13325 ) ;
  assign w13327 = w5005 & w13326 ;
  assign w13328 = w12857 | w12862 ;
  assign w13329 = w13145 & ~w13328 ;
  assign w13330 = w12860 ^ w13329 ;
  assign w13331 = ( ~w5005 & w13319 ) | ( ~w5005 & w13325 ) | ( w13319 & w13325 ) ;
  assign w13332 = ~w13319 & w13331 ;
  assign w13333 = w13330 | w13332 ;
  assign w13334 = ( w4727 & w13327 ) | ( w4727 & ~w13333 ) | ( w13327 & ~w13333 ) ;
  assign w13335 = w4727 & w13334 ;
  assign w13336 = w12865 | w12870 ;
  assign w13337 = w13145 & ~w13336 ;
  assign w13338 = w12868 ^ w13337 ;
  assign w13339 = ( ~w4727 & w13327 ) | ( ~w4727 & w13333 ) | ( w13327 & w13333 ) ;
  assign w13340 = ~w13327 & w13339 ;
  assign w13341 = w13338 | w13340 ;
  assign w13342 = ( w4457 & w13335 ) | ( w4457 & ~w13341 ) | ( w13335 & ~w13341 ) ;
  assign w13343 = w4457 & w13342 ;
  assign w13344 = w12873 | w12878 ;
  assign w13345 = w13145 & ~w13344 ;
  assign w13346 = w12876 ^ w13345 ;
  assign w13347 = ( ~w4457 & w13335 ) | ( ~w4457 & w13341 ) | ( w13335 & w13341 ) ;
  assign w13348 = ~w13335 & w13347 ;
  assign w13349 = w13346 | w13348 ;
  assign w13350 = ( w4195 & w13343 ) | ( w4195 & ~w13349 ) | ( w13343 & ~w13349 ) ;
  assign w13351 = w4195 & w13350 ;
  assign w13352 = w12881 | w12886 ;
  assign w13353 = w13145 & ~w13352 ;
  assign w13354 = w12884 ^ w13353 ;
  assign w13355 = ( ~w4195 & w13343 ) | ( ~w4195 & w13349 ) | ( w13343 & w13349 ) ;
  assign w13356 = ~w13343 & w13355 ;
  assign w13357 = w13354 | w13356 ;
  assign w13358 = ( w3941 & w13351 ) | ( w3941 & ~w13357 ) | ( w13351 & ~w13357 ) ;
  assign w13359 = w3941 & w13358 ;
  assign w13360 = w12889 | w12894 ;
  assign w13361 = w13145 & ~w13360 ;
  assign w13362 = w12892 ^ w13361 ;
  assign w13363 = ( ~w3941 & w13351 ) | ( ~w3941 & w13357 ) | ( w13351 & w13357 ) ;
  assign w13364 = ~w13351 & w13363 ;
  assign w13365 = w13362 | w13364 ;
  assign w13366 = ( w3695 & w13359 ) | ( w3695 & ~w13365 ) | ( w13359 & ~w13365 ) ;
  assign w13367 = w3695 & w13366 ;
  assign w13368 = w12897 | w12902 ;
  assign w13369 = w13145 & ~w13368 ;
  assign w13370 = w12900 ^ w13369 ;
  assign w13371 = ( ~w3695 & w13359 ) | ( ~w3695 & w13365 ) | ( w13359 & w13365 ) ;
  assign w13372 = ~w13359 & w13371 ;
  assign w13373 = w13370 | w13372 ;
  assign w13374 = ( w3457 & w13367 ) | ( w3457 & ~w13373 ) | ( w13367 & ~w13373 ) ;
  assign w13375 = w3457 & w13374 ;
  assign w13376 = w12905 | w12910 ;
  assign w13377 = w13145 & ~w13376 ;
  assign w13378 = w12908 ^ w13377 ;
  assign w13379 = ( ~w3457 & w13367 ) | ( ~w3457 & w13373 ) | ( w13367 & w13373 ) ;
  assign w13380 = ~w13367 & w13379 ;
  assign w13381 = w13378 | w13380 ;
  assign w13382 = ( w3227 & w13375 ) | ( w3227 & ~w13381 ) | ( w13375 & ~w13381 ) ;
  assign w13383 = w3227 & w13382 ;
  assign w13384 = w12913 | w12918 ;
  assign w13385 = w13145 & ~w13384 ;
  assign w13386 = w12916 ^ w13385 ;
  assign w13387 = ( ~w3227 & w13375 ) | ( ~w3227 & w13381 ) | ( w13375 & w13381 ) ;
  assign w13388 = ~w13375 & w13387 ;
  assign w13389 = w13386 | w13388 ;
  assign w13390 = ( w3005 & w13383 ) | ( w3005 & ~w13389 ) | ( w13383 & ~w13389 ) ;
  assign w13391 = w3005 & w13390 ;
  assign w13392 = w12921 | w12926 ;
  assign w13393 = w13145 & ~w13392 ;
  assign w13394 = w12924 ^ w13393 ;
  assign w13395 = ( ~w3005 & w13383 ) | ( ~w3005 & w13389 ) | ( w13383 & w13389 ) ;
  assign w13396 = ~w13383 & w13395 ;
  assign w13397 = w13394 | w13396 ;
  assign w13398 = ( w2791 & w13391 ) | ( w2791 & ~w13397 ) | ( w13391 & ~w13397 ) ;
  assign w13399 = w2791 & w13398 ;
  assign w13400 = w12929 | w12934 ;
  assign w13401 = w13145 & ~w13400 ;
  assign w13402 = w12932 ^ w13401 ;
  assign w13403 = ( ~w2791 & w13391 ) | ( ~w2791 & w13397 ) | ( w13391 & w13397 ) ;
  assign w13404 = ~w13391 & w13403 ;
  assign w13405 = w13402 | w13404 ;
  assign w13406 = ( w2585 & w13399 ) | ( w2585 & ~w13405 ) | ( w13399 & ~w13405 ) ;
  assign w13407 = w2585 & w13406 ;
  assign w13408 = w12937 | w12942 ;
  assign w13409 = w13145 & ~w13408 ;
  assign w13410 = w12940 ^ w13409 ;
  assign w13411 = ( ~w2585 & w13399 ) | ( ~w2585 & w13405 ) | ( w13399 & w13405 ) ;
  assign w13412 = ~w13399 & w13411 ;
  assign w13413 = w13410 | w13412 ;
  assign w13414 = ( w2387 & w13407 ) | ( w2387 & ~w13413 ) | ( w13407 & ~w13413 ) ;
  assign w13415 = w2387 & w13414 ;
  assign w13416 = w12945 | w12950 ;
  assign w13417 = w13145 & ~w13416 ;
  assign w13418 = w12948 ^ w13417 ;
  assign w13419 = ( ~w2387 & w13407 ) | ( ~w2387 & w13413 ) | ( w13407 & w13413 ) ;
  assign w13420 = ~w13407 & w13419 ;
  assign w13421 = w13418 | w13420 ;
  assign w13422 = ( w2197 & w13415 ) | ( w2197 & ~w13421 ) | ( w13415 & ~w13421 ) ;
  assign w13423 = w2197 & w13422 ;
  assign w13424 = w12953 | w12958 ;
  assign w13425 = w13145 & ~w13424 ;
  assign w13426 = w12956 ^ w13425 ;
  assign w13427 = ( ~w2197 & w13415 ) | ( ~w2197 & w13421 ) | ( w13415 & w13421 ) ;
  assign w13428 = ~w13415 & w13427 ;
  assign w13429 = w13426 | w13428 ;
  assign w13430 = ( w2015 & w13423 ) | ( w2015 & ~w13429 ) | ( w13423 & ~w13429 ) ;
  assign w13431 = w2015 & w13430 ;
  assign w13432 = w12961 | w12966 ;
  assign w13433 = w13145 & ~w13432 ;
  assign w13434 = w12964 ^ w13433 ;
  assign w13435 = ( ~w2015 & w13423 ) | ( ~w2015 & w13429 ) | ( w13423 & w13429 ) ;
  assign w13436 = ~w13423 & w13435 ;
  assign w13437 = w13434 | w13436 ;
  assign w13438 = ( w1841 & w13431 ) | ( w1841 & ~w13437 ) | ( w13431 & ~w13437 ) ;
  assign w13439 = w1841 & w13438 ;
  assign w13440 = w12969 | w12974 ;
  assign w13441 = w13145 & ~w13440 ;
  assign w13442 = w12972 ^ w13441 ;
  assign w13443 = ( ~w1841 & w13431 ) | ( ~w1841 & w13437 ) | ( w13431 & w13437 ) ;
  assign w13444 = ~w13431 & w13443 ;
  assign w13445 = w13442 | w13444 ;
  assign w13446 = ( w1675 & w13439 ) | ( w1675 & ~w13445 ) | ( w13439 & ~w13445 ) ;
  assign w13447 = w1675 & w13446 ;
  assign w13448 = w12977 | w12982 ;
  assign w13449 = w13145 & ~w13448 ;
  assign w13450 = w12980 ^ w13449 ;
  assign w13451 = ( ~w1675 & w13439 ) | ( ~w1675 & w13445 ) | ( w13439 & w13445 ) ;
  assign w13452 = ~w13439 & w13451 ;
  assign w13453 = w13450 | w13452 ;
  assign w13454 = ( w1517 & w13447 ) | ( w1517 & ~w13453 ) | ( w13447 & ~w13453 ) ;
  assign w13455 = w1517 & w13454 ;
  assign w13456 = w12985 | w12990 ;
  assign w13457 = w13145 & ~w13456 ;
  assign w13458 = w12988 ^ w13457 ;
  assign w13459 = ( ~w1517 & w13447 ) | ( ~w1517 & w13453 ) | ( w13447 & w13453 ) ;
  assign w13460 = ~w13447 & w13459 ;
  assign w13461 = w13458 | w13460 ;
  assign w13462 = ( w1367 & w13455 ) | ( w1367 & ~w13461 ) | ( w13455 & ~w13461 ) ;
  assign w13463 = w1367 & w13462 ;
  assign w13464 = w12993 | w12998 ;
  assign w13465 = w13145 & ~w13464 ;
  assign w13466 = w12996 ^ w13465 ;
  assign w13467 = ( ~w1367 & w13455 ) | ( ~w1367 & w13461 ) | ( w13455 & w13461 ) ;
  assign w13468 = ~w13455 & w13467 ;
  assign w13469 = w13466 | w13468 ;
  assign w13470 = ( w1225 & w13463 ) | ( w1225 & ~w13469 ) | ( w13463 & ~w13469 ) ;
  assign w13471 = w1225 & w13470 ;
  assign w13472 = w13001 | w13006 ;
  assign w13473 = w13145 & ~w13472 ;
  assign w13474 = w13004 ^ w13473 ;
  assign w13475 = ( ~w1225 & w13463 ) | ( ~w1225 & w13469 ) | ( w13463 & w13469 ) ;
  assign w13476 = ~w13463 & w13475 ;
  assign w13477 = w13474 | w13476 ;
  assign w13478 = ( w1091 & w13471 ) | ( w1091 & ~w13477 ) | ( w13471 & ~w13477 ) ;
  assign w13479 = w1091 & w13478 ;
  assign w13480 = w13009 | w13014 ;
  assign w13481 = w13145 & ~w13480 ;
  assign w13482 = w13012 ^ w13481 ;
  assign w13483 = ( ~w1091 & w13471 ) | ( ~w1091 & w13477 ) | ( w13471 & w13477 ) ;
  assign w13484 = ~w13471 & w13483 ;
  assign w13485 = w13482 | w13484 ;
  assign w13486 = ( w965 & w13479 ) | ( w965 & ~w13485 ) | ( w13479 & ~w13485 ) ;
  assign w13487 = w965 & w13486 ;
  assign w13488 = w13017 | w13022 ;
  assign w13489 = w13145 & ~w13488 ;
  assign w13490 = w13020 ^ w13489 ;
  assign w13491 = ( ~w965 & w13479 ) | ( ~w965 & w13485 ) | ( w13479 & w13485 ) ;
  assign w13492 = ~w13479 & w13491 ;
  assign w13493 = w13490 | w13492 ;
  assign w13494 = ( w847 & w13487 ) | ( w847 & ~w13493 ) | ( w13487 & ~w13493 ) ;
  assign w13495 = w847 & w13494 ;
  assign w13496 = w13025 | w13030 ;
  assign w13497 = w13145 & ~w13496 ;
  assign w13498 = w13028 ^ w13497 ;
  assign w13499 = ( ~w847 & w13487 ) | ( ~w847 & w13493 ) | ( w13487 & w13493 ) ;
  assign w13500 = ~w13487 & w13499 ;
  assign w13501 = w13498 | w13500 ;
  assign w13502 = ( w737 & w13495 ) | ( w737 & ~w13501 ) | ( w13495 & ~w13501 ) ;
  assign w13503 = w737 & w13502 ;
  assign w13504 = w13033 | w13038 ;
  assign w13505 = w13145 & ~w13504 ;
  assign w13506 = w13036 ^ w13505 ;
  assign w13507 = ( ~w737 & w13495 ) | ( ~w737 & w13501 ) | ( w13495 & w13501 ) ;
  assign w13508 = ~w13495 & w13507 ;
  assign w13509 = w13506 | w13508 ;
  assign w13510 = ( w635 & w13503 ) | ( w635 & ~w13509 ) | ( w13503 & ~w13509 ) ;
  assign w13511 = w635 & w13510 ;
  assign w13512 = w13041 | w13046 ;
  assign w13513 = w13145 & ~w13512 ;
  assign w13514 = w13044 ^ w13513 ;
  assign w13515 = ( ~w635 & w13503 ) | ( ~w635 & w13509 ) | ( w13503 & w13509 ) ;
  assign w13516 = ~w13503 & w13515 ;
  assign w13517 = w13514 | w13516 ;
  assign w13518 = ( w541 & w13511 ) | ( w541 & ~w13517 ) | ( w13511 & ~w13517 ) ;
  assign w13519 = w541 & w13518 ;
  assign w13520 = w13049 | w13054 ;
  assign w13521 = w13145 & ~w13520 ;
  assign w13522 = w13052 ^ w13521 ;
  assign w13523 = ( ~w541 & w13511 ) | ( ~w541 & w13517 ) | ( w13511 & w13517 ) ;
  assign w13524 = ~w13511 & w13523 ;
  assign w13525 = w13522 | w13524 ;
  assign w13526 = ( w455 & w13519 ) | ( w455 & ~w13525 ) | ( w13519 & ~w13525 ) ;
  assign w13527 = w455 & w13526 ;
  assign w13528 = ( ~w455 & w13519 ) | ( ~w455 & w13525 ) | ( w13519 & w13525 ) ;
  assign w13529 = ~w13519 & w13528 ;
  assign w13530 = w13057 | w13059 ;
  assign w13531 = w13145 & ~w13530 ;
  assign w13532 = w13062 ^ w13531 ;
  assign w13533 = w13529 | w13532 ;
  assign w13534 = ( w377 & w13527 ) | ( w377 & ~w13533 ) | ( w13527 & ~w13533 ) ;
  assign w13535 = w377 & w13534 ;
  assign w13536 = w13065 | w13070 ;
  assign w13537 = w13145 & ~w13536 ;
  assign w13538 = w13068 ^ w13537 ;
  assign w13539 = ( ~w377 & w13527 ) | ( ~w377 & w13533 ) | ( w13527 & w13533 ) ;
  assign w13540 = ~w13527 & w13539 ;
  assign w13541 = w13538 | w13540 ;
  assign w13542 = ( w307 & w13535 ) | ( w307 & ~w13541 ) | ( w13535 & ~w13541 ) ;
  assign w13543 = w307 & w13542 ;
  assign w13544 = w13073 | w13078 ;
  assign w13545 = w13145 & ~w13544 ;
  assign w13546 = w13076 ^ w13545 ;
  assign w13547 = ( ~w307 & w13535 ) | ( ~w307 & w13541 ) | ( w13535 & w13541 ) ;
  assign w13548 = ~w13535 & w13547 ;
  assign w13549 = w13546 | w13548 ;
  assign w13550 = ( w246 & w13543 ) | ( w246 & ~w13549 ) | ( w13543 & ~w13549 ) ;
  assign w13551 = w246 & w13550 ;
  assign w13552 = w13081 | w13086 ;
  assign w13553 = w13145 & ~w13552 ;
  assign w13554 = w13084 ^ w13553 ;
  assign w13555 = ( ~w246 & w13543 ) | ( ~w246 & w13549 ) | ( w13543 & w13549 ) ;
  assign w13556 = ~w13543 & w13555 ;
  assign w13557 = w13554 | w13556 ;
  assign w13558 = ( w185 & w13551 ) | ( w185 & ~w13557 ) | ( w13551 & ~w13557 ) ;
  assign w13559 = w185 & w13558 ;
  assign w13560 = w13089 | w13094 ;
  assign w13561 = w13145 & ~w13560 ;
  assign w13562 = w13092 ^ w13561 ;
  assign w13563 = ( ~w185 & w13551 ) | ( ~w185 & w13557 ) | ( w13551 & w13557 ) ;
  assign w13564 = ~w13551 & w13563 ;
  assign w13565 = w13562 | w13564 ;
  assign w13566 = ( w145 & w13559 ) | ( w145 & ~w13565 ) | ( w13559 & ~w13565 ) ;
  assign w13567 = w145 & w13566 ;
  assign w13568 = w13097 | w13102 ;
  assign w13569 = w13145 & ~w13568 ;
  assign w13570 = w13100 ^ w13569 ;
  assign w13571 = ( ~w145 & w13559 ) | ( ~w145 & w13565 ) | ( w13559 & w13565 ) ;
  assign w13572 = ~w13559 & w13571 ;
  assign w13573 = w13570 | w13572 ;
  assign w13574 = ( w132 & w13567 ) | ( w132 & ~w13573 ) | ( w13567 & ~w13573 ) ;
  assign w13575 = w132 & w13574 ;
  assign w13576 = w13105 | w13110 ;
  assign w13577 = w13145 & ~w13576 ;
  assign w13578 = w13108 ^ w13577 ;
  assign w13579 = ( ~w132 & w13567 ) | ( ~w132 & w13573 ) | ( w13567 & w13573 ) ;
  assign w13580 = ~w13567 & w13579 ;
  assign w13581 = w13578 | w13580 ;
  assign w13582 = ~w13575 & w13581 ;
  assign w13583 = w13113 | w13118 ;
  assign w13584 = w13145 & ~w13583 ;
  assign w13585 = w13116 ^ w13584 ;
  assign w13586 = ( ~w13131 & w13582 ) | ( ~w13131 & w13585 ) | ( w13582 & w13585 ) ;
  assign w13587 = w13120 & ~w13586 ;
  assign w13588 = ~w13123 & w13145 ;
  assign w13589 = ( w13586 & ~w13587 ) | ( w13586 & w13588 ) | ( ~w13587 & w13588 ) ;
  assign w13590 = w13131 | w13589 ;
  assign w13591 = ~w129 & w13590 ;
  assign w13592 = ( w13575 & w13581 ) | ( w13575 & w13585 ) | ( w13581 & w13585 ) ;
  assign w13593 = ~w13575 & w13592 ;
  assign w13594 = ( w129 & w13120 ) | ( w129 & w13123 ) | ( w13120 & w13123 ) ;
  assign w13595 = ( w13123 & ~w13145 ) | ( w13123 & w13594 ) | ( ~w13145 & w13594 ) ;
  assign w13596 = w13120 & w13595 ;
  assign w13597 = w13594 ^ w13596 ;
  assign w13598 = ( w12659 & w12664 ) | ( w12659 & w12691 ) | ( w12664 & w12691 ) ;
  assign w13599 = w12691 & ~w13598 ;
  assign w13600 = w12662 ^ w13599 ;
  assign w13601 = ( ~w13135 & w13142 ) | ( ~w13135 & w13600 ) | ( w13142 & w13600 ) ;
  assign w13602 = ~w13142 & w13601 ;
  assign w13603 = ( ~w13129 & w13131 ) | ( ~w13129 & w13602 ) | ( w13131 & w13602 ) ;
  assign w13604 = ~w13131 & w13603 ;
  assign w13605 = w13593 | w13604 ;
  assign w13606 = ( w13591 & ~w13593 ) | ( w13591 & w13597 ) | ( ~w13593 & w13597 ) ;
  assign w13607 = w13605 | w13606 ;
  assign w13608 = ( ~\pi015 & \pi016 ) | ( ~\pi015 & w13145 ) | ( \pi016 & w13145 ) ;
  assign w13609 = ( ~\pi014 & \pi016 ) | ( ~\pi014 & w13608 ) | ( \pi016 & w13608 ) ;
  assign w13610 = ( ~\pi016 & w13145 ) | ( ~\pi016 & w13607 ) | ( w13145 & w13607 ) ;
  assign w13611 = w13609 & w13610 ;
  assign w13612 = ( w13131 & w13135 ) | ( w13131 & ~w13142 ) | ( w13135 & ~w13142 ) ;
  assign w13613 = \pi015 & ~w13612 ;
  assign w13614 = \pi014 | \pi016 ;
  assign w13615 = ( ~w13612 & w13613 ) | ( ~w13612 & w13614 ) | ( w13613 & w13614 ) ;
  assign w13616 = ~w13142 & w13615 ;
  assign w13617 = ~w13129 & w13616 ;
  assign w13618 = ( \pi016 & w13607 ) | ( \pi016 & ~w13616 ) | ( w13607 & ~w13616 ) ;
  assign w13619 = w13617 & ~w13618 ;
  assign w13620 = ~\pi016 & w13607 ;
  assign w13621 = \pi017 ^ w13620 ;
  assign w13622 = w13619 | w13621 ;
  assign w13623 = ( w12691 & w13611 ) | ( w12691 & ~w13622 ) | ( w13611 & ~w13622 ) ;
  assign w13624 = w12691 & w13623 ;
  assign w13625 = ( ~w12691 & w13611 ) | ( ~w12691 & w13622 ) | ( w13611 & w13622 ) ;
  assign w13626 = ~w13611 & w13625 ;
  assign w13627 = w13145 & ~w13604 ;
  assign w13628 = ~w13593 & w13627 ;
  assign w13629 = ~w13606 & w13628 ;
  assign w13630 = \pi017 & w13607 ;
  assign w13631 = ( \pi016 & w13607 ) | ( \pi016 & ~w13630 ) | ( w13607 & ~w13630 ) ;
  assign w13632 = ( ~\pi016 & w13629 ) | ( ~\pi016 & w13631 ) | ( w13629 & w13631 ) ;
  assign w13633 = \pi018 ^ w13632 ;
  assign w13634 = w13626 | w13633 ;
  assign w13635 = ( w12245 & w13624 ) | ( w12245 & ~w13634 ) | ( w13624 & ~w13634 ) ;
  assign w13636 = w12245 & w13635 ;
  assign w13637 = ( w13149 & ~w13157 ) | ( w13149 & w13607 ) | ( ~w13157 & w13607 ) ;
  assign w13638 = ~w13149 & w13637 ;
  assign w13639 = \pi019 ^ w13638 ;
  assign w13640 = w13158 ^ w13639 ;
  assign w13641 = ( ~w12245 & w13624 ) | ( ~w12245 & w13634 ) | ( w13624 & w13634 ) ;
  assign w13642 = ~w13624 & w13641 ;
  assign w13643 = w13640 | w13642 ;
  assign w13644 = ( w11807 & w13636 ) | ( w11807 & ~w13643 ) | ( w13636 & ~w13643 ) ;
  assign w13645 = w11807 & w13644 ;
  assign w13646 = w13162 | w13164 ;
  assign w13647 = w13607 & ~w13646 ;
  assign w13648 = w13171 ^ w13647 ;
  assign w13649 = ( ~w11807 & w13636 ) | ( ~w11807 & w13643 ) | ( w13636 & w13643 ) ;
  assign w13650 = ~w13636 & w13649 ;
  assign w13651 = w13648 | w13650 ;
  assign w13652 = ( w11377 & w13645 ) | ( w11377 & ~w13651 ) | ( w13645 & ~w13651 ) ;
  assign w13653 = w11377 & w13652 ;
  assign w13654 = w13174 | w13180 ;
  assign w13655 = w13607 & ~w13654 ;
  assign w13656 = w13178 ^ w13655 ;
  assign w13657 = ( ~w11377 & w13645 ) | ( ~w11377 & w13651 ) | ( w13645 & w13651 ) ;
  assign w13658 = ~w13645 & w13657 ;
  assign w13659 = w13656 | w13658 ;
  assign w13660 = ( w10955 & w13653 ) | ( w10955 & ~w13659 ) | ( w13653 & ~w13659 ) ;
  assign w13661 = w10955 & w13660 ;
  assign w13662 = w13183 | w13188 ;
  assign w13663 = w13607 & ~w13662 ;
  assign w13664 = w13186 ^ w13663 ;
  assign w13665 = ( ~w10955 & w13653 ) | ( ~w10955 & w13659 ) | ( w13653 & w13659 ) ;
  assign w13666 = ~w13653 & w13665 ;
  assign w13667 = w13664 | w13666 ;
  assign w13668 = ( w10541 & w13661 ) | ( w10541 & ~w13667 ) | ( w13661 & ~w13667 ) ;
  assign w13669 = w10541 & w13668 ;
  assign w13670 = w13191 | w13196 ;
  assign w13671 = w13607 & ~w13670 ;
  assign w13672 = w13194 ^ w13671 ;
  assign w13673 = ( ~w10541 & w13661 ) | ( ~w10541 & w13667 ) | ( w13661 & w13667 ) ;
  assign w13674 = ~w13661 & w13673 ;
  assign w13675 = w13672 | w13674 ;
  assign w13676 = ( w10135 & w13669 ) | ( w10135 & ~w13675 ) | ( w13669 & ~w13675 ) ;
  assign w13677 = w10135 & w13676 ;
  assign w13678 = w13199 | w13204 ;
  assign w13679 = w13607 & ~w13678 ;
  assign w13680 = w13202 ^ w13679 ;
  assign w13681 = ( ~w10135 & w13669 ) | ( ~w10135 & w13675 ) | ( w13669 & w13675 ) ;
  assign w13682 = ~w13669 & w13681 ;
  assign w13683 = w13680 | w13682 ;
  assign w13684 = ( w9737 & w13677 ) | ( w9737 & ~w13683 ) | ( w13677 & ~w13683 ) ;
  assign w13685 = w9737 & w13684 ;
  assign w13686 = w13207 | w13212 ;
  assign w13687 = w13607 & ~w13686 ;
  assign w13688 = w13210 ^ w13687 ;
  assign w13689 = ( ~w9737 & w13677 ) | ( ~w9737 & w13683 ) | ( w13677 & w13683 ) ;
  assign w13690 = ~w13677 & w13689 ;
  assign w13691 = w13688 | w13690 ;
  assign w13692 = ( w9347 & w13685 ) | ( w9347 & ~w13691 ) | ( w13685 & ~w13691 ) ;
  assign w13693 = w9347 & w13692 ;
  assign w13694 = w13215 | w13220 ;
  assign w13695 = w13607 & ~w13694 ;
  assign w13696 = w13218 ^ w13695 ;
  assign w13697 = ( ~w9347 & w13685 ) | ( ~w9347 & w13691 ) | ( w13685 & w13691 ) ;
  assign w13698 = ~w13685 & w13697 ;
  assign w13699 = w13696 | w13698 ;
  assign w13700 = ( w8965 & w13693 ) | ( w8965 & ~w13699 ) | ( w13693 & ~w13699 ) ;
  assign w13701 = w8965 & w13700 ;
  assign w13702 = w13223 | w13228 ;
  assign w13703 = w13607 & ~w13702 ;
  assign w13704 = w13226 ^ w13703 ;
  assign w13705 = ( ~w8965 & w13693 ) | ( ~w8965 & w13699 ) | ( w13693 & w13699 ) ;
  assign w13706 = ~w13693 & w13705 ;
  assign w13707 = w13704 | w13706 ;
  assign w13708 = ( w8591 & w13701 ) | ( w8591 & ~w13707 ) | ( w13701 & ~w13707 ) ;
  assign w13709 = w8591 & w13708 ;
  assign w13710 = w13231 | w13236 ;
  assign w13711 = w13607 & ~w13710 ;
  assign w13712 = w13234 ^ w13711 ;
  assign w13713 = ( ~w8591 & w13701 ) | ( ~w8591 & w13707 ) | ( w13701 & w13707 ) ;
  assign w13714 = ~w13701 & w13713 ;
  assign w13715 = w13712 | w13714 ;
  assign w13716 = ( w8225 & w13709 ) | ( w8225 & ~w13715 ) | ( w13709 & ~w13715 ) ;
  assign w13717 = w8225 & w13716 ;
  assign w13718 = w13239 | w13244 ;
  assign w13719 = w13607 & ~w13718 ;
  assign w13720 = w13242 ^ w13719 ;
  assign w13721 = ( ~w8225 & w13709 ) | ( ~w8225 & w13715 ) | ( w13709 & w13715 ) ;
  assign w13722 = ~w13709 & w13721 ;
  assign w13723 = w13720 | w13722 ;
  assign w13724 = ( w7867 & w13717 ) | ( w7867 & ~w13723 ) | ( w13717 & ~w13723 ) ;
  assign w13725 = w7867 & w13724 ;
  assign w13726 = w13247 | w13252 ;
  assign w13727 = w13607 & ~w13726 ;
  assign w13728 = w13250 ^ w13727 ;
  assign w13729 = ( ~w7867 & w13717 ) | ( ~w7867 & w13723 ) | ( w13717 & w13723 ) ;
  assign w13730 = ~w13717 & w13729 ;
  assign w13731 = w13728 | w13730 ;
  assign w13732 = ( w7517 & w13725 ) | ( w7517 & ~w13731 ) | ( w13725 & ~w13731 ) ;
  assign w13733 = w7517 & w13732 ;
  assign w13734 = w13255 | w13260 ;
  assign w13735 = w13607 & ~w13734 ;
  assign w13736 = w13258 ^ w13735 ;
  assign w13737 = ( ~w7517 & w13725 ) | ( ~w7517 & w13731 ) | ( w13725 & w13731 ) ;
  assign w13738 = ~w13725 & w13737 ;
  assign w13739 = w13736 | w13738 ;
  assign w13740 = ( w7175 & w13733 ) | ( w7175 & ~w13739 ) | ( w13733 & ~w13739 ) ;
  assign w13741 = w7175 & w13740 ;
  assign w13742 = w13263 | w13268 ;
  assign w13743 = w13607 & ~w13742 ;
  assign w13744 = w13266 ^ w13743 ;
  assign w13745 = ( ~w7175 & w13733 ) | ( ~w7175 & w13739 ) | ( w13733 & w13739 ) ;
  assign w13746 = ~w13733 & w13745 ;
  assign w13747 = w13744 | w13746 ;
  assign w13748 = ( w6841 & w13741 ) | ( w6841 & ~w13747 ) | ( w13741 & ~w13747 ) ;
  assign w13749 = w6841 & w13748 ;
  assign w13750 = w13271 | w13276 ;
  assign w13751 = w13607 & ~w13750 ;
  assign w13752 = w13274 ^ w13751 ;
  assign w13753 = ( ~w6841 & w13741 ) | ( ~w6841 & w13747 ) | ( w13741 & w13747 ) ;
  assign w13754 = ~w13741 & w13753 ;
  assign w13755 = w13752 | w13754 ;
  assign w13756 = ( w6515 & w13749 ) | ( w6515 & ~w13755 ) | ( w13749 & ~w13755 ) ;
  assign w13757 = w6515 & w13756 ;
  assign w13758 = w13279 | w13284 ;
  assign w13759 = w13607 & ~w13758 ;
  assign w13760 = w13282 ^ w13759 ;
  assign w13761 = ( ~w6515 & w13749 ) | ( ~w6515 & w13755 ) | ( w13749 & w13755 ) ;
  assign w13762 = ~w13749 & w13761 ;
  assign w13763 = w13760 | w13762 ;
  assign w13764 = ( w6197 & w13757 ) | ( w6197 & ~w13763 ) | ( w13757 & ~w13763 ) ;
  assign w13765 = w6197 & w13764 ;
  assign w13766 = w13287 | w13292 ;
  assign w13767 = w13607 & ~w13766 ;
  assign w13768 = w13290 ^ w13767 ;
  assign w13769 = ( ~w6197 & w13757 ) | ( ~w6197 & w13763 ) | ( w13757 & w13763 ) ;
  assign w13770 = ~w13757 & w13769 ;
  assign w13771 = w13768 | w13770 ;
  assign w13772 = ( w5887 & w13765 ) | ( w5887 & ~w13771 ) | ( w13765 & ~w13771 ) ;
  assign w13773 = w5887 & w13772 ;
  assign w13774 = w13295 | w13300 ;
  assign w13775 = w13607 & ~w13774 ;
  assign w13776 = w13298 ^ w13775 ;
  assign w13777 = ( ~w5887 & w13765 ) | ( ~w5887 & w13771 ) | ( w13765 & w13771 ) ;
  assign w13778 = ~w13765 & w13777 ;
  assign w13779 = w13776 | w13778 ;
  assign w13780 = ( w5585 & w13773 ) | ( w5585 & ~w13779 ) | ( w13773 & ~w13779 ) ;
  assign w13781 = w5585 & w13780 ;
  assign w13782 = w13303 | w13308 ;
  assign w13783 = w13607 & ~w13782 ;
  assign w13784 = w13306 ^ w13783 ;
  assign w13785 = ( ~w5585 & w13773 ) | ( ~w5585 & w13779 ) | ( w13773 & w13779 ) ;
  assign w13786 = ~w13773 & w13785 ;
  assign w13787 = w13784 | w13786 ;
  assign w13788 = ( w5291 & w13781 ) | ( w5291 & ~w13787 ) | ( w13781 & ~w13787 ) ;
  assign w13789 = w5291 & w13788 ;
  assign w13790 = w13311 | w13316 ;
  assign w13791 = w13607 & ~w13790 ;
  assign w13792 = w13314 ^ w13791 ;
  assign w13793 = ( ~w5291 & w13781 ) | ( ~w5291 & w13787 ) | ( w13781 & w13787 ) ;
  assign w13794 = ~w13781 & w13793 ;
  assign w13795 = w13792 | w13794 ;
  assign w13796 = ( w5005 & w13789 ) | ( w5005 & ~w13795 ) | ( w13789 & ~w13795 ) ;
  assign w13797 = w5005 & w13796 ;
  assign w13798 = w13319 | w13324 ;
  assign w13799 = w13607 & ~w13798 ;
  assign w13800 = w13322 ^ w13799 ;
  assign w13801 = ( ~w5005 & w13789 ) | ( ~w5005 & w13795 ) | ( w13789 & w13795 ) ;
  assign w13802 = ~w13789 & w13801 ;
  assign w13803 = w13800 | w13802 ;
  assign w13804 = ( w4727 & w13797 ) | ( w4727 & ~w13803 ) | ( w13797 & ~w13803 ) ;
  assign w13805 = w4727 & w13804 ;
  assign w13806 = w13327 | w13332 ;
  assign w13807 = w13607 & ~w13806 ;
  assign w13808 = w13330 ^ w13807 ;
  assign w13809 = ( ~w4727 & w13797 ) | ( ~w4727 & w13803 ) | ( w13797 & w13803 ) ;
  assign w13810 = ~w13797 & w13809 ;
  assign w13811 = w13808 | w13810 ;
  assign w13812 = ( w4457 & w13805 ) | ( w4457 & ~w13811 ) | ( w13805 & ~w13811 ) ;
  assign w13813 = w4457 & w13812 ;
  assign w13814 = w13335 | w13340 ;
  assign w13815 = w13607 & ~w13814 ;
  assign w13816 = w13338 ^ w13815 ;
  assign w13817 = ( ~w4457 & w13805 ) | ( ~w4457 & w13811 ) | ( w13805 & w13811 ) ;
  assign w13818 = ~w13805 & w13817 ;
  assign w13819 = w13816 | w13818 ;
  assign w13820 = ( w4195 & w13813 ) | ( w4195 & ~w13819 ) | ( w13813 & ~w13819 ) ;
  assign w13821 = w4195 & w13820 ;
  assign w13822 = w13343 | w13348 ;
  assign w13823 = w13607 & ~w13822 ;
  assign w13824 = w13346 ^ w13823 ;
  assign w13825 = ( ~w4195 & w13813 ) | ( ~w4195 & w13819 ) | ( w13813 & w13819 ) ;
  assign w13826 = ~w13813 & w13825 ;
  assign w13827 = w13824 | w13826 ;
  assign w13828 = ( w3941 & w13821 ) | ( w3941 & ~w13827 ) | ( w13821 & ~w13827 ) ;
  assign w13829 = w3941 & w13828 ;
  assign w13830 = w13351 | w13356 ;
  assign w13831 = w13607 & ~w13830 ;
  assign w13832 = w13354 ^ w13831 ;
  assign w13833 = ( ~w3941 & w13821 ) | ( ~w3941 & w13827 ) | ( w13821 & w13827 ) ;
  assign w13834 = ~w13821 & w13833 ;
  assign w13835 = w13832 | w13834 ;
  assign w13836 = ( w3695 & w13829 ) | ( w3695 & ~w13835 ) | ( w13829 & ~w13835 ) ;
  assign w13837 = w3695 & w13836 ;
  assign w13838 = w13359 | w13364 ;
  assign w13839 = w13607 & ~w13838 ;
  assign w13840 = w13362 ^ w13839 ;
  assign w13841 = ( ~w3695 & w13829 ) | ( ~w3695 & w13835 ) | ( w13829 & w13835 ) ;
  assign w13842 = ~w13829 & w13841 ;
  assign w13843 = w13840 | w13842 ;
  assign w13844 = ( w3457 & w13837 ) | ( w3457 & ~w13843 ) | ( w13837 & ~w13843 ) ;
  assign w13845 = w3457 & w13844 ;
  assign w13846 = w13367 | w13372 ;
  assign w13847 = w13607 & ~w13846 ;
  assign w13848 = w13370 ^ w13847 ;
  assign w13849 = ( ~w3457 & w13837 ) | ( ~w3457 & w13843 ) | ( w13837 & w13843 ) ;
  assign w13850 = ~w13837 & w13849 ;
  assign w13851 = w13848 | w13850 ;
  assign w13852 = ( w3227 & w13845 ) | ( w3227 & ~w13851 ) | ( w13845 & ~w13851 ) ;
  assign w13853 = w3227 & w13852 ;
  assign w13854 = w13375 | w13380 ;
  assign w13855 = w13607 & ~w13854 ;
  assign w13856 = w13378 ^ w13855 ;
  assign w13857 = ( ~w3227 & w13845 ) | ( ~w3227 & w13851 ) | ( w13845 & w13851 ) ;
  assign w13858 = ~w13845 & w13857 ;
  assign w13859 = w13856 | w13858 ;
  assign w13860 = ( w3005 & w13853 ) | ( w3005 & ~w13859 ) | ( w13853 & ~w13859 ) ;
  assign w13861 = w3005 & w13860 ;
  assign w13862 = w13383 | w13388 ;
  assign w13863 = w13607 & ~w13862 ;
  assign w13864 = w13386 ^ w13863 ;
  assign w13865 = ( ~w3005 & w13853 ) | ( ~w3005 & w13859 ) | ( w13853 & w13859 ) ;
  assign w13866 = ~w13853 & w13865 ;
  assign w13867 = w13864 | w13866 ;
  assign w13868 = ( w2791 & w13861 ) | ( w2791 & ~w13867 ) | ( w13861 & ~w13867 ) ;
  assign w13869 = w2791 & w13868 ;
  assign w13870 = w13391 | w13396 ;
  assign w13871 = w13607 & ~w13870 ;
  assign w13872 = w13394 ^ w13871 ;
  assign w13873 = ( ~w2791 & w13861 ) | ( ~w2791 & w13867 ) | ( w13861 & w13867 ) ;
  assign w13874 = ~w13861 & w13873 ;
  assign w13875 = w13872 | w13874 ;
  assign w13876 = ( w2585 & w13869 ) | ( w2585 & ~w13875 ) | ( w13869 & ~w13875 ) ;
  assign w13877 = w2585 & w13876 ;
  assign w13878 = w13399 | w13404 ;
  assign w13879 = w13607 & ~w13878 ;
  assign w13880 = w13402 ^ w13879 ;
  assign w13881 = ( ~w2585 & w13869 ) | ( ~w2585 & w13875 ) | ( w13869 & w13875 ) ;
  assign w13882 = ~w13869 & w13881 ;
  assign w13883 = w13880 | w13882 ;
  assign w13884 = ( w2387 & w13877 ) | ( w2387 & ~w13883 ) | ( w13877 & ~w13883 ) ;
  assign w13885 = w2387 & w13884 ;
  assign w13886 = w13407 | w13412 ;
  assign w13887 = w13607 & ~w13886 ;
  assign w13888 = w13410 ^ w13887 ;
  assign w13889 = ( ~w2387 & w13877 ) | ( ~w2387 & w13883 ) | ( w13877 & w13883 ) ;
  assign w13890 = ~w13877 & w13889 ;
  assign w13891 = w13888 | w13890 ;
  assign w13892 = ( w2197 & w13885 ) | ( w2197 & ~w13891 ) | ( w13885 & ~w13891 ) ;
  assign w13893 = w2197 & w13892 ;
  assign w13894 = w13415 | w13420 ;
  assign w13895 = w13607 & ~w13894 ;
  assign w13896 = w13418 ^ w13895 ;
  assign w13897 = ( ~w2197 & w13885 ) | ( ~w2197 & w13891 ) | ( w13885 & w13891 ) ;
  assign w13898 = ~w13885 & w13897 ;
  assign w13899 = w13896 | w13898 ;
  assign w13900 = ( w2015 & w13893 ) | ( w2015 & ~w13899 ) | ( w13893 & ~w13899 ) ;
  assign w13901 = w2015 & w13900 ;
  assign w13902 = w13423 | w13428 ;
  assign w13903 = w13607 & ~w13902 ;
  assign w13904 = w13426 ^ w13903 ;
  assign w13905 = ( ~w2015 & w13893 ) | ( ~w2015 & w13899 ) | ( w13893 & w13899 ) ;
  assign w13906 = ~w13893 & w13905 ;
  assign w13907 = w13904 | w13906 ;
  assign w13908 = ( w1841 & w13901 ) | ( w1841 & ~w13907 ) | ( w13901 & ~w13907 ) ;
  assign w13909 = w1841 & w13908 ;
  assign w13910 = w13431 | w13436 ;
  assign w13911 = w13607 & ~w13910 ;
  assign w13912 = w13434 ^ w13911 ;
  assign w13913 = ( ~w1841 & w13901 ) | ( ~w1841 & w13907 ) | ( w13901 & w13907 ) ;
  assign w13914 = ~w13901 & w13913 ;
  assign w13915 = w13912 | w13914 ;
  assign w13916 = ( w1675 & w13909 ) | ( w1675 & ~w13915 ) | ( w13909 & ~w13915 ) ;
  assign w13917 = w1675 & w13916 ;
  assign w13918 = w13439 | w13444 ;
  assign w13919 = w13607 & ~w13918 ;
  assign w13920 = w13442 ^ w13919 ;
  assign w13921 = ( ~w1675 & w13909 ) | ( ~w1675 & w13915 ) | ( w13909 & w13915 ) ;
  assign w13922 = ~w13909 & w13921 ;
  assign w13923 = w13920 | w13922 ;
  assign w13924 = ( w1517 & w13917 ) | ( w1517 & ~w13923 ) | ( w13917 & ~w13923 ) ;
  assign w13925 = w1517 & w13924 ;
  assign w13926 = w13447 | w13452 ;
  assign w13927 = w13607 & ~w13926 ;
  assign w13928 = w13450 ^ w13927 ;
  assign w13929 = ( ~w1517 & w13917 ) | ( ~w1517 & w13923 ) | ( w13917 & w13923 ) ;
  assign w13930 = ~w13917 & w13929 ;
  assign w13931 = w13928 | w13930 ;
  assign w13932 = ( w1367 & w13925 ) | ( w1367 & ~w13931 ) | ( w13925 & ~w13931 ) ;
  assign w13933 = w1367 & w13932 ;
  assign w13934 = w13455 | w13460 ;
  assign w13935 = w13607 & ~w13934 ;
  assign w13936 = w13458 ^ w13935 ;
  assign w13937 = ( ~w1367 & w13925 ) | ( ~w1367 & w13931 ) | ( w13925 & w13931 ) ;
  assign w13938 = ~w13925 & w13937 ;
  assign w13939 = w13936 | w13938 ;
  assign w13940 = ( w1225 & w13933 ) | ( w1225 & ~w13939 ) | ( w13933 & ~w13939 ) ;
  assign w13941 = w1225 & w13940 ;
  assign w13942 = w13463 | w13468 ;
  assign w13943 = w13607 & ~w13942 ;
  assign w13944 = w13466 ^ w13943 ;
  assign w13945 = ( ~w1225 & w13933 ) | ( ~w1225 & w13939 ) | ( w13933 & w13939 ) ;
  assign w13946 = ~w13933 & w13945 ;
  assign w13947 = w13944 | w13946 ;
  assign w13948 = ( w1091 & w13941 ) | ( w1091 & ~w13947 ) | ( w13941 & ~w13947 ) ;
  assign w13949 = w1091 & w13948 ;
  assign w13950 = w13471 | w13476 ;
  assign w13951 = w13607 & ~w13950 ;
  assign w13952 = w13474 ^ w13951 ;
  assign w13953 = ( ~w1091 & w13941 ) | ( ~w1091 & w13947 ) | ( w13941 & w13947 ) ;
  assign w13954 = ~w13941 & w13953 ;
  assign w13955 = w13952 | w13954 ;
  assign w13956 = ( w965 & w13949 ) | ( w965 & ~w13955 ) | ( w13949 & ~w13955 ) ;
  assign w13957 = w965 & w13956 ;
  assign w13958 = w13479 | w13484 ;
  assign w13959 = w13607 & ~w13958 ;
  assign w13960 = w13482 ^ w13959 ;
  assign w13961 = ( ~w965 & w13949 ) | ( ~w965 & w13955 ) | ( w13949 & w13955 ) ;
  assign w13962 = ~w13949 & w13961 ;
  assign w13963 = w13960 | w13962 ;
  assign w13964 = ( w847 & w13957 ) | ( w847 & ~w13963 ) | ( w13957 & ~w13963 ) ;
  assign w13965 = w847 & w13964 ;
  assign w13966 = w13487 | w13492 ;
  assign w13967 = w13607 & ~w13966 ;
  assign w13968 = w13490 ^ w13967 ;
  assign w13969 = ( ~w847 & w13957 ) | ( ~w847 & w13963 ) | ( w13957 & w13963 ) ;
  assign w13970 = ~w13957 & w13969 ;
  assign w13971 = w13968 | w13970 ;
  assign w13972 = ( w737 & w13965 ) | ( w737 & ~w13971 ) | ( w13965 & ~w13971 ) ;
  assign w13973 = w737 & w13972 ;
  assign w13974 = w13495 | w13500 ;
  assign w13975 = w13607 & ~w13974 ;
  assign w13976 = w13498 ^ w13975 ;
  assign w13977 = ( ~w737 & w13965 ) | ( ~w737 & w13971 ) | ( w13965 & w13971 ) ;
  assign w13978 = ~w13965 & w13977 ;
  assign w13979 = w13976 | w13978 ;
  assign w13980 = ( w635 & w13973 ) | ( w635 & ~w13979 ) | ( w13973 & ~w13979 ) ;
  assign w13981 = w635 & w13980 ;
  assign w13982 = w13503 | w13508 ;
  assign w13983 = w13607 & ~w13982 ;
  assign w13984 = w13506 ^ w13983 ;
  assign w13985 = ( ~w635 & w13973 ) | ( ~w635 & w13979 ) | ( w13973 & w13979 ) ;
  assign w13986 = ~w13973 & w13985 ;
  assign w13987 = w13984 | w13986 ;
  assign w13988 = ( w541 & w13981 ) | ( w541 & ~w13987 ) | ( w13981 & ~w13987 ) ;
  assign w13989 = w541 & w13988 ;
  assign w13990 = w13511 | w13516 ;
  assign w13991 = w13607 & ~w13990 ;
  assign w13992 = w13514 ^ w13991 ;
  assign w13993 = ( ~w541 & w13981 ) | ( ~w541 & w13987 ) | ( w13981 & w13987 ) ;
  assign w13994 = ~w13981 & w13993 ;
  assign w13995 = w13992 | w13994 ;
  assign w13996 = ( w455 & w13989 ) | ( w455 & ~w13995 ) | ( w13989 & ~w13995 ) ;
  assign w13997 = w455 & w13996 ;
  assign w13998 = w13519 | w13524 ;
  assign w13999 = w13607 & ~w13998 ;
  assign w14000 = w13522 ^ w13999 ;
  assign w14001 = ( ~w455 & w13989 ) | ( ~w455 & w13995 ) | ( w13989 & w13995 ) ;
  assign w14002 = ~w13989 & w14001 ;
  assign w14003 = w14000 | w14002 ;
  assign w14004 = ( w377 & w13997 ) | ( w377 & ~w14003 ) | ( w13997 & ~w14003 ) ;
  assign w14005 = w377 & w14004 ;
  assign w14006 = ( ~w377 & w13997 ) | ( ~w377 & w14003 ) | ( w13997 & w14003 ) ;
  assign w14007 = ~w13997 & w14006 ;
  assign w14008 = w13527 | w13529 ;
  assign w14009 = w13607 & ~w14008 ;
  assign w14010 = w13532 ^ w14009 ;
  assign w14011 = w14007 | w14010 ;
  assign w14012 = ( w307 & w14005 ) | ( w307 & ~w14011 ) | ( w14005 & ~w14011 ) ;
  assign w14013 = w307 & w14012 ;
  assign w14014 = w13535 | w13540 ;
  assign w14015 = w13607 & ~w14014 ;
  assign w14016 = w13538 ^ w14015 ;
  assign w14017 = ( ~w307 & w14005 ) | ( ~w307 & w14011 ) | ( w14005 & w14011 ) ;
  assign w14018 = ~w14005 & w14017 ;
  assign w14019 = w14016 | w14018 ;
  assign w14020 = ( w246 & w14013 ) | ( w246 & ~w14019 ) | ( w14013 & ~w14019 ) ;
  assign w14021 = w246 & w14020 ;
  assign w14022 = w13543 | w13548 ;
  assign w14023 = w13607 & ~w14022 ;
  assign w14024 = w13546 ^ w14023 ;
  assign w14025 = ( ~w246 & w14013 ) | ( ~w246 & w14019 ) | ( w14013 & w14019 ) ;
  assign w14026 = ~w14013 & w14025 ;
  assign w14027 = w14024 | w14026 ;
  assign w14028 = ( w185 & w14021 ) | ( w185 & ~w14027 ) | ( w14021 & ~w14027 ) ;
  assign w14029 = w185 & w14028 ;
  assign w14030 = w13551 | w13556 ;
  assign w14031 = w13607 & ~w14030 ;
  assign w14032 = w13554 ^ w14031 ;
  assign w14033 = ( ~w185 & w14021 ) | ( ~w185 & w14027 ) | ( w14021 & w14027 ) ;
  assign w14034 = ~w14021 & w14033 ;
  assign w14035 = w14032 | w14034 ;
  assign w14036 = ( w145 & w14029 ) | ( w145 & ~w14035 ) | ( w14029 & ~w14035 ) ;
  assign w14037 = w145 & w14036 ;
  assign w14038 = w13559 | w13564 ;
  assign w14039 = w13607 & ~w14038 ;
  assign w14040 = w13562 ^ w14039 ;
  assign w14041 = ( ~w145 & w14029 ) | ( ~w145 & w14035 ) | ( w14029 & w14035 ) ;
  assign w14042 = ~w14029 & w14041 ;
  assign w14043 = w14040 | w14042 ;
  assign w14044 = ( w132 & w14037 ) | ( w132 & ~w14043 ) | ( w14037 & ~w14043 ) ;
  assign w14045 = w132 & w14044 ;
  assign w14046 = w13567 | w13572 ;
  assign w14047 = w13607 & ~w14046 ;
  assign w14048 = w13570 ^ w14047 ;
  assign w14049 = ( ~w132 & w14037 ) | ( ~w132 & w14043 ) | ( w14037 & w14043 ) ;
  assign w14050 = ~w14037 & w14049 ;
  assign w14051 = w14048 | w14050 ;
  assign w14052 = ~w14045 & w14051 ;
  assign w14053 = w13575 | w13580 ;
  assign w14054 = w13607 & ~w14053 ;
  assign w14055 = w13578 ^ w14054 ;
  assign w14056 = ( ~w13593 & w14052 ) | ( ~w13593 & w14055 ) | ( w14052 & w14055 ) ;
  assign w14057 = w13582 & ~w14056 ;
  assign w14058 = ~w13585 & w13607 ;
  assign w14059 = ( w14056 & ~w14057 ) | ( w14056 & w14058 ) | ( ~w14057 & w14058 ) ;
  assign w14060 = w13593 | w14059 ;
  assign w14061 = ~w129 & w14060 ;
  assign w14062 = ( w14045 & w14051 ) | ( w14045 & w14055 ) | ( w14051 & w14055 ) ;
  assign w14063 = ~w14045 & w14062 ;
  assign w14064 = ( w129 & w13582 ) | ( w129 & w13585 ) | ( w13582 & w13585 ) ;
  assign w14065 = ( w13585 & ~w13607 ) | ( w13585 & w14064 ) | ( ~w13607 & w14064 ) ;
  assign w14066 = w13582 & w14065 ;
  assign w14067 = w14064 ^ w14066 ;
  assign w14068 = ( w13113 & w13118 ) | ( w13113 & w13145 ) | ( w13118 & w13145 ) ;
  assign w14069 = w13145 & ~w14068 ;
  assign w14070 = w13116 ^ w14069 ;
  assign w14071 = ( ~w13597 & w13604 ) | ( ~w13597 & w14070 ) | ( w13604 & w14070 ) ;
  assign w14072 = ~w13604 & w14071 ;
  assign w14073 = ( ~w13591 & w13593 ) | ( ~w13591 & w14072 ) | ( w13593 & w14072 ) ;
  assign w14074 = ~w13593 & w14073 ;
  assign w14075 = w14063 | w14074 ;
  assign w14076 = ( w14061 & ~w14063 ) | ( w14061 & w14067 ) | ( ~w14063 & w14067 ) ;
  assign w14077 = w14075 | w14076 ;
  assign w14078 = ( ~\pi013 & \pi014 ) | ( ~\pi013 & w13607 ) | ( \pi014 & w13607 ) ;
  assign w14079 = ( ~\pi012 & \pi014 ) | ( ~\pi012 & w14078 ) | ( \pi014 & w14078 ) ;
  assign w14080 = ( ~\pi014 & w13607 ) | ( ~\pi014 & w14077 ) | ( w13607 & w14077 ) ;
  assign w14081 = w14079 & w14080 ;
  assign w14082 = ( w13593 & w13597 ) | ( w13593 & ~w13604 ) | ( w13597 & ~w13604 ) ;
  assign w14083 = \pi013 & ~w14082 ;
  assign w14084 = \pi012 | \pi014 ;
  assign w14085 = ( ~w14082 & w14083 ) | ( ~w14082 & w14084 ) | ( w14083 & w14084 ) ;
  assign w14086 = ~w13604 & w14085 ;
  assign w14087 = ~w13591 & w14086 ;
  assign w14088 = ( \pi014 & w14077 ) | ( \pi014 & ~w14086 ) | ( w14077 & ~w14086 ) ;
  assign w14089 = w14087 & ~w14088 ;
  assign w14090 = ~\pi014 & w14077 ;
  assign w14091 = \pi015 ^ w14090 ;
  assign w14092 = w14089 | w14091 ;
  assign w14093 = ( w13145 & w14081 ) | ( w13145 & ~w14092 ) | ( w14081 & ~w14092 ) ;
  assign w14094 = w13145 & w14093 ;
  assign w14095 = ( ~w13145 & w14081 ) | ( ~w13145 & w14092 ) | ( w14081 & w14092 ) ;
  assign w14096 = ~w14081 & w14095 ;
  assign w14097 = w13607 & ~w14074 ;
  assign w14098 = ~w14063 & w14097 ;
  assign w14099 = ~w14076 & w14098 ;
  assign w14100 = \pi015 & w14077 ;
  assign w14101 = ( \pi014 & w14077 ) | ( \pi014 & ~w14100 ) | ( w14077 & ~w14100 ) ;
  assign w14102 = ( ~\pi014 & w14099 ) | ( ~\pi014 & w14101 ) | ( w14099 & w14101 ) ;
  assign w14103 = \pi016 ^ w14102 ;
  assign w14104 = w14096 | w14103 ;
  assign w14105 = ( w12691 & w14094 ) | ( w12691 & ~w14104 ) | ( w14094 & ~w14104 ) ;
  assign w14106 = w12691 & w14105 ;
  assign w14107 = ( w13611 & ~w13619 ) | ( w13611 & w14077 ) | ( ~w13619 & w14077 ) ;
  assign w14108 = ~w13611 & w14107 ;
  assign w14109 = \pi017 ^ w14108 ;
  assign w14110 = w13620 ^ w14109 ;
  assign w14111 = ( ~w12691 & w14094 ) | ( ~w12691 & w14104 ) | ( w14094 & w14104 ) ;
  assign w14112 = ~w14094 & w14111 ;
  assign w14113 = w14110 | w14112 ;
  assign w14114 = ( w12245 & w14106 ) | ( w12245 & ~w14113 ) | ( w14106 & ~w14113 ) ;
  assign w14115 = w12245 & w14114 ;
  assign w14116 = w13624 | w13626 ;
  assign w14117 = w14077 & ~w14116 ;
  assign w14118 = w13633 ^ w14117 ;
  assign w14119 = ( ~w12245 & w14106 ) | ( ~w12245 & w14113 ) | ( w14106 & w14113 ) ;
  assign w14120 = ~w14106 & w14119 ;
  assign w14121 = w14118 | w14120 ;
  assign w14122 = ( w11807 & w14115 ) | ( w11807 & ~w14121 ) | ( w14115 & ~w14121 ) ;
  assign w14123 = w11807 & w14122 ;
  assign w14124 = w13636 | w13642 ;
  assign w14125 = w14077 & ~w14124 ;
  assign w14126 = w13640 ^ w14125 ;
  assign w14127 = ( ~w11807 & w14115 ) | ( ~w11807 & w14121 ) | ( w14115 & w14121 ) ;
  assign w14128 = ~w14115 & w14127 ;
  assign w14129 = w14126 | w14128 ;
  assign w14130 = ( w11377 & w14123 ) | ( w11377 & ~w14129 ) | ( w14123 & ~w14129 ) ;
  assign w14131 = w11377 & w14130 ;
  assign w14132 = w13645 | w13650 ;
  assign w14133 = w14077 & ~w14132 ;
  assign w14134 = w13648 ^ w14133 ;
  assign w14135 = ( ~w11377 & w14123 ) | ( ~w11377 & w14129 ) | ( w14123 & w14129 ) ;
  assign w14136 = ~w14123 & w14135 ;
  assign w14137 = w14134 | w14136 ;
  assign w14138 = ( w10955 & w14131 ) | ( w10955 & ~w14137 ) | ( w14131 & ~w14137 ) ;
  assign w14139 = w10955 & w14138 ;
  assign w14140 = w13653 | w13658 ;
  assign w14141 = w14077 & ~w14140 ;
  assign w14142 = w13656 ^ w14141 ;
  assign w14143 = ( ~w10955 & w14131 ) | ( ~w10955 & w14137 ) | ( w14131 & w14137 ) ;
  assign w14144 = ~w14131 & w14143 ;
  assign w14145 = w14142 | w14144 ;
  assign w14146 = ( w10541 & w14139 ) | ( w10541 & ~w14145 ) | ( w14139 & ~w14145 ) ;
  assign w14147 = w10541 & w14146 ;
  assign w14148 = w13661 | w13666 ;
  assign w14149 = w14077 & ~w14148 ;
  assign w14150 = w13664 ^ w14149 ;
  assign w14151 = ( ~w10541 & w14139 ) | ( ~w10541 & w14145 ) | ( w14139 & w14145 ) ;
  assign w14152 = ~w14139 & w14151 ;
  assign w14153 = w14150 | w14152 ;
  assign w14154 = ( w10135 & w14147 ) | ( w10135 & ~w14153 ) | ( w14147 & ~w14153 ) ;
  assign w14155 = w10135 & w14154 ;
  assign w14156 = w13669 | w13674 ;
  assign w14157 = w14077 & ~w14156 ;
  assign w14158 = w13672 ^ w14157 ;
  assign w14159 = ( ~w10135 & w14147 ) | ( ~w10135 & w14153 ) | ( w14147 & w14153 ) ;
  assign w14160 = ~w14147 & w14159 ;
  assign w14161 = w14158 | w14160 ;
  assign w14162 = ( w9737 & w14155 ) | ( w9737 & ~w14161 ) | ( w14155 & ~w14161 ) ;
  assign w14163 = w9737 & w14162 ;
  assign w14164 = w13677 | w13682 ;
  assign w14165 = w14077 & ~w14164 ;
  assign w14166 = w13680 ^ w14165 ;
  assign w14167 = ( ~w9737 & w14155 ) | ( ~w9737 & w14161 ) | ( w14155 & w14161 ) ;
  assign w14168 = ~w14155 & w14167 ;
  assign w14169 = w14166 | w14168 ;
  assign w14170 = ( w9347 & w14163 ) | ( w9347 & ~w14169 ) | ( w14163 & ~w14169 ) ;
  assign w14171 = w9347 & w14170 ;
  assign w14172 = w13685 | w13690 ;
  assign w14173 = w14077 & ~w14172 ;
  assign w14174 = w13688 ^ w14173 ;
  assign w14175 = ( ~w9347 & w14163 ) | ( ~w9347 & w14169 ) | ( w14163 & w14169 ) ;
  assign w14176 = ~w14163 & w14175 ;
  assign w14177 = w14174 | w14176 ;
  assign w14178 = ( w8965 & w14171 ) | ( w8965 & ~w14177 ) | ( w14171 & ~w14177 ) ;
  assign w14179 = w8965 & w14178 ;
  assign w14180 = w13693 | w13698 ;
  assign w14181 = w14077 & ~w14180 ;
  assign w14182 = w13696 ^ w14181 ;
  assign w14183 = ( ~w8965 & w14171 ) | ( ~w8965 & w14177 ) | ( w14171 & w14177 ) ;
  assign w14184 = ~w14171 & w14183 ;
  assign w14185 = w14182 | w14184 ;
  assign w14186 = ( w8591 & w14179 ) | ( w8591 & ~w14185 ) | ( w14179 & ~w14185 ) ;
  assign w14187 = w8591 & w14186 ;
  assign w14188 = w13701 | w13706 ;
  assign w14189 = w14077 & ~w14188 ;
  assign w14190 = w13704 ^ w14189 ;
  assign w14191 = ( ~w8591 & w14179 ) | ( ~w8591 & w14185 ) | ( w14179 & w14185 ) ;
  assign w14192 = ~w14179 & w14191 ;
  assign w14193 = w14190 | w14192 ;
  assign w14194 = ( w8225 & w14187 ) | ( w8225 & ~w14193 ) | ( w14187 & ~w14193 ) ;
  assign w14195 = w8225 & w14194 ;
  assign w14196 = w13709 | w13714 ;
  assign w14197 = w14077 & ~w14196 ;
  assign w14198 = w13712 ^ w14197 ;
  assign w14199 = ( ~w8225 & w14187 ) | ( ~w8225 & w14193 ) | ( w14187 & w14193 ) ;
  assign w14200 = ~w14187 & w14199 ;
  assign w14201 = w14198 | w14200 ;
  assign w14202 = ( w7867 & w14195 ) | ( w7867 & ~w14201 ) | ( w14195 & ~w14201 ) ;
  assign w14203 = w7867 & w14202 ;
  assign w14204 = w13717 | w13722 ;
  assign w14205 = w14077 & ~w14204 ;
  assign w14206 = w13720 ^ w14205 ;
  assign w14207 = ( ~w7867 & w14195 ) | ( ~w7867 & w14201 ) | ( w14195 & w14201 ) ;
  assign w14208 = ~w14195 & w14207 ;
  assign w14209 = w14206 | w14208 ;
  assign w14210 = ( w7517 & w14203 ) | ( w7517 & ~w14209 ) | ( w14203 & ~w14209 ) ;
  assign w14211 = w7517 & w14210 ;
  assign w14212 = w13725 | w13730 ;
  assign w14213 = w14077 & ~w14212 ;
  assign w14214 = w13728 ^ w14213 ;
  assign w14215 = ( ~w7517 & w14203 ) | ( ~w7517 & w14209 ) | ( w14203 & w14209 ) ;
  assign w14216 = ~w14203 & w14215 ;
  assign w14217 = w14214 | w14216 ;
  assign w14218 = ( w7175 & w14211 ) | ( w7175 & ~w14217 ) | ( w14211 & ~w14217 ) ;
  assign w14219 = w7175 & w14218 ;
  assign w14220 = w13733 | w13738 ;
  assign w14221 = w14077 & ~w14220 ;
  assign w14222 = w13736 ^ w14221 ;
  assign w14223 = ( ~w7175 & w14211 ) | ( ~w7175 & w14217 ) | ( w14211 & w14217 ) ;
  assign w14224 = ~w14211 & w14223 ;
  assign w14225 = w14222 | w14224 ;
  assign w14226 = ( w6841 & w14219 ) | ( w6841 & ~w14225 ) | ( w14219 & ~w14225 ) ;
  assign w14227 = w6841 & w14226 ;
  assign w14228 = w13741 | w13746 ;
  assign w14229 = w14077 & ~w14228 ;
  assign w14230 = w13744 ^ w14229 ;
  assign w14231 = ( ~w6841 & w14219 ) | ( ~w6841 & w14225 ) | ( w14219 & w14225 ) ;
  assign w14232 = ~w14219 & w14231 ;
  assign w14233 = w14230 | w14232 ;
  assign w14234 = ( w6515 & w14227 ) | ( w6515 & ~w14233 ) | ( w14227 & ~w14233 ) ;
  assign w14235 = w6515 & w14234 ;
  assign w14236 = w13749 | w13754 ;
  assign w14237 = w14077 & ~w14236 ;
  assign w14238 = w13752 ^ w14237 ;
  assign w14239 = ( ~w6515 & w14227 ) | ( ~w6515 & w14233 ) | ( w14227 & w14233 ) ;
  assign w14240 = ~w14227 & w14239 ;
  assign w14241 = w14238 | w14240 ;
  assign w14242 = ( w6197 & w14235 ) | ( w6197 & ~w14241 ) | ( w14235 & ~w14241 ) ;
  assign w14243 = w6197 & w14242 ;
  assign w14244 = w13757 | w13762 ;
  assign w14245 = w14077 & ~w14244 ;
  assign w14246 = w13760 ^ w14245 ;
  assign w14247 = ( ~w6197 & w14235 ) | ( ~w6197 & w14241 ) | ( w14235 & w14241 ) ;
  assign w14248 = ~w14235 & w14247 ;
  assign w14249 = w14246 | w14248 ;
  assign w14250 = ( w5887 & w14243 ) | ( w5887 & ~w14249 ) | ( w14243 & ~w14249 ) ;
  assign w14251 = w5887 & w14250 ;
  assign w14252 = w13765 | w13770 ;
  assign w14253 = w14077 & ~w14252 ;
  assign w14254 = w13768 ^ w14253 ;
  assign w14255 = ( ~w5887 & w14243 ) | ( ~w5887 & w14249 ) | ( w14243 & w14249 ) ;
  assign w14256 = ~w14243 & w14255 ;
  assign w14257 = w14254 | w14256 ;
  assign w14258 = ( w5585 & w14251 ) | ( w5585 & ~w14257 ) | ( w14251 & ~w14257 ) ;
  assign w14259 = w5585 & w14258 ;
  assign w14260 = w13773 | w13778 ;
  assign w14261 = w14077 & ~w14260 ;
  assign w14262 = w13776 ^ w14261 ;
  assign w14263 = ( ~w5585 & w14251 ) | ( ~w5585 & w14257 ) | ( w14251 & w14257 ) ;
  assign w14264 = ~w14251 & w14263 ;
  assign w14265 = w14262 | w14264 ;
  assign w14266 = ( w5291 & w14259 ) | ( w5291 & ~w14265 ) | ( w14259 & ~w14265 ) ;
  assign w14267 = w5291 & w14266 ;
  assign w14268 = w13781 | w13786 ;
  assign w14269 = w14077 & ~w14268 ;
  assign w14270 = w13784 ^ w14269 ;
  assign w14271 = ( ~w5291 & w14259 ) | ( ~w5291 & w14265 ) | ( w14259 & w14265 ) ;
  assign w14272 = ~w14259 & w14271 ;
  assign w14273 = w14270 | w14272 ;
  assign w14274 = ( w5005 & w14267 ) | ( w5005 & ~w14273 ) | ( w14267 & ~w14273 ) ;
  assign w14275 = w5005 & w14274 ;
  assign w14276 = w13789 | w13794 ;
  assign w14277 = w14077 & ~w14276 ;
  assign w14278 = w13792 ^ w14277 ;
  assign w14279 = ( ~w5005 & w14267 ) | ( ~w5005 & w14273 ) | ( w14267 & w14273 ) ;
  assign w14280 = ~w14267 & w14279 ;
  assign w14281 = w14278 | w14280 ;
  assign w14282 = ( w4727 & w14275 ) | ( w4727 & ~w14281 ) | ( w14275 & ~w14281 ) ;
  assign w14283 = w4727 & w14282 ;
  assign w14284 = w13797 | w13802 ;
  assign w14285 = w14077 & ~w14284 ;
  assign w14286 = w13800 ^ w14285 ;
  assign w14287 = ( ~w4727 & w14275 ) | ( ~w4727 & w14281 ) | ( w14275 & w14281 ) ;
  assign w14288 = ~w14275 & w14287 ;
  assign w14289 = w14286 | w14288 ;
  assign w14290 = ( w4457 & w14283 ) | ( w4457 & ~w14289 ) | ( w14283 & ~w14289 ) ;
  assign w14291 = w4457 & w14290 ;
  assign w14292 = w13805 | w13810 ;
  assign w14293 = w14077 & ~w14292 ;
  assign w14294 = w13808 ^ w14293 ;
  assign w14295 = ( ~w4457 & w14283 ) | ( ~w4457 & w14289 ) | ( w14283 & w14289 ) ;
  assign w14296 = ~w14283 & w14295 ;
  assign w14297 = w14294 | w14296 ;
  assign w14298 = ( w4195 & w14291 ) | ( w4195 & ~w14297 ) | ( w14291 & ~w14297 ) ;
  assign w14299 = w4195 & w14298 ;
  assign w14300 = w13813 | w13818 ;
  assign w14301 = w14077 & ~w14300 ;
  assign w14302 = w13816 ^ w14301 ;
  assign w14303 = ( ~w4195 & w14291 ) | ( ~w4195 & w14297 ) | ( w14291 & w14297 ) ;
  assign w14304 = ~w14291 & w14303 ;
  assign w14305 = w14302 | w14304 ;
  assign w14306 = ( w3941 & w14299 ) | ( w3941 & ~w14305 ) | ( w14299 & ~w14305 ) ;
  assign w14307 = w3941 & w14306 ;
  assign w14308 = w13821 | w13826 ;
  assign w14309 = w14077 & ~w14308 ;
  assign w14310 = w13824 ^ w14309 ;
  assign w14311 = ( ~w3941 & w14299 ) | ( ~w3941 & w14305 ) | ( w14299 & w14305 ) ;
  assign w14312 = ~w14299 & w14311 ;
  assign w14313 = w14310 | w14312 ;
  assign w14314 = ( w3695 & w14307 ) | ( w3695 & ~w14313 ) | ( w14307 & ~w14313 ) ;
  assign w14315 = w3695 & w14314 ;
  assign w14316 = w13829 | w13834 ;
  assign w14317 = w14077 & ~w14316 ;
  assign w14318 = w13832 ^ w14317 ;
  assign w14319 = ( ~w3695 & w14307 ) | ( ~w3695 & w14313 ) | ( w14307 & w14313 ) ;
  assign w14320 = ~w14307 & w14319 ;
  assign w14321 = w14318 | w14320 ;
  assign w14322 = ( w3457 & w14315 ) | ( w3457 & ~w14321 ) | ( w14315 & ~w14321 ) ;
  assign w14323 = w3457 & w14322 ;
  assign w14324 = w13837 | w13842 ;
  assign w14325 = w14077 & ~w14324 ;
  assign w14326 = w13840 ^ w14325 ;
  assign w14327 = ( ~w3457 & w14315 ) | ( ~w3457 & w14321 ) | ( w14315 & w14321 ) ;
  assign w14328 = ~w14315 & w14327 ;
  assign w14329 = w14326 | w14328 ;
  assign w14330 = ( w3227 & w14323 ) | ( w3227 & ~w14329 ) | ( w14323 & ~w14329 ) ;
  assign w14331 = w3227 & w14330 ;
  assign w14332 = w13845 | w13850 ;
  assign w14333 = w14077 & ~w14332 ;
  assign w14334 = w13848 ^ w14333 ;
  assign w14335 = ( ~w3227 & w14323 ) | ( ~w3227 & w14329 ) | ( w14323 & w14329 ) ;
  assign w14336 = ~w14323 & w14335 ;
  assign w14337 = w14334 | w14336 ;
  assign w14338 = ( w3005 & w14331 ) | ( w3005 & ~w14337 ) | ( w14331 & ~w14337 ) ;
  assign w14339 = w3005 & w14338 ;
  assign w14340 = w13853 | w13858 ;
  assign w14341 = w14077 & ~w14340 ;
  assign w14342 = w13856 ^ w14341 ;
  assign w14343 = ( ~w3005 & w14331 ) | ( ~w3005 & w14337 ) | ( w14331 & w14337 ) ;
  assign w14344 = ~w14331 & w14343 ;
  assign w14345 = w14342 | w14344 ;
  assign w14346 = ( w2791 & w14339 ) | ( w2791 & ~w14345 ) | ( w14339 & ~w14345 ) ;
  assign w14347 = w2791 & w14346 ;
  assign w14348 = w13861 | w13866 ;
  assign w14349 = w14077 & ~w14348 ;
  assign w14350 = w13864 ^ w14349 ;
  assign w14351 = ( ~w2791 & w14339 ) | ( ~w2791 & w14345 ) | ( w14339 & w14345 ) ;
  assign w14352 = ~w14339 & w14351 ;
  assign w14353 = w14350 | w14352 ;
  assign w14354 = ( w2585 & w14347 ) | ( w2585 & ~w14353 ) | ( w14347 & ~w14353 ) ;
  assign w14355 = w2585 & w14354 ;
  assign w14356 = w13869 | w13874 ;
  assign w14357 = w14077 & ~w14356 ;
  assign w14358 = w13872 ^ w14357 ;
  assign w14359 = ( ~w2585 & w14347 ) | ( ~w2585 & w14353 ) | ( w14347 & w14353 ) ;
  assign w14360 = ~w14347 & w14359 ;
  assign w14361 = w14358 | w14360 ;
  assign w14362 = ( w2387 & w14355 ) | ( w2387 & ~w14361 ) | ( w14355 & ~w14361 ) ;
  assign w14363 = w2387 & w14362 ;
  assign w14364 = w13877 | w13882 ;
  assign w14365 = w14077 & ~w14364 ;
  assign w14366 = w13880 ^ w14365 ;
  assign w14367 = ( ~w2387 & w14355 ) | ( ~w2387 & w14361 ) | ( w14355 & w14361 ) ;
  assign w14368 = ~w14355 & w14367 ;
  assign w14369 = w14366 | w14368 ;
  assign w14370 = ( w2197 & w14363 ) | ( w2197 & ~w14369 ) | ( w14363 & ~w14369 ) ;
  assign w14371 = w2197 & w14370 ;
  assign w14372 = w13885 | w13890 ;
  assign w14373 = w14077 & ~w14372 ;
  assign w14374 = w13888 ^ w14373 ;
  assign w14375 = ( ~w2197 & w14363 ) | ( ~w2197 & w14369 ) | ( w14363 & w14369 ) ;
  assign w14376 = ~w14363 & w14375 ;
  assign w14377 = w14374 | w14376 ;
  assign w14378 = ( w2015 & w14371 ) | ( w2015 & ~w14377 ) | ( w14371 & ~w14377 ) ;
  assign w14379 = w2015 & w14378 ;
  assign w14380 = w13893 | w13898 ;
  assign w14381 = w14077 & ~w14380 ;
  assign w14382 = w13896 ^ w14381 ;
  assign w14383 = ( ~w2015 & w14371 ) | ( ~w2015 & w14377 ) | ( w14371 & w14377 ) ;
  assign w14384 = ~w14371 & w14383 ;
  assign w14385 = w14382 | w14384 ;
  assign w14386 = ( w1841 & w14379 ) | ( w1841 & ~w14385 ) | ( w14379 & ~w14385 ) ;
  assign w14387 = w1841 & w14386 ;
  assign w14388 = w13901 | w13906 ;
  assign w14389 = w14077 & ~w14388 ;
  assign w14390 = w13904 ^ w14389 ;
  assign w14391 = ( ~w1841 & w14379 ) | ( ~w1841 & w14385 ) | ( w14379 & w14385 ) ;
  assign w14392 = ~w14379 & w14391 ;
  assign w14393 = w14390 | w14392 ;
  assign w14394 = ( w1675 & w14387 ) | ( w1675 & ~w14393 ) | ( w14387 & ~w14393 ) ;
  assign w14395 = w1675 & w14394 ;
  assign w14396 = w13909 | w13914 ;
  assign w14397 = w14077 & ~w14396 ;
  assign w14398 = w13912 ^ w14397 ;
  assign w14399 = ( ~w1675 & w14387 ) | ( ~w1675 & w14393 ) | ( w14387 & w14393 ) ;
  assign w14400 = ~w14387 & w14399 ;
  assign w14401 = w14398 | w14400 ;
  assign w14402 = ( w1517 & w14395 ) | ( w1517 & ~w14401 ) | ( w14395 & ~w14401 ) ;
  assign w14403 = w1517 & w14402 ;
  assign w14404 = w13917 | w13922 ;
  assign w14405 = w14077 & ~w14404 ;
  assign w14406 = w13920 ^ w14405 ;
  assign w14407 = ( ~w1517 & w14395 ) | ( ~w1517 & w14401 ) | ( w14395 & w14401 ) ;
  assign w14408 = ~w14395 & w14407 ;
  assign w14409 = w14406 | w14408 ;
  assign w14410 = ( w1367 & w14403 ) | ( w1367 & ~w14409 ) | ( w14403 & ~w14409 ) ;
  assign w14411 = w1367 & w14410 ;
  assign w14412 = w13925 | w13930 ;
  assign w14413 = w14077 & ~w14412 ;
  assign w14414 = w13928 ^ w14413 ;
  assign w14415 = ( ~w1367 & w14403 ) | ( ~w1367 & w14409 ) | ( w14403 & w14409 ) ;
  assign w14416 = ~w14403 & w14415 ;
  assign w14417 = w14414 | w14416 ;
  assign w14418 = ( w1225 & w14411 ) | ( w1225 & ~w14417 ) | ( w14411 & ~w14417 ) ;
  assign w14419 = w1225 & w14418 ;
  assign w14420 = w13933 | w13938 ;
  assign w14421 = w14077 & ~w14420 ;
  assign w14422 = w13936 ^ w14421 ;
  assign w14423 = ( ~w1225 & w14411 ) | ( ~w1225 & w14417 ) | ( w14411 & w14417 ) ;
  assign w14424 = ~w14411 & w14423 ;
  assign w14425 = w14422 | w14424 ;
  assign w14426 = ( w1091 & w14419 ) | ( w1091 & ~w14425 ) | ( w14419 & ~w14425 ) ;
  assign w14427 = w1091 & w14426 ;
  assign w14428 = w13941 | w13946 ;
  assign w14429 = w14077 & ~w14428 ;
  assign w14430 = w13944 ^ w14429 ;
  assign w14431 = ( ~w1091 & w14419 ) | ( ~w1091 & w14425 ) | ( w14419 & w14425 ) ;
  assign w14432 = ~w14419 & w14431 ;
  assign w14433 = w14430 | w14432 ;
  assign w14434 = ( w965 & w14427 ) | ( w965 & ~w14433 ) | ( w14427 & ~w14433 ) ;
  assign w14435 = w965 & w14434 ;
  assign w14436 = w13949 | w13954 ;
  assign w14437 = w14077 & ~w14436 ;
  assign w14438 = w13952 ^ w14437 ;
  assign w14439 = ( ~w965 & w14427 ) | ( ~w965 & w14433 ) | ( w14427 & w14433 ) ;
  assign w14440 = ~w14427 & w14439 ;
  assign w14441 = w14438 | w14440 ;
  assign w14442 = ( w847 & w14435 ) | ( w847 & ~w14441 ) | ( w14435 & ~w14441 ) ;
  assign w14443 = w847 & w14442 ;
  assign w14444 = w13957 | w13962 ;
  assign w14445 = w14077 & ~w14444 ;
  assign w14446 = w13960 ^ w14445 ;
  assign w14447 = ( ~w847 & w14435 ) | ( ~w847 & w14441 ) | ( w14435 & w14441 ) ;
  assign w14448 = ~w14435 & w14447 ;
  assign w14449 = w14446 | w14448 ;
  assign w14450 = ( w737 & w14443 ) | ( w737 & ~w14449 ) | ( w14443 & ~w14449 ) ;
  assign w14451 = w737 & w14450 ;
  assign w14452 = w13965 | w13970 ;
  assign w14453 = w14077 & ~w14452 ;
  assign w14454 = w13968 ^ w14453 ;
  assign w14455 = ( ~w737 & w14443 ) | ( ~w737 & w14449 ) | ( w14443 & w14449 ) ;
  assign w14456 = ~w14443 & w14455 ;
  assign w14457 = w14454 | w14456 ;
  assign w14458 = ( w635 & w14451 ) | ( w635 & ~w14457 ) | ( w14451 & ~w14457 ) ;
  assign w14459 = w635 & w14458 ;
  assign w14460 = w13973 | w13978 ;
  assign w14461 = w14077 & ~w14460 ;
  assign w14462 = w13976 ^ w14461 ;
  assign w14463 = ( ~w635 & w14451 ) | ( ~w635 & w14457 ) | ( w14451 & w14457 ) ;
  assign w14464 = ~w14451 & w14463 ;
  assign w14465 = w14462 | w14464 ;
  assign w14466 = ( w541 & w14459 ) | ( w541 & ~w14465 ) | ( w14459 & ~w14465 ) ;
  assign w14467 = w541 & w14466 ;
  assign w14468 = w13981 | w13986 ;
  assign w14469 = w14077 & ~w14468 ;
  assign w14470 = w13984 ^ w14469 ;
  assign w14471 = ( ~w541 & w14459 ) | ( ~w541 & w14465 ) | ( w14459 & w14465 ) ;
  assign w14472 = ~w14459 & w14471 ;
  assign w14473 = w14470 | w14472 ;
  assign w14474 = ( w455 & w14467 ) | ( w455 & ~w14473 ) | ( w14467 & ~w14473 ) ;
  assign w14475 = w455 & w14474 ;
  assign w14476 = w13989 | w13994 ;
  assign w14477 = w14077 & ~w14476 ;
  assign w14478 = w13992 ^ w14477 ;
  assign w14479 = ( ~w455 & w14467 ) | ( ~w455 & w14473 ) | ( w14467 & w14473 ) ;
  assign w14480 = ~w14467 & w14479 ;
  assign w14481 = w14478 | w14480 ;
  assign w14482 = ( w377 & w14475 ) | ( w377 & ~w14481 ) | ( w14475 & ~w14481 ) ;
  assign w14483 = w377 & w14482 ;
  assign w14484 = w13997 | w14002 ;
  assign w14485 = w14077 & ~w14484 ;
  assign w14486 = w14000 ^ w14485 ;
  assign w14487 = ( ~w377 & w14475 ) | ( ~w377 & w14481 ) | ( w14475 & w14481 ) ;
  assign w14488 = ~w14475 & w14487 ;
  assign w14489 = w14486 | w14488 ;
  assign w14490 = ( w307 & w14483 ) | ( w307 & ~w14489 ) | ( w14483 & ~w14489 ) ;
  assign w14491 = w307 & w14490 ;
  assign w14492 = ( ~w307 & w14483 ) | ( ~w307 & w14489 ) | ( w14483 & w14489 ) ;
  assign w14493 = ~w14483 & w14492 ;
  assign w14494 = w14005 | w14007 ;
  assign w14495 = w14077 & ~w14494 ;
  assign w14496 = w14010 ^ w14495 ;
  assign w14497 = w14493 | w14496 ;
  assign w14498 = ( w246 & w14491 ) | ( w246 & ~w14497 ) | ( w14491 & ~w14497 ) ;
  assign w14499 = w246 & w14498 ;
  assign w14500 = w14013 | w14018 ;
  assign w14501 = w14077 & ~w14500 ;
  assign w14502 = w14016 ^ w14501 ;
  assign w14503 = ( ~w246 & w14491 ) | ( ~w246 & w14497 ) | ( w14491 & w14497 ) ;
  assign w14504 = ~w14491 & w14503 ;
  assign w14505 = w14502 | w14504 ;
  assign w14506 = ( w185 & w14499 ) | ( w185 & ~w14505 ) | ( w14499 & ~w14505 ) ;
  assign w14507 = w185 & w14506 ;
  assign w14508 = w14021 | w14026 ;
  assign w14509 = w14077 & ~w14508 ;
  assign w14510 = w14024 ^ w14509 ;
  assign w14511 = ( ~w185 & w14499 ) | ( ~w185 & w14505 ) | ( w14499 & w14505 ) ;
  assign w14512 = ~w14499 & w14511 ;
  assign w14513 = w14510 | w14512 ;
  assign w14514 = ( w145 & w14507 ) | ( w145 & ~w14513 ) | ( w14507 & ~w14513 ) ;
  assign w14515 = w145 & w14514 ;
  assign w14516 = w14029 | w14034 ;
  assign w14517 = w14077 & ~w14516 ;
  assign w14518 = w14032 ^ w14517 ;
  assign w14519 = ( ~w145 & w14507 ) | ( ~w145 & w14513 ) | ( w14507 & w14513 ) ;
  assign w14520 = ~w14507 & w14519 ;
  assign w14521 = w14518 | w14520 ;
  assign w14522 = ( w132 & w14515 ) | ( w132 & ~w14521 ) | ( w14515 & ~w14521 ) ;
  assign w14523 = w132 & w14522 ;
  assign w14524 = w14037 | w14042 ;
  assign w14525 = w14077 & ~w14524 ;
  assign w14526 = w14040 ^ w14525 ;
  assign w14527 = ( ~w132 & w14515 ) | ( ~w132 & w14521 ) | ( w14515 & w14521 ) ;
  assign w14528 = ~w14515 & w14527 ;
  assign w14529 = w14526 | w14528 ;
  assign w14530 = ~w14523 & w14529 ;
  assign w14531 = w14045 | w14050 ;
  assign w14532 = w14077 & ~w14531 ;
  assign w14533 = w14048 ^ w14532 ;
  assign w14534 = ( ~w14063 & w14530 ) | ( ~w14063 & w14533 ) | ( w14530 & w14533 ) ;
  assign w14535 = w14052 & ~w14534 ;
  assign w14536 = ~w14055 & w14077 ;
  assign w14537 = ( w14534 & ~w14535 ) | ( w14534 & w14536 ) | ( ~w14535 & w14536 ) ;
  assign w14538 = w14063 | w14537 ;
  assign w14539 = ~w129 & w14538 ;
  assign w14540 = ( w14523 & w14529 ) | ( w14523 & w14533 ) | ( w14529 & w14533 ) ;
  assign w14541 = ~w14523 & w14540 ;
  assign w14542 = ( w129 & w14052 ) | ( w129 & w14055 ) | ( w14052 & w14055 ) ;
  assign w14543 = ( w14055 & ~w14077 ) | ( w14055 & w14542 ) | ( ~w14077 & w14542 ) ;
  assign w14544 = w14052 & w14543 ;
  assign w14545 = w14542 ^ w14544 ;
  assign w14546 = ( w13575 & w13580 ) | ( w13575 & w13607 ) | ( w13580 & w13607 ) ;
  assign w14547 = w13607 & ~w14546 ;
  assign w14548 = w13578 ^ w14547 ;
  assign w14549 = ( ~w14067 & w14074 ) | ( ~w14067 & w14548 ) | ( w14074 & w14548 ) ;
  assign w14550 = ~w14074 & w14549 ;
  assign w14551 = ( ~w14061 & w14063 ) | ( ~w14061 & w14550 ) | ( w14063 & w14550 ) ;
  assign w14552 = ~w14063 & w14551 ;
  assign w14553 = w14541 | w14552 ;
  assign w14554 = ( w14539 & ~w14541 ) | ( w14539 & w14545 ) | ( ~w14541 & w14545 ) ;
  assign w14555 = w14553 | w14554 ;
  assign w14556 = \pi010 | \pi011 ;
  assign w14557 = ( \pi012 & w14077 ) | ( \pi012 & ~w14556 ) | ( w14077 & ~w14556 ) ;
  assign w14558 = ( ~\pi012 & w14077 ) | ( ~\pi012 & w14555 ) | ( w14077 & w14555 ) ;
  assign w14559 = w14557 & w14558 ;
  assign w14560 = w14063 | w14067 ;
  assign w14561 = ( \pi012 & w14556 ) | ( \pi012 & ~w14560 ) | ( w14556 & ~w14560 ) ;
  assign w14562 = ( ~w14074 & w14560 ) | ( ~w14074 & w14561 ) | ( w14560 & w14561 ) ;
  assign w14563 = ~w14560 & w14562 ;
  assign w14564 = ~w14061 & w14563 ;
  assign w14565 = ( \pi012 & w14555 ) | ( \pi012 & ~w14563 ) | ( w14555 & ~w14563 ) ;
  assign w14566 = w14564 & ~w14565 ;
  assign w14567 = ~\pi012 & w14555 ;
  assign w14568 = \pi013 ^ w14567 ;
  assign w14569 = w14566 | w14568 ;
  assign w14570 = ( w13607 & w14559 ) | ( w13607 & ~w14569 ) | ( w14559 & ~w14569 ) ;
  assign w14571 = w13607 & w14570 ;
  assign w14572 = ( ~w13607 & w14559 ) | ( ~w13607 & w14569 ) | ( w14559 & w14569 ) ;
  assign w14573 = ~w14559 & w14572 ;
  assign w14574 = w14077 & ~w14552 ;
  assign w14575 = ~w14541 & w14574 ;
  assign w14576 = ~w14554 & w14575 ;
  assign w14577 = \pi013 & w14555 ;
  assign w14578 = ( \pi012 & w14555 ) | ( \pi012 & ~w14577 ) | ( w14555 & ~w14577 ) ;
  assign w14579 = ( ~\pi012 & w14576 ) | ( ~\pi012 & w14578 ) | ( w14576 & w14578 ) ;
  assign w14580 = \pi014 ^ w14579 ;
  assign w14581 = w14573 | w14580 ;
  assign w14582 = ( w13145 & w14571 ) | ( w13145 & ~w14581 ) | ( w14571 & ~w14581 ) ;
  assign w14583 = w13145 & w14582 ;
  assign w14584 = ( w14081 & ~w14089 ) | ( w14081 & w14555 ) | ( ~w14089 & w14555 ) ;
  assign w14585 = ~w14081 & w14584 ;
  assign w14586 = \pi015 ^ w14585 ;
  assign w14587 = w14090 ^ w14586 ;
  assign w14588 = ( ~w13145 & w14571 ) | ( ~w13145 & w14581 ) | ( w14571 & w14581 ) ;
  assign w14589 = ~w14571 & w14588 ;
  assign w14590 = w14587 | w14589 ;
  assign w14591 = ( w12691 & w14583 ) | ( w12691 & ~w14590 ) | ( w14583 & ~w14590 ) ;
  assign w14592 = w12691 & w14591 ;
  assign w14593 = w14094 | w14096 ;
  assign w14594 = w14555 & ~w14593 ;
  assign w14595 = w14103 ^ w14594 ;
  assign w14596 = ( ~w12691 & w14583 ) | ( ~w12691 & w14590 ) | ( w14583 & w14590 ) ;
  assign w14597 = ~w14583 & w14596 ;
  assign w14598 = w14595 | w14597 ;
  assign w14599 = ( w12245 & w14592 ) | ( w12245 & ~w14598 ) | ( w14592 & ~w14598 ) ;
  assign w14600 = w12245 & w14599 ;
  assign w14601 = w14106 | w14112 ;
  assign w14602 = w14555 & ~w14601 ;
  assign w14603 = w14110 ^ w14602 ;
  assign w14604 = ( ~w12245 & w14592 ) | ( ~w12245 & w14598 ) | ( w14592 & w14598 ) ;
  assign w14605 = ~w14592 & w14604 ;
  assign w14606 = w14603 | w14605 ;
  assign w14607 = ( w11807 & w14600 ) | ( w11807 & ~w14606 ) | ( w14600 & ~w14606 ) ;
  assign w14608 = w11807 & w14607 ;
  assign w14609 = w14115 | w14120 ;
  assign w14610 = w14555 & ~w14609 ;
  assign w14611 = w14118 ^ w14610 ;
  assign w14612 = ( ~w11807 & w14600 ) | ( ~w11807 & w14606 ) | ( w14600 & w14606 ) ;
  assign w14613 = ~w14600 & w14612 ;
  assign w14614 = w14611 | w14613 ;
  assign w14615 = ( w11377 & w14608 ) | ( w11377 & ~w14614 ) | ( w14608 & ~w14614 ) ;
  assign w14616 = w11377 & w14615 ;
  assign w14617 = w14123 | w14128 ;
  assign w14618 = w14555 & ~w14617 ;
  assign w14619 = w14126 ^ w14618 ;
  assign w14620 = ( ~w11377 & w14608 ) | ( ~w11377 & w14614 ) | ( w14608 & w14614 ) ;
  assign w14621 = ~w14608 & w14620 ;
  assign w14622 = w14619 | w14621 ;
  assign w14623 = ( w10955 & w14616 ) | ( w10955 & ~w14622 ) | ( w14616 & ~w14622 ) ;
  assign w14624 = w10955 & w14623 ;
  assign w14625 = w14131 | w14136 ;
  assign w14626 = w14555 & ~w14625 ;
  assign w14627 = w14134 ^ w14626 ;
  assign w14628 = ( ~w10955 & w14616 ) | ( ~w10955 & w14622 ) | ( w14616 & w14622 ) ;
  assign w14629 = ~w14616 & w14628 ;
  assign w14630 = w14627 | w14629 ;
  assign w14631 = ( w10541 & w14624 ) | ( w10541 & ~w14630 ) | ( w14624 & ~w14630 ) ;
  assign w14632 = w10541 & w14631 ;
  assign w14633 = w14139 | w14144 ;
  assign w14634 = w14555 & ~w14633 ;
  assign w14635 = w14142 ^ w14634 ;
  assign w14636 = ( ~w10541 & w14624 ) | ( ~w10541 & w14630 ) | ( w14624 & w14630 ) ;
  assign w14637 = ~w14624 & w14636 ;
  assign w14638 = w14635 | w14637 ;
  assign w14639 = ( w10135 & w14632 ) | ( w10135 & ~w14638 ) | ( w14632 & ~w14638 ) ;
  assign w14640 = w10135 & w14639 ;
  assign w14641 = w14147 | w14152 ;
  assign w14642 = w14555 & ~w14641 ;
  assign w14643 = w14150 ^ w14642 ;
  assign w14644 = ( ~w10135 & w14632 ) | ( ~w10135 & w14638 ) | ( w14632 & w14638 ) ;
  assign w14645 = ~w14632 & w14644 ;
  assign w14646 = w14643 | w14645 ;
  assign w14647 = ( w9737 & w14640 ) | ( w9737 & ~w14646 ) | ( w14640 & ~w14646 ) ;
  assign w14648 = w9737 & w14647 ;
  assign w14649 = w14155 | w14160 ;
  assign w14650 = w14555 & ~w14649 ;
  assign w14651 = w14158 ^ w14650 ;
  assign w14652 = ( ~w9737 & w14640 ) | ( ~w9737 & w14646 ) | ( w14640 & w14646 ) ;
  assign w14653 = ~w14640 & w14652 ;
  assign w14654 = w14651 | w14653 ;
  assign w14655 = ( w9347 & w14648 ) | ( w9347 & ~w14654 ) | ( w14648 & ~w14654 ) ;
  assign w14656 = w9347 & w14655 ;
  assign w14657 = w14163 | w14168 ;
  assign w14658 = w14555 & ~w14657 ;
  assign w14659 = w14166 ^ w14658 ;
  assign w14660 = ( ~w9347 & w14648 ) | ( ~w9347 & w14654 ) | ( w14648 & w14654 ) ;
  assign w14661 = ~w14648 & w14660 ;
  assign w14662 = w14659 | w14661 ;
  assign w14663 = ( w8965 & w14656 ) | ( w8965 & ~w14662 ) | ( w14656 & ~w14662 ) ;
  assign w14664 = w8965 & w14663 ;
  assign w14665 = w14171 | w14176 ;
  assign w14666 = w14555 & ~w14665 ;
  assign w14667 = w14174 ^ w14666 ;
  assign w14668 = ( ~w8965 & w14656 ) | ( ~w8965 & w14662 ) | ( w14656 & w14662 ) ;
  assign w14669 = ~w14656 & w14668 ;
  assign w14670 = w14667 | w14669 ;
  assign w14671 = ( w8591 & w14664 ) | ( w8591 & ~w14670 ) | ( w14664 & ~w14670 ) ;
  assign w14672 = w8591 & w14671 ;
  assign w14673 = w14179 | w14184 ;
  assign w14674 = w14555 & ~w14673 ;
  assign w14675 = w14182 ^ w14674 ;
  assign w14676 = ( ~w8591 & w14664 ) | ( ~w8591 & w14670 ) | ( w14664 & w14670 ) ;
  assign w14677 = ~w14664 & w14676 ;
  assign w14678 = w14675 | w14677 ;
  assign w14679 = ( w8225 & w14672 ) | ( w8225 & ~w14678 ) | ( w14672 & ~w14678 ) ;
  assign w14680 = w8225 & w14679 ;
  assign w14681 = w14187 | w14192 ;
  assign w14682 = w14555 & ~w14681 ;
  assign w14683 = w14190 ^ w14682 ;
  assign w14684 = ( ~w8225 & w14672 ) | ( ~w8225 & w14678 ) | ( w14672 & w14678 ) ;
  assign w14685 = ~w14672 & w14684 ;
  assign w14686 = w14683 | w14685 ;
  assign w14687 = ( w7867 & w14680 ) | ( w7867 & ~w14686 ) | ( w14680 & ~w14686 ) ;
  assign w14688 = w7867 & w14687 ;
  assign w14689 = w14195 | w14200 ;
  assign w14690 = w14555 & ~w14689 ;
  assign w14691 = w14198 ^ w14690 ;
  assign w14692 = ( ~w7867 & w14680 ) | ( ~w7867 & w14686 ) | ( w14680 & w14686 ) ;
  assign w14693 = ~w14680 & w14692 ;
  assign w14694 = w14691 | w14693 ;
  assign w14695 = ( w7517 & w14688 ) | ( w7517 & ~w14694 ) | ( w14688 & ~w14694 ) ;
  assign w14696 = w7517 & w14695 ;
  assign w14697 = w14203 | w14208 ;
  assign w14698 = w14555 & ~w14697 ;
  assign w14699 = w14206 ^ w14698 ;
  assign w14700 = ( ~w7517 & w14688 ) | ( ~w7517 & w14694 ) | ( w14688 & w14694 ) ;
  assign w14701 = ~w14688 & w14700 ;
  assign w14702 = w14699 | w14701 ;
  assign w14703 = ( w7175 & w14696 ) | ( w7175 & ~w14702 ) | ( w14696 & ~w14702 ) ;
  assign w14704 = w7175 & w14703 ;
  assign w14705 = w14211 | w14216 ;
  assign w14706 = w14555 & ~w14705 ;
  assign w14707 = w14214 ^ w14706 ;
  assign w14708 = ( ~w7175 & w14696 ) | ( ~w7175 & w14702 ) | ( w14696 & w14702 ) ;
  assign w14709 = ~w14696 & w14708 ;
  assign w14710 = w14707 | w14709 ;
  assign w14711 = ( w6841 & w14704 ) | ( w6841 & ~w14710 ) | ( w14704 & ~w14710 ) ;
  assign w14712 = w6841 & w14711 ;
  assign w14713 = w14219 | w14224 ;
  assign w14714 = w14555 & ~w14713 ;
  assign w14715 = w14222 ^ w14714 ;
  assign w14716 = ( ~w6841 & w14704 ) | ( ~w6841 & w14710 ) | ( w14704 & w14710 ) ;
  assign w14717 = ~w14704 & w14716 ;
  assign w14718 = w14715 | w14717 ;
  assign w14719 = ( w6515 & w14712 ) | ( w6515 & ~w14718 ) | ( w14712 & ~w14718 ) ;
  assign w14720 = w6515 & w14719 ;
  assign w14721 = w14227 | w14232 ;
  assign w14722 = w14555 & ~w14721 ;
  assign w14723 = w14230 ^ w14722 ;
  assign w14724 = ( ~w6515 & w14712 ) | ( ~w6515 & w14718 ) | ( w14712 & w14718 ) ;
  assign w14725 = ~w14712 & w14724 ;
  assign w14726 = w14723 | w14725 ;
  assign w14727 = ( w6197 & w14720 ) | ( w6197 & ~w14726 ) | ( w14720 & ~w14726 ) ;
  assign w14728 = w6197 & w14727 ;
  assign w14729 = w14235 | w14240 ;
  assign w14730 = w14555 & ~w14729 ;
  assign w14731 = w14238 ^ w14730 ;
  assign w14732 = ( ~w6197 & w14720 ) | ( ~w6197 & w14726 ) | ( w14720 & w14726 ) ;
  assign w14733 = ~w14720 & w14732 ;
  assign w14734 = w14731 | w14733 ;
  assign w14735 = ( w5887 & w14728 ) | ( w5887 & ~w14734 ) | ( w14728 & ~w14734 ) ;
  assign w14736 = w5887 & w14735 ;
  assign w14737 = w14243 | w14248 ;
  assign w14738 = w14555 & ~w14737 ;
  assign w14739 = w14246 ^ w14738 ;
  assign w14740 = ( ~w5887 & w14728 ) | ( ~w5887 & w14734 ) | ( w14728 & w14734 ) ;
  assign w14741 = ~w14728 & w14740 ;
  assign w14742 = w14739 | w14741 ;
  assign w14743 = ( w5585 & w14736 ) | ( w5585 & ~w14742 ) | ( w14736 & ~w14742 ) ;
  assign w14744 = w5585 & w14743 ;
  assign w14745 = w14251 | w14256 ;
  assign w14746 = w14555 & ~w14745 ;
  assign w14747 = w14254 ^ w14746 ;
  assign w14748 = ( ~w5585 & w14736 ) | ( ~w5585 & w14742 ) | ( w14736 & w14742 ) ;
  assign w14749 = ~w14736 & w14748 ;
  assign w14750 = w14747 | w14749 ;
  assign w14751 = ( w5291 & w14744 ) | ( w5291 & ~w14750 ) | ( w14744 & ~w14750 ) ;
  assign w14752 = w5291 & w14751 ;
  assign w14753 = w14259 | w14264 ;
  assign w14754 = w14555 & ~w14753 ;
  assign w14755 = w14262 ^ w14754 ;
  assign w14756 = ( ~w5291 & w14744 ) | ( ~w5291 & w14750 ) | ( w14744 & w14750 ) ;
  assign w14757 = ~w14744 & w14756 ;
  assign w14758 = w14755 | w14757 ;
  assign w14759 = ( w5005 & w14752 ) | ( w5005 & ~w14758 ) | ( w14752 & ~w14758 ) ;
  assign w14760 = w5005 & w14759 ;
  assign w14761 = w14267 | w14272 ;
  assign w14762 = w14555 & ~w14761 ;
  assign w14763 = w14270 ^ w14762 ;
  assign w14764 = ( ~w5005 & w14752 ) | ( ~w5005 & w14758 ) | ( w14752 & w14758 ) ;
  assign w14765 = ~w14752 & w14764 ;
  assign w14766 = w14763 | w14765 ;
  assign w14767 = ( w4727 & w14760 ) | ( w4727 & ~w14766 ) | ( w14760 & ~w14766 ) ;
  assign w14768 = w4727 & w14767 ;
  assign w14769 = w14275 | w14280 ;
  assign w14770 = w14555 & ~w14769 ;
  assign w14771 = w14278 ^ w14770 ;
  assign w14772 = ( ~w4727 & w14760 ) | ( ~w4727 & w14766 ) | ( w14760 & w14766 ) ;
  assign w14773 = ~w14760 & w14772 ;
  assign w14774 = w14771 | w14773 ;
  assign w14775 = ( w4457 & w14768 ) | ( w4457 & ~w14774 ) | ( w14768 & ~w14774 ) ;
  assign w14776 = w4457 & w14775 ;
  assign w14777 = w14283 | w14288 ;
  assign w14778 = w14555 & ~w14777 ;
  assign w14779 = w14286 ^ w14778 ;
  assign w14780 = ( ~w4457 & w14768 ) | ( ~w4457 & w14774 ) | ( w14768 & w14774 ) ;
  assign w14781 = ~w14768 & w14780 ;
  assign w14782 = w14779 | w14781 ;
  assign w14783 = ( w4195 & w14776 ) | ( w4195 & ~w14782 ) | ( w14776 & ~w14782 ) ;
  assign w14784 = w4195 & w14783 ;
  assign w14785 = w14291 | w14296 ;
  assign w14786 = w14555 & ~w14785 ;
  assign w14787 = w14294 ^ w14786 ;
  assign w14788 = ( ~w4195 & w14776 ) | ( ~w4195 & w14782 ) | ( w14776 & w14782 ) ;
  assign w14789 = ~w14776 & w14788 ;
  assign w14790 = w14787 | w14789 ;
  assign w14791 = ( w3941 & w14784 ) | ( w3941 & ~w14790 ) | ( w14784 & ~w14790 ) ;
  assign w14792 = w3941 & w14791 ;
  assign w14793 = w14299 | w14304 ;
  assign w14794 = w14555 & ~w14793 ;
  assign w14795 = w14302 ^ w14794 ;
  assign w14796 = ( ~w3941 & w14784 ) | ( ~w3941 & w14790 ) | ( w14784 & w14790 ) ;
  assign w14797 = ~w14784 & w14796 ;
  assign w14798 = w14795 | w14797 ;
  assign w14799 = ( w3695 & w14792 ) | ( w3695 & ~w14798 ) | ( w14792 & ~w14798 ) ;
  assign w14800 = w3695 & w14799 ;
  assign w14801 = w14307 | w14312 ;
  assign w14802 = w14555 & ~w14801 ;
  assign w14803 = w14310 ^ w14802 ;
  assign w14804 = ( ~w3695 & w14792 ) | ( ~w3695 & w14798 ) | ( w14792 & w14798 ) ;
  assign w14805 = ~w14792 & w14804 ;
  assign w14806 = w14803 | w14805 ;
  assign w14807 = ( w3457 & w14800 ) | ( w3457 & ~w14806 ) | ( w14800 & ~w14806 ) ;
  assign w14808 = w3457 & w14807 ;
  assign w14809 = w14315 | w14320 ;
  assign w14810 = w14555 & ~w14809 ;
  assign w14811 = w14318 ^ w14810 ;
  assign w14812 = ( ~w3457 & w14800 ) | ( ~w3457 & w14806 ) | ( w14800 & w14806 ) ;
  assign w14813 = ~w14800 & w14812 ;
  assign w14814 = w14811 | w14813 ;
  assign w14815 = ( w3227 & w14808 ) | ( w3227 & ~w14814 ) | ( w14808 & ~w14814 ) ;
  assign w14816 = w3227 & w14815 ;
  assign w14817 = w14323 | w14328 ;
  assign w14818 = w14555 & ~w14817 ;
  assign w14819 = w14326 ^ w14818 ;
  assign w14820 = ( ~w3227 & w14808 ) | ( ~w3227 & w14814 ) | ( w14808 & w14814 ) ;
  assign w14821 = ~w14808 & w14820 ;
  assign w14822 = w14819 | w14821 ;
  assign w14823 = ( w3005 & w14816 ) | ( w3005 & ~w14822 ) | ( w14816 & ~w14822 ) ;
  assign w14824 = w3005 & w14823 ;
  assign w14825 = w14331 | w14336 ;
  assign w14826 = w14555 & ~w14825 ;
  assign w14827 = w14334 ^ w14826 ;
  assign w14828 = ( ~w3005 & w14816 ) | ( ~w3005 & w14822 ) | ( w14816 & w14822 ) ;
  assign w14829 = ~w14816 & w14828 ;
  assign w14830 = w14827 | w14829 ;
  assign w14831 = ( w2791 & w14824 ) | ( w2791 & ~w14830 ) | ( w14824 & ~w14830 ) ;
  assign w14832 = w2791 & w14831 ;
  assign w14833 = w14339 | w14344 ;
  assign w14834 = w14555 & ~w14833 ;
  assign w14835 = w14342 ^ w14834 ;
  assign w14836 = ( ~w2791 & w14824 ) | ( ~w2791 & w14830 ) | ( w14824 & w14830 ) ;
  assign w14837 = ~w14824 & w14836 ;
  assign w14838 = w14835 | w14837 ;
  assign w14839 = ( w2585 & w14832 ) | ( w2585 & ~w14838 ) | ( w14832 & ~w14838 ) ;
  assign w14840 = w2585 & w14839 ;
  assign w14841 = w14347 | w14352 ;
  assign w14842 = w14555 & ~w14841 ;
  assign w14843 = w14350 ^ w14842 ;
  assign w14844 = ( ~w2585 & w14832 ) | ( ~w2585 & w14838 ) | ( w14832 & w14838 ) ;
  assign w14845 = ~w14832 & w14844 ;
  assign w14846 = w14843 | w14845 ;
  assign w14847 = ( w2387 & w14840 ) | ( w2387 & ~w14846 ) | ( w14840 & ~w14846 ) ;
  assign w14848 = w2387 & w14847 ;
  assign w14849 = w14355 | w14360 ;
  assign w14850 = w14555 & ~w14849 ;
  assign w14851 = w14358 ^ w14850 ;
  assign w14852 = ( ~w2387 & w14840 ) | ( ~w2387 & w14846 ) | ( w14840 & w14846 ) ;
  assign w14853 = ~w14840 & w14852 ;
  assign w14854 = w14851 | w14853 ;
  assign w14855 = ( w2197 & w14848 ) | ( w2197 & ~w14854 ) | ( w14848 & ~w14854 ) ;
  assign w14856 = w2197 & w14855 ;
  assign w14857 = w14363 | w14368 ;
  assign w14858 = w14555 & ~w14857 ;
  assign w14859 = w14366 ^ w14858 ;
  assign w14860 = ( ~w2197 & w14848 ) | ( ~w2197 & w14854 ) | ( w14848 & w14854 ) ;
  assign w14861 = ~w14848 & w14860 ;
  assign w14862 = w14859 | w14861 ;
  assign w14863 = ( w2015 & w14856 ) | ( w2015 & ~w14862 ) | ( w14856 & ~w14862 ) ;
  assign w14864 = w2015 & w14863 ;
  assign w14865 = w14371 | w14376 ;
  assign w14866 = w14555 & ~w14865 ;
  assign w14867 = w14374 ^ w14866 ;
  assign w14868 = ( ~w2015 & w14856 ) | ( ~w2015 & w14862 ) | ( w14856 & w14862 ) ;
  assign w14869 = ~w14856 & w14868 ;
  assign w14870 = w14867 | w14869 ;
  assign w14871 = ( w1841 & w14864 ) | ( w1841 & ~w14870 ) | ( w14864 & ~w14870 ) ;
  assign w14872 = w1841 & w14871 ;
  assign w14873 = w14379 | w14384 ;
  assign w14874 = w14555 & ~w14873 ;
  assign w14875 = w14382 ^ w14874 ;
  assign w14876 = ( ~w1841 & w14864 ) | ( ~w1841 & w14870 ) | ( w14864 & w14870 ) ;
  assign w14877 = ~w14864 & w14876 ;
  assign w14878 = w14875 | w14877 ;
  assign w14879 = ( w1675 & w14872 ) | ( w1675 & ~w14878 ) | ( w14872 & ~w14878 ) ;
  assign w14880 = w1675 & w14879 ;
  assign w14881 = w14387 | w14392 ;
  assign w14882 = w14555 & ~w14881 ;
  assign w14883 = w14390 ^ w14882 ;
  assign w14884 = ( ~w1675 & w14872 ) | ( ~w1675 & w14878 ) | ( w14872 & w14878 ) ;
  assign w14885 = ~w14872 & w14884 ;
  assign w14886 = w14883 | w14885 ;
  assign w14887 = ( w1517 & w14880 ) | ( w1517 & ~w14886 ) | ( w14880 & ~w14886 ) ;
  assign w14888 = w1517 & w14887 ;
  assign w14889 = w14395 | w14400 ;
  assign w14890 = w14555 & ~w14889 ;
  assign w14891 = w14398 ^ w14890 ;
  assign w14892 = ( ~w1517 & w14880 ) | ( ~w1517 & w14886 ) | ( w14880 & w14886 ) ;
  assign w14893 = ~w14880 & w14892 ;
  assign w14894 = w14891 | w14893 ;
  assign w14895 = ( w1367 & w14888 ) | ( w1367 & ~w14894 ) | ( w14888 & ~w14894 ) ;
  assign w14896 = w1367 & w14895 ;
  assign w14897 = w14403 | w14408 ;
  assign w14898 = w14555 & ~w14897 ;
  assign w14899 = w14406 ^ w14898 ;
  assign w14900 = ( ~w1367 & w14888 ) | ( ~w1367 & w14894 ) | ( w14888 & w14894 ) ;
  assign w14901 = ~w14888 & w14900 ;
  assign w14902 = w14899 | w14901 ;
  assign w14903 = ( w1225 & w14896 ) | ( w1225 & ~w14902 ) | ( w14896 & ~w14902 ) ;
  assign w14904 = w1225 & w14903 ;
  assign w14905 = w14411 | w14416 ;
  assign w14906 = w14555 & ~w14905 ;
  assign w14907 = w14414 ^ w14906 ;
  assign w14908 = ( ~w1225 & w14896 ) | ( ~w1225 & w14902 ) | ( w14896 & w14902 ) ;
  assign w14909 = ~w14896 & w14908 ;
  assign w14910 = w14907 | w14909 ;
  assign w14911 = ( w1091 & w14904 ) | ( w1091 & ~w14910 ) | ( w14904 & ~w14910 ) ;
  assign w14912 = w1091 & w14911 ;
  assign w14913 = w14419 | w14424 ;
  assign w14914 = w14555 & ~w14913 ;
  assign w14915 = w14422 ^ w14914 ;
  assign w14916 = ( ~w1091 & w14904 ) | ( ~w1091 & w14910 ) | ( w14904 & w14910 ) ;
  assign w14917 = ~w14904 & w14916 ;
  assign w14918 = w14915 | w14917 ;
  assign w14919 = ( w965 & w14912 ) | ( w965 & ~w14918 ) | ( w14912 & ~w14918 ) ;
  assign w14920 = w965 & w14919 ;
  assign w14921 = w14427 | w14432 ;
  assign w14922 = w14555 & ~w14921 ;
  assign w14923 = w14430 ^ w14922 ;
  assign w14924 = ( ~w965 & w14912 ) | ( ~w965 & w14918 ) | ( w14912 & w14918 ) ;
  assign w14925 = ~w14912 & w14924 ;
  assign w14926 = w14923 | w14925 ;
  assign w14927 = ( w847 & w14920 ) | ( w847 & ~w14926 ) | ( w14920 & ~w14926 ) ;
  assign w14928 = w847 & w14927 ;
  assign w14929 = w14435 | w14440 ;
  assign w14930 = w14555 & ~w14929 ;
  assign w14931 = w14438 ^ w14930 ;
  assign w14932 = ( ~w847 & w14920 ) | ( ~w847 & w14926 ) | ( w14920 & w14926 ) ;
  assign w14933 = ~w14920 & w14932 ;
  assign w14934 = w14931 | w14933 ;
  assign w14935 = ( w737 & w14928 ) | ( w737 & ~w14934 ) | ( w14928 & ~w14934 ) ;
  assign w14936 = w737 & w14935 ;
  assign w14937 = w14443 | w14448 ;
  assign w14938 = w14555 & ~w14937 ;
  assign w14939 = w14446 ^ w14938 ;
  assign w14940 = ( ~w737 & w14928 ) | ( ~w737 & w14934 ) | ( w14928 & w14934 ) ;
  assign w14941 = ~w14928 & w14940 ;
  assign w14942 = w14939 | w14941 ;
  assign w14943 = ( w635 & w14936 ) | ( w635 & ~w14942 ) | ( w14936 & ~w14942 ) ;
  assign w14944 = w635 & w14943 ;
  assign w14945 = w14451 | w14456 ;
  assign w14946 = w14555 & ~w14945 ;
  assign w14947 = w14454 ^ w14946 ;
  assign w14948 = ( ~w635 & w14936 ) | ( ~w635 & w14942 ) | ( w14936 & w14942 ) ;
  assign w14949 = ~w14936 & w14948 ;
  assign w14950 = w14947 | w14949 ;
  assign w14951 = ( w541 & w14944 ) | ( w541 & ~w14950 ) | ( w14944 & ~w14950 ) ;
  assign w14952 = w541 & w14951 ;
  assign w14953 = w14459 | w14464 ;
  assign w14954 = w14555 & ~w14953 ;
  assign w14955 = w14462 ^ w14954 ;
  assign w14956 = ( ~w541 & w14944 ) | ( ~w541 & w14950 ) | ( w14944 & w14950 ) ;
  assign w14957 = ~w14944 & w14956 ;
  assign w14958 = w14955 | w14957 ;
  assign w14959 = ( w455 & w14952 ) | ( w455 & ~w14958 ) | ( w14952 & ~w14958 ) ;
  assign w14960 = w455 & w14959 ;
  assign w14961 = w14467 | w14472 ;
  assign w14962 = w14555 & ~w14961 ;
  assign w14963 = w14470 ^ w14962 ;
  assign w14964 = ( ~w455 & w14952 ) | ( ~w455 & w14958 ) | ( w14952 & w14958 ) ;
  assign w14965 = ~w14952 & w14964 ;
  assign w14966 = w14963 | w14965 ;
  assign w14967 = ( w377 & w14960 ) | ( w377 & ~w14966 ) | ( w14960 & ~w14966 ) ;
  assign w14968 = w377 & w14967 ;
  assign w14969 = w14475 | w14480 ;
  assign w14970 = w14555 & ~w14969 ;
  assign w14971 = w14478 ^ w14970 ;
  assign w14972 = ( ~w377 & w14960 ) | ( ~w377 & w14966 ) | ( w14960 & w14966 ) ;
  assign w14973 = ~w14960 & w14972 ;
  assign w14974 = w14971 | w14973 ;
  assign w14975 = ( w307 & w14968 ) | ( w307 & ~w14974 ) | ( w14968 & ~w14974 ) ;
  assign w14976 = w307 & w14975 ;
  assign w14977 = w14483 | w14488 ;
  assign w14978 = w14555 & ~w14977 ;
  assign w14979 = w14486 ^ w14978 ;
  assign w14980 = ( ~w307 & w14968 ) | ( ~w307 & w14974 ) | ( w14968 & w14974 ) ;
  assign w14981 = ~w14968 & w14980 ;
  assign w14982 = w14979 | w14981 ;
  assign w14983 = ( w246 & w14976 ) | ( w246 & ~w14982 ) | ( w14976 & ~w14982 ) ;
  assign w14984 = w246 & w14983 ;
  assign w14985 = ( ~w246 & w14976 ) | ( ~w246 & w14982 ) | ( w14976 & w14982 ) ;
  assign w14986 = ~w14976 & w14985 ;
  assign w14987 = w14491 | w14493 ;
  assign w14988 = w14555 & ~w14987 ;
  assign w14989 = w14496 ^ w14988 ;
  assign w14990 = w14986 | w14989 ;
  assign w14991 = ( w185 & w14984 ) | ( w185 & ~w14990 ) | ( w14984 & ~w14990 ) ;
  assign w14992 = w185 & w14991 ;
  assign w14993 = w14499 | w14504 ;
  assign w14994 = w14555 & ~w14993 ;
  assign w14995 = w14502 ^ w14994 ;
  assign w14996 = ( ~w185 & w14984 ) | ( ~w185 & w14990 ) | ( w14984 & w14990 ) ;
  assign w14997 = ~w14984 & w14996 ;
  assign w14998 = w14995 | w14997 ;
  assign w14999 = ( w145 & w14992 ) | ( w145 & ~w14998 ) | ( w14992 & ~w14998 ) ;
  assign w15000 = w145 & w14999 ;
  assign w15001 = w14507 | w14512 ;
  assign w15002 = w14555 & ~w15001 ;
  assign w15003 = w14510 ^ w15002 ;
  assign w15004 = ( ~w145 & w14992 ) | ( ~w145 & w14998 ) | ( w14992 & w14998 ) ;
  assign w15005 = ~w14992 & w15004 ;
  assign w15006 = w15003 | w15005 ;
  assign w15007 = ( w132 & w15000 ) | ( w132 & ~w15006 ) | ( w15000 & ~w15006 ) ;
  assign w15008 = w132 & w15007 ;
  assign w15009 = w14515 | w14520 ;
  assign w15010 = w14555 & ~w15009 ;
  assign w15011 = w14518 ^ w15010 ;
  assign w15012 = ( ~w132 & w15000 ) | ( ~w132 & w15006 ) | ( w15000 & w15006 ) ;
  assign w15013 = ~w15000 & w15012 ;
  assign w15014 = w15011 | w15013 ;
  assign w15015 = ~w15008 & w15014 ;
  assign w15016 = w14523 | w14528 ;
  assign w15017 = w14555 & ~w15016 ;
  assign w15018 = w14526 ^ w15017 ;
  assign w15019 = ( ~w14541 & w15015 ) | ( ~w14541 & w15018 ) | ( w15015 & w15018 ) ;
  assign w15020 = w14530 & ~w15019 ;
  assign w15021 = ~w14533 & w14555 ;
  assign w15022 = ( w15019 & ~w15020 ) | ( w15019 & w15021 ) | ( ~w15020 & w15021 ) ;
  assign w15023 = w14541 | w15022 ;
  assign w15024 = ~w129 & w15023 ;
  assign w15025 = ( w15008 & w15014 ) | ( w15008 & w15018 ) | ( w15014 & w15018 ) ;
  assign w15026 = ~w15008 & w15025 ;
  assign w15027 = ( w129 & w14530 ) | ( w129 & w14533 ) | ( w14530 & w14533 ) ;
  assign w15028 = ( w14533 & ~w14555 ) | ( w14533 & w15027 ) | ( ~w14555 & w15027 ) ;
  assign w15029 = w14530 & w15028 ;
  assign w15030 = w15027 ^ w15029 ;
  assign w15031 = ( w15024 & ~w15026 ) | ( w15024 & w15030 ) | ( ~w15026 & w15030 ) ;
  assign w15032 = w15026 | w15031 ;
  assign w15033 = \pi008 | \pi009 ;
  assign w15034 = ( \pi010 & w14555 ) | ( \pi010 & ~w15033 ) | ( w14555 & ~w15033 ) ;
  assign w15035 = ( ~\pi010 & w14555 ) | ( ~\pi010 & w15032 ) | ( w14555 & w15032 ) ;
  assign w15036 = w15034 & w15035 ;
  assign w15037 = w14541 | w14545 ;
  assign w15038 = ( \pi010 & w15033 ) | ( \pi010 & ~w15037 ) | ( w15033 & ~w15037 ) ;
  assign w15039 = ( ~w14552 & w15037 ) | ( ~w14552 & w15038 ) | ( w15037 & w15038 ) ;
  assign w15040 = ~w15037 & w15039 ;
  assign w15041 = ~w14539 & w15040 ;
  assign w15042 = ( \pi010 & w15032 ) | ( \pi010 & ~w15040 ) | ( w15032 & ~w15040 ) ;
  assign w15043 = w15041 & ~w15042 ;
  assign w15044 = ~\pi010 & w15032 ;
  assign w15045 = \pi011 ^ w15044 ;
  assign w15046 = w15043 | w15045 ;
  assign w15047 = ( w14077 & w15036 ) | ( w14077 & ~w15046 ) | ( w15036 & ~w15046 ) ;
  assign w15048 = w14077 & w15047 ;
  assign w15049 = ( ~w14077 & w15036 ) | ( ~w14077 & w15046 ) | ( w15036 & w15046 ) ;
  assign w15050 = ~w15036 & w15049 ;
  assign w15051 = w15024 | w15026 ;
  assign w15052 = w15030 | w15051 ;
  assign w15053 = w14555 ^ w15052 ;
  assign w15054 = ( w14555 & ~w14556 ) | ( w14555 & w15053 ) | ( ~w14556 & w15053 ) ;
  assign w15055 = \pi012 ^ w15054 ;
  assign w15056 = w15050 | w15055 ;
  assign w15057 = ( w13607 & w15048 ) | ( w13607 & ~w15056 ) | ( w15048 & ~w15056 ) ;
  assign w15058 = w13607 & w15057 ;
  assign w15059 = ( w14559 & ~w14566 ) | ( w14559 & w15032 ) | ( ~w14566 & w15032 ) ;
  assign w15060 = ~w14559 & w15059 ;
  assign w15061 = \pi013 ^ w15060 ;
  assign w15062 = w14567 ^ w15061 ;
  assign w15063 = ( ~w13607 & w15048 ) | ( ~w13607 & w15056 ) | ( w15048 & w15056 ) ;
  assign w15064 = ~w15048 & w15063 ;
  assign w15065 = w15062 | w15064 ;
  assign w15066 = ( w13145 & w15058 ) | ( w13145 & ~w15065 ) | ( w15058 & ~w15065 ) ;
  assign w15067 = w13145 & w15066 ;
  assign w15068 = w14571 | w14573 ;
  assign w15069 = w15032 & ~w15068 ;
  assign w15070 = w14580 ^ w15069 ;
  assign w15071 = ( ~w13145 & w15058 ) | ( ~w13145 & w15065 ) | ( w15058 & w15065 ) ;
  assign w15072 = ~w15058 & w15071 ;
  assign w15073 = w15070 | w15072 ;
  assign w15074 = ( w12691 & w15067 ) | ( w12691 & ~w15073 ) | ( w15067 & ~w15073 ) ;
  assign w15075 = w12691 & w15074 ;
  assign w15076 = w14583 | w14589 ;
  assign w15077 = w15032 & ~w15076 ;
  assign w15078 = w14587 ^ w15077 ;
  assign w15079 = ( ~w12691 & w15067 ) | ( ~w12691 & w15073 ) | ( w15067 & w15073 ) ;
  assign w15080 = ~w15067 & w15079 ;
  assign w15081 = w15078 | w15080 ;
  assign w15082 = ( w12245 & w15075 ) | ( w12245 & ~w15081 ) | ( w15075 & ~w15081 ) ;
  assign w15083 = w12245 & w15082 ;
  assign w15084 = w14592 | w14597 ;
  assign w15085 = w15032 & ~w15084 ;
  assign w15086 = w14595 ^ w15085 ;
  assign w15087 = ( ~w12245 & w15075 ) | ( ~w12245 & w15081 ) | ( w15075 & w15081 ) ;
  assign w15088 = ~w15075 & w15087 ;
  assign w15089 = w15086 | w15088 ;
  assign w15090 = ( w11807 & w15083 ) | ( w11807 & ~w15089 ) | ( w15083 & ~w15089 ) ;
  assign w15091 = w11807 & w15090 ;
  assign w15092 = w14600 | w14605 ;
  assign w15093 = w15032 & ~w15092 ;
  assign w15094 = w14603 ^ w15093 ;
  assign w15095 = ( ~w11807 & w15083 ) | ( ~w11807 & w15089 ) | ( w15083 & w15089 ) ;
  assign w15096 = ~w15083 & w15095 ;
  assign w15097 = w15094 | w15096 ;
  assign w15098 = ( w11377 & w15091 ) | ( w11377 & ~w15097 ) | ( w15091 & ~w15097 ) ;
  assign w15099 = w11377 & w15098 ;
  assign w15100 = w14608 | w14613 ;
  assign w15101 = w15032 & ~w15100 ;
  assign w15102 = w14611 ^ w15101 ;
  assign w15103 = ( ~w11377 & w15091 ) | ( ~w11377 & w15097 ) | ( w15091 & w15097 ) ;
  assign w15104 = ~w15091 & w15103 ;
  assign w15105 = w15102 | w15104 ;
  assign w15106 = ( w10955 & w15099 ) | ( w10955 & ~w15105 ) | ( w15099 & ~w15105 ) ;
  assign w15107 = w10955 & w15106 ;
  assign w15108 = w14616 | w14621 ;
  assign w15109 = w15032 & ~w15108 ;
  assign w15110 = w14619 ^ w15109 ;
  assign w15111 = ( ~w10955 & w15099 ) | ( ~w10955 & w15105 ) | ( w15099 & w15105 ) ;
  assign w15112 = ~w15099 & w15111 ;
  assign w15113 = w15110 | w15112 ;
  assign w15114 = ( w10541 & w15107 ) | ( w10541 & ~w15113 ) | ( w15107 & ~w15113 ) ;
  assign w15115 = w10541 & w15114 ;
  assign w15116 = w14624 | w14629 ;
  assign w15117 = w15032 & ~w15116 ;
  assign w15118 = w14627 ^ w15117 ;
  assign w15119 = ( ~w10541 & w15107 ) | ( ~w10541 & w15113 ) | ( w15107 & w15113 ) ;
  assign w15120 = ~w15107 & w15119 ;
  assign w15121 = w15118 | w15120 ;
  assign w15122 = ( w10135 & w15115 ) | ( w10135 & ~w15121 ) | ( w15115 & ~w15121 ) ;
  assign w15123 = w10135 & w15122 ;
  assign w15124 = w14632 | w14637 ;
  assign w15125 = w15032 & ~w15124 ;
  assign w15126 = w14635 ^ w15125 ;
  assign w15127 = ( ~w10135 & w15115 ) | ( ~w10135 & w15121 ) | ( w15115 & w15121 ) ;
  assign w15128 = ~w15115 & w15127 ;
  assign w15129 = w15126 | w15128 ;
  assign w15130 = ( w9737 & w15123 ) | ( w9737 & ~w15129 ) | ( w15123 & ~w15129 ) ;
  assign w15131 = w9737 & w15130 ;
  assign w15132 = w14640 | w14645 ;
  assign w15133 = w15032 & ~w15132 ;
  assign w15134 = w14643 ^ w15133 ;
  assign w15135 = ( ~w9737 & w15123 ) | ( ~w9737 & w15129 ) | ( w15123 & w15129 ) ;
  assign w15136 = ~w15123 & w15135 ;
  assign w15137 = w15134 | w15136 ;
  assign w15138 = ( w9347 & w15131 ) | ( w9347 & ~w15137 ) | ( w15131 & ~w15137 ) ;
  assign w15139 = w9347 & w15138 ;
  assign w15140 = w14648 | w14653 ;
  assign w15141 = w15032 & ~w15140 ;
  assign w15142 = w14651 ^ w15141 ;
  assign w15143 = ( ~w9347 & w15131 ) | ( ~w9347 & w15137 ) | ( w15131 & w15137 ) ;
  assign w15144 = ~w15131 & w15143 ;
  assign w15145 = w15142 | w15144 ;
  assign w15146 = ( w8965 & w15139 ) | ( w8965 & ~w15145 ) | ( w15139 & ~w15145 ) ;
  assign w15147 = w8965 & w15146 ;
  assign w15148 = w14656 | w14661 ;
  assign w15149 = w15032 & ~w15148 ;
  assign w15150 = w14659 ^ w15149 ;
  assign w15151 = ( ~w8965 & w15139 ) | ( ~w8965 & w15145 ) | ( w15139 & w15145 ) ;
  assign w15152 = ~w15139 & w15151 ;
  assign w15153 = w15150 | w15152 ;
  assign w15154 = ( w8591 & w15147 ) | ( w8591 & ~w15153 ) | ( w15147 & ~w15153 ) ;
  assign w15155 = w8591 & w15154 ;
  assign w15156 = w14664 | w14669 ;
  assign w15157 = w15032 & ~w15156 ;
  assign w15158 = w14667 ^ w15157 ;
  assign w15159 = ( ~w8591 & w15147 ) | ( ~w8591 & w15153 ) | ( w15147 & w15153 ) ;
  assign w15160 = ~w15147 & w15159 ;
  assign w15161 = w15158 | w15160 ;
  assign w15162 = ( w8225 & w15155 ) | ( w8225 & ~w15161 ) | ( w15155 & ~w15161 ) ;
  assign w15163 = w8225 & w15162 ;
  assign w15164 = w14672 | w14677 ;
  assign w15165 = w15032 & ~w15164 ;
  assign w15166 = w14675 ^ w15165 ;
  assign w15167 = ( ~w8225 & w15155 ) | ( ~w8225 & w15161 ) | ( w15155 & w15161 ) ;
  assign w15168 = ~w15155 & w15167 ;
  assign w15169 = w15166 | w15168 ;
  assign w15170 = ( w7867 & w15163 ) | ( w7867 & ~w15169 ) | ( w15163 & ~w15169 ) ;
  assign w15171 = w7867 & w15170 ;
  assign w15172 = w14680 | w14685 ;
  assign w15173 = w15032 & ~w15172 ;
  assign w15174 = w14683 ^ w15173 ;
  assign w15175 = ( ~w7867 & w15163 ) | ( ~w7867 & w15169 ) | ( w15163 & w15169 ) ;
  assign w15176 = ~w15163 & w15175 ;
  assign w15177 = w15174 | w15176 ;
  assign w15178 = ( w7517 & w15171 ) | ( w7517 & ~w15177 ) | ( w15171 & ~w15177 ) ;
  assign w15179 = w7517 & w15178 ;
  assign w15180 = w14688 | w14693 ;
  assign w15181 = w15032 & ~w15180 ;
  assign w15182 = w14691 ^ w15181 ;
  assign w15183 = ( ~w7517 & w15171 ) | ( ~w7517 & w15177 ) | ( w15171 & w15177 ) ;
  assign w15184 = ~w15171 & w15183 ;
  assign w15185 = w15182 | w15184 ;
  assign w15186 = ( w7175 & w15179 ) | ( w7175 & ~w15185 ) | ( w15179 & ~w15185 ) ;
  assign w15187 = w7175 & w15186 ;
  assign w15188 = w14696 | w14701 ;
  assign w15189 = w15032 & ~w15188 ;
  assign w15190 = w14699 ^ w15189 ;
  assign w15191 = ( ~w7175 & w15179 ) | ( ~w7175 & w15185 ) | ( w15179 & w15185 ) ;
  assign w15192 = ~w15179 & w15191 ;
  assign w15193 = w15190 | w15192 ;
  assign w15194 = ( w6841 & w15187 ) | ( w6841 & ~w15193 ) | ( w15187 & ~w15193 ) ;
  assign w15195 = w6841 & w15194 ;
  assign w15196 = w14704 | w14709 ;
  assign w15197 = w15032 & ~w15196 ;
  assign w15198 = w14707 ^ w15197 ;
  assign w15199 = ( ~w6841 & w15187 ) | ( ~w6841 & w15193 ) | ( w15187 & w15193 ) ;
  assign w15200 = ~w15187 & w15199 ;
  assign w15201 = w15198 | w15200 ;
  assign w15202 = ( w6515 & w15195 ) | ( w6515 & ~w15201 ) | ( w15195 & ~w15201 ) ;
  assign w15203 = w6515 & w15202 ;
  assign w15204 = w14712 | w14717 ;
  assign w15205 = w15032 & ~w15204 ;
  assign w15206 = w14715 ^ w15205 ;
  assign w15207 = ( ~w6515 & w15195 ) | ( ~w6515 & w15201 ) | ( w15195 & w15201 ) ;
  assign w15208 = ~w15195 & w15207 ;
  assign w15209 = w15206 | w15208 ;
  assign w15210 = ( w6197 & w15203 ) | ( w6197 & ~w15209 ) | ( w15203 & ~w15209 ) ;
  assign w15211 = w6197 & w15210 ;
  assign w15212 = w14720 | w14725 ;
  assign w15213 = w15032 & ~w15212 ;
  assign w15214 = w14723 ^ w15213 ;
  assign w15215 = ( ~w6197 & w15203 ) | ( ~w6197 & w15209 ) | ( w15203 & w15209 ) ;
  assign w15216 = ~w15203 & w15215 ;
  assign w15217 = w15214 | w15216 ;
  assign w15218 = ( w5887 & w15211 ) | ( w5887 & ~w15217 ) | ( w15211 & ~w15217 ) ;
  assign w15219 = w5887 & w15218 ;
  assign w15220 = w14728 | w14733 ;
  assign w15221 = w15032 & ~w15220 ;
  assign w15222 = w14731 ^ w15221 ;
  assign w15223 = ( ~w5887 & w15211 ) | ( ~w5887 & w15217 ) | ( w15211 & w15217 ) ;
  assign w15224 = ~w15211 & w15223 ;
  assign w15225 = w15222 | w15224 ;
  assign w15226 = ( w5585 & w15219 ) | ( w5585 & ~w15225 ) | ( w15219 & ~w15225 ) ;
  assign w15227 = w5585 & w15226 ;
  assign w15228 = w14736 | w14741 ;
  assign w15229 = w15032 & ~w15228 ;
  assign w15230 = w14739 ^ w15229 ;
  assign w15231 = ( ~w5585 & w15219 ) | ( ~w5585 & w15225 ) | ( w15219 & w15225 ) ;
  assign w15232 = ~w15219 & w15231 ;
  assign w15233 = w15230 | w15232 ;
  assign w15234 = ( w5291 & w15227 ) | ( w5291 & ~w15233 ) | ( w15227 & ~w15233 ) ;
  assign w15235 = w5291 & w15234 ;
  assign w15236 = w14744 | w14749 ;
  assign w15237 = w15032 & ~w15236 ;
  assign w15238 = w14747 ^ w15237 ;
  assign w15239 = ( ~w5291 & w15227 ) | ( ~w5291 & w15233 ) | ( w15227 & w15233 ) ;
  assign w15240 = ~w15227 & w15239 ;
  assign w15241 = w15238 | w15240 ;
  assign w15242 = ( w5005 & w15235 ) | ( w5005 & ~w15241 ) | ( w15235 & ~w15241 ) ;
  assign w15243 = w5005 & w15242 ;
  assign w15244 = w14752 | w14757 ;
  assign w15245 = w15032 & ~w15244 ;
  assign w15246 = w14755 ^ w15245 ;
  assign w15247 = ( ~w5005 & w15235 ) | ( ~w5005 & w15241 ) | ( w15235 & w15241 ) ;
  assign w15248 = ~w15235 & w15247 ;
  assign w15249 = w15246 | w15248 ;
  assign w15250 = ( w4727 & w15243 ) | ( w4727 & ~w15249 ) | ( w15243 & ~w15249 ) ;
  assign w15251 = w4727 & w15250 ;
  assign w15252 = w14760 | w14765 ;
  assign w15253 = w15032 & ~w15252 ;
  assign w15254 = w14763 ^ w15253 ;
  assign w15255 = ( ~w4727 & w15243 ) | ( ~w4727 & w15249 ) | ( w15243 & w15249 ) ;
  assign w15256 = ~w15243 & w15255 ;
  assign w15257 = w15254 | w15256 ;
  assign w15258 = ( w4457 & w15251 ) | ( w4457 & ~w15257 ) | ( w15251 & ~w15257 ) ;
  assign w15259 = w4457 & w15258 ;
  assign w15260 = w14768 | w14773 ;
  assign w15261 = w15032 & ~w15260 ;
  assign w15262 = w14771 ^ w15261 ;
  assign w15263 = ( ~w4457 & w15251 ) | ( ~w4457 & w15257 ) | ( w15251 & w15257 ) ;
  assign w15264 = ~w15251 & w15263 ;
  assign w15265 = w15262 | w15264 ;
  assign w15266 = ( w4195 & w15259 ) | ( w4195 & ~w15265 ) | ( w15259 & ~w15265 ) ;
  assign w15267 = w4195 & w15266 ;
  assign w15268 = w14776 | w14781 ;
  assign w15269 = w15032 & ~w15268 ;
  assign w15270 = w14779 ^ w15269 ;
  assign w15271 = ( ~w4195 & w15259 ) | ( ~w4195 & w15265 ) | ( w15259 & w15265 ) ;
  assign w15272 = ~w15259 & w15271 ;
  assign w15273 = w15270 | w15272 ;
  assign w15274 = ( w3941 & w15267 ) | ( w3941 & ~w15273 ) | ( w15267 & ~w15273 ) ;
  assign w15275 = w3941 & w15274 ;
  assign w15276 = w14784 | w14789 ;
  assign w15277 = w15032 & ~w15276 ;
  assign w15278 = w14787 ^ w15277 ;
  assign w15279 = ( ~w3941 & w15267 ) | ( ~w3941 & w15273 ) | ( w15267 & w15273 ) ;
  assign w15280 = ~w15267 & w15279 ;
  assign w15281 = w15278 | w15280 ;
  assign w15282 = ( w3695 & w15275 ) | ( w3695 & ~w15281 ) | ( w15275 & ~w15281 ) ;
  assign w15283 = w3695 & w15282 ;
  assign w15284 = w14792 | w14797 ;
  assign w15285 = w15032 & ~w15284 ;
  assign w15286 = w14795 ^ w15285 ;
  assign w15287 = ( ~w3695 & w15275 ) | ( ~w3695 & w15281 ) | ( w15275 & w15281 ) ;
  assign w15288 = ~w15275 & w15287 ;
  assign w15289 = w15286 | w15288 ;
  assign w15290 = ( w3457 & w15283 ) | ( w3457 & ~w15289 ) | ( w15283 & ~w15289 ) ;
  assign w15291 = w3457 & w15290 ;
  assign w15292 = w14800 | w14805 ;
  assign w15293 = w15032 & ~w15292 ;
  assign w15294 = w14803 ^ w15293 ;
  assign w15295 = ( ~w3457 & w15283 ) | ( ~w3457 & w15289 ) | ( w15283 & w15289 ) ;
  assign w15296 = ~w15283 & w15295 ;
  assign w15297 = w15294 | w15296 ;
  assign w15298 = ( w3227 & w15291 ) | ( w3227 & ~w15297 ) | ( w15291 & ~w15297 ) ;
  assign w15299 = w3227 & w15298 ;
  assign w15300 = w14808 | w14813 ;
  assign w15301 = w15032 & ~w15300 ;
  assign w15302 = w14811 ^ w15301 ;
  assign w15303 = ( ~w3227 & w15291 ) | ( ~w3227 & w15297 ) | ( w15291 & w15297 ) ;
  assign w15304 = ~w15291 & w15303 ;
  assign w15305 = w15302 | w15304 ;
  assign w15306 = ( w3005 & w15299 ) | ( w3005 & ~w15305 ) | ( w15299 & ~w15305 ) ;
  assign w15307 = w3005 & w15306 ;
  assign w15308 = w14816 | w14821 ;
  assign w15309 = w15032 & ~w15308 ;
  assign w15310 = w14819 ^ w15309 ;
  assign w15311 = ( ~w3005 & w15299 ) | ( ~w3005 & w15305 ) | ( w15299 & w15305 ) ;
  assign w15312 = ~w15299 & w15311 ;
  assign w15313 = w15310 | w15312 ;
  assign w15314 = ( w2791 & w15307 ) | ( w2791 & ~w15313 ) | ( w15307 & ~w15313 ) ;
  assign w15315 = w2791 & w15314 ;
  assign w15316 = w14824 | w14829 ;
  assign w15317 = w15032 & ~w15316 ;
  assign w15318 = w14827 ^ w15317 ;
  assign w15319 = ( ~w2791 & w15307 ) | ( ~w2791 & w15313 ) | ( w15307 & w15313 ) ;
  assign w15320 = ~w15307 & w15319 ;
  assign w15321 = w15318 | w15320 ;
  assign w15322 = ( w2585 & w15315 ) | ( w2585 & ~w15321 ) | ( w15315 & ~w15321 ) ;
  assign w15323 = w2585 & w15322 ;
  assign w15324 = w14832 | w14837 ;
  assign w15325 = w15032 & ~w15324 ;
  assign w15326 = w14835 ^ w15325 ;
  assign w15327 = ( ~w2585 & w15315 ) | ( ~w2585 & w15321 ) | ( w15315 & w15321 ) ;
  assign w15328 = ~w15315 & w15327 ;
  assign w15329 = w15326 | w15328 ;
  assign w15330 = ( w2387 & w15323 ) | ( w2387 & ~w15329 ) | ( w15323 & ~w15329 ) ;
  assign w15331 = w2387 & w15330 ;
  assign w15332 = w14840 | w14845 ;
  assign w15333 = w15032 & ~w15332 ;
  assign w15334 = w14843 ^ w15333 ;
  assign w15335 = ( ~w2387 & w15323 ) | ( ~w2387 & w15329 ) | ( w15323 & w15329 ) ;
  assign w15336 = ~w15323 & w15335 ;
  assign w15337 = w15334 | w15336 ;
  assign w15338 = ( w2197 & w15331 ) | ( w2197 & ~w15337 ) | ( w15331 & ~w15337 ) ;
  assign w15339 = w2197 & w15338 ;
  assign w15340 = w14848 | w14853 ;
  assign w15341 = w15032 & ~w15340 ;
  assign w15342 = w14851 ^ w15341 ;
  assign w15343 = ( ~w2197 & w15331 ) | ( ~w2197 & w15337 ) | ( w15331 & w15337 ) ;
  assign w15344 = ~w15331 & w15343 ;
  assign w15345 = w15342 | w15344 ;
  assign w15346 = ( w2015 & w15339 ) | ( w2015 & ~w15345 ) | ( w15339 & ~w15345 ) ;
  assign w15347 = w2015 & w15346 ;
  assign w15348 = w14856 | w14861 ;
  assign w15349 = w15032 & ~w15348 ;
  assign w15350 = w14859 ^ w15349 ;
  assign w15351 = ( ~w2015 & w15339 ) | ( ~w2015 & w15345 ) | ( w15339 & w15345 ) ;
  assign w15352 = ~w15339 & w15351 ;
  assign w15353 = w15350 | w15352 ;
  assign w15354 = ( w1841 & w15347 ) | ( w1841 & ~w15353 ) | ( w15347 & ~w15353 ) ;
  assign w15355 = w1841 & w15354 ;
  assign w15356 = w14864 | w14869 ;
  assign w15357 = w15032 & ~w15356 ;
  assign w15358 = w14867 ^ w15357 ;
  assign w15359 = ( ~w1841 & w15347 ) | ( ~w1841 & w15353 ) | ( w15347 & w15353 ) ;
  assign w15360 = ~w15347 & w15359 ;
  assign w15361 = w15358 | w15360 ;
  assign w15362 = ( w1675 & w15355 ) | ( w1675 & ~w15361 ) | ( w15355 & ~w15361 ) ;
  assign w15363 = w1675 & w15362 ;
  assign w15364 = w14872 | w14877 ;
  assign w15365 = w15032 & ~w15364 ;
  assign w15366 = w14875 ^ w15365 ;
  assign w15367 = ( ~w1675 & w15355 ) | ( ~w1675 & w15361 ) | ( w15355 & w15361 ) ;
  assign w15368 = ~w15355 & w15367 ;
  assign w15369 = w15366 | w15368 ;
  assign w15370 = ( w1517 & w15363 ) | ( w1517 & ~w15369 ) | ( w15363 & ~w15369 ) ;
  assign w15371 = w1517 & w15370 ;
  assign w15372 = w14880 | w14885 ;
  assign w15373 = w15032 & ~w15372 ;
  assign w15374 = w14883 ^ w15373 ;
  assign w15375 = ( ~w1517 & w15363 ) | ( ~w1517 & w15369 ) | ( w15363 & w15369 ) ;
  assign w15376 = ~w15363 & w15375 ;
  assign w15377 = w15374 | w15376 ;
  assign w15378 = ( w1367 & w15371 ) | ( w1367 & ~w15377 ) | ( w15371 & ~w15377 ) ;
  assign w15379 = w1367 & w15378 ;
  assign w15380 = w14888 | w14893 ;
  assign w15381 = w15032 & ~w15380 ;
  assign w15382 = w14891 ^ w15381 ;
  assign w15383 = ( ~w1367 & w15371 ) | ( ~w1367 & w15377 ) | ( w15371 & w15377 ) ;
  assign w15384 = ~w15371 & w15383 ;
  assign w15385 = w15382 | w15384 ;
  assign w15386 = ( w1225 & w15379 ) | ( w1225 & ~w15385 ) | ( w15379 & ~w15385 ) ;
  assign w15387 = w1225 & w15386 ;
  assign w15388 = w14896 | w14901 ;
  assign w15389 = w15032 & ~w15388 ;
  assign w15390 = w14899 ^ w15389 ;
  assign w15391 = ( ~w1225 & w15379 ) | ( ~w1225 & w15385 ) | ( w15379 & w15385 ) ;
  assign w15392 = ~w15379 & w15391 ;
  assign w15393 = w15390 | w15392 ;
  assign w15394 = ( w1091 & w15387 ) | ( w1091 & ~w15393 ) | ( w15387 & ~w15393 ) ;
  assign w15395 = w1091 & w15394 ;
  assign w15396 = w14904 | w14909 ;
  assign w15397 = w15032 & ~w15396 ;
  assign w15398 = w14907 ^ w15397 ;
  assign w15399 = ( ~w1091 & w15387 ) | ( ~w1091 & w15393 ) | ( w15387 & w15393 ) ;
  assign w15400 = ~w15387 & w15399 ;
  assign w15401 = w15398 | w15400 ;
  assign w15402 = ( w965 & w15395 ) | ( w965 & ~w15401 ) | ( w15395 & ~w15401 ) ;
  assign w15403 = w965 & w15402 ;
  assign w15404 = w14912 | w14917 ;
  assign w15405 = w15032 & ~w15404 ;
  assign w15406 = w14915 ^ w15405 ;
  assign w15407 = ( ~w965 & w15395 ) | ( ~w965 & w15401 ) | ( w15395 & w15401 ) ;
  assign w15408 = ~w15395 & w15407 ;
  assign w15409 = w15406 | w15408 ;
  assign w15410 = ( w847 & w15403 ) | ( w847 & ~w15409 ) | ( w15403 & ~w15409 ) ;
  assign w15411 = w847 & w15410 ;
  assign w15412 = w14920 | w14925 ;
  assign w15413 = w15032 & ~w15412 ;
  assign w15414 = w14923 ^ w15413 ;
  assign w15415 = ( ~w847 & w15403 ) | ( ~w847 & w15409 ) | ( w15403 & w15409 ) ;
  assign w15416 = ~w15403 & w15415 ;
  assign w15417 = w15414 | w15416 ;
  assign w15418 = ( w737 & w15411 ) | ( w737 & ~w15417 ) | ( w15411 & ~w15417 ) ;
  assign w15419 = w737 & w15418 ;
  assign w15420 = w14928 | w14933 ;
  assign w15421 = w15032 & ~w15420 ;
  assign w15422 = w14931 ^ w15421 ;
  assign w15423 = ( ~w737 & w15411 ) | ( ~w737 & w15417 ) | ( w15411 & w15417 ) ;
  assign w15424 = ~w15411 & w15423 ;
  assign w15425 = w15422 | w15424 ;
  assign w15426 = ( w635 & w15419 ) | ( w635 & ~w15425 ) | ( w15419 & ~w15425 ) ;
  assign w15427 = w635 & w15426 ;
  assign w15428 = w14936 | w14941 ;
  assign w15429 = w15032 & ~w15428 ;
  assign w15430 = w14939 ^ w15429 ;
  assign w15431 = ( ~w635 & w15419 ) | ( ~w635 & w15425 ) | ( w15419 & w15425 ) ;
  assign w15432 = ~w15419 & w15431 ;
  assign w15433 = w15430 | w15432 ;
  assign w15434 = ( w541 & w15427 ) | ( w541 & ~w15433 ) | ( w15427 & ~w15433 ) ;
  assign w15435 = w541 & w15434 ;
  assign w15436 = w14944 | w14949 ;
  assign w15437 = w15032 & ~w15436 ;
  assign w15438 = w14947 ^ w15437 ;
  assign w15439 = ( ~w541 & w15427 ) | ( ~w541 & w15433 ) | ( w15427 & w15433 ) ;
  assign w15440 = ~w15427 & w15439 ;
  assign w15441 = w15438 | w15440 ;
  assign w15442 = ( w455 & w15435 ) | ( w455 & ~w15441 ) | ( w15435 & ~w15441 ) ;
  assign w15443 = w455 & w15442 ;
  assign w15444 = w14952 | w14957 ;
  assign w15445 = w15032 & ~w15444 ;
  assign w15446 = w14955 ^ w15445 ;
  assign w15447 = ( ~w455 & w15435 ) | ( ~w455 & w15441 ) | ( w15435 & w15441 ) ;
  assign w15448 = ~w15435 & w15447 ;
  assign w15449 = w15446 | w15448 ;
  assign w15450 = ( w377 & w15443 ) | ( w377 & ~w15449 ) | ( w15443 & ~w15449 ) ;
  assign w15451 = w377 & w15450 ;
  assign w15452 = w14960 | w14965 ;
  assign w15453 = w15032 & ~w15452 ;
  assign w15454 = w14963 ^ w15453 ;
  assign w15455 = ( ~w377 & w15443 ) | ( ~w377 & w15449 ) | ( w15443 & w15449 ) ;
  assign w15456 = ~w15443 & w15455 ;
  assign w15457 = w15454 | w15456 ;
  assign w15458 = ( w307 & w15451 ) | ( w307 & ~w15457 ) | ( w15451 & ~w15457 ) ;
  assign w15459 = w307 & w15458 ;
  assign w15460 = w14968 | w14973 ;
  assign w15461 = w15032 & ~w15460 ;
  assign w15462 = w14971 ^ w15461 ;
  assign w15463 = ( ~w307 & w15451 ) | ( ~w307 & w15457 ) | ( w15451 & w15457 ) ;
  assign w15464 = ~w15451 & w15463 ;
  assign w15465 = w15462 | w15464 ;
  assign w15466 = ( w246 & w15459 ) | ( w246 & ~w15465 ) | ( w15459 & ~w15465 ) ;
  assign w15467 = w246 & w15466 ;
  assign w15468 = w14976 | w14981 ;
  assign w15469 = w15032 & ~w15468 ;
  assign w15470 = w14979 ^ w15469 ;
  assign w15471 = ( ~w246 & w15459 ) | ( ~w246 & w15465 ) | ( w15459 & w15465 ) ;
  assign w15472 = ~w15459 & w15471 ;
  assign w15473 = w15470 | w15472 ;
  assign w15474 = ( w185 & w15467 ) | ( w185 & ~w15473 ) | ( w15467 & ~w15473 ) ;
  assign w15475 = w185 & w15474 ;
  assign w15476 = ( ~w185 & w15467 ) | ( ~w185 & w15473 ) | ( w15467 & w15473 ) ;
  assign w15477 = ~w15467 & w15476 ;
  assign w15478 = w14984 | w14986 ;
  assign w15479 = w15032 & ~w15478 ;
  assign w15480 = w14989 ^ w15479 ;
  assign w15481 = w15477 | w15480 ;
  assign w15482 = ( w145 & w15475 ) | ( w145 & ~w15481 ) | ( w15475 & ~w15481 ) ;
  assign w15483 = w145 & w15482 ;
  assign w15484 = w14992 | w14997 ;
  assign w15485 = w15032 & ~w15484 ;
  assign w15486 = w14995 ^ w15485 ;
  assign w15487 = ( ~w145 & w15475 ) | ( ~w145 & w15481 ) | ( w15475 & w15481 ) ;
  assign w15488 = ~w15475 & w15487 ;
  assign w15489 = w15486 | w15488 ;
  assign w15490 = ( w132 & w15483 ) | ( w132 & ~w15489 ) | ( w15483 & ~w15489 ) ;
  assign w15491 = w132 & w15490 ;
  assign w15492 = w15000 | w15005 ;
  assign w15493 = w15032 & ~w15492 ;
  assign w15494 = w15003 ^ w15493 ;
  assign w15495 = ( ~w132 & w15483 ) | ( ~w132 & w15489 ) | ( w15483 & w15489 ) ;
  assign w15496 = ~w15483 & w15495 ;
  assign w15497 = w15494 | w15496 ;
  assign w15498 = ~w15491 & w15497 ;
  assign w15499 = w15008 | w15013 ;
  assign w15500 = w15032 & ~w15499 ;
  assign w15501 = w15011 ^ w15500 ;
  assign w15502 = ( ~w15026 & w15498 ) | ( ~w15026 & w15501 ) | ( w15498 & w15501 ) ;
  assign w15503 = w15015 & ~w15502 ;
  assign w15504 = ~w15018 & w15032 ;
  assign w15505 = ( w15502 & ~w15503 ) | ( w15502 & w15504 ) | ( ~w15503 & w15504 ) ;
  assign w15506 = w15026 | w15505 ;
  assign w15507 = ~w129 & w15506 ;
  assign w15508 = ( w15491 & w15497 ) | ( w15491 & w15501 ) | ( w15497 & w15501 ) ;
  assign w15509 = ~w15491 & w15508 ;
  assign w15510 = ( w129 & w15015 ) | ( w129 & w15018 ) | ( w15015 & w15018 ) ;
  assign w15511 = ( w15018 & ~w15032 ) | ( w15018 & w15510 ) | ( ~w15032 & w15510 ) ;
  assign w15512 = w15015 & w15511 ;
  assign w15513 = w15510 ^ w15512 ;
  assign w15514 = ( w15507 & ~w15509 ) | ( w15507 & w15513 ) | ( ~w15509 & w15513 ) ;
  assign w15515 = w15509 | w15514 ;
  assign w15516 = \pi006 | \pi007 ;
  assign w15517 = ( \pi008 & w15032 ) | ( \pi008 & ~w15516 ) | ( w15032 & ~w15516 ) ;
  assign w15518 = ( ~\pi008 & w15032 ) | ( ~\pi008 & w15515 ) | ( w15032 & w15515 ) ;
  assign w15519 = w15517 & w15518 ;
  assign w15520 = \pi008 & ~w15515 ;
  assign w15521 = ( ~\pi008 & w15024 ) | ( ~\pi008 & w15516 ) | ( w15024 & w15516 ) ;
  assign w15522 = ( ~w15024 & w15026 ) | ( ~w15024 & w15030 ) | ( w15026 & w15030 ) ;
  assign w15523 = ( w15520 & w15521 ) | ( w15520 & ~w15522 ) | ( w15521 & ~w15522 ) ;
  assign w15524 = ~w15024 & w15523 ;
  assign w15525 = ~\pi008 & w15515 ;
  assign w15526 = \pi009 ^ w15525 ;
  assign w15527 = w15524 | w15526 ;
  assign w15528 = ( w14555 & w15519 ) | ( w14555 & ~w15527 ) | ( w15519 & ~w15527 ) ;
  assign w15529 = w14555 & w15528 ;
  assign w15530 = ( ~w14555 & w15519 ) | ( ~w14555 & w15527 ) | ( w15519 & w15527 ) ;
  assign w15531 = ~w15519 & w15530 ;
  assign w15532 = w15507 | w15509 ;
  assign w15533 = w15513 | w15532 ;
  assign w15534 = w15032 ^ w15533 ;
  assign w15535 = ( w15032 & ~w15033 ) | ( w15032 & w15534 ) | ( ~w15033 & w15534 ) ;
  assign w15536 = \pi010 ^ w15535 ;
  assign w15537 = w15531 | w15536 ;
  assign w15538 = ( w14077 & w15529 ) | ( w14077 & ~w15537 ) | ( w15529 & ~w15537 ) ;
  assign w15539 = w14077 & w15538 ;
  assign w15540 = ( w15036 & ~w15043 ) | ( w15036 & w15515 ) | ( ~w15043 & w15515 ) ;
  assign w15541 = ~w15036 & w15540 ;
  assign w15542 = \pi011 ^ w15541 ;
  assign w15543 = w15044 ^ w15542 ;
  assign w15544 = ( ~w14077 & w15529 ) | ( ~w14077 & w15537 ) | ( w15529 & w15537 ) ;
  assign w15545 = ~w15529 & w15544 ;
  assign w15546 = w15543 | w15545 ;
  assign w15547 = ( w13607 & w15539 ) | ( w13607 & ~w15546 ) | ( w15539 & ~w15546 ) ;
  assign w15548 = w13607 & w15547 ;
  assign w15549 = w15048 | w15050 ;
  assign w15550 = w15515 & ~w15549 ;
  assign w15551 = w15055 ^ w15550 ;
  assign w15552 = ( ~w13607 & w15539 ) | ( ~w13607 & w15546 ) | ( w15539 & w15546 ) ;
  assign w15553 = ~w15539 & w15552 ;
  assign w15554 = w15551 | w15553 ;
  assign w15555 = ( w13145 & w15548 ) | ( w13145 & ~w15554 ) | ( w15548 & ~w15554 ) ;
  assign w15556 = w13145 & w15555 ;
  assign w15557 = w15058 | w15064 ;
  assign w15558 = w15515 & ~w15557 ;
  assign w15559 = w15062 ^ w15558 ;
  assign w15560 = ( ~w13145 & w15548 ) | ( ~w13145 & w15554 ) | ( w15548 & w15554 ) ;
  assign w15561 = ~w15548 & w15560 ;
  assign w15562 = w15559 | w15561 ;
  assign w15563 = ( w12691 & w15556 ) | ( w12691 & ~w15562 ) | ( w15556 & ~w15562 ) ;
  assign w15564 = w12691 & w15563 ;
  assign w15565 = w15067 | w15072 ;
  assign w15566 = w15515 & ~w15565 ;
  assign w15567 = w15070 ^ w15566 ;
  assign w15568 = ( ~w12691 & w15556 ) | ( ~w12691 & w15562 ) | ( w15556 & w15562 ) ;
  assign w15569 = ~w15556 & w15568 ;
  assign w15570 = w15567 | w15569 ;
  assign w15571 = ( w12245 & w15564 ) | ( w12245 & ~w15570 ) | ( w15564 & ~w15570 ) ;
  assign w15572 = w12245 & w15571 ;
  assign w15573 = w15075 | w15080 ;
  assign w15574 = w15515 & ~w15573 ;
  assign w15575 = w15078 ^ w15574 ;
  assign w15576 = ( ~w12245 & w15564 ) | ( ~w12245 & w15570 ) | ( w15564 & w15570 ) ;
  assign w15577 = ~w15564 & w15576 ;
  assign w15578 = w15575 | w15577 ;
  assign w15579 = ( w11807 & w15572 ) | ( w11807 & ~w15578 ) | ( w15572 & ~w15578 ) ;
  assign w15580 = w11807 & w15579 ;
  assign w15581 = w15083 | w15088 ;
  assign w15582 = w15515 & ~w15581 ;
  assign w15583 = w15086 ^ w15582 ;
  assign w15584 = ( ~w11807 & w15572 ) | ( ~w11807 & w15578 ) | ( w15572 & w15578 ) ;
  assign w15585 = ~w15572 & w15584 ;
  assign w15586 = w15583 | w15585 ;
  assign w15587 = ( w11377 & w15580 ) | ( w11377 & ~w15586 ) | ( w15580 & ~w15586 ) ;
  assign w15588 = w11377 & w15587 ;
  assign w15589 = w15091 | w15096 ;
  assign w15590 = w15515 & ~w15589 ;
  assign w15591 = w15094 ^ w15590 ;
  assign w15592 = ( ~w11377 & w15580 ) | ( ~w11377 & w15586 ) | ( w15580 & w15586 ) ;
  assign w15593 = ~w15580 & w15592 ;
  assign w15594 = w15591 | w15593 ;
  assign w15595 = ( w10955 & w15588 ) | ( w10955 & ~w15594 ) | ( w15588 & ~w15594 ) ;
  assign w15596 = w10955 & w15595 ;
  assign w15597 = w15099 | w15104 ;
  assign w15598 = w15515 & ~w15597 ;
  assign w15599 = w15102 ^ w15598 ;
  assign w15600 = ( ~w10955 & w15588 ) | ( ~w10955 & w15594 ) | ( w15588 & w15594 ) ;
  assign w15601 = ~w15588 & w15600 ;
  assign w15602 = w15599 | w15601 ;
  assign w15603 = ( w10541 & w15596 ) | ( w10541 & ~w15602 ) | ( w15596 & ~w15602 ) ;
  assign w15604 = w10541 & w15603 ;
  assign w15605 = w15107 | w15112 ;
  assign w15606 = w15515 & ~w15605 ;
  assign w15607 = w15110 ^ w15606 ;
  assign w15608 = ( ~w10541 & w15596 ) | ( ~w10541 & w15602 ) | ( w15596 & w15602 ) ;
  assign w15609 = ~w15596 & w15608 ;
  assign w15610 = w15607 | w15609 ;
  assign w15611 = ( w10135 & w15604 ) | ( w10135 & ~w15610 ) | ( w15604 & ~w15610 ) ;
  assign w15612 = w10135 & w15611 ;
  assign w15613 = w15115 | w15120 ;
  assign w15614 = w15515 & ~w15613 ;
  assign w15615 = w15118 ^ w15614 ;
  assign w15616 = ( ~w10135 & w15604 ) | ( ~w10135 & w15610 ) | ( w15604 & w15610 ) ;
  assign w15617 = ~w15604 & w15616 ;
  assign w15618 = w15615 | w15617 ;
  assign w15619 = ( w9737 & w15612 ) | ( w9737 & ~w15618 ) | ( w15612 & ~w15618 ) ;
  assign w15620 = w9737 & w15619 ;
  assign w15621 = w15123 | w15128 ;
  assign w15622 = w15515 & ~w15621 ;
  assign w15623 = w15126 ^ w15622 ;
  assign w15624 = ( ~w9737 & w15612 ) | ( ~w9737 & w15618 ) | ( w15612 & w15618 ) ;
  assign w15625 = ~w15612 & w15624 ;
  assign w15626 = w15623 | w15625 ;
  assign w15627 = ( w9347 & w15620 ) | ( w9347 & ~w15626 ) | ( w15620 & ~w15626 ) ;
  assign w15628 = w9347 & w15627 ;
  assign w15629 = w15131 | w15136 ;
  assign w15630 = w15515 & ~w15629 ;
  assign w15631 = w15134 ^ w15630 ;
  assign w15632 = ( ~w9347 & w15620 ) | ( ~w9347 & w15626 ) | ( w15620 & w15626 ) ;
  assign w15633 = ~w15620 & w15632 ;
  assign w15634 = w15631 | w15633 ;
  assign w15635 = ( w8965 & w15628 ) | ( w8965 & ~w15634 ) | ( w15628 & ~w15634 ) ;
  assign w15636 = w8965 & w15635 ;
  assign w15637 = w15139 | w15144 ;
  assign w15638 = w15515 & ~w15637 ;
  assign w15639 = w15142 ^ w15638 ;
  assign w15640 = ( ~w8965 & w15628 ) | ( ~w8965 & w15634 ) | ( w15628 & w15634 ) ;
  assign w15641 = ~w15628 & w15640 ;
  assign w15642 = w15639 | w15641 ;
  assign w15643 = ( w8591 & w15636 ) | ( w8591 & ~w15642 ) | ( w15636 & ~w15642 ) ;
  assign w15644 = w8591 & w15643 ;
  assign w15645 = w15147 | w15152 ;
  assign w15646 = w15515 & ~w15645 ;
  assign w15647 = w15150 ^ w15646 ;
  assign w15648 = ( ~w8591 & w15636 ) | ( ~w8591 & w15642 ) | ( w15636 & w15642 ) ;
  assign w15649 = ~w15636 & w15648 ;
  assign w15650 = w15647 | w15649 ;
  assign w15651 = ( w8225 & w15644 ) | ( w8225 & ~w15650 ) | ( w15644 & ~w15650 ) ;
  assign w15652 = w8225 & w15651 ;
  assign w15653 = w15155 | w15160 ;
  assign w15654 = w15515 & ~w15653 ;
  assign w15655 = w15158 ^ w15654 ;
  assign w15656 = ( ~w8225 & w15644 ) | ( ~w8225 & w15650 ) | ( w15644 & w15650 ) ;
  assign w15657 = ~w15644 & w15656 ;
  assign w15658 = w15655 | w15657 ;
  assign w15659 = ( w7867 & w15652 ) | ( w7867 & ~w15658 ) | ( w15652 & ~w15658 ) ;
  assign w15660 = w7867 & w15659 ;
  assign w15661 = w15163 | w15168 ;
  assign w15662 = w15515 & ~w15661 ;
  assign w15663 = w15166 ^ w15662 ;
  assign w15664 = ( ~w7867 & w15652 ) | ( ~w7867 & w15658 ) | ( w15652 & w15658 ) ;
  assign w15665 = ~w15652 & w15664 ;
  assign w15666 = w15663 | w15665 ;
  assign w15667 = ( w7517 & w15660 ) | ( w7517 & ~w15666 ) | ( w15660 & ~w15666 ) ;
  assign w15668 = w7517 & w15667 ;
  assign w15669 = w15171 | w15176 ;
  assign w15670 = w15515 & ~w15669 ;
  assign w15671 = w15174 ^ w15670 ;
  assign w15672 = ( ~w7517 & w15660 ) | ( ~w7517 & w15666 ) | ( w15660 & w15666 ) ;
  assign w15673 = ~w15660 & w15672 ;
  assign w15674 = w15671 | w15673 ;
  assign w15675 = ( w7175 & w15668 ) | ( w7175 & ~w15674 ) | ( w15668 & ~w15674 ) ;
  assign w15676 = w7175 & w15675 ;
  assign w15677 = w15179 | w15184 ;
  assign w15678 = w15515 & ~w15677 ;
  assign w15679 = w15182 ^ w15678 ;
  assign w15680 = ( ~w7175 & w15668 ) | ( ~w7175 & w15674 ) | ( w15668 & w15674 ) ;
  assign w15681 = ~w15668 & w15680 ;
  assign w15682 = w15679 | w15681 ;
  assign w15683 = ( w6841 & w15676 ) | ( w6841 & ~w15682 ) | ( w15676 & ~w15682 ) ;
  assign w15684 = w6841 & w15683 ;
  assign w15685 = w15187 | w15192 ;
  assign w15686 = w15515 & ~w15685 ;
  assign w15687 = w15190 ^ w15686 ;
  assign w15688 = ( ~w6841 & w15676 ) | ( ~w6841 & w15682 ) | ( w15676 & w15682 ) ;
  assign w15689 = ~w15676 & w15688 ;
  assign w15690 = w15687 | w15689 ;
  assign w15691 = ( w6515 & w15684 ) | ( w6515 & ~w15690 ) | ( w15684 & ~w15690 ) ;
  assign w15692 = w6515 & w15691 ;
  assign w15693 = w15195 | w15200 ;
  assign w15694 = w15515 & ~w15693 ;
  assign w15695 = w15198 ^ w15694 ;
  assign w15696 = ( ~w6515 & w15684 ) | ( ~w6515 & w15690 ) | ( w15684 & w15690 ) ;
  assign w15697 = ~w15684 & w15696 ;
  assign w15698 = w15695 | w15697 ;
  assign w15699 = ( w6197 & w15692 ) | ( w6197 & ~w15698 ) | ( w15692 & ~w15698 ) ;
  assign w15700 = w6197 & w15699 ;
  assign w15701 = w15203 | w15208 ;
  assign w15702 = w15515 & ~w15701 ;
  assign w15703 = w15206 ^ w15702 ;
  assign w15704 = ( ~w6197 & w15692 ) | ( ~w6197 & w15698 ) | ( w15692 & w15698 ) ;
  assign w15705 = ~w15692 & w15704 ;
  assign w15706 = w15703 | w15705 ;
  assign w15707 = ( w5887 & w15700 ) | ( w5887 & ~w15706 ) | ( w15700 & ~w15706 ) ;
  assign w15708 = w5887 & w15707 ;
  assign w15709 = w15211 | w15216 ;
  assign w15710 = w15515 & ~w15709 ;
  assign w15711 = w15214 ^ w15710 ;
  assign w15712 = ( ~w5887 & w15700 ) | ( ~w5887 & w15706 ) | ( w15700 & w15706 ) ;
  assign w15713 = ~w15700 & w15712 ;
  assign w15714 = w15711 | w15713 ;
  assign w15715 = ( w5585 & w15708 ) | ( w5585 & ~w15714 ) | ( w15708 & ~w15714 ) ;
  assign w15716 = w5585 & w15715 ;
  assign w15717 = w15219 | w15224 ;
  assign w15718 = w15515 & ~w15717 ;
  assign w15719 = w15222 ^ w15718 ;
  assign w15720 = ( ~w5585 & w15708 ) | ( ~w5585 & w15714 ) | ( w15708 & w15714 ) ;
  assign w15721 = ~w15708 & w15720 ;
  assign w15722 = w15719 | w15721 ;
  assign w15723 = ( w5291 & w15716 ) | ( w5291 & ~w15722 ) | ( w15716 & ~w15722 ) ;
  assign w15724 = w5291 & w15723 ;
  assign w15725 = w15227 | w15232 ;
  assign w15726 = w15515 & ~w15725 ;
  assign w15727 = w15230 ^ w15726 ;
  assign w15728 = ( ~w5291 & w15716 ) | ( ~w5291 & w15722 ) | ( w15716 & w15722 ) ;
  assign w15729 = ~w15716 & w15728 ;
  assign w15730 = w15727 | w15729 ;
  assign w15731 = ( w5005 & w15724 ) | ( w5005 & ~w15730 ) | ( w15724 & ~w15730 ) ;
  assign w15732 = w5005 & w15731 ;
  assign w15733 = w15235 | w15240 ;
  assign w15734 = w15515 & ~w15733 ;
  assign w15735 = w15238 ^ w15734 ;
  assign w15736 = ( ~w5005 & w15724 ) | ( ~w5005 & w15730 ) | ( w15724 & w15730 ) ;
  assign w15737 = ~w15724 & w15736 ;
  assign w15738 = w15735 | w15737 ;
  assign w15739 = ( w4727 & w15732 ) | ( w4727 & ~w15738 ) | ( w15732 & ~w15738 ) ;
  assign w15740 = w4727 & w15739 ;
  assign w15741 = w15243 | w15248 ;
  assign w15742 = w15515 & ~w15741 ;
  assign w15743 = w15246 ^ w15742 ;
  assign w15744 = ( ~w4727 & w15732 ) | ( ~w4727 & w15738 ) | ( w15732 & w15738 ) ;
  assign w15745 = ~w15732 & w15744 ;
  assign w15746 = w15743 | w15745 ;
  assign w15747 = ( w4457 & w15740 ) | ( w4457 & ~w15746 ) | ( w15740 & ~w15746 ) ;
  assign w15748 = w4457 & w15747 ;
  assign w15749 = w15251 | w15256 ;
  assign w15750 = w15515 & ~w15749 ;
  assign w15751 = w15254 ^ w15750 ;
  assign w15752 = ( ~w4457 & w15740 ) | ( ~w4457 & w15746 ) | ( w15740 & w15746 ) ;
  assign w15753 = ~w15740 & w15752 ;
  assign w15754 = w15751 | w15753 ;
  assign w15755 = ( w4195 & w15748 ) | ( w4195 & ~w15754 ) | ( w15748 & ~w15754 ) ;
  assign w15756 = w4195 & w15755 ;
  assign w15757 = w15259 | w15264 ;
  assign w15758 = w15515 & ~w15757 ;
  assign w15759 = w15262 ^ w15758 ;
  assign w15760 = ( ~w4195 & w15748 ) | ( ~w4195 & w15754 ) | ( w15748 & w15754 ) ;
  assign w15761 = ~w15748 & w15760 ;
  assign w15762 = w15759 | w15761 ;
  assign w15763 = ( w3941 & w15756 ) | ( w3941 & ~w15762 ) | ( w15756 & ~w15762 ) ;
  assign w15764 = w3941 & w15763 ;
  assign w15765 = w15267 | w15272 ;
  assign w15766 = w15515 & ~w15765 ;
  assign w15767 = w15270 ^ w15766 ;
  assign w15768 = ( ~w3941 & w15756 ) | ( ~w3941 & w15762 ) | ( w15756 & w15762 ) ;
  assign w15769 = ~w15756 & w15768 ;
  assign w15770 = w15767 | w15769 ;
  assign w15771 = ( w3695 & w15764 ) | ( w3695 & ~w15770 ) | ( w15764 & ~w15770 ) ;
  assign w15772 = w3695 & w15771 ;
  assign w15773 = w15275 | w15280 ;
  assign w15774 = w15515 & ~w15773 ;
  assign w15775 = w15278 ^ w15774 ;
  assign w15776 = ( ~w3695 & w15764 ) | ( ~w3695 & w15770 ) | ( w15764 & w15770 ) ;
  assign w15777 = ~w15764 & w15776 ;
  assign w15778 = w15775 | w15777 ;
  assign w15779 = ( w3457 & w15772 ) | ( w3457 & ~w15778 ) | ( w15772 & ~w15778 ) ;
  assign w15780 = w3457 & w15779 ;
  assign w15781 = w15283 | w15288 ;
  assign w15782 = w15515 & ~w15781 ;
  assign w15783 = w15286 ^ w15782 ;
  assign w15784 = ( ~w3457 & w15772 ) | ( ~w3457 & w15778 ) | ( w15772 & w15778 ) ;
  assign w15785 = ~w15772 & w15784 ;
  assign w15786 = w15783 | w15785 ;
  assign w15787 = ( w3227 & w15780 ) | ( w3227 & ~w15786 ) | ( w15780 & ~w15786 ) ;
  assign w15788 = w3227 & w15787 ;
  assign w15789 = w15291 | w15296 ;
  assign w15790 = w15515 & ~w15789 ;
  assign w15791 = w15294 ^ w15790 ;
  assign w15792 = ( ~w3227 & w15780 ) | ( ~w3227 & w15786 ) | ( w15780 & w15786 ) ;
  assign w15793 = ~w15780 & w15792 ;
  assign w15794 = w15791 | w15793 ;
  assign w15795 = ( w3005 & w15788 ) | ( w3005 & ~w15794 ) | ( w15788 & ~w15794 ) ;
  assign w15796 = w3005 & w15795 ;
  assign w15797 = w15299 | w15304 ;
  assign w15798 = w15515 & ~w15797 ;
  assign w15799 = w15302 ^ w15798 ;
  assign w15800 = ( ~w3005 & w15788 ) | ( ~w3005 & w15794 ) | ( w15788 & w15794 ) ;
  assign w15801 = ~w15788 & w15800 ;
  assign w15802 = w15799 | w15801 ;
  assign w15803 = ( w2791 & w15796 ) | ( w2791 & ~w15802 ) | ( w15796 & ~w15802 ) ;
  assign w15804 = w2791 & w15803 ;
  assign w15805 = w15307 | w15312 ;
  assign w15806 = w15515 & ~w15805 ;
  assign w15807 = w15310 ^ w15806 ;
  assign w15808 = ( ~w2791 & w15796 ) | ( ~w2791 & w15802 ) | ( w15796 & w15802 ) ;
  assign w15809 = ~w15796 & w15808 ;
  assign w15810 = w15807 | w15809 ;
  assign w15811 = ( w2585 & w15804 ) | ( w2585 & ~w15810 ) | ( w15804 & ~w15810 ) ;
  assign w15812 = w2585 & w15811 ;
  assign w15813 = w15315 | w15320 ;
  assign w15814 = w15515 & ~w15813 ;
  assign w15815 = w15318 ^ w15814 ;
  assign w15816 = ( ~w2585 & w15804 ) | ( ~w2585 & w15810 ) | ( w15804 & w15810 ) ;
  assign w15817 = ~w15804 & w15816 ;
  assign w15818 = w15815 | w15817 ;
  assign w15819 = ( w2387 & w15812 ) | ( w2387 & ~w15818 ) | ( w15812 & ~w15818 ) ;
  assign w15820 = w2387 & w15819 ;
  assign w15821 = w15323 | w15328 ;
  assign w15822 = w15515 & ~w15821 ;
  assign w15823 = w15326 ^ w15822 ;
  assign w15824 = ( ~w2387 & w15812 ) | ( ~w2387 & w15818 ) | ( w15812 & w15818 ) ;
  assign w15825 = ~w15812 & w15824 ;
  assign w15826 = w15823 | w15825 ;
  assign w15827 = ( w2197 & w15820 ) | ( w2197 & ~w15826 ) | ( w15820 & ~w15826 ) ;
  assign w15828 = w2197 & w15827 ;
  assign w15829 = w15331 | w15336 ;
  assign w15830 = w15515 & ~w15829 ;
  assign w15831 = w15334 ^ w15830 ;
  assign w15832 = ( ~w2197 & w15820 ) | ( ~w2197 & w15826 ) | ( w15820 & w15826 ) ;
  assign w15833 = ~w15820 & w15832 ;
  assign w15834 = w15831 | w15833 ;
  assign w15835 = ( w2015 & w15828 ) | ( w2015 & ~w15834 ) | ( w15828 & ~w15834 ) ;
  assign w15836 = w2015 & w15835 ;
  assign w15837 = w15339 | w15344 ;
  assign w15838 = w15515 & ~w15837 ;
  assign w15839 = w15342 ^ w15838 ;
  assign w15840 = ( ~w2015 & w15828 ) | ( ~w2015 & w15834 ) | ( w15828 & w15834 ) ;
  assign w15841 = ~w15828 & w15840 ;
  assign w15842 = w15839 | w15841 ;
  assign w15843 = ( w1841 & w15836 ) | ( w1841 & ~w15842 ) | ( w15836 & ~w15842 ) ;
  assign w15844 = w1841 & w15843 ;
  assign w15845 = w15347 | w15352 ;
  assign w15846 = w15515 & ~w15845 ;
  assign w15847 = w15350 ^ w15846 ;
  assign w15848 = ( ~w1841 & w15836 ) | ( ~w1841 & w15842 ) | ( w15836 & w15842 ) ;
  assign w15849 = ~w15836 & w15848 ;
  assign w15850 = w15847 | w15849 ;
  assign w15851 = ( w1675 & w15844 ) | ( w1675 & ~w15850 ) | ( w15844 & ~w15850 ) ;
  assign w15852 = w1675 & w15851 ;
  assign w15853 = w15355 | w15360 ;
  assign w15854 = w15515 & ~w15853 ;
  assign w15855 = w15358 ^ w15854 ;
  assign w15856 = ( ~w1675 & w15844 ) | ( ~w1675 & w15850 ) | ( w15844 & w15850 ) ;
  assign w15857 = ~w15844 & w15856 ;
  assign w15858 = w15855 | w15857 ;
  assign w15859 = ( w1517 & w15852 ) | ( w1517 & ~w15858 ) | ( w15852 & ~w15858 ) ;
  assign w15860 = w1517 & w15859 ;
  assign w15861 = w15363 | w15368 ;
  assign w15862 = w15515 & ~w15861 ;
  assign w15863 = w15366 ^ w15862 ;
  assign w15864 = ( ~w1517 & w15852 ) | ( ~w1517 & w15858 ) | ( w15852 & w15858 ) ;
  assign w15865 = ~w15852 & w15864 ;
  assign w15866 = w15863 | w15865 ;
  assign w15867 = ( w1367 & w15860 ) | ( w1367 & ~w15866 ) | ( w15860 & ~w15866 ) ;
  assign w15868 = w1367 & w15867 ;
  assign w15869 = w15371 | w15376 ;
  assign w15870 = w15515 & ~w15869 ;
  assign w15871 = w15374 ^ w15870 ;
  assign w15872 = ( ~w1367 & w15860 ) | ( ~w1367 & w15866 ) | ( w15860 & w15866 ) ;
  assign w15873 = ~w15860 & w15872 ;
  assign w15874 = w15871 | w15873 ;
  assign w15875 = ( w1225 & w15868 ) | ( w1225 & ~w15874 ) | ( w15868 & ~w15874 ) ;
  assign w15876 = w1225 & w15875 ;
  assign w15877 = w15379 | w15384 ;
  assign w15878 = w15515 & ~w15877 ;
  assign w15879 = w15382 ^ w15878 ;
  assign w15880 = ( ~w1225 & w15868 ) | ( ~w1225 & w15874 ) | ( w15868 & w15874 ) ;
  assign w15881 = ~w15868 & w15880 ;
  assign w15882 = w15879 | w15881 ;
  assign w15883 = ( w1091 & w15876 ) | ( w1091 & ~w15882 ) | ( w15876 & ~w15882 ) ;
  assign w15884 = w1091 & w15883 ;
  assign w15885 = w15387 | w15392 ;
  assign w15886 = w15515 & ~w15885 ;
  assign w15887 = w15390 ^ w15886 ;
  assign w15888 = ( ~w1091 & w15876 ) | ( ~w1091 & w15882 ) | ( w15876 & w15882 ) ;
  assign w15889 = ~w15876 & w15888 ;
  assign w15890 = w15887 | w15889 ;
  assign w15891 = ( w965 & w15884 ) | ( w965 & ~w15890 ) | ( w15884 & ~w15890 ) ;
  assign w15892 = w965 & w15891 ;
  assign w15893 = w15395 | w15400 ;
  assign w15894 = w15515 & ~w15893 ;
  assign w15895 = w15398 ^ w15894 ;
  assign w15896 = ( ~w965 & w15884 ) | ( ~w965 & w15890 ) | ( w15884 & w15890 ) ;
  assign w15897 = ~w15884 & w15896 ;
  assign w15898 = w15895 | w15897 ;
  assign w15899 = ( w847 & w15892 ) | ( w847 & ~w15898 ) | ( w15892 & ~w15898 ) ;
  assign w15900 = w847 & w15899 ;
  assign w15901 = w15403 | w15408 ;
  assign w15902 = w15515 & ~w15901 ;
  assign w15903 = w15406 ^ w15902 ;
  assign w15904 = ( ~w847 & w15892 ) | ( ~w847 & w15898 ) | ( w15892 & w15898 ) ;
  assign w15905 = ~w15892 & w15904 ;
  assign w15906 = w15903 | w15905 ;
  assign w15907 = ( w737 & w15900 ) | ( w737 & ~w15906 ) | ( w15900 & ~w15906 ) ;
  assign w15908 = w737 & w15907 ;
  assign w15909 = w15411 | w15416 ;
  assign w15910 = w15515 & ~w15909 ;
  assign w15911 = w15414 ^ w15910 ;
  assign w15912 = ( ~w737 & w15900 ) | ( ~w737 & w15906 ) | ( w15900 & w15906 ) ;
  assign w15913 = ~w15900 & w15912 ;
  assign w15914 = w15911 | w15913 ;
  assign w15915 = ( w635 & w15908 ) | ( w635 & ~w15914 ) | ( w15908 & ~w15914 ) ;
  assign w15916 = w635 & w15915 ;
  assign w15917 = w15419 | w15424 ;
  assign w15918 = w15515 & ~w15917 ;
  assign w15919 = w15422 ^ w15918 ;
  assign w15920 = ( ~w635 & w15908 ) | ( ~w635 & w15914 ) | ( w15908 & w15914 ) ;
  assign w15921 = ~w15908 & w15920 ;
  assign w15922 = w15919 | w15921 ;
  assign w15923 = ( w541 & w15916 ) | ( w541 & ~w15922 ) | ( w15916 & ~w15922 ) ;
  assign w15924 = w541 & w15923 ;
  assign w15925 = w15427 | w15432 ;
  assign w15926 = w15515 & ~w15925 ;
  assign w15927 = w15430 ^ w15926 ;
  assign w15928 = ( ~w541 & w15916 ) | ( ~w541 & w15922 ) | ( w15916 & w15922 ) ;
  assign w15929 = ~w15916 & w15928 ;
  assign w15930 = w15927 | w15929 ;
  assign w15931 = ( w455 & w15924 ) | ( w455 & ~w15930 ) | ( w15924 & ~w15930 ) ;
  assign w15932 = w455 & w15931 ;
  assign w15933 = w15435 | w15440 ;
  assign w15934 = w15515 & ~w15933 ;
  assign w15935 = w15438 ^ w15934 ;
  assign w15936 = ( ~w455 & w15924 ) | ( ~w455 & w15930 ) | ( w15924 & w15930 ) ;
  assign w15937 = ~w15924 & w15936 ;
  assign w15938 = w15935 | w15937 ;
  assign w15939 = ( w377 & w15932 ) | ( w377 & ~w15938 ) | ( w15932 & ~w15938 ) ;
  assign w15940 = w377 & w15939 ;
  assign w15941 = w15443 | w15448 ;
  assign w15942 = w15515 & ~w15941 ;
  assign w15943 = w15446 ^ w15942 ;
  assign w15944 = ( ~w377 & w15932 ) | ( ~w377 & w15938 ) | ( w15932 & w15938 ) ;
  assign w15945 = ~w15932 & w15944 ;
  assign w15946 = w15943 | w15945 ;
  assign w15947 = ( w307 & w15940 ) | ( w307 & ~w15946 ) | ( w15940 & ~w15946 ) ;
  assign w15948 = w307 & w15947 ;
  assign w15949 = w15451 | w15456 ;
  assign w15950 = w15515 & ~w15949 ;
  assign w15951 = w15454 ^ w15950 ;
  assign w15952 = ( ~w307 & w15940 ) | ( ~w307 & w15946 ) | ( w15940 & w15946 ) ;
  assign w15953 = ~w15940 & w15952 ;
  assign w15954 = w15951 | w15953 ;
  assign w15955 = ( w246 & w15948 ) | ( w246 & ~w15954 ) | ( w15948 & ~w15954 ) ;
  assign w15956 = w246 & w15955 ;
  assign w15957 = w15459 | w15464 ;
  assign w15958 = w15515 & ~w15957 ;
  assign w15959 = w15462 ^ w15958 ;
  assign w15960 = ( ~w246 & w15948 ) | ( ~w246 & w15954 ) | ( w15948 & w15954 ) ;
  assign w15961 = ~w15948 & w15960 ;
  assign w15962 = w15959 | w15961 ;
  assign w15963 = ( w185 & w15956 ) | ( w185 & ~w15962 ) | ( w15956 & ~w15962 ) ;
  assign w15964 = w185 & w15963 ;
  assign w15965 = w15467 | w15472 ;
  assign w15966 = w15515 & ~w15965 ;
  assign w15967 = w15470 ^ w15966 ;
  assign w15968 = ( ~w185 & w15956 ) | ( ~w185 & w15962 ) | ( w15956 & w15962 ) ;
  assign w15969 = ~w15956 & w15968 ;
  assign w15970 = w15967 | w15969 ;
  assign w15971 = ( w145 & w15964 ) | ( w145 & ~w15970 ) | ( w15964 & ~w15970 ) ;
  assign w15972 = w145 & w15971 ;
  assign w15973 = ( ~w145 & w15964 ) | ( ~w145 & w15970 ) | ( w15964 & w15970 ) ;
  assign w15974 = ~w15964 & w15973 ;
  assign w15975 = w15475 | w15477 ;
  assign w15976 = w15515 & ~w15975 ;
  assign w15977 = w15480 ^ w15976 ;
  assign w15978 = w15974 | w15977 ;
  assign w15979 = ( w132 & w15972 ) | ( w132 & ~w15978 ) | ( w15972 & ~w15978 ) ;
  assign w15980 = w132 & w15979 ;
  assign w15981 = w15483 | w15488 ;
  assign w15982 = w15515 & ~w15981 ;
  assign w15983 = w15486 ^ w15982 ;
  assign w15984 = ( ~w132 & w15972 ) | ( ~w132 & w15978 ) | ( w15972 & w15978 ) ;
  assign w15985 = ~w15972 & w15984 ;
  assign w15986 = w15983 | w15985 ;
  assign w15987 = ~w15980 & w15986 ;
  assign w15988 = w15491 | w15496 ;
  assign w15989 = w15515 & ~w15988 ;
  assign w15990 = w15494 ^ w15989 ;
  assign w15991 = ( ~w15509 & w15987 ) | ( ~w15509 & w15990 ) | ( w15987 & w15990 ) ;
  assign w15992 = w15498 & ~w15991 ;
  assign w15993 = ~w15501 & w15515 ;
  assign w15994 = ( w15991 & ~w15992 ) | ( w15991 & w15993 ) | ( ~w15992 & w15993 ) ;
  assign w15995 = w15509 | w15994 ;
  assign w15996 = ~w129 & w15995 ;
  assign w15997 = ( w15980 & w15986 ) | ( w15980 & w15990 ) | ( w15986 & w15990 ) ;
  assign w15998 = ~w15980 & w15997 ;
  assign w15999 = ( w129 & w15498 ) | ( w129 & w15501 ) | ( w15498 & w15501 ) ;
  assign w16000 = ( w15501 & ~w15515 ) | ( w15501 & w15999 ) | ( ~w15515 & w15999 ) ;
  assign w16001 = w15498 & w16000 ;
  assign w16002 = w15999 ^ w16001 ;
  assign w16003 = ( w15996 & ~w15998 ) | ( w15996 & w16002 ) | ( ~w15998 & w16002 ) ;
  assign w16004 = w15998 | w16003 ;
  assign w16005 = \pi004 | \pi005 ;
  assign w16006 = ( \pi006 & w15515 ) | ( \pi006 & ~w16005 ) | ( w15515 & ~w16005 ) ;
  assign w16007 = ( ~\pi006 & w15515 ) | ( ~\pi006 & w16004 ) | ( w15515 & w16004 ) ;
  assign w16008 = w16006 & w16007 ;
  assign w16009 = \pi006 & ~w16004 ;
  assign w16010 = ( ~\pi006 & w15507 ) | ( ~\pi006 & w16005 ) | ( w15507 & w16005 ) ;
  assign w16011 = ( ~w15507 & w15509 ) | ( ~w15507 & w15513 ) | ( w15509 & w15513 ) ;
  assign w16012 = ( w16009 & w16010 ) | ( w16009 & ~w16011 ) | ( w16010 & ~w16011 ) ;
  assign w16013 = ~w15507 & w16012 ;
  assign w16014 = ~\pi006 & w16004 ;
  assign w16015 = \pi007 ^ w16014 ;
  assign w16016 = w16013 | w16015 ;
  assign w16017 = ( w15032 & w16008 ) | ( w15032 & ~w16016 ) | ( w16008 & ~w16016 ) ;
  assign w16018 = w15032 & w16017 ;
  assign w16019 = ( ~w15032 & w16008 ) | ( ~w15032 & w16016 ) | ( w16008 & w16016 ) ;
  assign w16020 = ~w16008 & w16019 ;
  assign w16021 = w15996 | w15998 ;
  assign w16022 = w16002 | w16021 ;
  assign w16023 = w15515 ^ w16022 ;
  assign w16024 = ( w15515 & ~w15516 ) | ( w15515 & w16023 ) | ( ~w15516 & w16023 ) ;
  assign w16025 = \pi008 ^ w16024 ;
  assign w16026 = w16020 | w16025 ;
  assign w16027 = ( w14555 & w16018 ) | ( w14555 & ~w16026 ) | ( w16018 & ~w16026 ) ;
  assign w16028 = w14555 & w16027 ;
  assign w16029 = ( w15519 & ~w15524 ) | ( w15519 & w16004 ) | ( ~w15524 & w16004 ) ;
  assign w16030 = ~w15519 & w16029 ;
  assign w16031 = \pi009 ^ w16030 ;
  assign w16032 = w15525 ^ w16031 ;
  assign w16033 = ( ~w14555 & w16018 ) | ( ~w14555 & w16026 ) | ( w16018 & w16026 ) ;
  assign w16034 = ~w16018 & w16033 ;
  assign w16035 = w16032 | w16034 ;
  assign w16036 = ( w14077 & w16028 ) | ( w14077 & ~w16035 ) | ( w16028 & ~w16035 ) ;
  assign w16037 = w14077 & w16036 ;
  assign w16038 = w15529 | w15531 ;
  assign w16039 = w16004 & ~w16038 ;
  assign w16040 = w15536 ^ w16039 ;
  assign w16041 = ( ~w14077 & w16028 ) | ( ~w14077 & w16035 ) | ( w16028 & w16035 ) ;
  assign w16042 = ~w16028 & w16041 ;
  assign w16043 = w16040 | w16042 ;
  assign w16044 = ( w13607 & w16037 ) | ( w13607 & ~w16043 ) | ( w16037 & ~w16043 ) ;
  assign w16045 = w13607 & w16044 ;
  assign w16046 = w15539 | w15545 ;
  assign w16047 = w16004 & ~w16046 ;
  assign w16048 = w15543 ^ w16047 ;
  assign w16049 = ( ~w13607 & w16037 ) | ( ~w13607 & w16043 ) | ( w16037 & w16043 ) ;
  assign w16050 = ~w16037 & w16049 ;
  assign w16051 = w16048 | w16050 ;
  assign w16052 = ( w13145 & w16045 ) | ( w13145 & ~w16051 ) | ( w16045 & ~w16051 ) ;
  assign w16053 = w13145 & w16052 ;
  assign w16054 = w15548 | w15553 ;
  assign w16055 = w16004 & ~w16054 ;
  assign w16056 = w15551 ^ w16055 ;
  assign w16057 = ( ~w13145 & w16045 ) | ( ~w13145 & w16051 ) | ( w16045 & w16051 ) ;
  assign w16058 = ~w16045 & w16057 ;
  assign w16059 = w16056 | w16058 ;
  assign w16060 = ( w12691 & w16053 ) | ( w12691 & ~w16059 ) | ( w16053 & ~w16059 ) ;
  assign w16061 = w12691 & w16060 ;
  assign w16062 = w15556 | w15561 ;
  assign w16063 = w16004 & ~w16062 ;
  assign w16064 = w15559 ^ w16063 ;
  assign w16065 = ( ~w12691 & w16053 ) | ( ~w12691 & w16059 ) | ( w16053 & w16059 ) ;
  assign w16066 = ~w16053 & w16065 ;
  assign w16067 = w16064 | w16066 ;
  assign w16068 = ( w12245 & w16061 ) | ( w12245 & ~w16067 ) | ( w16061 & ~w16067 ) ;
  assign w16069 = w12245 & w16068 ;
  assign w16070 = w15564 | w15569 ;
  assign w16071 = w16004 & ~w16070 ;
  assign w16072 = w15567 ^ w16071 ;
  assign w16073 = ( ~w12245 & w16061 ) | ( ~w12245 & w16067 ) | ( w16061 & w16067 ) ;
  assign w16074 = ~w16061 & w16073 ;
  assign w16075 = w16072 | w16074 ;
  assign w16076 = ( w11807 & w16069 ) | ( w11807 & ~w16075 ) | ( w16069 & ~w16075 ) ;
  assign w16077 = w11807 & w16076 ;
  assign w16078 = w15572 | w15577 ;
  assign w16079 = w16004 & ~w16078 ;
  assign w16080 = w15575 ^ w16079 ;
  assign w16081 = ( ~w11807 & w16069 ) | ( ~w11807 & w16075 ) | ( w16069 & w16075 ) ;
  assign w16082 = ~w16069 & w16081 ;
  assign w16083 = w16080 | w16082 ;
  assign w16084 = ( w11377 & w16077 ) | ( w11377 & ~w16083 ) | ( w16077 & ~w16083 ) ;
  assign w16085 = w11377 & w16084 ;
  assign w16086 = w15580 | w15585 ;
  assign w16087 = w16004 & ~w16086 ;
  assign w16088 = w15583 ^ w16087 ;
  assign w16089 = ( ~w11377 & w16077 ) | ( ~w11377 & w16083 ) | ( w16077 & w16083 ) ;
  assign w16090 = ~w16077 & w16089 ;
  assign w16091 = w16088 | w16090 ;
  assign w16092 = ( w10955 & w16085 ) | ( w10955 & ~w16091 ) | ( w16085 & ~w16091 ) ;
  assign w16093 = w10955 & w16092 ;
  assign w16094 = w15588 | w15593 ;
  assign w16095 = w16004 & ~w16094 ;
  assign w16096 = w15591 ^ w16095 ;
  assign w16097 = ( ~w10955 & w16085 ) | ( ~w10955 & w16091 ) | ( w16085 & w16091 ) ;
  assign w16098 = ~w16085 & w16097 ;
  assign w16099 = w16096 | w16098 ;
  assign w16100 = ( w10541 & w16093 ) | ( w10541 & ~w16099 ) | ( w16093 & ~w16099 ) ;
  assign w16101 = w10541 & w16100 ;
  assign w16102 = w15596 | w15601 ;
  assign w16103 = w16004 & ~w16102 ;
  assign w16104 = w15599 ^ w16103 ;
  assign w16105 = ( ~w10541 & w16093 ) | ( ~w10541 & w16099 ) | ( w16093 & w16099 ) ;
  assign w16106 = ~w16093 & w16105 ;
  assign w16107 = w16104 | w16106 ;
  assign w16108 = ( w10135 & w16101 ) | ( w10135 & ~w16107 ) | ( w16101 & ~w16107 ) ;
  assign w16109 = w10135 & w16108 ;
  assign w16110 = w15604 | w15609 ;
  assign w16111 = w16004 & ~w16110 ;
  assign w16112 = w15607 ^ w16111 ;
  assign w16113 = ( ~w10135 & w16101 ) | ( ~w10135 & w16107 ) | ( w16101 & w16107 ) ;
  assign w16114 = ~w16101 & w16113 ;
  assign w16115 = w16112 | w16114 ;
  assign w16116 = ( w9737 & w16109 ) | ( w9737 & ~w16115 ) | ( w16109 & ~w16115 ) ;
  assign w16117 = w9737 & w16116 ;
  assign w16118 = w15612 | w15617 ;
  assign w16119 = w16004 & ~w16118 ;
  assign w16120 = w15615 ^ w16119 ;
  assign w16121 = ( ~w9737 & w16109 ) | ( ~w9737 & w16115 ) | ( w16109 & w16115 ) ;
  assign w16122 = ~w16109 & w16121 ;
  assign w16123 = w16120 | w16122 ;
  assign w16124 = ( w9347 & w16117 ) | ( w9347 & ~w16123 ) | ( w16117 & ~w16123 ) ;
  assign w16125 = w9347 & w16124 ;
  assign w16126 = w15620 | w15625 ;
  assign w16127 = w16004 & ~w16126 ;
  assign w16128 = w15623 ^ w16127 ;
  assign w16129 = ( ~w9347 & w16117 ) | ( ~w9347 & w16123 ) | ( w16117 & w16123 ) ;
  assign w16130 = ~w16117 & w16129 ;
  assign w16131 = w16128 | w16130 ;
  assign w16132 = ( w8965 & w16125 ) | ( w8965 & ~w16131 ) | ( w16125 & ~w16131 ) ;
  assign w16133 = w8965 & w16132 ;
  assign w16134 = w15628 | w15633 ;
  assign w16135 = w16004 & ~w16134 ;
  assign w16136 = w15631 ^ w16135 ;
  assign w16137 = ( ~w8965 & w16125 ) | ( ~w8965 & w16131 ) | ( w16125 & w16131 ) ;
  assign w16138 = ~w16125 & w16137 ;
  assign w16139 = w16136 | w16138 ;
  assign w16140 = ( w8591 & w16133 ) | ( w8591 & ~w16139 ) | ( w16133 & ~w16139 ) ;
  assign w16141 = w8591 & w16140 ;
  assign w16142 = w15636 | w15641 ;
  assign w16143 = w16004 & ~w16142 ;
  assign w16144 = w15639 ^ w16143 ;
  assign w16145 = ( ~w8591 & w16133 ) | ( ~w8591 & w16139 ) | ( w16133 & w16139 ) ;
  assign w16146 = ~w16133 & w16145 ;
  assign w16147 = w16144 | w16146 ;
  assign w16148 = ( w8225 & w16141 ) | ( w8225 & ~w16147 ) | ( w16141 & ~w16147 ) ;
  assign w16149 = w8225 & w16148 ;
  assign w16150 = w15644 | w15649 ;
  assign w16151 = w16004 & ~w16150 ;
  assign w16152 = w15647 ^ w16151 ;
  assign w16153 = ( ~w8225 & w16141 ) | ( ~w8225 & w16147 ) | ( w16141 & w16147 ) ;
  assign w16154 = ~w16141 & w16153 ;
  assign w16155 = w16152 | w16154 ;
  assign w16156 = ( w7867 & w16149 ) | ( w7867 & ~w16155 ) | ( w16149 & ~w16155 ) ;
  assign w16157 = w7867 & w16156 ;
  assign w16158 = w15652 | w15657 ;
  assign w16159 = w16004 & ~w16158 ;
  assign w16160 = w15655 ^ w16159 ;
  assign w16161 = ( ~w7867 & w16149 ) | ( ~w7867 & w16155 ) | ( w16149 & w16155 ) ;
  assign w16162 = ~w16149 & w16161 ;
  assign w16163 = w16160 | w16162 ;
  assign w16164 = ( w7517 & w16157 ) | ( w7517 & ~w16163 ) | ( w16157 & ~w16163 ) ;
  assign w16165 = w7517 & w16164 ;
  assign w16166 = w15660 | w15665 ;
  assign w16167 = w16004 & ~w16166 ;
  assign w16168 = w15663 ^ w16167 ;
  assign w16169 = ( ~w7517 & w16157 ) | ( ~w7517 & w16163 ) | ( w16157 & w16163 ) ;
  assign w16170 = ~w16157 & w16169 ;
  assign w16171 = w16168 | w16170 ;
  assign w16172 = ( w7175 & w16165 ) | ( w7175 & ~w16171 ) | ( w16165 & ~w16171 ) ;
  assign w16173 = w7175 & w16172 ;
  assign w16174 = w15668 | w15673 ;
  assign w16175 = w16004 & ~w16174 ;
  assign w16176 = w15671 ^ w16175 ;
  assign w16177 = ( ~w7175 & w16165 ) | ( ~w7175 & w16171 ) | ( w16165 & w16171 ) ;
  assign w16178 = ~w16165 & w16177 ;
  assign w16179 = w16176 | w16178 ;
  assign w16180 = ( w6841 & w16173 ) | ( w6841 & ~w16179 ) | ( w16173 & ~w16179 ) ;
  assign w16181 = w6841 & w16180 ;
  assign w16182 = w15676 | w15681 ;
  assign w16183 = w16004 & ~w16182 ;
  assign w16184 = w15679 ^ w16183 ;
  assign w16185 = ( ~w6841 & w16173 ) | ( ~w6841 & w16179 ) | ( w16173 & w16179 ) ;
  assign w16186 = ~w16173 & w16185 ;
  assign w16187 = w16184 | w16186 ;
  assign w16188 = ( w6515 & w16181 ) | ( w6515 & ~w16187 ) | ( w16181 & ~w16187 ) ;
  assign w16189 = w6515 & w16188 ;
  assign w16190 = w15684 | w15689 ;
  assign w16191 = w16004 & ~w16190 ;
  assign w16192 = w15687 ^ w16191 ;
  assign w16193 = ( ~w6515 & w16181 ) | ( ~w6515 & w16187 ) | ( w16181 & w16187 ) ;
  assign w16194 = ~w16181 & w16193 ;
  assign w16195 = w16192 | w16194 ;
  assign w16196 = ( w6197 & w16189 ) | ( w6197 & ~w16195 ) | ( w16189 & ~w16195 ) ;
  assign w16197 = w6197 & w16196 ;
  assign w16198 = w15692 | w15697 ;
  assign w16199 = w16004 & ~w16198 ;
  assign w16200 = w15695 ^ w16199 ;
  assign w16201 = ( ~w6197 & w16189 ) | ( ~w6197 & w16195 ) | ( w16189 & w16195 ) ;
  assign w16202 = ~w16189 & w16201 ;
  assign w16203 = w16200 | w16202 ;
  assign w16204 = ( w5887 & w16197 ) | ( w5887 & ~w16203 ) | ( w16197 & ~w16203 ) ;
  assign w16205 = w5887 & w16204 ;
  assign w16206 = w15700 | w15705 ;
  assign w16207 = w16004 & ~w16206 ;
  assign w16208 = w15703 ^ w16207 ;
  assign w16209 = ( ~w5887 & w16197 ) | ( ~w5887 & w16203 ) | ( w16197 & w16203 ) ;
  assign w16210 = ~w16197 & w16209 ;
  assign w16211 = w16208 | w16210 ;
  assign w16212 = ( w5585 & w16205 ) | ( w5585 & ~w16211 ) | ( w16205 & ~w16211 ) ;
  assign w16213 = w5585 & w16212 ;
  assign w16214 = w15708 | w15713 ;
  assign w16215 = w16004 & ~w16214 ;
  assign w16216 = w15711 ^ w16215 ;
  assign w16217 = ( ~w5585 & w16205 ) | ( ~w5585 & w16211 ) | ( w16205 & w16211 ) ;
  assign w16218 = ~w16205 & w16217 ;
  assign w16219 = w16216 | w16218 ;
  assign w16220 = ( w5291 & w16213 ) | ( w5291 & ~w16219 ) | ( w16213 & ~w16219 ) ;
  assign w16221 = w5291 & w16220 ;
  assign w16222 = w15716 | w15721 ;
  assign w16223 = w16004 & ~w16222 ;
  assign w16224 = w15719 ^ w16223 ;
  assign w16225 = ( ~w5291 & w16213 ) | ( ~w5291 & w16219 ) | ( w16213 & w16219 ) ;
  assign w16226 = ~w16213 & w16225 ;
  assign w16227 = w16224 | w16226 ;
  assign w16228 = ( w5005 & w16221 ) | ( w5005 & ~w16227 ) | ( w16221 & ~w16227 ) ;
  assign w16229 = w5005 & w16228 ;
  assign w16230 = w15724 | w15729 ;
  assign w16231 = w16004 & ~w16230 ;
  assign w16232 = w15727 ^ w16231 ;
  assign w16233 = ( ~w5005 & w16221 ) | ( ~w5005 & w16227 ) | ( w16221 & w16227 ) ;
  assign w16234 = ~w16221 & w16233 ;
  assign w16235 = w16232 | w16234 ;
  assign w16236 = ( w4727 & w16229 ) | ( w4727 & ~w16235 ) | ( w16229 & ~w16235 ) ;
  assign w16237 = w4727 & w16236 ;
  assign w16238 = w15732 | w15737 ;
  assign w16239 = w16004 & ~w16238 ;
  assign w16240 = w15735 ^ w16239 ;
  assign w16241 = ( ~w4727 & w16229 ) | ( ~w4727 & w16235 ) | ( w16229 & w16235 ) ;
  assign w16242 = ~w16229 & w16241 ;
  assign w16243 = w16240 | w16242 ;
  assign w16244 = ( w4457 & w16237 ) | ( w4457 & ~w16243 ) | ( w16237 & ~w16243 ) ;
  assign w16245 = w4457 & w16244 ;
  assign w16246 = w15740 | w15745 ;
  assign w16247 = w16004 & ~w16246 ;
  assign w16248 = w15743 ^ w16247 ;
  assign w16249 = ( ~w4457 & w16237 ) | ( ~w4457 & w16243 ) | ( w16237 & w16243 ) ;
  assign w16250 = ~w16237 & w16249 ;
  assign w16251 = w16248 | w16250 ;
  assign w16252 = ( w4195 & w16245 ) | ( w4195 & ~w16251 ) | ( w16245 & ~w16251 ) ;
  assign w16253 = w4195 & w16252 ;
  assign w16254 = w15748 | w15753 ;
  assign w16255 = w16004 & ~w16254 ;
  assign w16256 = w15751 ^ w16255 ;
  assign w16257 = ( ~w4195 & w16245 ) | ( ~w4195 & w16251 ) | ( w16245 & w16251 ) ;
  assign w16258 = ~w16245 & w16257 ;
  assign w16259 = w16256 | w16258 ;
  assign w16260 = ( w3941 & w16253 ) | ( w3941 & ~w16259 ) | ( w16253 & ~w16259 ) ;
  assign w16261 = w3941 & w16260 ;
  assign w16262 = w15756 | w15761 ;
  assign w16263 = w16004 & ~w16262 ;
  assign w16264 = w15759 ^ w16263 ;
  assign w16265 = ( ~w3941 & w16253 ) | ( ~w3941 & w16259 ) | ( w16253 & w16259 ) ;
  assign w16266 = ~w16253 & w16265 ;
  assign w16267 = w16264 | w16266 ;
  assign w16268 = ( w3695 & w16261 ) | ( w3695 & ~w16267 ) | ( w16261 & ~w16267 ) ;
  assign w16269 = w3695 & w16268 ;
  assign w16270 = w15764 | w15769 ;
  assign w16271 = w16004 & ~w16270 ;
  assign w16272 = w15767 ^ w16271 ;
  assign w16273 = ( ~w3695 & w16261 ) | ( ~w3695 & w16267 ) | ( w16261 & w16267 ) ;
  assign w16274 = ~w16261 & w16273 ;
  assign w16275 = w16272 | w16274 ;
  assign w16276 = ( w3457 & w16269 ) | ( w3457 & ~w16275 ) | ( w16269 & ~w16275 ) ;
  assign w16277 = w3457 & w16276 ;
  assign w16278 = w15772 | w15777 ;
  assign w16279 = w16004 & ~w16278 ;
  assign w16280 = w15775 ^ w16279 ;
  assign w16281 = ( ~w3457 & w16269 ) | ( ~w3457 & w16275 ) | ( w16269 & w16275 ) ;
  assign w16282 = ~w16269 & w16281 ;
  assign w16283 = w16280 | w16282 ;
  assign w16284 = ( w3227 & w16277 ) | ( w3227 & ~w16283 ) | ( w16277 & ~w16283 ) ;
  assign w16285 = w3227 & w16284 ;
  assign w16286 = w15780 | w15785 ;
  assign w16287 = w16004 & ~w16286 ;
  assign w16288 = w15783 ^ w16287 ;
  assign w16289 = ( ~w3227 & w16277 ) | ( ~w3227 & w16283 ) | ( w16277 & w16283 ) ;
  assign w16290 = ~w16277 & w16289 ;
  assign w16291 = w16288 | w16290 ;
  assign w16292 = ( w3005 & w16285 ) | ( w3005 & ~w16291 ) | ( w16285 & ~w16291 ) ;
  assign w16293 = w3005 & w16292 ;
  assign w16294 = w15788 | w15793 ;
  assign w16295 = w16004 & ~w16294 ;
  assign w16296 = w15791 ^ w16295 ;
  assign w16297 = ( ~w3005 & w16285 ) | ( ~w3005 & w16291 ) | ( w16285 & w16291 ) ;
  assign w16298 = ~w16285 & w16297 ;
  assign w16299 = w16296 | w16298 ;
  assign w16300 = ( w2791 & w16293 ) | ( w2791 & ~w16299 ) | ( w16293 & ~w16299 ) ;
  assign w16301 = w2791 & w16300 ;
  assign w16302 = w15796 | w15801 ;
  assign w16303 = w16004 & ~w16302 ;
  assign w16304 = w15799 ^ w16303 ;
  assign w16305 = ( ~w2791 & w16293 ) | ( ~w2791 & w16299 ) | ( w16293 & w16299 ) ;
  assign w16306 = ~w16293 & w16305 ;
  assign w16307 = w16304 | w16306 ;
  assign w16308 = ( w2585 & w16301 ) | ( w2585 & ~w16307 ) | ( w16301 & ~w16307 ) ;
  assign w16309 = w2585 & w16308 ;
  assign w16310 = w15804 | w15809 ;
  assign w16311 = w16004 & ~w16310 ;
  assign w16312 = w15807 ^ w16311 ;
  assign w16313 = ( ~w2585 & w16301 ) | ( ~w2585 & w16307 ) | ( w16301 & w16307 ) ;
  assign w16314 = ~w16301 & w16313 ;
  assign w16315 = w16312 | w16314 ;
  assign w16316 = ( w2387 & w16309 ) | ( w2387 & ~w16315 ) | ( w16309 & ~w16315 ) ;
  assign w16317 = w2387 & w16316 ;
  assign w16318 = w15812 | w15817 ;
  assign w16319 = w16004 & ~w16318 ;
  assign w16320 = w15815 ^ w16319 ;
  assign w16321 = ( ~w2387 & w16309 ) | ( ~w2387 & w16315 ) | ( w16309 & w16315 ) ;
  assign w16322 = ~w16309 & w16321 ;
  assign w16323 = w16320 | w16322 ;
  assign w16324 = ( w2197 & w16317 ) | ( w2197 & ~w16323 ) | ( w16317 & ~w16323 ) ;
  assign w16325 = w2197 & w16324 ;
  assign w16326 = w15820 | w15825 ;
  assign w16327 = w16004 & ~w16326 ;
  assign w16328 = w15823 ^ w16327 ;
  assign w16329 = ( ~w2197 & w16317 ) | ( ~w2197 & w16323 ) | ( w16317 & w16323 ) ;
  assign w16330 = ~w16317 & w16329 ;
  assign w16331 = w16328 | w16330 ;
  assign w16332 = ( w2015 & w16325 ) | ( w2015 & ~w16331 ) | ( w16325 & ~w16331 ) ;
  assign w16333 = w2015 & w16332 ;
  assign w16334 = w15828 | w15833 ;
  assign w16335 = w16004 & ~w16334 ;
  assign w16336 = w15831 ^ w16335 ;
  assign w16337 = ( ~w2015 & w16325 ) | ( ~w2015 & w16331 ) | ( w16325 & w16331 ) ;
  assign w16338 = ~w16325 & w16337 ;
  assign w16339 = w16336 | w16338 ;
  assign w16340 = ( w1841 & w16333 ) | ( w1841 & ~w16339 ) | ( w16333 & ~w16339 ) ;
  assign w16341 = w1841 & w16340 ;
  assign w16342 = w15836 | w15841 ;
  assign w16343 = w16004 & ~w16342 ;
  assign w16344 = w15839 ^ w16343 ;
  assign w16345 = ( ~w1841 & w16333 ) | ( ~w1841 & w16339 ) | ( w16333 & w16339 ) ;
  assign w16346 = ~w16333 & w16345 ;
  assign w16347 = w16344 | w16346 ;
  assign w16348 = ( w1675 & w16341 ) | ( w1675 & ~w16347 ) | ( w16341 & ~w16347 ) ;
  assign w16349 = w1675 & w16348 ;
  assign w16350 = w15844 | w15849 ;
  assign w16351 = w16004 & ~w16350 ;
  assign w16352 = w15847 ^ w16351 ;
  assign w16353 = ( ~w1675 & w16341 ) | ( ~w1675 & w16347 ) | ( w16341 & w16347 ) ;
  assign w16354 = ~w16341 & w16353 ;
  assign w16355 = w16352 | w16354 ;
  assign w16356 = ( w1517 & w16349 ) | ( w1517 & ~w16355 ) | ( w16349 & ~w16355 ) ;
  assign w16357 = w1517 & w16356 ;
  assign w16358 = w15852 | w15857 ;
  assign w16359 = w16004 & ~w16358 ;
  assign w16360 = w15855 ^ w16359 ;
  assign w16361 = ( ~w1517 & w16349 ) | ( ~w1517 & w16355 ) | ( w16349 & w16355 ) ;
  assign w16362 = ~w16349 & w16361 ;
  assign w16363 = w16360 | w16362 ;
  assign w16364 = ( w1367 & w16357 ) | ( w1367 & ~w16363 ) | ( w16357 & ~w16363 ) ;
  assign w16365 = w1367 & w16364 ;
  assign w16366 = w15860 | w15865 ;
  assign w16367 = w16004 & ~w16366 ;
  assign w16368 = w15863 ^ w16367 ;
  assign w16369 = ( ~w1367 & w16357 ) | ( ~w1367 & w16363 ) | ( w16357 & w16363 ) ;
  assign w16370 = ~w16357 & w16369 ;
  assign w16371 = w16368 | w16370 ;
  assign w16372 = ( w1225 & w16365 ) | ( w1225 & ~w16371 ) | ( w16365 & ~w16371 ) ;
  assign w16373 = w1225 & w16372 ;
  assign w16374 = w15868 | w15873 ;
  assign w16375 = w16004 & ~w16374 ;
  assign w16376 = w15871 ^ w16375 ;
  assign w16377 = ( ~w1225 & w16365 ) | ( ~w1225 & w16371 ) | ( w16365 & w16371 ) ;
  assign w16378 = ~w16365 & w16377 ;
  assign w16379 = w16376 | w16378 ;
  assign w16380 = ( w1091 & w16373 ) | ( w1091 & ~w16379 ) | ( w16373 & ~w16379 ) ;
  assign w16381 = w1091 & w16380 ;
  assign w16382 = w15876 | w15881 ;
  assign w16383 = w16004 & ~w16382 ;
  assign w16384 = w15879 ^ w16383 ;
  assign w16385 = ( ~w1091 & w16373 ) | ( ~w1091 & w16379 ) | ( w16373 & w16379 ) ;
  assign w16386 = ~w16373 & w16385 ;
  assign w16387 = w16384 | w16386 ;
  assign w16388 = ( w965 & w16381 ) | ( w965 & ~w16387 ) | ( w16381 & ~w16387 ) ;
  assign w16389 = w965 & w16388 ;
  assign w16390 = w15884 | w15889 ;
  assign w16391 = w16004 & ~w16390 ;
  assign w16392 = w15887 ^ w16391 ;
  assign w16393 = ( ~w965 & w16381 ) | ( ~w965 & w16387 ) | ( w16381 & w16387 ) ;
  assign w16394 = ~w16381 & w16393 ;
  assign w16395 = w16392 | w16394 ;
  assign w16396 = ( w847 & w16389 ) | ( w847 & ~w16395 ) | ( w16389 & ~w16395 ) ;
  assign w16397 = w847 & w16396 ;
  assign w16398 = w15892 | w15897 ;
  assign w16399 = w16004 & ~w16398 ;
  assign w16400 = w15895 ^ w16399 ;
  assign w16401 = ( ~w847 & w16389 ) | ( ~w847 & w16395 ) | ( w16389 & w16395 ) ;
  assign w16402 = ~w16389 & w16401 ;
  assign w16403 = w16400 | w16402 ;
  assign w16404 = ( w737 & w16397 ) | ( w737 & ~w16403 ) | ( w16397 & ~w16403 ) ;
  assign w16405 = w737 & w16404 ;
  assign w16406 = w15900 | w15905 ;
  assign w16407 = w16004 & ~w16406 ;
  assign w16408 = w15903 ^ w16407 ;
  assign w16409 = ( ~w737 & w16397 ) | ( ~w737 & w16403 ) | ( w16397 & w16403 ) ;
  assign w16410 = ~w16397 & w16409 ;
  assign w16411 = w16408 | w16410 ;
  assign w16412 = ( w635 & w16405 ) | ( w635 & ~w16411 ) | ( w16405 & ~w16411 ) ;
  assign w16413 = w635 & w16412 ;
  assign w16414 = w15908 | w15913 ;
  assign w16415 = w16004 & ~w16414 ;
  assign w16416 = w15911 ^ w16415 ;
  assign w16417 = ( ~w635 & w16405 ) | ( ~w635 & w16411 ) | ( w16405 & w16411 ) ;
  assign w16418 = ~w16405 & w16417 ;
  assign w16419 = w16416 | w16418 ;
  assign w16420 = ( w541 & w16413 ) | ( w541 & ~w16419 ) | ( w16413 & ~w16419 ) ;
  assign w16421 = w541 & w16420 ;
  assign w16422 = w15916 | w15921 ;
  assign w16423 = w16004 & ~w16422 ;
  assign w16424 = w15919 ^ w16423 ;
  assign w16425 = ( ~w541 & w16413 ) | ( ~w541 & w16419 ) | ( w16413 & w16419 ) ;
  assign w16426 = ~w16413 & w16425 ;
  assign w16427 = w16424 | w16426 ;
  assign w16428 = ( w455 & w16421 ) | ( w455 & ~w16427 ) | ( w16421 & ~w16427 ) ;
  assign w16429 = w455 & w16428 ;
  assign w16430 = w15924 | w15929 ;
  assign w16431 = w16004 & ~w16430 ;
  assign w16432 = w15927 ^ w16431 ;
  assign w16433 = ( ~w455 & w16421 ) | ( ~w455 & w16427 ) | ( w16421 & w16427 ) ;
  assign w16434 = ~w16421 & w16433 ;
  assign w16435 = w16432 | w16434 ;
  assign w16436 = ( w377 & w16429 ) | ( w377 & ~w16435 ) | ( w16429 & ~w16435 ) ;
  assign w16437 = w377 & w16436 ;
  assign w16438 = w15932 | w15937 ;
  assign w16439 = w16004 & ~w16438 ;
  assign w16440 = w15935 ^ w16439 ;
  assign w16441 = ( ~w377 & w16429 ) | ( ~w377 & w16435 ) | ( w16429 & w16435 ) ;
  assign w16442 = ~w16429 & w16441 ;
  assign w16443 = w16440 | w16442 ;
  assign w16444 = ( w307 & w16437 ) | ( w307 & ~w16443 ) | ( w16437 & ~w16443 ) ;
  assign w16445 = w307 & w16444 ;
  assign w16446 = w15940 | w15945 ;
  assign w16447 = w16004 & ~w16446 ;
  assign w16448 = w15943 ^ w16447 ;
  assign w16449 = ( ~w307 & w16437 ) | ( ~w307 & w16443 ) | ( w16437 & w16443 ) ;
  assign w16450 = ~w16437 & w16449 ;
  assign w16451 = w16448 | w16450 ;
  assign w16452 = ( w246 & w16445 ) | ( w246 & ~w16451 ) | ( w16445 & ~w16451 ) ;
  assign w16453 = w246 & w16452 ;
  assign w16454 = w15948 | w15953 ;
  assign w16455 = w16004 & ~w16454 ;
  assign w16456 = w15951 ^ w16455 ;
  assign w16457 = ( ~w246 & w16445 ) | ( ~w246 & w16451 ) | ( w16445 & w16451 ) ;
  assign w16458 = ~w16445 & w16457 ;
  assign w16459 = w16456 | w16458 ;
  assign w16460 = ( w185 & w16453 ) | ( w185 & ~w16459 ) | ( w16453 & ~w16459 ) ;
  assign w16461 = w185 & w16460 ;
  assign w16462 = w15956 | w15961 ;
  assign w16463 = w16004 & ~w16462 ;
  assign w16464 = w15959 ^ w16463 ;
  assign w16465 = ( ~w185 & w16453 ) | ( ~w185 & w16459 ) | ( w16453 & w16459 ) ;
  assign w16466 = ~w16453 & w16465 ;
  assign w16467 = w16464 | w16466 ;
  assign w16468 = ( w145 & w16461 ) | ( w145 & ~w16467 ) | ( w16461 & ~w16467 ) ;
  assign w16469 = w145 & w16468 ;
  assign w16470 = w15964 | w15969 ;
  assign w16471 = w16004 & ~w16470 ;
  assign w16472 = w15967 ^ w16471 ;
  assign w16473 = ( ~w145 & w16461 ) | ( ~w145 & w16467 ) | ( w16461 & w16467 ) ;
  assign w16474 = ~w16461 & w16473 ;
  assign w16475 = w16472 | w16474 ;
  assign w16476 = ( w132 & w16469 ) | ( w132 & ~w16475 ) | ( w16469 & ~w16475 ) ;
  assign w16477 = w132 & w16476 ;
  assign w16478 = ( ~w132 & w16469 ) | ( ~w132 & w16475 ) | ( w16469 & w16475 ) ;
  assign w16479 = ~w16469 & w16478 ;
  assign w16480 = w15972 | w15974 ;
  assign w16481 = w16004 & ~w16480 ;
  assign w16482 = w15977 ^ w16481 ;
  assign w16483 = w16479 | w16482 ;
  assign w16484 = ~w16477 & w16483 ;
  assign w16485 = w15980 | w15985 ;
  assign w16486 = w16004 & ~w16485 ;
  assign w16487 = w15983 ^ w16486 ;
  assign w16488 = ( ~w15998 & w16484 ) | ( ~w15998 & w16487 ) | ( w16484 & w16487 ) ;
  assign w16489 = w15987 & ~w16488 ;
  assign w16490 = ~w15990 & w16004 ;
  assign w16491 = ( w16488 & ~w16489 ) | ( w16488 & w16490 ) | ( ~w16489 & w16490 ) ;
  assign w16492 = w15998 | w16491 ;
  assign w16493 = ~w129 & w16492 ;
  assign w16494 = ( w16477 & w16483 ) | ( w16477 & w16487 ) | ( w16483 & w16487 ) ;
  assign w16495 = ~w16477 & w16494 ;
  assign w16496 = ( w129 & w15987 ) | ( w129 & w15990 ) | ( w15987 & w15990 ) ;
  assign w16497 = ( w15990 & ~w16004 ) | ( w15990 & w16496 ) | ( ~w16004 & w16496 ) ;
  assign w16498 = w15987 & w16497 ;
  assign w16499 = w16496 ^ w16498 ;
  assign w16500 = ( w16493 & ~w16495 ) | ( w16493 & w16499 ) | ( ~w16495 & w16499 ) ;
  assign w16501 = w16495 | w16500 ;
  assign w16502 = w16461 | w16466 ;
  assign w16503 = w16501 & ~w16502 ;
  assign w16504 = w16464 ^ w16503 ;
  assign w16505 = \pi002 | \pi003 ;
  assign w16506 = ( \pi004 & w16004 ) | ( \pi004 & ~w16505 ) | ( w16004 & ~w16505 ) ;
  assign w16507 = ( ~\pi004 & w16004 ) | ( ~\pi004 & w16501 ) | ( w16004 & w16501 ) ;
  assign w16508 = w16506 & w16507 ;
  assign w16509 = \pi004 & ~w16501 ;
  assign w16510 = ( ~\pi004 & w15996 ) | ( ~\pi004 & w16505 ) | ( w15996 & w16505 ) ;
  assign w16511 = ( ~w15996 & w15998 ) | ( ~w15996 & w16002 ) | ( w15998 & w16002 ) ;
  assign w16512 = ( w16509 & w16510 ) | ( w16509 & ~w16511 ) | ( w16510 & ~w16511 ) ;
  assign w16513 = ~w15996 & w16512 ;
  assign w16514 = ~\pi004 & w16501 ;
  assign w16515 = \pi005 ^ w16514 ;
  assign w16516 = w16513 | w16515 ;
  assign w16517 = ( w15515 & w16508 ) | ( w15515 & ~w16516 ) | ( w16508 & ~w16516 ) ;
  assign w16518 = w15515 & w16517 ;
  assign w16519 = ( ~w15515 & w16508 ) | ( ~w15515 & w16516 ) | ( w16508 & w16516 ) ;
  assign w16520 = ~w16508 & w16519 ;
  assign w16521 = w16493 | w16495 ;
  assign w16522 = w16499 | w16521 ;
  assign w16523 = w16004 ^ w16522 ;
  assign w16524 = ( w16004 & ~w16005 ) | ( w16004 & w16523 ) | ( ~w16005 & w16523 ) ;
  assign w16525 = \pi006 ^ w16524 ;
  assign w16526 = w16520 | w16525 ;
  assign w16527 = ( w15032 & w16518 ) | ( w15032 & ~w16526 ) | ( w16518 & ~w16526 ) ;
  assign w16528 = w15032 & w16527 ;
  assign w16529 = ( w16008 & ~w16013 ) | ( w16008 & w16501 ) | ( ~w16013 & w16501 ) ;
  assign w16530 = ~w16008 & w16529 ;
  assign w16531 = \pi007 ^ w16530 ;
  assign w16532 = w16014 ^ w16531 ;
  assign w16533 = ( ~w15032 & w16518 ) | ( ~w15032 & w16526 ) | ( w16518 & w16526 ) ;
  assign w16534 = ~w16518 & w16533 ;
  assign w16535 = w16532 | w16534 ;
  assign w16536 = ( w14555 & w16528 ) | ( w14555 & ~w16535 ) | ( w16528 & ~w16535 ) ;
  assign w16537 = w14555 & w16536 ;
  assign w16538 = w16018 | w16020 ;
  assign w16539 = w16501 & ~w16538 ;
  assign w16540 = w16025 ^ w16539 ;
  assign w16541 = ( ~w14555 & w16528 ) | ( ~w14555 & w16535 ) | ( w16528 & w16535 ) ;
  assign w16542 = ~w16528 & w16541 ;
  assign w16543 = w16540 | w16542 ;
  assign w16544 = ( w14077 & w16537 ) | ( w14077 & ~w16543 ) | ( w16537 & ~w16543 ) ;
  assign w16545 = w14077 & w16544 ;
  assign w16546 = w16028 | w16034 ;
  assign w16547 = w16501 & ~w16546 ;
  assign w16548 = w16032 ^ w16547 ;
  assign w16549 = ( ~w14077 & w16537 ) | ( ~w14077 & w16543 ) | ( w16537 & w16543 ) ;
  assign w16550 = ~w16537 & w16549 ;
  assign w16551 = w16548 | w16550 ;
  assign w16552 = ( w13607 & w16545 ) | ( w13607 & ~w16551 ) | ( w16545 & ~w16551 ) ;
  assign w16553 = w13607 & w16552 ;
  assign w16554 = w16037 | w16042 ;
  assign w16555 = w16501 & ~w16554 ;
  assign w16556 = w16040 ^ w16555 ;
  assign w16557 = ( ~w13607 & w16545 ) | ( ~w13607 & w16551 ) | ( w16545 & w16551 ) ;
  assign w16558 = ~w16545 & w16557 ;
  assign w16559 = w16556 | w16558 ;
  assign w16560 = ( w13145 & w16553 ) | ( w13145 & ~w16559 ) | ( w16553 & ~w16559 ) ;
  assign w16561 = w13145 & w16560 ;
  assign w16562 = w16045 | w16050 ;
  assign w16563 = w16501 & ~w16562 ;
  assign w16564 = w16048 ^ w16563 ;
  assign w16565 = ( ~w13145 & w16553 ) | ( ~w13145 & w16559 ) | ( w16553 & w16559 ) ;
  assign w16566 = ~w16553 & w16565 ;
  assign w16567 = w16564 | w16566 ;
  assign w16568 = ( w12691 & w16561 ) | ( w12691 & ~w16567 ) | ( w16561 & ~w16567 ) ;
  assign w16569 = w12691 & w16568 ;
  assign w16570 = w16053 | w16058 ;
  assign w16571 = w16501 & ~w16570 ;
  assign w16572 = w16056 ^ w16571 ;
  assign w16573 = ( ~w12691 & w16561 ) | ( ~w12691 & w16567 ) | ( w16561 & w16567 ) ;
  assign w16574 = ~w16561 & w16573 ;
  assign w16575 = w16572 | w16574 ;
  assign w16576 = ( w12245 & w16569 ) | ( w12245 & ~w16575 ) | ( w16569 & ~w16575 ) ;
  assign w16577 = w12245 & w16576 ;
  assign w16578 = w16061 | w16066 ;
  assign w16579 = w16501 & ~w16578 ;
  assign w16580 = w16064 ^ w16579 ;
  assign w16581 = ( ~w12245 & w16569 ) | ( ~w12245 & w16575 ) | ( w16569 & w16575 ) ;
  assign w16582 = ~w16569 & w16581 ;
  assign w16583 = w16580 | w16582 ;
  assign w16584 = ( w11807 & w16577 ) | ( w11807 & ~w16583 ) | ( w16577 & ~w16583 ) ;
  assign w16585 = w11807 & w16584 ;
  assign w16586 = w16069 | w16074 ;
  assign w16587 = w16501 & ~w16586 ;
  assign w16588 = w16072 ^ w16587 ;
  assign w16589 = ( ~w11807 & w16577 ) | ( ~w11807 & w16583 ) | ( w16577 & w16583 ) ;
  assign w16590 = ~w16577 & w16589 ;
  assign w16591 = w16588 | w16590 ;
  assign w16592 = ( w11377 & w16585 ) | ( w11377 & ~w16591 ) | ( w16585 & ~w16591 ) ;
  assign w16593 = w11377 & w16592 ;
  assign w16594 = w16077 | w16082 ;
  assign w16595 = w16501 & ~w16594 ;
  assign w16596 = w16080 ^ w16595 ;
  assign w16597 = ( ~w11377 & w16585 ) | ( ~w11377 & w16591 ) | ( w16585 & w16591 ) ;
  assign w16598 = ~w16585 & w16597 ;
  assign w16599 = w16596 | w16598 ;
  assign w16600 = ( w10955 & w16593 ) | ( w10955 & ~w16599 ) | ( w16593 & ~w16599 ) ;
  assign w16601 = w10955 & w16600 ;
  assign w16602 = w16085 | w16090 ;
  assign w16603 = w16501 & ~w16602 ;
  assign w16604 = w16088 ^ w16603 ;
  assign w16605 = ( ~w10955 & w16593 ) | ( ~w10955 & w16599 ) | ( w16593 & w16599 ) ;
  assign w16606 = ~w16593 & w16605 ;
  assign w16607 = w16604 | w16606 ;
  assign w16608 = ( w10541 & w16601 ) | ( w10541 & ~w16607 ) | ( w16601 & ~w16607 ) ;
  assign w16609 = w10541 & w16608 ;
  assign w16610 = w16093 | w16098 ;
  assign w16611 = w16501 & ~w16610 ;
  assign w16612 = w16096 ^ w16611 ;
  assign w16613 = ( ~w10541 & w16601 ) | ( ~w10541 & w16607 ) | ( w16601 & w16607 ) ;
  assign w16614 = ~w16601 & w16613 ;
  assign w16615 = w16612 | w16614 ;
  assign w16616 = ( w10135 & w16609 ) | ( w10135 & ~w16615 ) | ( w16609 & ~w16615 ) ;
  assign w16617 = w10135 & w16616 ;
  assign w16618 = w16101 | w16106 ;
  assign w16619 = w16501 & ~w16618 ;
  assign w16620 = w16104 ^ w16619 ;
  assign w16621 = ( ~w10135 & w16609 ) | ( ~w10135 & w16615 ) | ( w16609 & w16615 ) ;
  assign w16622 = ~w16609 & w16621 ;
  assign w16623 = w16620 | w16622 ;
  assign w16624 = ( w9737 & w16617 ) | ( w9737 & ~w16623 ) | ( w16617 & ~w16623 ) ;
  assign w16625 = w9737 & w16624 ;
  assign w16626 = w16109 | w16114 ;
  assign w16627 = w16501 & ~w16626 ;
  assign w16628 = w16112 ^ w16627 ;
  assign w16629 = ( ~w9737 & w16617 ) | ( ~w9737 & w16623 ) | ( w16617 & w16623 ) ;
  assign w16630 = ~w16617 & w16629 ;
  assign w16631 = w16628 | w16630 ;
  assign w16632 = ( w9347 & w16625 ) | ( w9347 & ~w16631 ) | ( w16625 & ~w16631 ) ;
  assign w16633 = w9347 & w16632 ;
  assign w16634 = w16117 | w16122 ;
  assign w16635 = w16501 & ~w16634 ;
  assign w16636 = w16120 ^ w16635 ;
  assign w16637 = ( ~w9347 & w16625 ) | ( ~w9347 & w16631 ) | ( w16625 & w16631 ) ;
  assign w16638 = ~w16625 & w16637 ;
  assign w16639 = w16636 | w16638 ;
  assign w16640 = ( w8965 & w16633 ) | ( w8965 & ~w16639 ) | ( w16633 & ~w16639 ) ;
  assign w16641 = w8965 & w16640 ;
  assign w16642 = w16125 | w16130 ;
  assign w16643 = w16501 & ~w16642 ;
  assign w16644 = w16128 ^ w16643 ;
  assign w16645 = ( ~w8965 & w16633 ) | ( ~w8965 & w16639 ) | ( w16633 & w16639 ) ;
  assign w16646 = ~w16633 & w16645 ;
  assign w16647 = w16644 | w16646 ;
  assign w16648 = ( w8591 & w16641 ) | ( w8591 & ~w16647 ) | ( w16641 & ~w16647 ) ;
  assign w16649 = w8591 & w16648 ;
  assign w16650 = w16133 | w16138 ;
  assign w16651 = w16501 & ~w16650 ;
  assign w16652 = w16136 ^ w16651 ;
  assign w16653 = ( ~w8591 & w16641 ) | ( ~w8591 & w16647 ) | ( w16641 & w16647 ) ;
  assign w16654 = ~w16641 & w16653 ;
  assign w16655 = w16652 | w16654 ;
  assign w16656 = ( w8225 & w16649 ) | ( w8225 & ~w16655 ) | ( w16649 & ~w16655 ) ;
  assign w16657 = w8225 & w16656 ;
  assign w16658 = w16141 | w16146 ;
  assign w16659 = w16501 & ~w16658 ;
  assign w16660 = w16144 ^ w16659 ;
  assign w16661 = ( ~w8225 & w16649 ) | ( ~w8225 & w16655 ) | ( w16649 & w16655 ) ;
  assign w16662 = ~w16649 & w16661 ;
  assign w16663 = w16660 | w16662 ;
  assign w16664 = ( w7867 & w16657 ) | ( w7867 & ~w16663 ) | ( w16657 & ~w16663 ) ;
  assign w16665 = w7867 & w16664 ;
  assign w16666 = w16149 | w16154 ;
  assign w16667 = w16501 & ~w16666 ;
  assign w16668 = w16152 ^ w16667 ;
  assign w16669 = ( ~w7867 & w16657 ) | ( ~w7867 & w16663 ) | ( w16657 & w16663 ) ;
  assign w16670 = ~w16657 & w16669 ;
  assign w16671 = w16668 | w16670 ;
  assign w16672 = ( w7517 & w16665 ) | ( w7517 & ~w16671 ) | ( w16665 & ~w16671 ) ;
  assign w16673 = w7517 & w16672 ;
  assign w16674 = w16157 | w16162 ;
  assign w16675 = w16501 & ~w16674 ;
  assign w16676 = w16160 ^ w16675 ;
  assign w16677 = ( ~w7517 & w16665 ) | ( ~w7517 & w16671 ) | ( w16665 & w16671 ) ;
  assign w16678 = ~w16665 & w16677 ;
  assign w16679 = w16676 | w16678 ;
  assign w16680 = ( w7175 & w16673 ) | ( w7175 & ~w16679 ) | ( w16673 & ~w16679 ) ;
  assign w16681 = w7175 & w16680 ;
  assign w16682 = w16165 | w16170 ;
  assign w16683 = w16501 & ~w16682 ;
  assign w16684 = w16168 ^ w16683 ;
  assign w16685 = ( ~w7175 & w16673 ) | ( ~w7175 & w16679 ) | ( w16673 & w16679 ) ;
  assign w16686 = ~w16673 & w16685 ;
  assign w16687 = w16684 | w16686 ;
  assign w16688 = ( w6841 & w16681 ) | ( w6841 & ~w16687 ) | ( w16681 & ~w16687 ) ;
  assign w16689 = w6841 & w16688 ;
  assign w16690 = w16173 | w16178 ;
  assign w16691 = w16501 & ~w16690 ;
  assign w16692 = w16176 ^ w16691 ;
  assign w16693 = ( ~w6841 & w16681 ) | ( ~w6841 & w16687 ) | ( w16681 & w16687 ) ;
  assign w16694 = ~w16681 & w16693 ;
  assign w16695 = w16692 | w16694 ;
  assign w16696 = ( w6515 & w16689 ) | ( w6515 & ~w16695 ) | ( w16689 & ~w16695 ) ;
  assign w16697 = w6515 & w16696 ;
  assign w16698 = w16181 | w16186 ;
  assign w16699 = w16501 & ~w16698 ;
  assign w16700 = w16184 ^ w16699 ;
  assign w16701 = ( ~w6515 & w16689 ) | ( ~w6515 & w16695 ) | ( w16689 & w16695 ) ;
  assign w16702 = ~w16689 & w16701 ;
  assign w16703 = w16700 | w16702 ;
  assign w16704 = ( w6197 & w16697 ) | ( w6197 & ~w16703 ) | ( w16697 & ~w16703 ) ;
  assign w16705 = w6197 & w16704 ;
  assign w16706 = w16189 | w16194 ;
  assign w16707 = w16501 & ~w16706 ;
  assign w16708 = w16192 ^ w16707 ;
  assign w16709 = ( ~w6197 & w16697 ) | ( ~w6197 & w16703 ) | ( w16697 & w16703 ) ;
  assign w16710 = ~w16697 & w16709 ;
  assign w16711 = w16708 | w16710 ;
  assign w16712 = ( w5887 & w16705 ) | ( w5887 & ~w16711 ) | ( w16705 & ~w16711 ) ;
  assign w16713 = w5887 & w16712 ;
  assign w16714 = w16197 | w16202 ;
  assign w16715 = w16501 & ~w16714 ;
  assign w16716 = w16200 ^ w16715 ;
  assign w16717 = ( ~w5887 & w16705 ) | ( ~w5887 & w16711 ) | ( w16705 & w16711 ) ;
  assign w16718 = ~w16705 & w16717 ;
  assign w16719 = w16716 | w16718 ;
  assign w16720 = ( w5585 & w16713 ) | ( w5585 & ~w16719 ) | ( w16713 & ~w16719 ) ;
  assign w16721 = w5585 & w16720 ;
  assign w16722 = w16205 | w16210 ;
  assign w16723 = w16501 & ~w16722 ;
  assign w16724 = w16208 ^ w16723 ;
  assign w16725 = ( ~w5585 & w16713 ) | ( ~w5585 & w16719 ) | ( w16713 & w16719 ) ;
  assign w16726 = ~w16713 & w16725 ;
  assign w16727 = w16724 | w16726 ;
  assign w16728 = ( w5291 & w16721 ) | ( w5291 & ~w16727 ) | ( w16721 & ~w16727 ) ;
  assign w16729 = w5291 & w16728 ;
  assign w16730 = w16213 | w16218 ;
  assign w16731 = w16501 & ~w16730 ;
  assign w16732 = w16216 ^ w16731 ;
  assign w16733 = ( ~w5291 & w16721 ) | ( ~w5291 & w16727 ) | ( w16721 & w16727 ) ;
  assign w16734 = ~w16721 & w16733 ;
  assign w16735 = w16732 | w16734 ;
  assign w16736 = ( w5005 & w16729 ) | ( w5005 & ~w16735 ) | ( w16729 & ~w16735 ) ;
  assign w16737 = w5005 & w16736 ;
  assign w16738 = w16221 | w16226 ;
  assign w16739 = w16501 & ~w16738 ;
  assign w16740 = w16224 ^ w16739 ;
  assign w16741 = ( ~w5005 & w16729 ) | ( ~w5005 & w16735 ) | ( w16729 & w16735 ) ;
  assign w16742 = ~w16729 & w16741 ;
  assign w16743 = w16740 | w16742 ;
  assign w16744 = ( w4727 & w16737 ) | ( w4727 & ~w16743 ) | ( w16737 & ~w16743 ) ;
  assign w16745 = w4727 & w16744 ;
  assign w16746 = w16229 | w16234 ;
  assign w16747 = w16501 & ~w16746 ;
  assign w16748 = w16232 ^ w16747 ;
  assign w16749 = ( ~w4727 & w16737 ) | ( ~w4727 & w16743 ) | ( w16737 & w16743 ) ;
  assign w16750 = ~w16737 & w16749 ;
  assign w16751 = w16748 | w16750 ;
  assign w16752 = ( w4457 & w16745 ) | ( w4457 & ~w16751 ) | ( w16745 & ~w16751 ) ;
  assign w16753 = w4457 & w16752 ;
  assign w16754 = w16237 | w16242 ;
  assign w16755 = w16501 & ~w16754 ;
  assign w16756 = w16240 ^ w16755 ;
  assign w16757 = ( ~w4457 & w16745 ) | ( ~w4457 & w16751 ) | ( w16745 & w16751 ) ;
  assign w16758 = ~w16745 & w16757 ;
  assign w16759 = w16756 | w16758 ;
  assign w16760 = ( w4195 & w16753 ) | ( w4195 & ~w16759 ) | ( w16753 & ~w16759 ) ;
  assign w16761 = w4195 & w16760 ;
  assign w16762 = w16245 | w16250 ;
  assign w16763 = w16501 & ~w16762 ;
  assign w16764 = w16248 ^ w16763 ;
  assign w16765 = ( ~w4195 & w16753 ) | ( ~w4195 & w16759 ) | ( w16753 & w16759 ) ;
  assign w16766 = ~w16753 & w16765 ;
  assign w16767 = w16764 | w16766 ;
  assign w16768 = ( w3941 & w16761 ) | ( w3941 & ~w16767 ) | ( w16761 & ~w16767 ) ;
  assign w16769 = w3941 & w16768 ;
  assign w16770 = w16253 | w16258 ;
  assign w16771 = w16501 & ~w16770 ;
  assign w16772 = w16256 ^ w16771 ;
  assign w16773 = ( ~w3941 & w16761 ) | ( ~w3941 & w16767 ) | ( w16761 & w16767 ) ;
  assign w16774 = ~w16761 & w16773 ;
  assign w16775 = w16772 | w16774 ;
  assign w16776 = ( w3695 & w16769 ) | ( w3695 & ~w16775 ) | ( w16769 & ~w16775 ) ;
  assign w16777 = w3695 & w16776 ;
  assign w16778 = w16261 | w16266 ;
  assign w16779 = w16501 & ~w16778 ;
  assign w16780 = w16264 ^ w16779 ;
  assign w16781 = ( ~w3695 & w16769 ) | ( ~w3695 & w16775 ) | ( w16769 & w16775 ) ;
  assign w16782 = ~w16769 & w16781 ;
  assign w16783 = w16780 | w16782 ;
  assign w16784 = ( w3457 & w16777 ) | ( w3457 & ~w16783 ) | ( w16777 & ~w16783 ) ;
  assign w16785 = w3457 & w16784 ;
  assign w16786 = w16269 | w16274 ;
  assign w16787 = w16501 & ~w16786 ;
  assign w16788 = w16272 ^ w16787 ;
  assign w16789 = ( ~w3457 & w16777 ) | ( ~w3457 & w16783 ) | ( w16777 & w16783 ) ;
  assign w16790 = ~w16777 & w16789 ;
  assign w16791 = w16788 | w16790 ;
  assign w16792 = ( w3227 & w16785 ) | ( w3227 & ~w16791 ) | ( w16785 & ~w16791 ) ;
  assign w16793 = w3227 & w16792 ;
  assign w16794 = w16277 | w16282 ;
  assign w16795 = w16501 & ~w16794 ;
  assign w16796 = w16280 ^ w16795 ;
  assign w16797 = ( ~w3227 & w16785 ) | ( ~w3227 & w16791 ) | ( w16785 & w16791 ) ;
  assign w16798 = ~w16785 & w16797 ;
  assign w16799 = w16796 | w16798 ;
  assign w16800 = ( w3005 & w16793 ) | ( w3005 & ~w16799 ) | ( w16793 & ~w16799 ) ;
  assign w16801 = w3005 & w16800 ;
  assign w16802 = w16285 | w16290 ;
  assign w16803 = w16501 & ~w16802 ;
  assign w16804 = w16288 ^ w16803 ;
  assign w16805 = ( ~w3005 & w16793 ) | ( ~w3005 & w16799 ) | ( w16793 & w16799 ) ;
  assign w16806 = ~w16793 & w16805 ;
  assign w16807 = w16804 | w16806 ;
  assign w16808 = ( w2791 & w16801 ) | ( w2791 & ~w16807 ) | ( w16801 & ~w16807 ) ;
  assign w16809 = w2791 & w16808 ;
  assign w16810 = w16293 | w16298 ;
  assign w16811 = w16501 & ~w16810 ;
  assign w16812 = w16296 ^ w16811 ;
  assign w16813 = ( ~w2791 & w16801 ) | ( ~w2791 & w16807 ) | ( w16801 & w16807 ) ;
  assign w16814 = ~w16801 & w16813 ;
  assign w16815 = w16812 | w16814 ;
  assign w16816 = ( w2585 & w16809 ) | ( w2585 & ~w16815 ) | ( w16809 & ~w16815 ) ;
  assign w16817 = w2585 & w16816 ;
  assign w16818 = w16301 | w16306 ;
  assign w16819 = w16501 & ~w16818 ;
  assign w16820 = w16304 ^ w16819 ;
  assign w16821 = ( ~w2585 & w16809 ) | ( ~w2585 & w16815 ) | ( w16809 & w16815 ) ;
  assign w16822 = ~w16809 & w16821 ;
  assign w16823 = w16820 | w16822 ;
  assign w16824 = ( w2387 & w16817 ) | ( w2387 & ~w16823 ) | ( w16817 & ~w16823 ) ;
  assign w16825 = w2387 & w16824 ;
  assign w16826 = w16309 | w16314 ;
  assign w16827 = w16501 & ~w16826 ;
  assign w16828 = w16312 ^ w16827 ;
  assign w16829 = ( ~w2387 & w16817 ) | ( ~w2387 & w16823 ) | ( w16817 & w16823 ) ;
  assign w16830 = ~w16817 & w16829 ;
  assign w16831 = w16828 | w16830 ;
  assign w16832 = ( w2197 & w16825 ) | ( w2197 & ~w16831 ) | ( w16825 & ~w16831 ) ;
  assign w16833 = w2197 & w16832 ;
  assign w16834 = w16317 | w16322 ;
  assign w16835 = w16501 & ~w16834 ;
  assign w16836 = w16320 ^ w16835 ;
  assign w16837 = ( ~w2197 & w16825 ) | ( ~w2197 & w16831 ) | ( w16825 & w16831 ) ;
  assign w16838 = ~w16825 & w16837 ;
  assign w16839 = w16836 | w16838 ;
  assign w16840 = ( w2015 & w16833 ) | ( w2015 & ~w16839 ) | ( w16833 & ~w16839 ) ;
  assign w16841 = w2015 & w16840 ;
  assign w16842 = w16325 | w16330 ;
  assign w16843 = w16501 & ~w16842 ;
  assign w16844 = w16328 ^ w16843 ;
  assign w16845 = ( ~w2015 & w16833 ) | ( ~w2015 & w16839 ) | ( w16833 & w16839 ) ;
  assign w16846 = ~w16833 & w16845 ;
  assign w16847 = w16844 | w16846 ;
  assign w16848 = ( w1841 & w16841 ) | ( w1841 & ~w16847 ) | ( w16841 & ~w16847 ) ;
  assign w16849 = w1841 & w16848 ;
  assign w16850 = w16333 | w16338 ;
  assign w16851 = w16501 & ~w16850 ;
  assign w16852 = w16336 ^ w16851 ;
  assign w16853 = ( ~w1841 & w16841 ) | ( ~w1841 & w16847 ) | ( w16841 & w16847 ) ;
  assign w16854 = ~w16841 & w16853 ;
  assign w16855 = w16852 | w16854 ;
  assign w16856 = ( w1675 & w16849 ) | ( w1675 & ~w16855 ) | ( w16849 & ~w16855 ) ;
  assign w16857 = w1675 & w16856 ;
  assign w16858 = w16341 | w16346 ;
  assign w16859 = w16501 & ~w16858 ;
  assign w16860 = w16344 ^ w16859 ;
  assign w16861 = ( ~w1675 & w16849 ) | ( ~w1675 & w16855 ) | ( w16849 & w16855 ) ;
  assign w16862 = ~w16849 & w16861 ;
  assign w16863 = w16860 | w16862 ;
  assign w16864 = ( w1517 & w16857 ) | ( w1517 & ~w16863 ) | ( w16857 & ~w16863 ) ;
  assign w16865 = w1517 & w16864 ;
  assign w16866 = w16349 | w16354 ;
  assign w16867 = w16501 & ~w16866 ;
  assign w16868 = w16352 ^ w16867 ;
  assign w16869 = ( ~w1517 & w16857 ) | ( ~w1517 & w16863 ) | ( w16857 & w16863 ) ;
  assign w16870 = ~w16857 & w16869 ;
  assign w16871 = w16868 | w16870 ;
  assign w16872 = ( w1367 & w16865 ) | ( w1367 & ~w16871 ) | ( w16865 & ~w16871 ) ;
  assign w16873 = w1367 & w16872 ;
  assign w16874 = w16357 | w16362 ;
  assign w16875 = w16501 & ~w16874 ;
  assign w16876 = w16360 ^ w16875 ;
  assign w16877 = ( ~w1367 & w16865 ) | ( ~w1367 & w16871 ) | ( w16865 & w16871 ) ;
  assign w16878 = ~w16865 & w16877 ;
  assign w16879 = w16876 | w16878 ;
  assign w16880 = ( w1225 & w16873 ) | ( w1225 & ~w16879 ) | ( w16873 & ~w16879 ) ;
  assign w16881 = w1225 & w16880 ;
  assign w16882 = w16365 | w16370 ;
  assign w16883 = w16501 & ~w16882 ;
  assign w16884 = w16368 ^ w16883 ;
  assign w16885 = ( ~w1225 & w16873 ) | ( ~w1225 & w16879 ) | ( w16873 & w16879 ) ;
  assign w16886 = ~w16873 & w16885 ;
  assign w16887 = w16884 | w16886 ;
  assign w16888 = ( w1091 & w16881 ) | ( w1091 & ~w16887 ) | ( w16881 & ~w16887 ) ;
  assign w16889 = w1091 & w16888 ;
  assign w16890 = w16373 | w16378 ;
  assign w16891 = w16501 & ~w16890 ;
  assign w16892 = w16376 ^ w16891 ;
  assign w16893 = ( ~w1091 & w16881 ) | ( ~w1091 & w16887 ) | ( w16881 & w16887 ) ;
  assign w16894 = ~w16881 & w16893 ;
  assign w16895 = w16892 | w16894 ;
  assign w16896 = ( w965 & w16889 ) | ( w965 & ~w16895 ) | ( w16889 & ~w16895 ) ;
  assign w16897 = w965 & w16896 ;
  assign w16898 = w16381 | w16386 ;
  assign w16899 = w16501 & ~w16898 ;
  assign w16900 = w16384 ^ w16899 ;
  assign w16901 = ( ~w965 & w16889 ) | ( ~w965 & w16895 ) | ( w16889 & w16895 ) ;
  assign w16902 = ~w16889 & w16901 ;
  assign w16903 = w16900 | w16902 ;
  assign w16904 = ( w847 & w16897 ) | ( w847 & ~w16903 ) | ( w16897 & ~w16903 ) ;
  assign w16905 = w847 & w16904 ;
  assign w16906 = w16389 | w16394 ;
  assign w16907 = w16501 & ~w16906 ;
  assign w16908 = w16392 ^ w16907 ;
  assign w16909 = ( ~w847 & w16897 ) | ( ~w847 & w16903 ) | ( w16897 & w16903 ) ;
  assign w16910 = ~w16897 & w16909 ;
  assign w16911 = w16908 | w16910 ;
  assign w16912 = ( w737 & w16905 ) | ( w737 & ~w16911 ) | ( w16905 & ~w16911 ) ;
  assign w16913 = w737 & w16912 ;
  assign w16914 = w16397 | w16402 ;
  assign w16915 = w16501 & ~w16914 ;
  assign w16916 = w16400 ^ w16915 ;
  assign w16917 = ( ~w737 & w16905 ) | ( ~w737 & w16911 ) | ( w16905 & w16911 ) ;
  assign w16918 = ~w16905 & w16917 ;
  assign w16919 = w16916 | w16918 ;
  assign w16920 = ( w635 & w16913 ) | ( w635 & ~w16919 ) | ( w16913 & ~w16919 ) ;
  assign w16921 = w635 & w16920 ;
  assign w16922 = w16405 | w16410 ;
  assign w16923 = w16501 & ~w16922 ;
  assign w16924 = w16408 ^ w16923 ;
  assign w16925 = ( ~w635 & w16913 ) | ( ~w635 & w16919 ) | ( w16913 & w16919 ) ;
  assign w16926 = ~w16913 & w16925 ;
  assign w16927 = w16924 | w16926 ;
  assign w16928 = ( w541 & w16921 ) | ( w541 & ~w16927 ) | ( w16921 & ~w16927 ) ;
  assign w16929 = w541 & w16928 ;
  assign w16930 = w16413 | w16418 ;
  assign w16931 = w16501 & ~w16930 ;
  assign w16932 = w16416 ^ w16931 ;
  assign w16933 = ( ~w541 & w16921 ) | ( ~w541 & w16927 ) | ( w16921 & w16927 ) ;
  assign w16934 = ~w16921 & w16933 ;
  assign w16935 = w16932 | w16934 ;
  assign w16936 = ( w455 & w16929 ) | ( w455 & ~w16935 ) | ( w16929 & ~w16935 ) ;
  assign w16937 = w455 & w16936 ;
  assign w16938 = w16421 | w16426 ;
  assign w16939 = w16501 & ~w16938 ;
  assign w16940 = w16424 ^ w16939 ;
  assign w16941 = ( ~w455 & w16929 ) | ( ~w455 & w16935 ) | ( w16929 & w16935 ) ;
  assign w16942 = ~w16929 & w16941 ;
  assign w16943 = w16940 | w16942 ;
  assign w16944 = ( w377 & w16937 ) | ( w377 & ~w16943 ) | ( w16937 & ~w16943 ) ;
  assign w16945 = w377 & w16944 ;
  assign w16946 = w16429 | w16434 ;
  assign w16947 = w16501 & ~w16946 ;
  assign w16948 = w16432 ^ w16947 ;
  assign w16949 = ( ~w377 & w16937 ) | ( ~w377 & w16943 ) | ( w16937 & w16943 ) ;
  assign w16950 = ~w16937 & w16949 ;
  assign w16951 = w16948 | w16950 ;
  assign w16952 = ( w307 & w16945 ) | ( w307 & ~w16951 ) | ( w16945 & ~w16951 ) ;
  assign w16953 = w307 & w16952 ;
  assign w16954 = w16437 | w16442 ;
  assign w16955 = w16501 & ~w16954 ;
  assign w16956 = w16440 ^ w16955 ;
  assign w16957 = ( ~w307 & w16945 ) | ( ~w307 & w16951 ) | ( w16945 & w16951 ) ;
  assign w16958 = ~w16945 & w16957 ;
  assign w16959 = w16956 | w16958 ;
  assign w16960 = ( w246 & w16953 ) | ( w246 & ~w16959 ) | ( w16953 & ~w16959 ) ;
  assign w16961 = w246 & w16960 ;
  assign w16962 = w16445 | w16450 ;
  assign w16963 = w16501 & ~w16962 ;
  assign w16964 = w16448 ^ w16963 ;
  assign w16965 = ( ~w246 & w16953 ) | ( ~w246 & w16959 ) | ( w16953 & w16959 ) ;
  assign w16966 = ~w16953 & w16965 ;
  assign w16967 = w16964 | w16966 ;
  assign w16968 = ( w185 & w16961 ) | ( w185 & ~w16967 ) | ( w16961 & ~w16967 ) ;
  assign w16969 = w185 & w16968 ;
  assign w16970 = w16453 | w16458 ;
  assign w16971 = w16501 & ~w16970 ;
  assign w16972 = w16456 ^ w16971 ;
  assign w16973 = ( ~w185 & w16961 ) | ( ~w185 & w16967 ) | ( w16961 & w16967 ) ;
  assign w16974 = ~w16961 & w16973 ;
  assign w16975 = w16972 | w16974 ;
  assign w16976 = ( w145 & w16969 ) | ( w145 & ~w16975 ) | ( w16969 & ~w16975 ) ;
  assign w16977 = w145 & w16976 ;
  assign w16978 = ( ~w145 & w16969 ) | ( ~w145 & w16975 ) | ( w16969 & w16975 ) ;
  assign w16979 = ~w16969 & w16978 ;
  assign w16980 = w16504 | w16979 ;
  assign w16981 = ( w132 & w16977 ) | ( w132 & ~w16980 ) | ( w16977 & ~w16980 ) ;
  assign w16982 = w132 & w16981 ;
  assign w16983 = w16469 | w16474 ;
  assign w16984 = w16501 & ~w16983 ;
  assign w16985 = w16472 ^ w16984 ;
  assign w16986 = ( ~w132 & w16977 ) | ( ~w132 & w16980 ) | ( w16977 & w16980 ) ;
  assign w16987 = ~w16977 & w16986 ;
  assign w16988 = w16985 | w16987 ;
  assign w16989 = ~w16982 & w16988 ;
  assign w16990 = w16477 | w16479 ;
  assign w16991 = w16501 & ~w16990 ;
  assign w16992 = w16482 ^ w16991 ;
  assign w16993 = ( ~w16495 & w16989 ) | ( ~w16495 & w16992 ) | ( w16989 & w16992 ) ;
  assign w16994 = w16484 & ~w16993 ;
  assign w16995 = ~w16487 & w16501 ;
  assign w16996 = ( w16993 & ~w16994 ) | ( w16993 & w16995 ) | ( ~w16994 & w16995 ) ;
  assign w16997 = w16495 | w16996 ;
  assign w16998 = ~w129 & w16997 ;
  assign w16999 = ( w16982 & w16988 ) | ( w16982 & w16992 ) | ( w16988 & w16992 ) ;
  assign w17000 = ~w16982 & w16999 ;
  assign w17001 = ( w129 & w16484 ) | ( w129 & w16487 ) | ( w16484 & w16487 ) ;
  assign w17002 = ( w16487 & ~w16501 ) | ( w16487 & w17001 ) | ( ~w16501 & w17001 ) ;
  assign w17003 = w16484 & w17002 ;
  assign w17004 = w17001 ^ w17003 ;
  assign w17005 = ( w16998 & ~w17000 ) | ( w16998 & w17004 ) | ( ~w17000 & w17004 ) ;
  assign w17006 = w17000 | w17005 ;
  assign w17007 = w16977 | w16979 ;
  assign w17008 = w17006 & ~w17007 ;
  assign w17009 = w16504 ^ w17008 ;
  assign w17010 = w16961 | w16966 ;
  assign w17011 = w17006 & ~w17010 ;
  assign w17012 = w16964 ^ w17011 ;
  assign w17013 = w16945 | w16950 ;
  assign w17014 = w17006 & ~w17013 ;
  assign w17015 = w16948 ^ w17014 ;
  assign w17016 = w16929 | w16934 ;
  assign w17017 = w17006 & ~w17016 ;
  assign w17018 = w16932 ^ w17017 ;
  assign w17019 = w16913 | w16918 ;
  assign w17020 = w17006 & ~w17019 ;
  assign w17021 = w16916 ^ w17020 ;
  assign w17022 = w16897 | w16902 ;
  assign w17023 = w17006 & ~w17022 ;
  assign w17024 = w16900 ^ w17023 ;
  assign w17025 = w16881 | w16886 ;
  assign w17026 = w17006 & ~w17025 ;
  assign w17027 = w16884 ^ w17026 ;
  assign w17028 = w16865 | w16870 ;
  assign w17029 = w17006 & ~w17028 ;
  assign w17030 = w16868 ^ w17029 ;
  assign w17031 = w16849 | w16854 ;
  assign w17032 = w17006 & ~w17031 ;
  assign w17033 = w16852 ^ w17032 ;
  assign w17034 = w16833 | w16838 ;
  assign w17035 = w17006 & ~w17034 ;
  assign w17036 = w16836 ^ w17035 ;
  assign w17037 = w16817 | w16822 ;
  assign w17038 = w17006 & ~w17037 ;
  assign w17039 = w16820 ^ w17038 ;
  assign w17040 = w16801 | w16806 ;
  assign w17041 = w17006 & ~w17040 ;
  assign w17042 = w16804 ^ w17041 ;
  assign w17043 = w16785 | w16790 ;
  assign w17044 = w17006 & ~w17043 ;
  assign w17045 = w16788 ^ w17044 ;
  assign w17046 = w16769 | w16774 ;
  assign w17047 = w17006 & ~w17046 ;
  assign w17048 = w16772 ^ w17047 ;
  assign w17049 = w16753 | w16758 ;
  assign w17050 = w17006 & ~w17049 ;
  assign w17051 = w16756 ^ w17050 ;
  assign w17052 = w16737 | w16742 ;
  assign w17053 = w17006 & ~w17052 ;
  assign w17054 = w16740 ^ w17053 ;
  assign w17055 = w16721 | w16726 ;
  assign w17056 = w17006 & ~w17055 ;
  assign w17057 = w16724 ^ w17056 ;
  assign w17058 = w16705 | w16710 ;
  assign w17059 = w17006 & ~w17058 ;
  assign w17060 = w16708 ^ w17059 ;
  assign w17061 = w16689 | w16694 ;
  assign w17062 = w17006 & ~w17061 ;
  assign w17063 = w16692 ^ w17062 ;
  assign w17064 = w16673 | w16678 ;
  assign w17065 = w17006 & ~w17064 ;
  assign w17066 = w16676 ^ w17065 ;
  assign w17067 = w16657 | w16662 ;
  assign w17068 = w17006 & ~w17067 ;
  assign w17069 = w16660 ^ w17068 ;
  assign w17070 = w16641 | w16646 ;
  assign w17071 = w17006 & ~w17070 ;
  assign w17072 = w16644 ^ w17071 ;
  assign w17073 = w16625 | w16630 ;
  assign w17074 = w17006 & ~w17073 ;
  assign w17075 = w16628 ^ w17074 ;
  assign w17076 = w16609 | w16614 ;
  assign w17077 = w17006 & ~w17076 ;
  assign w17078 = w16612 ^ w17077 ;
  assign w17079 = w16593 | w16598 ;
  assign w17080 = w17006 & ~w17079 ;
  assign w17081 = w16596 ^ w17080 ;
  assign w17082 = w16577 | w16582 ;
  assign w17083 = w17006 & ~w17082 ;
  assign w17084 = w16580 ^ w17083 ;
  assign w17085 = w16561 | w16566 ;
  assign w17086 = w17006 & ~w17085 ;
  assign w17087 = w16564 ^ w17086 ;
  assign w17088 = w16545 | w16550 ;
  assign w17089 = w17006 & ~w17088 ;
  assign w17090 = w16548 ^ w17089 ;
  assign w17091 = w16528 | w16534 ;
  assign w17092 = w17006 & ~w17091 ;
  assign w17093 = w16532 ^ w17092 ;
  assign w17094 = ( w16508 & ~w16513 ) | ( w16508 & w17006 ) | ( ~w16513 & w17006 ) ;
  assign w17095 = ~w16508 & w17094 ;
  assign w17096 = \pi005 ^ w17095 ;
  assign w17097 = w16514 ^ w17096 ;
  assign w17098 = w16998 | w17000 ;
  assign w17099 = w17004 | w17098 ;
  assign w17100 = w16501 ^ w17099 ;
  assign w17101 = ( w16501 & ~w16505 ) | ( w16501 & w17100 ) | ( ~w16505 & w17100 ) ;
  assign w17102 = \pi004 ^ w17101 ;
  assign w17103 = \pi000 | \pi001 ;
  assign w17104 = \pi002 ^ w17103 ;
  assign w17105 = ( w16998 & w17000 ) | ( w16998 & ~w17004 ) | ( w17000 & ~w17004 ) ;
  assign w17106 = w17004 | w17105 ;
  assign w17107 = ( w17103 & w17104 ) | ( w17103 & ~w17106 ) | ( w17104 & ~w17106 ) ;
  assign w17108 = ~\pi002 & w17006 ;
  assign w17109 = \pi003 ^ w17108 ;
  assign w17110 = ( ~w16501 & w17107 ) | ( ~w16501 & w17109 ) | ( w17107 & w17109 ) ;
  assign w17111 = ( ~w16004 & w17102 ) | ( ~w16004 & w17110 ) | ( w17102 & w17110 ) ;
  assign w17112 = w17097 & w17111 ;
  assign w17113 = ~w15515 & w17097 ;
  assign w17114 = ( ~w15515 & w17111 ) | ( ~w15515 & w17113 ) | ( w17111 & w17113 ) ;
  assign w17115 = w16518 | w16520 ;
  assign w17116 = w17006 & ~w17115 ;
  assign w17117 = w16525 ^ w17116 ;
  assign w17118 = w17112 & ~w17114 ;
  assign w17119 = ( w17114 & w17117 ) | ( w17114 & ~w17118 ) | ( w17117 & ~w17118 ) ;
  assign w17120 = ( ~w15032 & w17118 ) | ( ~w15032 & w17119 ) | ( w17118 & w17119 ) ;
  assign w17121 = ( w17112 & w17114 ) | ( w17112 & w17117 ) | ( w17114 & w17117 ) ;
  assign w17122 = w17117 & w17121 ;
  assign w17123 = w16537 | w16542 ;
  assign w17124 = w17006 & ~w17123 ;
  assign w17125 = w16540 ^ w17124 ;
  assign w17126 = ~w14077 & w17125 ;
  assign w17127 = ( w17120 & w17122 ) | ( w17120 & ~w17126 ) | ( w17122 & ~w17126 ) ;
  assign w17128 = ( ~w14555 & w17093 ) | ( ~w14555 & w17127 ) | ( w17093 & w17127 ) ;
  assign w17129 = ( ~w14077 & w17126 ) | ( ~w14077 & w17128 ) | ( w17126 & w17128 ) ;
  assign w17130 = w17120 | w17122 ;
  assign w17131 = ( ~w14555 & w17093 ) | ( ~w14555 & w17130 ) | ( w17093 & w17130 ) ;
  assign w17132 = w17125 & w17131 ;
  assign w17133 = ( w17090 & w17129 ) | ( w17090 & w17132 ) | ( w17129 & w17132 ) ;
  assign w17134 = w17090 & w17133 ;
  assign w17135 = w17129 & ~w17132 ;
  assign w17136 = ( w17090 & w17132 ) | ( w17090 & ~w17135 ) | ( w17132 & ~w17135 ) ;
  assign w17137 = ( ~w13607 & w17135 ) | ( ~w13607 & w17136 ) | ( w17135 & w17136 ) ;
  assign w17138 = w16553 | w16558 ;
  assign w17139 = w17006 & ~w17138 ;
  assign w17140 = w16556 ^ w17139 ;
  assign w17141 = w17134 & ~w17137 ;
  assign w17142 = ( w17137 & w17140 ) | ( w17137 & ~w17141 ) | ( w17140 & ~w17141 ) ;
  assign w17143 = ( ~w13145 & w17141 ) | ( ~w13145 & w17142 ) | ( w17141 & w17142 ) ;
  assign w17144 = ( w17134 & w17137 ) | ( w17134 & w17140 ) | ( w17137 & w17140 ) ;
  assign w17145 = w17140 & w17144 ;
  assign w17146 = ( w17087 & w17143 ) | ( w17087 & w17145 ) | ( w17143 & w17145 ) ;
  assign w17147 = w17087 & w17146 ;
  assign w17148 = w17143 & ~w17145 ;
  assign w17149 = ( w17087 & w17145 ) | ( w17087 & ~w17148 ) | ( w17145 & ~w17148 ) ;
  assign w17150 = ( ~w12691 & w17148 ) | ( ~w12691 & w17149 ) | ( w17148 & w17149 ) ;
  assign w17151 = w16569 | w16574 ;
  assign w17152 = w17006 & ~w17151 ;
  assign w17153 = w16572 ^ w17152 ;
  assign w17154 = w17147 & ~w17150 ;
  assign w17155 = ( w17150 & w17153 ) | ( w17150 & ~w17154 ) | ( w17153 & ~w17154 ) ;
  assign w17156 = ( ~w12245 & w17154 ) | ( ~w12245 & w17155 ) | ( w17154 & w17155 ) ;
  assign w17157 = ( w17147 & w17150 ) | ( w17147 & w17153 ) | ( w17150 & w17153 ) ;
  assign w17158 = w17153 & w17157 ;
  assign w17159 = ( w17084 & w17156 ) | ( w17084 & w17158 ) | ( w17156 & w17158 ) ;
  assign w17160 = w17084 & w17159 ;
  assign w17161 = w17156 & ~w17158 ;
  assign w17162 = ( w17084 & w17158 ) | ( w17084 & ~w17161 ) | ( w17158 & ~w17161 ) ;
  assign w17163 = ( ~w11807 & w17161 ) | ( ~w11807 & w17162 ) | ( w17161 & w17162 ) ;
  assign w17164 = w16585 | w16590 ;
  assign w17165 = w17006 & ~w17164 ;
  assign w17166 = w16588 ^ w17165 ;
  assign w17167 = w17160 & ~w17163 ;
  assign w17168 = ( w17163 & w17166 ) | ( w17163 & ~w17167 ) | ( w17166 & ~w17167 ) ;
  assign w17169 = ( ~w11377 & w17167 ) | ( ~w11377 & w17168 ) | ( w17167 & w17168 ) ;
  assign w17170 = ( w17160 & w17163 ) | ( w17160 & w17166 ) | ( w17163 & w17166 ) ;
  assign w17171 = w17166 & w17170 ;
  assign w17172 = ( w17081 & w17169 ) | ( w17081 & w17171 ) | ( w17169 & w17171 ) ;
  assign w17173 = w17081 & w17172 ;
  assign w17174 = w17169 & ~w17171 ;
  assign w17175 = ( w17081 & w17171 ) | ( w17081 & ~w17174 ) | ( w17171 & ~w17174 ) ;
  assign w17176 = ( ~w10955 & w17174 ) | ( ~w10955 & w17175 ) | ( w17174 & w17175 ) ;
  assign w17177 = w16601 | w16606 ;
  assign w17178 = w17006 & ~w17177 ;
  assign w17179 = w16604 ^ w17178 ;
  assign w17180 = w17173 & ~w17176 ;
  assign w17181 = ( w17176 & w17179 ) | ( w17176 & ~w17180 ) | ( w17179 & ~w17180 ) ;
  assign w17182 = ( ~w10541 & w17180 ) | ( ~w10541 & w17181 ) | ( w17180 & w17181 ) ;
  assign w17183 = ( w17173 & w17176 ) | ( w17173 & w17179 ) | ( w17176 & w17179 ) ;
  assign w17184 = w17179 & w17183 ;
  assign w17185 = ( w17078 & w17182 ) | ( w17078 & w17184 ) | ( w17182 & w17184 ) ;
  assign w17186 = w17078 & w17185 ;
  assign w17187 = w17182 & ~w17184 ;
  assign w17188 = ( w17078 & w17184 ) | ( w17078 & ~w17187 ) | ( w17184 & ~w17187 ) ;
  assign w17189 = ( ~w10135 & w17187 ) | ( ~w10135 & w17188 ) | ( w17187 & w17188 ) ;
  assign w17190 = w16617 | w16622 ;
  assign w17191 = w17006 & ~w17190 ;
  assign w17192 = w16620 ^ w17191 ;
  assign w17193 = w17186 & ~w17189 ;
  assign w17194 = ( w17189 & w17192 ) | ( w17189 & ~w17193 ) | ( w17192 & ~w17193 ) ;
  assign w17195 = ( ~w9737 & w17193 ) | ( ~w9737 & w17194 ) | ( w17193 & w17194 ) ;
  assign w17196 = ( w17186 & w17189 ) | ( w17186 & w17192 ) | ( w17189 & w17192 ) ;
  assign w17197 = w17192 & w17196 ;
  assign w17198 = ( w17075 & w17195 ) | ( w17075 & w17197 ) | ( w17195 & w17197 ) ;
  assign w17199 = w17075 & w17198 ;
  assign w17200 = w17195 & ~w17197 ;
  assign w17201 = ( w17075 & w17197 ) | ( w17075 & ~w17200 ) | ( w17197 & ~w17200 ) ;
  assign w17202 = ( ~w9347 & w17200 ) | ( ~w9347 & w17201 ) | ( w17200 & w17201 ) ;
  assign w17203 = w16633 | w16638 ;
  assign w17204 = w17006 & ~w17203 ;
  assign w17205 = w16636 ^ w17204 ;
  assign w17206 = w17199 & ~w17202 ;
  assign w17207 = ( w17202 & w17205 ) | ( w17202 & ~w17206 ) | ( w17205 & ~w17206 ) ;
  assign w17208 = ( ~w8965 & w17206 ) | ( ~w8965 & w17207 ) | ( w17206 & w17207 ) ;
  assign w17209 = ( w17199 & w17202 ) | ( w17199 & w17205 ) | ( w17202 & w17205 ) ;
  assign w17210 = w17205 & w17209 ;
  assign w17211 = ( w17072 & w17208 ) | ( w17072 & w17210 ) | ( w17208 & w17210 ) ;
  assign w17212 = w17072 & w17211 ;
  assign w17213 = w17208 & ~w17210 ;
  assign w17214 = ( w17072 & w17210 ) | ( w17072 & ~w17213 ) | ( w17210 & ~w17213 ) ;
  assign w17215 = ( ~w8591 & w17213 ) | ( ~w8591 & w17214 ) | ( w17213 & w17214 ) ;
  assign w17216 = w16649 | w16654 ;
  assign w17217 = w17006 & ~w17216 ;
  assign w17218 = w16652 ^ w17217 ;
  assign w17219 = w17212 & ~w17215 ;
  assign w17220 = ( w17215 & w17218 ) | ( w17215 & ~w17219 ) | ( w17218 & ~w17219 ) ;
  assign w17221 = ( ~w8225 & w17219 ) | ( ~w8225 & w17220 ) | ( w17219 & w17220 ) ;
  assign w17222 = ( w17212 & w17215 ) | ( w17212 & w17218 ) | ( w17215 & w17218 ) ;
  assign w17223 = w17218 & w17222 ;
  assign w17224 = ( w17069 & w17221 ) | ( w17069 & w17223 ) | ( w17221 & w17223 ) ;
  assign w17225 = w17069 & w17224 ;
  assign w17226 = w17221 & ~w17223 ;
  assign w17227 = ( w17069 & w17223 ) | ( w17069 & ~w17226 ) | ( w17223 & ~w17226 ) ;
  assign w17228 = ( ~w7867 & w17226 ) | ( ~w7867 & w17227 ) | ( w17226 & w17227 ) ;
  assign w17229 = w16665 | w16670 ;
  assign w17230 = w17006 & ~w17229 ;
  assign w17231 = w16668 ^ w17230 ;
  assign w17232 = w17225 & ~w17228 ;
  assign w17233 = ( w17228 & w17231 ) | ( w17228 & ~w17232 ) | ( w17231 & ~w17232 ) ;
  assign w17234 = ( ~w7517 & w17232 ) | ( ~w7517 & w17233 ) | ( w17232 & w17233 ) ;
  assign w17235 = ( w17225 & w17228 ) | ( w17225 & w17231 ) | ( w17228 & w17231 ) ;
  assign w17236 = w17231 & w17235 ;
  assign w17237 = ( w17066 & w17234 ) | ( w17066 & w17236 ) | ( w17234 & w17236 ) ;
  assign w17238 = w17066 & w17237 ;
  assign w17239 = w17234 & ~w17236 ;
  assign w17240 = ( w17066 & w17236 ) | ( w17066 & ~w17239 ) | ( w17236 & ~w17239 ) ;
  assign w17241 = ( ~w7175 & w17239 ) | ( ~w7175 & w17240 ) | ( w17239 & w17240 ) ;
  assign w17242 = w16681 | w16686 ;
  assign w17243 = w17006 & ~w17242 ;
  assign w17244 = w16684 ^ w17243 ;
  assign w17245 = w17238 & ~w17241 ;
  assign w17246 = ( w17241 & w17244 ) | ( w17241 & ~w17245 ) | ( w17244 & ~w17245 ) ;
  assign w17247 = ( ~w6841 & w17245 ) | ( ~w6841 & w17246 ) | ( w17245 & w17246 ) ;
  assign w17248 = ( w17238 & w17241 ) | ( w17238 & w17244 ) | ( w17241 & w17244 ) ;
  assign w17249 = w17244 & w17248 ;
  assign w17250 = ( w17063 & w17247 ) | ( w17063 & w17249 ) | ( w17247 & w17249 ) ;
  assign w17251 = w17063 & w17250 ;
  assign w17252 = w17247 & ~w17249 ;
  assign w17253 = ( w17063 & w17249 ) | ( w17063 & ~w17252 ) | ( w17249 & ~w17252 ) ;
  assign w17254 = ( ~w6515 & w17252 ) | ( ~w6515 & w17253 ) | ( w17252 & w17253 ) ;
  assign w17255 = w16697 | w16702 ;
  assign w17256 = w17006 & ~w17255 ;
  assign w17257 = w16700 ^ w17256 ;
  assign w17258 = w17251 & ~w17254 ;
  assign w17259 = ( w17254 & w17257 ) | ( w17254 & ~w17258 ) | ( w17257 & ~w17258 ) ;
  assign w17260 = ( ~w6197 & w17258 ) | ( ~w6197 & w17259 ) | ( w17258 & w17259 ) ;
  assign w17261 = ( w17251 & w17254 ) | ( w17251 & w17257 ) | ( w17254 & w17257 ) ;
  assign w17262 = w17257 & w17261 ;
  assign w17263 = ( w17060 & w17260 ) | ( w17060 & w17262 ) | ( w17260 & w17262 ) ;
  assign w17264 = w17060 & w17263 ;
  assign w17265 = w17260 & ~w17262 ;
  assign w17266 = ( w17060 & w17262 ) | ( w17060 & ~w17265 ) | ( w17262 & ~w17265 ) ;
  assign w17267 = ( ~w5887 & w17265 ) | ( ~w5887 & w17266 ) | ( w17265 & w17266 ) ;
  assign w17268 = w16713 | w16718 ;
  assign w17269 = w17006 & ~w17268 ;
  assign w17270 = w16716 ^ w17269 ;
  assign w17271 = w17264 & ~w17267 ;
  assign w17272 = ( w17267 & w17270 ) | ( w17267 & ~w17271 ) | ( w17270 & ~w17271 ) ;
  assign w17273 = ( ~w5585 & w17271 ) | ( ~w5585 & w17272 ) | ( w17271 & w17272 ) ;
  assign w17274 = ( w17264 & w17267 ) | ( w17264 & w17270 ) | ( w17267 & w17270 ) ;
  assign w17275 = w17270 & w17274 ;
  assign w17276 = ( w17057 & w17273 ) | ( w17057 & w17275 ) | ( w17273 & w17275 ) ;
  assign w17277 = w17057 & w17276 ;
  assign w17278 = w17273 & ~w17275 ;
  assign w17279 = ( w17057 & w17275 ) | ( w17057 & ~w17278 ) | ( w17275 & ~w17278 ) ;
  assign w17280 = ( ~w5291 & w17278 ) | ( ~w5291 & w17279 ) | ( w17278 & w17279 ) ;
  assign w17281 = w16729 | w16734 ;
  assign w17282 = w17006 & ~w17281 ;
  assign w17283 = w16732 ^ w17282 ;
  assign w17284 = w17277 & ~w17280 ;
  assign w17285 = ( w17280 & w17283 ) | ( w17280 & ~w17284 ) | ( w17283 & ~w17284 ) ;
  assign w17286 = ( ~w5005 & w17284 ) | ( ~w5005 & w17285 ) | ( w17284 & w17285 ) ;
  assign w17287 = ( w17277 & w17280 ) | ( w17277 & w17283 ) | ( w17280 & w17283 ) ;
  assign w17288 = w17283 & w17287 ;
  assign w17289 = ( w17054 & w17286 ) | ( w17054 & w17288 ) | ( w17286 & w17288 ) ;
  assign w17290 = w17054 & w17289 ;
  assign w17291 = w17286 & ~w17288 ;
  assign w17292 = ( w17054 & w17288 ) | ( w17054 & ~w17291 ) | ( w17288 & ~w17291 ) ;
  assign w17293 = ( ~w4727 & w17291 ) | ( ~w4727 & w17292 ) | ( w17291 & w17292 ) ;
  assign w17294 = w16745 | w16750 ;
  assign w17295 = w17006 & ~w17294 ;
  assign w17296 = w16748 ^ w17295 ;
  assign w17297 = w17290 & ~w17293 ;
  assign w17298 = ( w17293 & w17296 ) | ( w17293 & ~w17297 ) | ( w17296 & ~w17297 ) ;
  assign w17299 = ( ~w4457 & w17297 ) | ( ~w4457 & w17298 ) | ( w17297 & w17298 ) ;
  assign w17300 = ( w17290 & w17293 ) | ( w17290 & w17296 ) | ( w17293 & w17296 ) ;
  assign w17301 = w17296 & w17300 ;
  assign w17302 = ( w17051 & w17299 ) | ( w17051 & w17301 ) | ( w17299 & w17301 ) ;
  assign w17303 = w17051 & w17302 ;
  assign w17304 = w17299 & ~w17301 ;
  assign w17305 = ( w17051 & w17301 ) | ( w17051 & ~w17304 ) | ( w17301 & ~w17304 ) ;
  assign w17306 = ( ~w4195 & w17304 ) | ( ~w4195 & w17305 ) | ( w17304 & w17305 ) ;
  assign w17307 = w16761 | w16766 ;
  assign w17308 = w17006 & ~w17307 ;
  assign w17309 = w16764 ^ w17308 ;
  assign w17310 = w17303 & ~w17306 ;
  assign w17311 = ( w17306 & w17309 ) | ( w17306 & ~w17310 ) | ( w17309 & ~w17310 ) ;
  assign w17312 = ( ~w3941 & w17310 ) | ( ~w3941 & w17311 ) | ( w17310 & w17311 ) ;
  assign w17313 = ( w17303 & w17306 ) | ( w17303 & w17309 ) | ( w17306 & w17309 ) ;
  assign w17314 = w17309 & w17313 ;
  assign w17315 = ( w17048 & w17312 ) | ( w17048 & w17314 ) | ( w17312 & w17314 ) ;
  assign w17316 = w17048 & w17315 ;
  assign w17317 = w17312 & ~w17314 ;
  assign w17318 = ( w17048 & w17314 ) | ( w17048 & ~w17317 ) | ( w17314 & ~w17317 ) ;
  assign w17319 = ( ~w3695 & w17317 ) | ( ~w3695 & w17318 ) | ( w17317 & w17318 ) ;
  assign w17320 = w16777 | w16782 ;
  assign w17321 = w17006 & ~w17320 ;
  assign w17322 = w16780 ^ w17321 ;
  assign w17323 = w17316 & ~w17319 ;
  assign w17324 = ( w17319 & w17322 ) | ( w17319 & ~w17323 ) | ( w17322 & ~w17323 ) ;
  assign w17325 = ( ~w3457 & w17323 ) | ( ~w3457 & w17324 ) | ( w17323 & w17324 ) ;
  assign w17326 = ( w17316 & w17319 ) | ( w17316 & w17322 ) | ( w17319 & w17322 ) ;
  assign w17327 = w17322 & w17326 ;
  assign w17328 = ( w17045 & w17325 ) | ( w17045 & w17327 ) | ( w17325 & w17327 ) ;
  assign w17329 = w17045 & w17328 ;
  assign w17330 = w17325 & ~w17327 ;
  assign w17331 = ( w17045 & w17327 ) | ( w17045 & ~w17330 ) | ( w17327 & ~w17330 ) ;
  assign w17332 = ( ~w3227 & w17330 ) | ( ~w3227 & w17331 ) | ( w17330 & w17331 ) ;
  assign w17333 = w16793 | w16798 ;
  assign w17334 = w17006 & ~w17333 ;
  assign w17335 = w16796 ^ w17334 ;
  assign w17336 = w17329 & ~w17332 ;
  assign w17337 = ( w17332 & w17335 ) | ( w17332 & ~w17336 ) | ( w17335 & ~w17336 ) ;
  assign w17338 = ( ~w3005 & w17336 ) | ( ~w3005 & w17337 ) | ( w17336 & w17337 ) ;
  assign w17339 = ( w17329 & w17332 ) | ( w17329 & w17335 ) | ( w17332 & w17335 ) ;
  assign w17340 = w17335 & w17339 ;
  assign w17341 = ( w17042 & w17338 ) | ( w17042 & w17340 ) | ( w17338 & w17340 ) ;
  assign w17342 = w17042 & w17341 ;
  assign w17343 = w17338 & ~w17340 ;
  assign w17344 = ( w17042 & w17340 ) | ( w17042 & ~w17343 ) | ( w17340 & ~w17343 ) ;
  assign w17345 = ( ~w2791 & w17343 ) | ( ~w2791 & w17344 ) | ( w17343 & w17344 ) ;
  assign w17346 = w16809 | w16814 ;
  assign w17347 = w17006 & ~w17346 ;
  assign w17348 = w16812 ^ w17347 ;
  assign w17349 = w17342 & ~w17345 ;
  assign w17350 = ( w17345 & w17348 ) | ( w17345 & ~w17349 ) | ( w17348 & ~w17349 ) ;
  assign w17351 = ( ~w2585 & w17349 ) | ( ~w2585 & w17350 ) | ( w17349 & w17350 ) ;
  assign w17352 = ( w17342 & w17345 ) | ( w17342 & w17348 ) | ( w17345 & w17348 ) ;
  assign w17353 = w17348 & w17352 ;
  assign w17354 = ( w17039 & w17351 ) | ( w17039 & w17353 ) | ( w17351 & w17353 ) ;
  assign w17355 = w17039 & w17354 ;
  assign w17356 = w17351 & ~w17353 ;
  assign w17357 = ( w17039 & w17353 ) | ( w17039 & ~w17356 ) | ( w17353 & ~w17356 ) ;
  assign w17358 = ( ~w2387 & w17356 ) | ( ~w2387 & w17357 ) | ( w17356 & w17357 ) ;
  assign w17359 = w16825 | w16830 ;
  assign w17360 = w17006 & ~w17359 ;
  assign w17361 = w16828 ^ w17360 ;
  assign w17362 = w17355 & ~w17358 ;
  assign w17363 = ( w17358 & w17361 ) | ( w17358 & ~w17362 ) | ( w17361 & ~w17362 ) ;
  assign w17364 = ( ~w2197 & w17362 ) | ( ~w2197 & w17363 ) | ( w17362 & w17363 ) ;
  assign w17365 = ( w17355 & w17358 ) | ( w17355 & w17361 ) | ( w17358 & w17361 ) ;
  assign w17366 = w17361 & w17365 ;
  assign w17367 = ( w17036 & w17364 ) | ( w17036 & w17366 ) | ( w17364 & w17366 ) ;
  assign w17368 = w17036 & w17367 ;
  assign w17369 = w17364 & ~w17366 ;
  assign w17370 = ( w17036 & w17366 ) | ( w17036 & ~w17369 ) | ( w17366 & ~w17369 ) ;
  assign w17371 = ( ~w2015 & w17369 ) | ( ~w2015 & w17370 ) | ( w17369 & w17370 ) ;
  assign w17372 = w16841 | w16846 ;
  assign w17373 = w17006 & ~w17372 ;
  assign w17374 = w16844 ^ w17373 ;
  assign w17375 = w17368 & ~w17371 ;
  assign w17376 = ( w17371 & w17374 ) | ( w17371 & ~w17375 ) | ( w17374 & ~w17375 ) ;
  assign w17377 = ( ~w1841 & w17375 ) | ( ~w1841 & w17376 ) | ( w17375 & w17376 ) ;
  assign w17378 = ( w17368 & w17371 ) | ( w17368 & w17374 ) | ( w17371 & w17374 ) ;
  assign w17379 = w17374 & w17378 ;
  assign w17380 = ( w17033 & w17377 ) | ( w17033 & w17379 ) | ( w17377 & w17379 ) ;
  assign w17381 = w17033 & w17380 ;
  assign w17382 = w17377 & ~w17379 ;
  assign w17383 = ( w17033 & w17379 ) | ( w17033 & ~w17382 ) | ( w17379 & ~w17382 ) ;
  assign w17384 = ( ~w1675 & w17382 ) | ( ~w1675 & w17383 ) | ( w17382 & w17383 ) ;
  assign w17385 = w16857 | w16862 ;
  assign w17386 = w17006 & ~w17385 ;
  assign w17387 = w16860 ^ w17386 ;
  assign w17388 = w17381 & ~w17384 ;
  assign w17389 = ( w17384 & w17387 ) | ( w17384 & ~w17388 ) | ( w17387 & ~w17388 ) ;
  assign w17390 = ( ~w1517 & w17388 ) | ( ~w1517 & w17389 ) | ( w17388 & w17389 ) ;
  assign w17391 = ( w17381 & w17384 ) | ( w17381 & w17387 ) | ( w17384 & w17387 ) ;
  assign w17392 = w17387 & w17391 ;
  assign w17393 = ( w17030 & w17390 ) | ( w17030 & w17392 ) | ( w17390 & w17392 ) ;
  assign w17394 = w17030 & w17393 ;
  assign w17395 = w17390 & ~w17392 ;
  assign w17396 = ( w17030 & w17392 ) | ( w17030 & ~w17395 ) | ( w17392 & ~w17395 ) ;
  assign w17397 = ( ~w1367 & w17395 ) | ( ~w1367 & w17396 ) | ( w17395 & w17396 ) ;
  assign w17398 = w16873 | w16878 ;
  assign w17399 = w17006 & ~w17398 ;
  assign w17400 = w16876 ^ w17399 ;
  assign w17401 = w17394 & ~w17397 ;
  assign w17402 = ( w17397 & w17400 ) | ( w17397 & ~w17401 ) | ( w17400 & ~w17401 ) ;
  assign w17403 = ( ~w1225 & w17401 ) | ( ~w1225 & w17402 ) | ( w17401 & w17402 ) ;
  assign w17404 = ( w17394 & w17397 ) | ( w17394 & w17400 ) | ( w17397 & w17400 ) ;
  assign w17405 = w17400 & w17404 ;
  assign w17406 = ( w17027 & w17403 ) | ( w17027 & w17405 ) | ( w17403 & w17405 ) ;
  assign w17407 = w17027 & w17406 ;
  assign w17408 = w17403 & ~w17405 ;
  assign w17409 = ( w17027 & w17405 ) | ( w17027 & ~w17408 ) | ( w17405 & ~w17408 ) ;
  assign w17410 = ( ~w1091 & w17408 ) | ( ~w1091 & w17409 ) | ( w17408 & w17409 ) ;
  assign w17411 = w16889 | w16894 ;
  assign w17412 = w17006 & ~w17411 ;
  assign w17413 = w16892 ^ w17412 ;
  assign w17414 = w17407 & ~w17410 ;
  assign w17415 = ( w17410 & w17413 ) | ( w17410 & ~w17414 ) | ( w17413 & ~w17414 ) ;
  assign w17416 = ( ~w965 & w17414 ) | ( ~w965 & w17415 ) | ( w17414 & w17415 ) ;
  assign w17417 = ( w17407 & w17410 ) | ( w17407 & w17413 ) | ( w17410 & w17413 ) ;
  assign w17418 = w17413 & w17417 ;
  assign w17419 = ( w17024 & w17416 ) | ( w17024 & w17418 ) | ( w17416 & w17418 ) ;
  assign w17420 = w17024 & w17419 ;
  assign w17421 = w17416 & ~w17418 ;
  assign w17422 = ( w17024 & w17418 ) | ( w17024 & ~w17421 ) | ( w17418 & ~w17421 ) ;
  assign w17423 = ( ~w847 & w17421 ) | ( ~w847 & w17422 ) | ( w17421 & w17422 ) ;
  assign w17424 = w16905 | w16910 ;
  assign w17425 = w17006 & ~w17424 ;
  assign w17426 = w16908 ^ w17425 ;
  assign w17427 = w17420 & ~w17423 ;
  assign w17428 = ( w17423 & w17426 ) | ( w17423 & ~w17427 ) | ( w17426 & ~w17427 ) ;
  assign w17429 = ( ~w737 & w17427 ) | ( ~w737 & w17428 ) | ( w17427 & w17428 ) ;
  assign w17430 = ( w17420 & w17423 ) | ( w17420 & w17426 ) | ( w17423 & w17426 ) ;
  assign w17431 = w17426 & w17430 ;
  assign w17432 = ( w17021 & w17429 ) | ( w17021 & w17431 ) | ( w17429 & w17431 ) ;
  assign w17433 = w17021 & w17432 ;
  assign w17434 = w17429 & ~w17431 ;
  assign w17435 = ( w17021 & w17431 ) | ( w17021 & ~w17434 ) | ( w17431 & ~w17434 ) ;
  assign w17436 = ( ~w635 & w17434 ) | ( ~w635 & w17435 ) | ( w17434 & w17435 ) ;
  assign w17437 = w16921 | w16926 ;
  assign w17438 = w17006 & ~w17437 ;
  assign w17439 = w16924 ^ w17438 ;
  assign w17440 = w17433 & ~w17436 ;
  assign w17441 = ( w17436 & w17439 ) | ( w17436 & ~w17440 ) | ( w17439 & ~w17440 ) ;
  assign w17442 = ( ~w541 & w17440 ) | ( ~w541 & w17441 ) | ( w17440 & w17441 ) ;
  assign w17443 = ( w17433 & w17436 ) | ( w17433 & w17439 ) | ( w17436 & w17439 ) ;
  assign w17444 = w17439 & w17443 ;
  assign w17445 = ( w17018 & w17442 ) | ( w17018 & w17444 ) | ( w17442 & w17444 ) ;
  assign w17446 = w17018 & w17445 ;
  assign w17447 = w17442 & ~w17444 ;
  assign w17448 = ( w17018 & w17444 ) | ( w17018 & ~w17447 ) | ( w17444 & ~w17447 ) ;
  assign w17449 = ( ~w455 & w17447 ) | ( ~w455 & w17448 ) | ( w17447 & w17448 ) ;
  assign w17450 = w16937 | w16942 ;
  assign w17451 = w17006 & ~w17450 ;
  assign w17452 = w16940 ^ w17451 ;
  assign w17453 = w17446 & ~w17449 ;
  assign w17454 = ( w17449 & w17452 ) | ( w17449 & ~w17453 ) | ( w17452 & ~w17453 ) ;
  assign w17455 = ( ~w377 & w17453 ) | ( ~w377 & w17454 ) | ( w17453 & w17454 ) ;
  assign w17456 = ( w17446 & w17449 ) | ( w17446 & w17452 ) | ( w17449 & w17452 ) ;
  assign w17457 = w17452 & w17456 ;
  assign w17458 = w16953 | w16958 ;
  assign w17459 = w17006 & ~w17458 ;
  assign w17460 = w16956 ^ w17459 ;
  assign w17461 = ~w246 & w17460 ;
  assign w17462 = ( w17455 & w17457 ) | ( w17455 & ~w17461 ) | ( w17457 & ~w17461 ) ;
  assign w17463 = ( ~w307 & w17015 ) | ( ~w307 & w17462 ) | ( w17015 & w17462 ) ;
  assign w17464 = ( ~w246 & w17461 ) | ( ~w246 & w17463 ) | ( w17461 & w17463 ) ;
  assign w17465 = w17455 | w17457 ;
  assign w17466 = ( ~w307 & w17015 ) | ( ~w307 & w17465 ) | ( w17015 & w17465 ) ;
  assign w17467 = w17460 & w17466 ;
  assign w17468 = w16969 | w16974 ;
  assign w17469 = w17006 & ~w17468 ;
  assign w17470 = w16972 ^ w17469 ;
  assign w17471 = ~w145 & w17470 ;
  assign w17472 = ( w17464 & w17467 ) | ( w17464 & ~w17471 ) | ( w17467 & ~w17471 ) ;
  assign w17473 = ( ~w185 & w17012 ) | ( ~w185 & w17472 ) | ( w17012 & w17472 ) ;
  assign w17474 = ( ~w145 & w17471 ) | ( ~w145 & w17473 ) | ( w17471 & w17473 ) ;
  assign w17475 = w17464 | w17467 ;
  assign w17476 = ( ~w185 & w17012 ) | ( ~w185 & w17475 ) | ( w17012 & w17475 ) ;
  assign w17477 = w17470 & w17476 ;
  assign w17478 = ( w17009 & w17474 ) | ( w17009 & w17477 ) | ( w17474 & w17477 ) ;
  assign w17479 = w17009 & w17478 ;
  assign w17480 = w17474 & ~w17477 ;
  assign w17481 = ( w17009 & w17477 ) | ( w17009 & ~w17480 ) | ( w17477 & ~w17480 ) ;
  assign w17482 = ( ~w132 & w17480 ) | ( ~w132 & w17481 ) | ( w17480 & w17481 ) ;
  assign w17483 = w16982 | w16987 ;
  assign w17484 = w17006 & ~w17483 ;
  assign w17485 = w16985 ^ w17484 ;
  assign w17486 = w16989 | w17006 ;
  assign w17487 = ( w16989 & w16992 ) | ( w16989 & w17486 ) | ( w16992 & w17486 ) ;
  assign w17488 = ( w17000 & w17486 ) | ( w17000 & ~w17487 ) | ( w17486 & ~w17487 ) ;
  assign w17489 = ( w129 & w16989 ) | ( w129 & w16992 ) | ( w16989 & w16992 ) ;
  assign w17490 = ( w16992 & ~w17006 ) | ( w16992 & w17489 ) | ( ~w17006 & w17489 ) ;
  assign w17491 = w16989 & w17490 ;
  assign w17492 = w17489 ^ w17491 ;
  assign w17493 = ~w129 & w17488 ;
  assign w17494 = ( w17479 & w17482 ) | ( w17479 & ~w17492 ) | ( w17482 & ~w17492 ) ;
  assign w17495 = ( ~w129 & w17485 ) | ( ~w129 & w17494 ) | ( w17485 & w17494 ) ;
  assign w17496 = w17492 | w17495 ;
  assign w17497 = w17493 | w17496 ;
  assign \po00 = w17497 ;
  assign \po01 = w17006 ;
  assign \po02 = w16501 ;
  assign \po03 = w16004 ;
  assign \po04 = w15515 ;
  assign \po05 = w15032 ;
  assign \po06 = w14555 ;
  assign \po07 = w14077 ;
  assign \po08 = w13607 ;
  assign \po09 = w13145 ;
  assign \po10 = w12691 ;
  assign \po11 = w12245 ;
  assign \po12 = w11807 ;
  assign \po13 = w11377 ;
  assign \po14 = w10955 ;
  assign \po15 = w10541 ;
  assign \po16 = w10135 ;
  assign \po17 = w9737 ;
  assign \po18 = w9347 ;
  assign \po19 = w8965 ;
  assign \po20 = w8591 ;
  assign \po21 = w8225 ;
  assign \po22 = w7867 ;
  assign \po23 = w7517 ;
  assign \po24 = w7175 ;
  assign \po25 = w6841 ;
  assign \po26 = w6515 ;
  assign \po27 = w6197 ;
  assign \po28 = w5887 ;
  assign \po29 = w5585 ;
  assign \po30 = w5291 ;
  assign \po31 = w5005 ;
  assign \po32 = w4727 ;
  assign \po33 = w4457 ;
  assign \po34 = w4195 ;
  assign \po35 = w3941 ;
  assign \po36 = w3695 ;
  assign \po37 = w3457 ;
  assign \po38 = w3227 ;
  assign \po39 = w3005 ;
  assign \po40 = w2791 ;
  assign \po41 = w2585 ;
  assign \po42 = w2387 ;
  assign \po43 = w2197 ;
  assign \po44 = w2015 ;
  assign \po45 = w1841 ;
  assign \po46 = w1675 ;
  assign \po47 = w1517 ;
  assign \po48 = w1367 ;
  assign \po49 = w1225 ;
  assign \po50 = w1091 ;
  assign \po51 = w965 ;
  assign \po52 = w847 ;
  assign \po53 = w737 ;
  assign \po54 = w635 ;
  assign \po55 = w541 ;
  assign \po56 = w455 ;
  assign \po57 = w377 ;
  assign \po58 = w307 ;
  assign \po59 = w246 ;
  assign \po60 = w185 ;
  assign \po61 = w145 ;
  assign \po62 = w132 ;
  assign \po63 = w129 ;
endmodule
