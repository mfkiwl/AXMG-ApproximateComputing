module square( \pi00 , \pi01 , \pi02 , \pi03 , \pi04 , \pi05 , \pi06 , \pi07 , \pi08 , \pi09 , \pi10 , \pi11 , \pi12 , \pi13 , \pi14 , \pi15 , \pi16 , \pi17 , \pi18 , \pi19 , \pi20 , \pi21 , \pi22 , \pi23 , \pi24 , \pi25 , \pi26 , \pi27 , \pi28 , \pi29 , \pi30 , \pi31 , \pi32 , \pi33 , \pi34 , \pi35 , \pi36 , \pi37 , \pi38 , \pi39 , \pi40 , \pi41 , \pi42 , \pi43 , \pi44 , \pi45 , \pi46 , \pi47 , \pi48 , \pi49 , \pi50 , \pi51 , \pi52 , \pi53 , \pi54 , \pi55 , \pi56 , \pi57 , \pi58 , \pi59 , \pi60 , \pi61 , \pi62 , \pi63 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 );
  input \pi00 , \pi01 , \pi02 , \pi03 , \pi04 , \pi05 , \pi06 , \pi07 , \pi08 , \pi09 , \pi10 , \pi11 , \pi12 , \pi13 , \pi14 , \pi15 , \pi16 , \pi17 , \pi18 , \pi19 , \pi20 , \pi21 , \pi22 , \pi23 , \pi24 , \pi25 , \pi26 , \pi27 , \pi28 , \pi29 , \pi30 , \pi31 , \pi32 , \pi33 , \pi34 , \pi35 , \pi36 , \pi37 , \pi38 , \pi39 , \pi40 , \pi41 , \pi42 , \pi43 , \pi44 , \pi45 , \pi46 , \pi47 , \pi48 , \pi49 , \pi50 , \pi51 , \pi52 , \pi53 , \pi54 , \pi55 , \pi56 , \pi57 , \pi58 , \pi59 , \pi60 , \pi61 , \pi62 , \pi63 ;
  output \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 ;
  wire zero , w65 , w66 , w67 , w68 , w69 , w70 , w71 , w72 , w73 , w74 , w75 , w76 , w77 , w78 , w79 , w80 , w81 , w82 , w83 , w84 , w85 , w86 , w87 , w88 , w89 , w90 , w91 , w92 , w93 , w94 , w95 , w96 , w97 , w98 , w99 , w100 , w101 , w102 , w103 , w104 , w105 , w106 , w107 , w108 , w109 , w110 , w111 , w112 , w113 , w114 , w115 , w116 , w117 , w118 , w119 , w120 , w121 , w122 , w123 , w124 , w125 , w126 , w127 , w128 , w129 , w130 , w131 , w132 , w133 , w134 , w135 , w136 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w146 , w147 , w148 , w149 , w150 , w151 , w152 , w153 , w154 , w155 , w156 , w157 , w158 , w159 , w160 , w161 , w162 , w163 , w164 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w174 , w175 , w176 , w177 , w178 , w179 , w180 , w181 , w182 , w183 , w184 , w185 , w186 , w187 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w203 , w204 , w205 , w206 , w207 , w208 , w209 , w210 , w211 , w212 , w213 , w214 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w224 , w225 , w226 , w227 , w228 , w229 , w230 , w231 , w232 , w233 , w234 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w250 , w251 , w252 , w253 , w254 , w255 , w256 , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 , w2495 , w2496 , w2497 , w2498 , w2499 , w2500 , w2501 , w2502 , w2503 , w2504 , w2505 , w2506 , w2507 , w2508 , w2509 , w2510 , w2511 , w2512 , w2513 , w2514 , w2515 , w2516 , w2517 , w2518 , w2519 , w2520 , w2521 , w2522 , w2523 , w2524 , w2525 , w2526 , w2527 , w2528 , w2529 , w2530 , w2531 , w2532 , w2533 , w2534 , w2535 , w2536 , w2537 , w2538 , w2539 , w2540 , w2541 , w2542 , w2543 , w2544 , w2545 , w2546 , w2547 , w2548 , w2549 , w2550 , w2551 , w2552 , w2553 , w2554 , w2555 , w2556 , w2557 , w2558 , w2559 , w2560 , w2561 , w2562 , w2563 , w2564 , w2565 , w2566 , w2567 , w2568 , w2569 , w2570 , w2571 , w2572 , w2573 , w2574 , w2575 , w2576 , w2577 , w2578 , w2579 , w2580 , w2581 , w2582 , w2583 , w2584 , w2585 , w2586 , w2587 , w2588 , w2589 , w2590 , w2591 , w2592 , w2593 , w2594 , w2595 , w2596 , w2597 , w2598 , w2599 , w2600 , w2601 , w2602 , w2603 , w2604 , w2605 , w2606 , w2607 , w2608 , w2609 , w2610 , w2611 , w2612 , w2613 , w2614 , w2615 , w2616 , w2617 , w2618 , w2619 , w2620 , w2621 , w2622 , w2623 , w2624 , w2625 , w2626 , w2627 , w2628 , w2629 , w2630 , w2631 , w2632 , w2633 , w2634 , w2635 , w2636 , w2637 , w2638 , w2639 , w2640 , w2641 , w2642 , w2643 , w2644 , w2645 , w2646 , w2647 , w2648 , w2649 , w2650 , w2651 , w2652 , w2653 , w2654 , w2655 , w2656 , w2657 , w2658 , w2659 , w2660 , w2661 , w2662 , w2663 , w2664 , w2665 , w2666 , w2667 , w2668 , w2669 , w2670 , w2671 , w2672 , w2673 , w2674 , w2675 , w2676 , w2677 , w2678 , w2679 , w2680 , w2681 , w2682 , w2683 , w2684 , w2685 , w2686 , w2687 , w2688 , w2689 , w2690 , w2691 , w2692 , w2693 , w2694 , w2695 , w2696 , w2697 , w2698 , w2699 , w2700 , w2701 , w2702 , w2703 , w2704 , w2705 , w2706 , w2707 , w2708 , w2709 , w2710 , w2711 , w2712 , w2713 , w2714 , w2715 , w2716 , w2717 , w2718 , w2719 , w2720 , w2721 , w2722 , w2723 , w2724 , w2725 , w2726 , w2727 , w2728 , w2729 , w2730 , w2731 , w2732 , w2733 , w2734 , w2735 , w2736 , w2737 , w2738 , w2739 , w2740 , w2741 , w2742 , w2743 , w2744 , w2745 , w2746 , w2747 , w2748 , w2749 , w2750 , w2751 , w2752 , w2753 , w2754 , w2755 , w2756 , w2757 , w2758 , w2759 , w2760 , w2761 , w2762 , w2763 , w2764 , w2765 , w2766 , w2767 , w2768 , w2769 , w2770 , w2771 , w2772 , w2773 , w2774 , w2775 , w2776 , w2777 , w2778 , w2779 , w2780 , w2781 , w2782 , w2783 , w2784 , w2785 , w2786 , w2787 , w2788 , w2789 , w2790 , w2791 , w2792 , w2793 , w2794 , w2795 , w2796 , w2797 , w2798 , w2799 , w2800 , w2801 , w2802 , w2803 , w2804 , w2805 , w2806 , w2807 , w2808 , w2809 , w2810 , w2811 , w2812 , w2813 , w2814 , w2815 , w2816 , w2817 , w2818 , w2819 , w2820 , w2821 , w2822 , w2823 , w2824 , w2825 , w2826 , w2827 , w2828 , w2829 , w2830 , w2831 , w2832 , w2833 , w2834 , w2835 , w2836 , w2837 , w2838 , w2839 , w2840 , w2841 , w2842 , w2843 , w2844 , w2845 , w2846 , w2847 , w2848 , w2849 , w2850 , w2851 , w2852 , w2853 , w2854 , w2855 , w2856 , w2857 , w2858 , w2859 , w2860 , w2861 , w2862 , w2863 , w2864 , w2865 , w2866 , w2867 , w2868 , w2869 , w2870 , w2871 , w2872 , w2873 , w2874 , w2875 , w2876 , w2877 , w2878 , w2879 , w2880 , w2881 , w2882 , w2883 , w2884 , w2885 , w2886 , w2887 , w2888 , w2889 , w2890 , w2891 , w2892 , w2893 , w2894 , w2895 , w2896 , w2897 , w2898 , w2899 , w2900 , w2901 , w2902 , w2903 , w2904 , w2905 , w2906 , w2907 , w2908 , w2909 , w2910 , w2911 , w2912 , w2913 , w2914 , w2915 , w2916 , w2917 , w2918 , w2919 , w2920 , w2921 , w2922 , w2923 , w2924 , w2925 , w2926 , w2927 , w2928 , w2929 , w2930 , w2931 , w2932 , w2933 , w2934 , w2935 , w2936 , w2937 , w2938 , w2939 , w2940 , w2941 , w2942 , w2943 , w2944 , w2945 , w2946 , w2947 , w2948 , w2949 , w2950 , w2951 , w2952 , w2953 , w2954 , w2955 , w2956 , w2957 , w2958 , w2959 , w2960 , w2961 , w2962 , w2963 , w2964 , w2965 , w2966 , w2967 , w2968 , w2969 , w2970 , w2971 , w2972 , w2973 , w2974 , w2975 , w2976 , w2977 , w2978 , w2979 , w2980 , w2981 , w2982 , w2983 , w2984 , w2985 , w2986 , w2987 , w2988 , w2989 , w2990 , w2991 , w2992 , w2993 , w2994 , w2995 , w2996 , w2997 , w2998 , w2999 , w3000 , w3001 , w3002 , w3003 , w3004 , w3005 , w3006 , w3007 , w3008 , w3009 , w3010 , w3011 , w3012 , w3013 , w3014 , w3015 , w3016 , w3017 , w3018 , w3019 , w3020 , w3021 , w3022 , w3023 , w3024 , w3025 , w3026 , w3027 , w3028 , w3029 , w3030 , w3031 , w3032 , w3033 , w3034 , w3035 , w3036 , w3037 , w3038 , w3039 , w3040 , w3041 , w3042 , w3043 , w3044 , w3045 , w3046 , w3047 , w3048 , w3049 , w3050 , w3051 , w3052 , w3053 , w3054 , w3055 , w3056 , w3057 , w3058 , w3059 , w3060 , w3061 , w3062 , w3063 , w3064 , w3065 , w3066 , w3067 , w3068 , w3069 , w3070 , w3071 , w3072 , w3073 , w3074 , w3075 , w3076 , w3077 , w3078 , w3079 , w3080 , w3081 , w3082 , w3083 , w3084 , w3085 , w3086 , w3087 , w3088 , w3089 , w3090 , w3091 , w3092 , w3093 , w3094 , w3095 , w3096 , w3097 , w3098 , w3099 , w3100 , w3101 , w3102 , w3103 , w3104 , w3105 , w3106 , w3107 , w3108 , w3109 , w3110 , w3111 , w3112 , w3113 , w3114 , w3115 , w3116 , w3117 , w3118 , w3119 , w3120 , w3121 , w3122 , w3123 , w3124 , w3125 , w3126 , w3127 , w3128 , w3129 , w3130 , w3131 , w3132 , w3133 , w3134 , w3135 , w3136 , w3137 , w3138 , w3139 , w3140 , w3141 , w3142 , w3143 , w3144 , w3145 , w3146 , w3147 , w3148 , w3149 , w3150 , w3151 , w3152 , w3153 , w3154 , w3155 , w3156 , w3157 , w3158 , w3159 , w3160 , w3161 , w3162 , w3163 , w3164 , w3165 , w3166 , w3167 , w3168 , w3169 , w3170 , w3171 , w3172 , w3173 , w3174 , w3175 , w3176 , w3177 , w3178 , w3179 , w3180 , w3181 , w3182 , w3183 , w3184 , w3185 , w3186 , w3187 , w3188 , w3189 , w3190 , w3191 , w3192 , w3193 , w3194 , w3195 , w3196 , w3197 , w3198 , w3199 , w3200 , w3201 , w3202 , w3203 , w3204 , w3205 , w3206 , w3207 , w3208 , w3209 , w3210 , w3211 , w3212 , w3213 , w3214 , w3215 , w3216 , w3217 , w3218 , w3219 , w3220 , w3221 , w3222 , w3223 , w3224 , w3225 , w3226 , w3227 , w3228 , w3229 , w3230 , w3231 , w3232 , w3233 , w3234 , w3235 , w3236 , w3237 , w3238 , w3239 , w3240 , w3241 , w3242 , w3243 , w3244 , w3245 , w3246 , w3247 , w3248 , w3249 , w3250 , w3251 , w3252 , w3253 , w3254 , w3255 , w3256 , w3257 , w3258 , w3259 , w3260 , w3261 , w3262 , w3263 , w3264 , w3265 , w3266 , w3267 , w3268 , w3269 , w3270 , w3271 , w3272 , w3273 , w3274 , w3275 , w3276 , w3277 , w3278 , w3279 , w3280 , w3281 , w3282 , w3283 , w3284 , w3285 , w3286 , w3287 , w3288 , w3289 , w3290 , w3291 , w3292 , w3293 , w3294 , w3295 , w3296 , w3297 , w3298 , w3299 , w3300 , w3301 , w3302 , w3303 , w3304 , w3305 , w3306 , w3307 , w3308 , w3309 , w3310 , w3311 , w3312 , w3313 , w3314 , w3315 , w3316 , w3317 , w3318 , w3319 , w3320 , w3321 , w3322 , w3323 , w3324 , w3325 , w3326 , w3327 , w3328 , w3329 , w3330 , w3331 , w3332 , w3333 , w3334 , w3335 , w3336 , w3337 , w3338 , w3339 , w3340 , w3341 , w3342 , w3343 , w3344 , w3345 , w3346 , w3347 , w3348 , w3349 , w3350 , w3351 , w3352 , w3353 , w3354 , w3355 , w3356 , w3357 , w3358 , w3359 , w3360 , w3361 , w3362 , w3363 , w3364 , w3365 , w3366 , w3367 , w3368 , w3369 , w3370 , w3371 , w3372 , w3373 , w3374 , w3375 , w3376 , w3377 , w3378 , w3379 , w3380 , w3381 , w3382 , w3383 , w3384 , w3385 , w3386 , w3387 , w3388 , w3389 , w3390 , w3391 , w3392 , w3393 , w3394 , w3395 , w3396 , w3397 , w3398 , w3399 , w3400 , w3401 , w3402 , w3403 , w3404 , w3405 , w3406 , w3407 , w3408 , w3409 , w3410 , w3411 , w3412 , w3413 , w3414 , w3415 , w3416 , w3417 , w3418 , w3419 , w3420 , w3421 , w3422 , w3423 , w3424 , w3425 , w3426 , w3427 , w3428 , w3429 , w3430 , w3431 , w3432 , w3433 , w3434 , w3435 , w3436 , w3437 , w3438 , w3439 , w3440 , w3441 , w3442 , w3443 , w3444 , w3445 , w3446 , w3447 , w3448 , w3449 , w3450 , w3451 , w3452 , w3453 , w3454 , w3455 , w3456 , w3457 , w3458 , w3459 , w3460 , w3461 , w3462 , w3463 , w3464 , w3465 , w3466 , w3467 , w3468 , w3469 , w3470 , w3471 , w3472 , w3473 , w3474 , w3475 , w3476 , w3477 , w3478 , w3479 , w3480 , w3481 , w3482 , w3483 , w3484 , w3485 , w3486 , w3487 , w3488 , w3489 , w3490 , w3491 , w3492 , w3493 , w3494 , w3495 , w3496 , w3497 , w3498 , w3499 , w3500 , w3501 , w3502 , w3503 , w3504 , w3505 , w3506 , w3507 , w3508 , w3509 , w3510 , w3511 , w3512 , w3513 , w3514 , w3515 , w3516 , w3517 , w3518 , w3519 , w3520 , w3521 , w3522 , w3523 , w3524 , w3525 , w3526 , w3527 , w3528 , w3529 , w3530 , w3531 , w3532 , w3533 , w3534 , w3535 , w3536 , w3537 , w3538 , w3539 , w3540 , w3541 , w3542 , w3543 , w3544 , w3545 , w3546 , w3547 , w3548 , w3549 , w3550 , w3551 , w3552 , w3553 , w3554 , w3555 , w3556 , w3557 , w3558 , w3559 , w3560 , w3561 , w3562 , w3563 , w3564 , w3565 , w3566 , w3567 , w3568 , w3569 , w3570 , w3571 , w3572 , w3573 , w3574 , w3575 , w3576 , w3577 , w3578 , w3579 , w3580 , w3581 , w3582 , w3583 , w3584 , w3585 , w3586 , w3587 , w3588 , w3589 , w3590 , w3591 , w3592 , w3593 , w3594 , w3595 , w3596 , w3597 , w3598 , w3599 , w3600 , w3601 , w3602 , w3603 , w3604 , w3605 , w3606 , w3607 , w3608 , w3609 , w3610 , w3611 , w3612 , w3613 , w3614 , w3615 , w3616 , w3617 , w3618 , w3619 , w3620 , w3621 , w3622 , w3623 , w3624 , w3625 , w3626 , w3627 , w3628 , w3629 , w3630 , w3631 , w3632 , w3633 , w3634 , w3635 , w3636 , w3637 , w3638 , w3639 , w3640 , w3641 , w3642 , w3643 , w3644 , w3645 , w3646 , w3647 , w3648 , w3649 , w3650 , w3651 , w3652 , w3653 , w3654 , w3655 , w3656 , w3657 , w3658 , w3659 , w3660 , w3661 , w3662 , w3663 , w3664 , w3665 , w3666 , w3667 , w3668 , w3669 , w3670 , w3671 , w3672 , w3673 , w3674 , w3675 , w3676 , w3677 , w3678 , w3679 , w3680 , w3681 , w3682 , w3683 , w3684 , w3685 , w3686 , w3687 , w3688 , w3689 , w3690 , w3691 , w3692 , w3693 , w3694 , w3695 , w3696 , w3697 , w3698 , w3699 , w3700 , w3701 , w3702 , w3703 , w3704 , w3705 , w3706 , w3707 , w3708 , w3709 , w3710 , w3711 , w3712 , w3713 , w3714 , w3715 , w3716 , w3717 , w3718 , w3719 , w3720 , w3721 , w3722 , w3723 , w3724 , w3725 , w3726 , w3727 , w3728 , w3729 , w3730 , w3731 , w3732 , w3733 , w3734 , w3735 , w3736 , w3737 , w3738 , w3739 , w3740 , w3741 , w3742 , w3743 , w3744 , w3745 , w3746 , w3747 , w3748 , w3749 , w3750 , w3751 , w3752 , w3753 , w3754 , w3755 , w3756 , w3757 , w3758 , w3759 , w3760 , w3761 , w3762 , w3763 , w3764 , w3765 , w3766 , w3767 , w3768 , w3769 , w3770 , w3771 , w3772 , w3773 , w3774 , w3775 , w3776 , w3777 , w3778 , w3779 , w3780 , w3781 , w3782 , w3783 , w3784 , w3785 , w3786 , w3787 , w3788 , w3789 , w3790 , w3791 , w3792 , w3793 , w3794 , w3795 , w3796 , w3797 , w3798 , w3799 , w3800 , w3801 , w3802 , w3803 , w3804 , w3805 , w3806 , w3807 , w3808 , w3809 , w3810 , w3811 , w3812 , w3813 , w3814 , w3815 , w3816 , w3817 , w3818 , w3819 , w3820 , w3821 , w3822 , w3823 , w3824 , w3825 , w3826 , w3827 , w3828 , w3829 , w3830 , w3831 , w3832 , w3833 , w3834 , w3835 , w3836 , w3837 , w3838 , w3839 , w3840 , w3841 , w3842 , w3843 , w3844 , w3845 , w3846 , w3847 , w3848 , w3849 , w3850 , w3851 , w3852 , w3853 , w3854 , w3855 , w3856 , w3857 , w3858 , w3859 , w3860 , w3861 , w3862 , w3863 , w3864 , w3865 , w3866 , w3867 , w3868 , w3869 , w3870 , w3871 , w3872 , w3873 , w3874 , w3875 , w3876 , w3877 , w3878 , w3879 , w3880 , w3881 , w3882 , w3883 , w3884 , w3885 , w3886 , w3887 , w3888 , w3889 , w3890 , w3891 , w3892 , w3893 , w3894 , w3895 , w3896 , w3897 , w3898 , w3899 , w3900 , w3901 , w3902 , w3903 , w3904 , w3905 , w3906 , w3907 , w3908 , w3909 , w3910 , w3911 , w3912 , w3913 , w3914 , w3915 , w3916 , w3917 , w3918 , w3919 , w3920 , w3921 , w3922 , w3923 , w3924 , w3925 , w3926 , w3927 , w3928 , w3929 , w3930 , w3931 , w3932 , w3933 , w3934 , w3935 , w3936 , w3937 , w3938 , w3939 , w3940 , w3941 , w3942 , w3943 , w3944 , w3945 , w3946 , w3947 , w3948 , w3949 , w3950 , w3951 , w3952 , w3953 , w3954 , w3955 , w3956 , w3957 , w3958 , w3959 , w3960 , w3961 , w3962 , w3963 , w3964 , w3965 , w3966 , w3967 , w3968 , w3969 , w3970 , w3971 , w3972 , w3973 , w3974 , w3975 , w3976 , w3977 , w3978 , w3979 , w3980 , w3981 , w3982 , w3983 , w3984 , w3985 , w3986 , w3987 , w3988 , w3989 , w3990 , w3991 , w3992 , w3993 , w3994 , w3995 , w3996 , w3997 , w3998 , w3999 , w4000 , w4001 , w4002 , w4003 , w4004 , w4005 , w4006 , w4007 , w4008 , w4009 , w4010 , w4011 , w4012 , w4013 , w4014 , w4015 , w4016 , w4017 , w4018 , w4019 , w4020 , w4021 , w4022 , w4023 , w4024 , w4025 , w4026 , w4027 , w4028 , w4029 , w4030 , w4031 , w4032 , w4033 , w4034 , w4035 , w4036 , w4037 , w4038 , w4039 , w4040 , w4041 , w4042 , w4043 , w4044 , w4045 , w4046 , w4047 , w4048 , w4049 , w4050 , w4051 , w4052 , w4053 , w4054 , w4055 , w4056 , w4057 , w4058 , w4059 , w4060 , w4061 , w4062 , w4063 , w4064 , w4065 , w4066 , w4067 , w4068 , w4069 , w4070 , w4071 , w4072 , w4073 , w4074 , w4075 , w4076 , w4077 , w4078 , w4079 , w4080 , w4081 , w4082 , w4083 , w4084 , w4085 , w4086 , w4087 , w4088 , w4089 , w4090 , w4091 , w4092 , w4093 , w4094 , w4095 , w4096 , w4097 , w4098 , w4099 , w4100 , w4101 , w4102 , w4103 , w4104 , w4105 , w4106 , w4107 , w4108 , w4109 , w4110 , w4111 , w4112 , w4113 , w4114 , w4115 , w4116 , w4117 , w4118 , w4119 , w4120 , w4121 , w4122 , w4123 , w4124 , w4125 , w4126 , w4127 , w4128 , w4129 , w4130 , w4131 , w4132 , w4133 , w4134 , w4135 , w4136 , w4137 , w4138 , w4139 , w4140 , w4141 , w4142 , w4143 , w4144 , w4145 , w4146 , w4147 , w4148 , w4149 , w4150 , w4151 , w4152 , w4153 , w4154 , w4155 , w4156 , w4157 , w4158 , w4159 , w4160 , w4161 , w4162 , w4163 , w4164 , w4165 , w4166 , w4167 , w4168 , w4169 , w4170 , w4171 , w4172 , w4173 , w4174 , w4175 , w4176 , w4177 , w4178 , w4179 , w4180 , w4181 , w4182 , w4183 , w4184 , w4185 , w4186 , w4187 , w4188 , w4189 , w4190 , w4191 , w4192 , w4193 , w4194 , w4195 , w4196 , w4197 , w4198 , w4199 , w4200 , w4201 , w4202 , w4203 , w4204 , w4205 , w4206 , w4207 , w4208 , w4209 , w4210 , w4211 , w4212 , w4213 , w4214 , w4215 , w4216 , w4217 , w4218 , w4219 , w4220 , w4221 , w4222 , w4223 , w4224 , w4225 , w4226 , w4227 , w4228 , w4229 , w4230 , w4231 , w4232 , w4233 , w4234 , w4235 , w4236 , w4237 , w4238 , w4239 , w4240 , w4241 , w4242 , w4243 , w4244 , w4245 , w4246 , w4247 , w4248 , w4249 , w4250 , w4251 , w4252 , w4253 , w4254 , w4255 , w4256 , w4257 , w4258 , w4259 , w4260 , w4261 , w4262 , w4263 , w4264 , w4265 , w4266 , w4267 , w4268 , w4269 , w4270 , w4271 , w4272 , w4273 , w4274 , w4275 , w4276 , w4277 , w4278 , w4279 , w4280 , w4281 , w4282 , w4283 , w4284 , w4285 , w4286 , w4287 , w4288 , w4289 , w4290 , w4291 , w4292 , w4293 , w4294 , w4295 , w4296 , w4297 , w4298 , w4299 , w4300 , w4301 , w4302 , w4303 , w4304 , w4305 , w4306 , w4307 , w4308 , w4309 , w4310 , w4311 , w4312 , w4313 , w4314 , w4315 , w4316 , w4317 , w4318 , w4319 , w4320 , w4321 , w4322 , w4323 , w4324 , w4325 , w4326 , w4327 , w4328 , w4329 , w4330 , w4331 , w4332 , w4333 , w4334 , w4335 , w4336 , w4337 , w4338 , w4339 , w4340 , w4341 , w4342 , w4343 , w4344 , w4345 , w4346 , w4347 , w4348 , w4349 , w4350 , w4351 , w4352 , w4353 , w4354 , w4355 , w4356 , w4357 , w4358 , w4359 , w4360 , w4361 , w4362 , w4363 , w4364 , w4365 , w4366 , w4367 , w4368 , w4369 , w4370 , w4371 , w4372 , w4373 , w4374 , w4375 , w4376 , w4377 , w4378 , w4379 , w4380 , w4381 , w4382 , w4383 , w4384 , w4385 , w4386 , w4387 , w4388 , w4389 , w4390 , w4391 , w4392 , w4393 , w4394 , w4395 , w4396 , w4397 , w4398 , w4399 , w4400 , w4401 , w4402 , w4403 , w4404 , w4405 , w4406 , w4407 , w4408 , w4409 , w4410 , w4411 , w4412 , w4413 , w4414 , w4415 , w4416 , w4417 , w4418 , w4419 , w4420 , w4421 , w4422 , w4423 , w4424 , w4425 , w4426 , w4427 , w4428 , w4429 , w4430 , w4431 , w4432 , w4433 , w4434 , w4435 , w4436 , w4437 , w4438 , w4439 , w4440 , w4441 , w4442 , w4443 , w4444 , w4445 , w4446 , w4447 , w4448 , w4449 , w4450 , w4451 , w4452 , w4453 , w4454 , w4455 , w4456 , w4457 , w4458 , w4459 , w4460 , w4461 , w4462 , w4463 , w4464 , w4465 , w4466 , w4467 , w4468 , w4469 , w4470 , w4471 , w4472 , w4473 , w4474 , w4475 , w4476 , w4477 , w4478 , w4479 , w4480 , w4481 , w4482 , w4483 , w4484 , w4485 , w4486 , w4487 , w4488 , w4489 , w4490 , w4491 , w4492 , w4493 , w4494 , w4495 , w4496 , w4497 , w4498 , w4499 , w4500 , w4501 , w4502 , w4503 , w4504 , w4505 , w4506 , w4507 , w4508 , w4509 , w4510 , w4511 , w4512 , w4513 , w4514 , w4515 , w4516 , w4517 , w4518 , w4519 , w4520 , w4521 , w4522 , w4523 , w4524 , w4525 , w4526 , w4527 , w4528 , w4529 , w4530 , w4531 , w4532 , w4533 , w4534 , w4535 , w4536 , w4537 , w4538 , w4539 , w4540 , w4541 , w4542 , w4543 , w4544 , w4545 , w4546 , w4547 , w4548 , w4549 , w4550 , w4551 , w4552 , w4553 , w4554 , w4555 , w4556 , w4557 , w4558 , w4559 , w4560 , w4561 , w4562 , w4563 , w4564 , w4565 , w4566 , w4567 , w4568 , w4569 , w4570 , w4571 , w4572 , w4573 , w4574 , w4575 , w4576 , w4577 , w4578 , w4579 , w4580 , w4581 , w4582 , w4583 , w4584 , w4585 , w4586 , w4587 , w4588 , w4589 , w4590 , w4591 , w4592 , w4593 , w4594 , w4595 , w4596 , w4597 , w4598 , w4599 , w4600 , w4601 , w4602 , w4603 , w4604 , w4605 , w4606 , w4607 , w4608 , w4609 , w4610 , w4611 , w4612 , w4613 , w4614 , w4615 , w4616 , w4617 , w4618 , w4619 , w4620 , w4621 , w4622 , w4623 , w4624 , w4625 , w4626 , w4627 , w4628 , w4629 , w4630 , w4631 , w4632 , w4633 , w4634 , w4635 , w4636 , w4637 , w4638 , w4639 , w4640 , w4641 , w4642 , w4643 , w4644 , w4645 , w4646 , w4647 , w4648 , w4649 , w4650 , w4651 , w4652 , w4653 , w4654 , w4655 , w4656 , w4657 , w4658 , w4659 , w4660 , w4661 , w4662 , w4663 , w4664 , w4665 , w4666 , w4667 , w4668 , w4669 , w4670 , w4671 , w4672 , w4673 , w4674 , w4675 , w4676 , w4677 , w4678 , w4679 , w4680 , w4681 , w4682 , w4683 , w4684 , w4685 , w4686 , w4687 , w4688 , w4689 , w4690 , w4691 , w4692 , w4693 , w4694 , w4695 , w4696 , w4697 , w4698 , w4699 , w4700 , w4701 , w4702 , w4703 , w4704 , w4705 , w4706 , w4707 , w4708 , w4709 , w4710 , w4711 , w4712 , w4713 , w4714 , w4715 , w4716 , w4717 , w4718 , w4719 , w4720 , w4721 , w4722 , w4723 , w4724 , w4725 , w4726 , w4727 , w4728 , w4729 , w4730 , w4731 , w4732 , w4733 , w4734 , w4735 , w4736 , w4737 , w4738 , w4739 , w4740 , w4741 , w4742 , w4743 , w4744 , w4745 , w4746 , w4747 , w4748 , w4749 , w4750 , w4751 , w4752 , w4753 , w4754 , w4755 , w4756 , w4757 , w4758 , w4759 , w4760 , w4761 , w4762 , w4763 , w4764 , w4765 , w4766 , w4767 , w4768 , w4769 , w4770 , w4771 , w4772 , w4773 , w4774 , w4775 , w4776 , w4777 , w4778 , w4779 , w4780 , w4781 , w4782 , w4783 , w4784 , w4785 , w4786 , w4787 , w4788 , w4789 , w4790 , w4791 , w4792 , w4793 , w4794 , w4795 , w4796 , w4797 , w4798 , w4799 , w4800 , w4801 , w4802 , w4803 , w4804 , w4805 , w4806 , w4807 , w4808 , w4809 , w4810 , w4811 , w4812 , w4813 , w4814 , w4815 , w4816 , w4817 , w4818 , w4819 , w4820 , w4821 , w4822 , w4823 , w4824 , w4825 , w4826 , w4827 , w4828 , w4829 , w4830 , w4831 , w4832 , w4833 , w4834 , w4835 , w4836 , w4837 , w4838 , w4839 , w4840 , w4841 , w4842 , w4843 , w4844 , w4845 , w4846 , w4847 , w4848 , w4849 , w4850 , w4851 , w4852 , w4853 , w4854 , w4855 , w4856 , w4857 , w4858 , w4859 , w4860 , w4861 , w4862 , w4863 , w4864 , w4865 , w4866 , w4867 , w4868 , w4869 , w4870 , w4871 , w4872 , w4873 , w4874 , w4875 , w4876 , w4877 , w4878 , w4879 , w4880 , w4881 , w4882 , w4883 , w4884 , w4885 , w4886 , w4887 , w4888 , w4889 , w4890 , w4891 , w4892 , w4893 , w4894 , w4895 , w4896 , w4897 , w4898 , w4899 , w4900 , w4901 , w4902 , w4903 , w4904 , w4905 , w4906 , w4907 , w4908 , w4909 , w4910 , w4911 , w4912 , w4913 , w4914 , w4915 , w4916 , w4917 , w4918 , w4919 , w4920 , w4921 , w4922 , w4923 , w4924 , w4925 , w4926 , w4927 , w4928 , w4929 , w4930 , w4931 , w4932 , w4933 , w4934 , w4935 , w4936 , w4937 , w4938 , w4939 , w4940 , w4941 , w4942 , w4943 , w4944 , w4945 , w4946 , w4947 , w4948 , w4949 , w4950 , w4951 , w4952 , w4953 , w4954 , w4955 , w4956 , w4957 , w4958 , w4959 , w4960 , w4961 , w4962 , w4963 , w4964 , w4965 , w4966 , w4967 , w4968 , w4969 , w4970 , w4971 , w4972 , w4973 , w4974 , w4975 , w4976 , w4977 , w4978 , w4979 , w4980 , w4981 , w4982 , w4983 , w4984 , w4985 , w4986 , w4987 , w4988 , w4989 , w4990 , w4991 , w4992 , w4993 , w4994 , w4995 , w4996 , w4997 , w4998 , w4999 , w5000 , w5001 , w5002 , w5003 , w5004 , w5005 , w5006 , w5007 , w5008 , w5009 , w5010 , w5011 , w5012 , w5013 , w5014 , w5015 , w5016 , w5017 , w5018 , w5019 , w5020 , w5021 , w5022 , w5023 , w5024 , w5025 , w5026 , w5027 , w5028 , w5029 , w5030 , w5031 , w5032 , w5033 , w5034 , w5035 , w5036 , w5037 , w5038 , w5039 , w5040 , w5041 , w5042 , w5043 , w5044 , w5045 , w5046 , w5047 , w5048 , w5049 , w5050 , w5051 , w5052 , w5053 , w5054 , w5055 , w5056 , w5057 , w5058 , w5059 , w5060 , w5061 , w5062 , w5063 , w5064 , w5065 , w5066 , w5067 , w5068 , w5069 , w5070 , w5071 , w5072 , w5073 , w5074 , w5075 , w5076 , w5077 , w5078 , w5079 , w5080 , w5081 , w5082 , w5083 , w5084 , w5085 , w5086 , w5087 , w5088 , w5089 , w5090 , w5091 , w5092 , w5093 , w5094 , w5095 , w5096 , w5097 , w5098 , w5099 , w5100 , w5101 , w5102 , w5103 , w5104 , w5105 , w5106 , w5107 , w5108 , w5109 , w5110 , w5111 , w5112 , w5113 , w5114 , w5115 , w5116 , w5117 , w5118 , w5119 , w5120 , w5121 , w5122 , w5123 , w5124 , w5125 , w5126 , w5127 , w5128 , w5129 , w5130 , w5131 , w5132 , w5133 , w5134 , w5135 , w5136 , w5137 , w5138 , w5139 , w5140 , w5141 , w5142 , w5143 , w5144 , w5145 , w5146 , w5147 , w5148 , w5149 , w5150 , w5151 , w5152 , w5153 , w5154 , w5155 , w5156 , w5157 , w5158 , w5159 , w5160 , w5161 , w5162 , w5163 , w5164 , w5165 , w5166 , w5167 , w5168 , w5169 , w5170 , w5171 , w5172 , w5173 , w5174 , w5175 , w5176 , w5177 , w5178 , w5179 , w5180 , w5181 , w5182 , w5183 , w5184 , w5185 , w5186 , w5187 , w5188 , w5189 , w5190 , w5191 , w5192 , w5193 , w5194 , w5195 , w5196 , w5197 , w5198 , w5199 , w5200 , w5201 , w5202 , w5203 , w5204 , w5205 , w5206 , w5207 , w5208 , w5209 , w5210 , w5211 , w5212 , w5213 , w5214 , w5215 , w5216 , w5217 , w5218 , w5219 , w5220 , w5221 , w5222 , w5223 , w5224 , w5225 , w5226 , w5227 , w5228 , w5229 , w5230 , w5231 , w5232 , w5233 , w5234 , w5235 , w5236 , w5237 , w5238 , w5239 , w5240 , w5241 , w5242 , w5243 , w5244 , w5245 , w5246 , w5247 , w5248 , w5249 , w5250 , w5251 , w5252 , w5253 , w5254 , w5255 , w5256 , w5257 , w5258 , w5259 , w5260 , w5261 , w5262 , w5263 , w5264 , w5265 , w5266 , w5267 , w5268 , w5269 , w5270 , w5271 , w5272 , w5273 , w5274 , w5275 , w5276 , w5277 , w5278 , w5279 , w5280 , w5281 , w5282 , w5283 , w5284 , w5285 , w5286 , w5287 , w5288 , w5289 , w5290 , w5291 , w5292 , w5293 , w5294 , w5295 , w5296 , w5297 , w5298 , w5299 , w5300 , w5301 , w5302 , w5303 , w5304 , w5305 , w5306 , w5307 , w5308 , w5309 , w5310 , w5311 , w5312 , w5313 , w5314 , w5315 , w5316 , w5317 , w5318 , w5319 , w5320 , w5321 , w5322 , w5323 , w5324 , w5325 , w5326 , w5327 , w5328 , w5329 , w5330 , w5331 , w5332 , w5333 , w5334 , w5335 , w5336 , w5337 , w5338 , w5339 , w5340 , w5341 , w5342 , w5343 , w5344 , w5345 , w5346 , w5347 , w5348 , w5349 , w5350 , w5351 , w5352 , w5353 , w5354 , w5355 , w5356 , w5357 , w5358 , w5359 , w5360 , w5361 , w5362 , w5363 , w5364 , w5365 , w5366 , w5367 , w5368 , w5369 , w5370 , w5371 , w5372 , w5373 , w5374 , w5375 , w5376 , w5377 , w5378 , w5379 , w5380 , w5381 , w5382 , w5383 , w5384 , w5385 , w5386 , w5387 , w5388 , w5389 , w5390 , w5391 , w5392 , w5393 , w5394 , w5395 , w5396 , w5397 , w5398 , w5399 , w5400 , w5401 , w5402 , w5403 , w5404 , w5405 , w5406 , w5407 , w5408 , w5409 , w5410 , w5411 , w5412 , w5413 , w5414 , w5415 , w5416 , w5417 , w5418 , w5419 , w5420 , w5421 , w5422 , w5423 , w5424 , w5425 , w5426 , w5427 , w5428 , w5429 , w5430 , w5431 , w5432 , w5433 , w5434 , w5435 , w5436 , w5437 , w5438 , w5439 , w5440 , w5441 , w5442 , w5443 , w5444 , w5445 , w5446 , w5447 , w5448 , w5449 , w5450 , w5451 , w5452 , w5453 , w5454 , w5455 , w5456 , w5457 , w5458 , w5459 , w5460 , w5461 , w5462 , w5463 , w5464 , w5465 , w5466 , w5467 , w5468 , w5469 , w5470 , w5471 , w5472 , w5473 , w5474 , w5475 , w5476 , w5477 , w5478 , w5479 , w5480 , w5481 , w5482 , w5483 , w5484 , w5485 , w5486 , w5487 , w5488 , w5489 , w5490 , w5491 , w5492 , w5493 , w5494 , w5495 , w5496 , w5497 , w5498 , w5499 , w5500 , w5501 , w5502 , w5503 , w5504 , w5505 , w5506 , w5507 , w5508 , w5509 , w5510 , w5511 , w5512 , w5513 , w5514 , w5515 , w5516 , w5517 , w5518 , w5519 , w5520 , w5521 , w5522 , w5523 , w5524 , w5525 , w5526 , w5527 , w5528 , w5529 , w5530 , w5531 , w5532 , w5533 , w5534 , w5535 , w5536 , w5537 , w5538 , w5539 , w5540 , w5541 , w5542 , w5543 , w5544 , w5545 , w5546 , w5547 , w5548 , w5549 , w5550 , w5551 , w5552 , w5553 , w5554 , w5555 , w5556 , w5557 , w5558 , w5559 , w5560 , w5561 , w5562 , w5563 , w5564 , w5565 , w5566 , w5567 , w5568 , w5569 , w5570 , w5571 , w5572 , w5573 , w5574 , w5575 , w5576 , w5577 , w5578 , w5579 , w5580 , w5581 , w5582 , w5583 , w5584 , w5585 , w5586 , w5587 , w5588 , w5589 , w5590 , w5591 , w5592 , w5593 , w5594 , w5595 , w5596 , w5597 , w5598 , w5599 , w5600 , w5601 , w5602 , w5603 , w5604 , w5605 , w5606 , w5607 , w5608 , w5609 , w5610 , w5611 , w5612 , w5613 , w5614 , w5615 , w5616 , w5617 , w5618 , w5619 , w5620 , w5621 , w5622 , w5623 , w5624 , w5625 , w5626 , w5627 , w5628 , w5629 , w5630 , w5631 , w5632 , w5633 , w5634 , w5635 , w5636 , w5637 , w5638 , w5639 , w5640 , w5641 , w5642 , w5643 , w5644 , w5645 , w5646 , w5647 , w5648 , w5649 , w5650 , w5651 , w5652 , w5653 , w5654 , w5655 , w5656 , w5657 , w5658 , w5659 , w5660 , w5661 , w5662 , w5663 , w5664 , w5665 , w5666 , w5667 , w5668 , w5669 , w5670 , w5671 , w5672 , w5673 , w5674 , w5675 , w5676 , w5677 , w5678 , w5679 , w5680 , w5681 , w5682 , w5683 , w5684 , w5685 , w5686 , w5687 , w5688 , w5689 , w5690 , w5691 , w5692 , w5693 , w5694 , w5695 , w5696 , w5697 , w5698 , w5699 , w5700 , w5701 , w5702 , w5703 , w5704 , w5705 , w5706 , w5707 , w5708 , w5709 , w5710 , w5711 , w5712 , w5713 , w5714 , w5715 , w5716 , w5717 , w5718 , w5719 , w5720 , w5721 , w5722 , w5723 , w5724 , w5725 , w5726 , w5727 , w5728 , w5729 , w5730 , w5731 , w5732 , w5733 , w5734 , w5735 , w5736 , w5737 , w5738 , w5739 , w5740 , w5741 , w5742 , w5743 , w5744 , w5745 , w5746 , w5747 , w5748 , w5749 , w5750 , w5751 , w5752 , w5753 , w5754 , w5755 , w5756 , w5757 , w5758 , w5759 , w5760 , w5761 , w5762 , w5763 , w5764 , w5765 , w5766 , w5767 , w5768 , w5769 , w5770 , w5771 , w5772 , w5773 , w5774 , w5775 , w5776 , w5777 , w5778 , w5779 , w5780 , w5781 , w5782 , w5783 , w5784 , w5785 , w5786 , w5787 , w5788 , w5789 , w5790 , w5791 , w5792 , w5793 , w5794 , w5795 , w5796 , w5797 , w5798 , w5799 , w5800 , w5801 , w5802 , w5803 , w5804 , w5805 , w5806 , w5807 , w5808 , w5809 , w5810 , w5811 , w5812 , w5813 , w5814 , w5815 , w5816 , w5817 , w5818 , w5819 , w5820 , w5821 , w5822 , w5823 , w5824 , w5825 , w5826 , w5827 , w5828 , w5829 , w5830 , w5831 , w5832 , w5833 , w5834 , w5835 , w5836 , w5837 , w5838 , w5839 , w5840 , w5841 , w5842 , w5843 , w5844 , w5845 , w5846 , w5847 , w5848 , w5849 , w5850 , w5851 , w5852 , w5853 , w5854 , w5855 , w5856 , w5857 , w5858 , w5859 , w5860 , w5861 , w5862 , w5863 , w5864 , w5865 , w5866 , w5867 , w5868 , w5869 , w5870 , w5871 , w5872 , w5873 , w5874 , w5875 , w5876 , w5877 , w5878 , w5879 , w5880 , w5881 , w5882 , w5883 , w5884 , w5885 , w5886 , w5887 , w5888 , w5889 , w5890 , w5891 , w5892 , w5893 , w5894 , w5895 , w5896 , w5897 , w5898 , w5899 , w5900 , w5901 , w5902 , w5903 , w5904 , w5905 , w5906 , w5907 , w5908 , w5909 , w5910 , w5911 , w5912 , w5913 , w5914 , w5915 , w5916 , w5917 , w5918 , w5919 , w5920 , w5921 , w5922 , w5923 , w5924 , w5925 , w5926 , w5927 , w5928 , w5929 , w5930 , w5931 , w5932 , w5933 , w5934 , w5935 , w5936 , w5937 , w5938 , w5939 , w5940 , w5941 , w5942 , w5943 , w5944 , w5945 , w5946 , w5947 , w5948 , w5949 , w5950 , w5951 , w5952 , w5953 , w5954 , w5955 , w5956 , w5957 , w5958 , w5959 , w5960 , w5961 , w5962 , w5963 , w5964 , w5965 , w5966 , w5967 , w5968 , w5969 , w5970 , w5971 , w5972 , w5973 , w5974 , w5975 , w5976 , w5977 , w5978 , w5979 , w5980 , w5981 , w5982 , w5983 , w5984 , w5985 , w5986 , w5987 , w5988 , w5989 , w5990 , w5991 , w5992 , w5993 , w5994 , w5995 , w5996 , w5997 , w5998 , w5999 , w6000 , w6001 , w6002 , w6003 , w6004 , w6005 , w6006 , w6007 , w6008 , w6009 , w6010 , w6011 , w6012 , w6013 , w6014 , w6015 , w6016 , w6017 , w6018 , w6019 , w6020 , w6021 , w6022 , w6023 , w6024 , w6025 , w6026 , w6027 , w6028 , w6029 , w6030 , w6031 , w6032 , w6033 , w6034 , w6035 , w6036 , w6037 , w6038 , w6039 , w6040 , w6041 , w6042 , w6043 , w6044 , w6045 , w6046 , w6047 , w6048 , w6049 , w6050 , w6051 , w6052 , w6053 , w6054 , w6055 , w6056 , w6057 , w6058 , w6059 , w6060 , w6061 , w6062 , w6063 , w6064 , w6065 , w6066 , w6067 , w6068 , w6069 , w6070 , w6071 , w6072 , w6073 , w6074 , w6075 , w6076 , w6077 , w6078 , w6079 , w6080 , w6081 , w6082 , w6083 , w6084 , w6085 , w6086 , w6087 , w6088 , w6089 , w6090 , w6091 , w6092 , w6093 , w6094 , w6095 , w6096 , w6097 , w6098 , w6099 , w6100 , w6101 , w6102 , w6103 , w6104 , w6105 , w6106 , w6107 , w6108 , w6109 , w6110 , w6111 , w6112 , w6113 , w6114 , w6115 , w6116 , w6117 , w6118 , w6119 , w6120 , w6121 , w6122 , w6123 , w6124 , w6125 , w6126 , w6127 , w6128 , w6129 , w6130 , w6131 , w6132 , w6133 , w6134 , w6135 , w6136 , w6137 , w6138 , w6139 , w6140 , w6141 , w6142 , w6143 , w6144 , w6145 , w6146 , w6147 , w6148 , w6149 , w6150 , w6151 , w6152 , w6153 , w6154 , w6155 , w6156 , w6157 , w6158 , w6159 , w6160 , w6161 , w6162 , w6163 , w6164 , w6165 , w6166 , w6167 , w6168 , w6169 , w6170 , w6171 , w6172 , w6173 , w6174 , w6175 , w6176 , w6177 , w6178 , w6179 , w6180 , w6181 , w6182 , w6183 , w6184 , w6185 , w6186 , w6187 , w6188 , w6189 , w6190 , w6191 , w6192 , w6193 , w6194 , w6195 , w6196 , w6197 , w6198 , w6199 , w6200 , w6201 , w6202 , w6203 , w6204 , w6205 , w6206 , w6207 , w6208 , w6209 , w6210 , w6211 , w6212 , w6213 , w6214 , w6215 , w6216 , w6217 , w6218 , w6219 , w6220 , w6221 , w6222 , w6223 , w6224 , w6225 , w6226 , w6227 , w6228 , w6229 , w6230 , w6231 , w6232 , w6233 , w6234 , w6235 , w6236 , w6237 , w6238 , w6239 , w6240 , w6241 , w6242 , w6243 , w6244 , w6245 , w6246 , w6247 , w6248 , w6249 , w6250 , w6251 , w6252 , w6253 , w6254 , w6255 , w6256 , w6257 , w6258 , w6259 , w6260 , w6261 , w6262 , w6263 , w6264 , w6265 , w6266 , w6267 , w6268 , w6269 , w6270 , w6271 , w6272 , w6273 , w6274 , w6275 , w6276 , w6277 , w6278 , w6279 , w6280 , w6281 , w6282 , w6283 , w6284 , w6285 , w6286 , w6287 , w6288 , w6289 , w6290 , w6291 , w6292 , w6293 , w6294 , w6295 , w6296 , w6297 , w6298 , w6299 , w6300 , w6301 , w6302 , w6303 , w6304 , w6305 , w6306 , w6307 , w6308 , w6309 , w6310 , w6311 , w6312 , w6313 , w6314 , w6315 , w6316 , w6317 , w6318 , w6319 , w6320 , w6321 , w6322 , w6323 , w6324 , w6325 , w6326 , w6327 , w6328 , w6329 , w6330 , w6331 , w6332 , w6333 , w6334 , w6335 , w6336 , w6337 , w6338 , w6339 , w6340 , w6341 , w6342 , w6343 , w6344 , w6345 , w6346 , w6347 , w6348 , w6349 , w6350 , w6351 , w6352 , w6353 , w6354 , w6355 , w6356 , w6357 , w6358 , w6359 , w6360 , w6361 , w6362 , w6363 , w6364 , w6365 , w6366 , w6367 , w6368 , w6369 , w6370 , w6371 , w6372 , w6373 , w6374 , w6375 , w6376 , w6377 , w6378 , w6379 , w6380 , w6381 , w6382 , w6383 , w6384 , w6385 , w6386 , w6387 , w6388 , w6389 , w6390 , w6391 , w6392 , w6393 , w6394 , w6395 , w6396 , w6397 , w6398 , w6399 , w6400 , w6401 , w6402 , w6403 , w6404 , w6405 , w6406 , w6407 , w6408 , w6409 , w6410 , w6411 , w6412 , w6413 , w6414 , w6415 , w6416 , w6417 , w6418 , w6419 , w6420 , w6421 , w6422 , w6423 , w6424 , w6425 , w6426 , w6427 , w6428 , w6429 , w6430 , w6431 , w6432 , w6433 , w6434 , w6435 , w6436 , w6437 , w6438 , w6439 , w6440 , w6441 , w6442 , w6443 , w6444 , w6445 , w6446 , w6447 , w6448 , w6449 , w6450 , w6451 , w6452 , w6453 , w6454 , w6455 , w6456 , w6457 , w6458 , w6459 , w6460 , w6461 , w6462 , w6463 , w6464 , w6465 , w6466 , w6467 , w6468 , w6469 , w6470 , w6471 , w6472 , w6473 , w6474 , w6475 , w6476 , w6477 , w6478 , w6479 , w6480 , w6481 , w6482 , w6483 , w6484 , w6485 , w6486 , w6487 , w6488 , w6489 , w6490 , w6491 , w6492 , w6493 , w6494 , w6495 , w6496 , w6497 , w6498 , w6499 , w6500 , w6501 , w6502 , w6503 , w6504 , w6505 , w6506 , w6507 , w6508 , w6509 , w6510 , w6511 , w6512 , w6513 , w6514 , w6515 , w6516 , w6517 , w6518 , w6519 , w6520 , w6521 , w6522 , w6523 , w6524 , w6525 , w6526 , w6527 , w6528 , w6529 , w6530 , w6531 , w6532 , w6533 , w6534 , w6535 , w6536 , w6537 , w6538 , w6539 , w6540 , w6541 , w6542 , w6543 , w6544 , w6545 , w6546 , w6547 , w6548 , w6549 , w6550 , w6551 , w6552 , w6553 , w6554 , w6555 , w6556 , w6557 , w6558 , w6559 , w6560 , w6561 , w6562 , w6563 , w6564 , w6565 , w6566 , w6567 , w6568 , w6569 , w6570 , w6571 , w6572 , w6573 , w6574 , w6575 , w6576 , w6577 , w6578 , w6579 , w6580 , w6581 , w6582 , w6583 , w6584 , w6585 , w6586 , w6587 , w6588 , w6589 , w6590 , w6591 , w6592 , w6593 , w6594 , w6595 , w6596 , w6597 , w6598 , w6599 , w6600 , w6601 , w6602 , w6603 , w6604 , w6605 , w6606 , w6607 , w6608 , w6609 , w6610 , w6611 , w6612 , w6613 , w6614 , w6615 , w6616 , w6617 , w6618 , w6619 , w6620 , w6621 , w6622 , w6623 , w6624 , w6625 , w6626 , w6627 , w6628 , w6629 , w6630 , w6631 , w6632 , w6633 , w6634 , w6635 , w6636 , w6637 , w6638 , w6639 , w6640 , w6641 , w6642 , w6643 , w6644 , w6645 , w6646 , w6647 , w6648 , w6649 , w6650 , w6651 , w6652 , w6653 , w6654 , w6655 , w6656 , w6657 , w6658 , w6659 , w6660 , w6661 , w6662 , w6663 , w6664 , w6665 , w6666 , w6667 , w6668 , w6669 , w6670 , w6671 , w6672 , w6673 , w6674 , w6675 , w6676 , w6677 , w6678 , w6679 , w6680 , w6681 , w6682 , w6683 , w6684 , w6685 , w6686 , w6687 , w6688 , w6689 , w6690 , w6691 , w6692 , w6693 , w6694 , w6695 , w6696 , w6697 , w6698 , w6699 , w6700 , w6701 , w6702 , w6703 , w6704 , w6705 , w6706 , w6707 , w6708 , w6709 , w6710 , w6711 , w6712 , w6713 , w6714 , w6715 , w6716 , w6717 , w6718 , w6719 , w6720 , w6721 , w6722 , w6723 , w6724 , w6725 , w6726 , w6727 , w6728 , w6729 , w6730 , w6731 , w6732 , w6733 , w6734 , w6735 , w6736 , w6737 , w6738 , w6739 , w6740 , w6741 , w6742 , w6743 , w6744 , w6745 , w6746 , w6747 , w6748 , w6749 , w6750 , w6751 , w6752 , w6753 , w6754 , w6755 , w6756 , w6757 , w6758 , w6759 , w6760 , w6761 , w6762 , w6763 , w6764 , w6765 , w6766 , w6767 , w6768 , w6769 , w6770 , w6771 , w6772 , w6773 , w6774 , w6775 , w6776 , w6777 , w6778 , w6779 , w6780 , w6781 , w6782 , w6783 , w6784 , w6785 , w6786 , w6787 , w6788 , w6789 , w6790 , w6791 , w6792 , w6793 , w6794 , w6795 , w6796 , w6797 , w6798 , w6799 , w6800 , w6801 , w6802 , w6803 , w6804 , w6805 , w6806 , w6807 , w6808 , w6809 , w6810 , w6811 , w6812 , w6813 , w6814 , w6815 , w6816 , w6817 , w6818 , w6819 , w6820 , w6821 , w6822 , w6823 , w6824 , w6825 , w6826 , w6827 , w6828 , w6829 , w6830 , w6831 , w6832 , w6833 , w6834 , w6835 , w6836 , w6837 , w6838 , w6839 , w6840 , w6841 , w6842 , w6843 , w6844 , w6845 , w6846 , w6847 , w6848 , w6849 , w6850 , w6851 , w6852 , w6853 , w6854 , w6855 , w6856 , w6857 , w6858 , w6859 , w6860 , w6861 , w6862 , w6863 , w6864 , w6865 , w6866 , w6867 , w6868 , w6869 , w6870 , w6871 , w6872 , w6873 , w6874 , w6875 , w6876 , w6877 , w6878 , w6879 , w6880 , w6881 , w6882 , w6883 , w6884 , w6885 , w6886 , w6887 , w6888 , w6889 , w6890 , w6891 , w6892 , w6893 , w6894 , w6895 , w6896 , w6897 , w6898 , w6899 , w6900 , w6901 , w6902 , w6903 , w6904 , w6905 , w6906 , w6907 , w6908 , w6909 , w6910 , w6911 , w6912 , w6913 , w6914 , w6915 , w6916 , w6917 , w6918 , w6919 , w6920 , w6921 , w6922 , w6923 , w6924 , w6925 , w6926 , w6927 , w6928 , w6929 , w6930 , w6931 , w6932 , w6933 , w6934 , w6935 , w6936 , w6937 , w6938 , w6939 , w6940 , w6941 , w6942 , w6943 , w6944 , w6945 , w6946 , w6947 , w6948 , w6949 , w6950 , w6951 , w6952 , w6953 , w6954 , w6955 , w6956 , w6957 , w6958 , w6959 , w6960 , w6961 , w6962 , w6963 , w6964 , w6965 , w6966 , w6967 , w6968 , w6969 , w6970 , w6971 , w6972 , w6973 , w6974 , w6975 , w6976 , w6977 , w6978 , w6979 , w6980 , w6981 , w6982 , w6983 , w6984 , w6985 , w6986 , w6987 , w6988 , w6989 , w6990 , w6991 , w6992 , w6993 , w6994 , w6995 , w6996 , w6997 , w6998 , w6999 , w7000 , w7001 , w7002 , w7003 , w7004 , w7005 , w7006 , w7007 , w7008 , w7009 , w7010 , w7011 , w7012 , w7013 , w7014 , w7015 , w7016 , w7017 , w7018 , w7019 , w7020 , w7021 , w7022 , w7023 , w7024 , w7025 , w7026 , w7027 , w7028 , w7029 , w7030 , w7031 , w7032 , w7033 , w7034 , w7035 , w7036 , w7037 , w7038 , w7039 , w7040 , w7041 , w7042 , w7043 , w7044 , w7045 , w7046 , w7047 , w7048 , w7049 , w7050 , w7051 , w7052 , w7053 , w7054 , w7055 , w7056 , w7057 , w7058 , w7059 , w7060 , w7061 , w7062 , w7063 , w7064 , w7065 , w7066 , w7067 , w7068 , w7069 , w7070 , w7071 , w7072 , w7073 , w7074 , w7075 , w7076 , w7077 , w7078 , w7079 , w7080 , w7081 , w7082 , w7083 , w7084 , w7085 , w7086 , w7087 , w7088 , w7089 , w7090 , w7091 , w7092 , w7093 , w7094 , w7095 , w7096 , w7097 , w7098 , w7099 , w7100 , w7101 , w7102 , w7103 , w7104 , w7105 , w7106 , w7107 , w7108 , w7109 , w7110 , w7111 , w7112 , w7113 , w7114 , w7115 , w7116 , w7117 , w7118 , w7119 , w7120 , w7121 , w7122 , w7123 , w7124 , w7125 , w7126 , w7127 , w7128 , w7129 , w7130 , w7131 , w7132 , w7133 , w7134 , w7135 , w7136 , w7137 , w7138 , w7139 , w7140 , w7141 , w7142 , w7143 , w7144 , w7145 , w7146 , w7147 , w7148 , w7149 , w7150 , w7151 , w7152 , w7153 , w7154 , w7155 , w7156 , w7157 , w7158 , w7159 , w7160 , w7161 , w7162 , w7163 , w7164 , w7165 , w7166 , w7167 , w7168 , w7169 , w7170 , w7171 , w7172 , w7173 , w7174 , w7175 , w7176 , w7177 , w7178 , w7179 , w7180 , w7181 , w7182 , w7183 , w7184 , w7185 , w7186 , w7187 , w7188 , w7189 , w7190 , w7191 , w7192 , w7193 , w7194 , w7195 , w7196 , w7197 , w7198 , w7199 , w7200 , w7201 , w7202 , w7203 , w7204 , w7205 , w7206 , w7207 , w7208 , w7209 , w7210 , w7211 , w7212 , w7213 , w7214 , w7215 , w7216 , w7217 , w7218 , w7219 , w7220 , w7221 , w7222 , w7223 , w7224 , w7225 , w7226 , w7227 , w7228 , w7229 , w7230 , w7231 , w7232 , w7233 , w7234 , w7235 , w7236 , w7237 , w7238 , w7239 , w7240 , w7241 , w7242 , w7243 , w7244 , w7245 , w7246 , w7247 , w7248 , w7249 , w7250 , w7251 , w7252 , w7253 , w7254 , w7255 , w7256 , w7257 , w7258 , w7259 , w7260 , w7261 , w7262 , w7263 , w7264 , w7265 , w7266 , w7267 , w7268 , w7269 , w7270 , w7271 , w7272 , w7273 , w7274 , w7275 , w7276 , w7277 , w7278 , w7279 , w7280 , w7281 , w7282 , w7283 , w7284 , w7285 , w7286 , w7287 , w7288 , w7289 , w7290 , w7291 , w7292 , w7293 , w7294 , w7295 , w7296 , w7297 , w7298 , w7299 , w7300 , w7301 , w7302 , w7303 , w7304 , w7305 , w7306 , w7307 , w7308 , w7309 , w7310 , w7311 , w7312 , w7313 , w7314 , w7315 , w7316 , w7317 , w7318 , w7319 , w7320 , w7321 , w7322 , w7323 , w7324 , w7325 , w7326 , w7327 , w7328 , w7329 , w7330 , w7331 , w7332 , w7333 , w7334 , w7335 , w7336 , w7337 , w7338 , w7339 , w7340 , w7341 , w7342 , w7343 , w7344 , w7345 , w7346 , w7347 , w7348 , w7349 , w7350 , w7351 , w7352 , w7353 , w7354 , w7355 , w7356 , w7357 , w7358 , w7359 , w7360 , w7361 , w7362 , w7363 , w7364 , w7365 , w7366 , w7367 , w7368 , w7369 , w7370 , w7371 , w7372 , w7373 , w7374 , w7375 , w7376 , w7377 , w7378 , w7379 , w7380 , w7381 , w7382 , w7383 , w7384 , w7385 , w7386 , w7387 , w7388 , w7389 , w7390 , w7391 , w7392 , w7393 , w7394 , w7395 , w7396 , w7397 , w7398 , w7399 , w7400 , w7401 , w7402 , w7403 , w7404 , w7405 , w7406 , w7407 , w7408 , w7409 , w7410 , w7411 , w7412 , w7413 , w7414 , w7415 , w7416 , w7417 , w7418 , w7419 , w7420 , w7421 , w7422 , w7423 , w7424 , w7425 , w7426 , w7427 , w7428 , w7429 , w7430 , w7431 , w7432 , w7433 , w7434 , w7435 , w7436 , w7437 , w7438 , w7439 , w7440 , w7441 , w7442 , w7443 , w7444 , w7445 , w7446 , w7447 , w7448 , w7449 , w7450 , w7451 , w7452 , w7453 , w7454 , w7455 , w7456 , w7457 , w7458 , w7459 , w7460 , w7461 , w7462 , w7463 , w7464 , w7465 , w7466 , w7467 , w7468 , w7469 , w7470 , w7471 , w7472 , w7473 , w7474 , w7475 , w7476 , w7477 , w7478 , w7479 , w7480 , w7481 , w7482 , w7483 , w7484 , w7485 , w7486 , w7487 , w7488 , w7489 , w7490 , w7491 , w7492 , w7493 , w7494 , w7495 , w7496 , w7497 , w7498 , w7499 , w7500 , w7501 , w7502 , w7503 , w7504 , w7505 , w7506 , w7507 , w7508 , w7509 , w7510 , w7511 , w7512 , w7513 , w7514 , w7515 , w7516 , w7517 , w7518 , w7519 , w7520 , w7521 , w7522 , w7523 , w7524 , w7525 , w7526 , w7527 , w7528 , w7529 , w7530 , w7531 , w7532 , w7533 , w7534 , w7535 , w7536 , w7537 , w7538 , w7539 , w7540 , w7541 , w7542 , w7543 , w7544 , w7545 , w7546 , w7547 , w7548 , w7549 , w7550 , w7551 , w7552 , w7553 , w7554 , w7555 , w7556 , w7557 , w7558 , w7559 , w7560 , w7561 , w7562 , w7563 , w7564 , w7565 , w7566 , w7567 , w7568 , w7569 , w7570 , w7571 , w7572 , w7573 , w7574 , w7575 , w7576 , w7577 , w7578 , w7579 , w7580 , w7581 , w7582 , w7583 , w7584 , w7585 , w7586 , w7587 , w7588 , w7589 , w7590 , w7591 , w7592 , w7593 , w7594 , w7595 , w7596 , w7597 , w7598 , w7599 , w7600 , w7601 , w7602 , w7603 , w7604 , w7605 , w7606 , w7607 , w7608 , w7609 , w7610 , w7611 , w7612 , w7613 , w7614 , w7615 , w7616 , w7617 , w7618 , w7619 , w7620 , w7621 , w7622 , w7623 , w7624 , w7625 , w7626 , w7627 , w7628 , w7629 , w7630 , w7631 , w7632 , w7633 , w7634 , w7635 , w7636 , w7637 , w7638 , w7639 , w7640 , w7641 , w7642 , w7643 , w7644 , w7645 , w7646 , w7647 , w7648 , w7649 , w7650 , w7651 , w7652 , w7653 , w7654 , w7655 , w7656 , w7657 , w7658 , w7659 , w7660 , w7661 , w7662 , w7663 , w7664 , w7665 , w7666 , w7667 , w7668 , w7669 , w7670 , w7671 , w7672 , w7673 , w7674 , w7675 , w7676 , w7677 , w7678 , w7679 , w7680 , w7681 , w7682 , w7683 , w7684 , w7685 , w7686 , w7687 , w7688 , w7689 , w7690 , w7691 , w7692 , w7693 , w7694 , w7695 , w7696 , w7697 , w7698 , w7699 , w7700 , w7701 , w7702 , w7703 , w7704 , w7705 , w7706 , w7707 , w7708 , w7709 , w7710 , w7711 , w7712 , w7713 , w7714 , w7715 , w7716 , w7717 , w7718 , w7719 , w7720 , w7721 , w7722 , w7723 , w7724 , w7725 , w7726 , w7727 , w7728 , w7729 , w7730 , w7731 , w7732 , w7733 , w7734 , w7735 , w7736 , w7737 , w7738 , w7739 , w7740 , w7741 , w7742 , w7743 , w7744 , w7745 , w7746 , w7747 , w7748 , w7749 , w7750 , w7751 , w7752 , w7753 , w7754 , w7755 , w7756 , w7757 , w7758 , w7759 , w7760 , w7761 , w7762 , w7763 , w7764 , w7765 , w7766 , w7767 , w7768 , w7769 , w7770 , w7771 , w7772 , w7773 , w7774 , w7775 , w7776 , w7777 , w7778 , w7779 , w7780 , w7781 , w7782 , w7783 , w7784 , w7785 , w7786 , w7787 , w7788 , w7789 , w7790 , w7791 , w7792 , w7793 , w7794 , w7795 , w7796 , w7797 , w7798 , w7799 , w7800 , w7801 , w7802 , w7803 , w7804 , w7805 , w7806 , w7807 , w7808 , w7809 , w7810 , w7811 , w7812 , w7813 , w7814 , w7815 , w7816 , w7817 , w7818 , w7819 , w7820 , w7821 , w7822 , w7823 , w7824 , w7825 , w7826 , w7827 , w7828 , w7829 , w7830 , w7831 , w7832 , w7833 , w7834 , w7835 , w7836 , w7837 , w7838 , w7839 , w7840 , w7841 , w7842 , w7843 , w7844 , w7845 , w7846 , w7847 , w7848 , w7849 , w7850 , w7851 , w7852 , w7853 , w7854 , w7855 , w7856 , w7857 , w7858 , w7859 , w7860 , w7861 , w7862 , w7863 , w7864 , w7865 , w7866 , w7867 , w7868 , w7869 , w7870 , w7871 , w7872 , w7873 , w7874 , w7875 , w7876 , w7877 , w7878 , w7879 , w7880 , w7881 , w7882 , w7883 , w7884 , w7885 , w7886 , w7887 , w7888 , w7889 , w7890 , w7891 , w7892 , w7893 , w7894 , w7895 , w7896 , w7897 , w7898 , w7899 , w7900 , w7901 , w7902 , w7903 , w7904 , w7905 , w7906 , w7907 , w7908 , w7909 , w7910 , w7911 , w7912 , w7913 , w7914 , w7915 , w7916 , w7917 , w7918 , w7919 , w7920 , w7921 , w7922 , w7923 , w7924 , w7925 , w7926 , w7927 , w7928 , w7929 , w7930 , w7931 , w7932 , w7933 , w7934 , w7935 , w7936 , w7937 , w7938 , w7939 , w7940 , w7941 , w7942 , w7943 , w7944 , w7945 , w7946 , w7947 , w7948 , w7949 , w7950 , w7951 , w7952 , w7953 , w7954 , w7955 , w7956 , w7957 , w7958 , w7959 , w7960 , w7961 , w7962 , w7963 , w7964 , w7965 , w7966 , w7967 , w7968 , w7969 , w7970 , w7971 , w7972 , w7973 , w7974 , w7975 , w7976 , w7977 , w7978 , w7979 , w7980 , w7981 , w7982 , w7983 , w7984 , w7985 , w7986 , w7987 , w7988 , w7989 , w7990 , w7991 , w7992 , w7993 , w7994 , w7995 , w7996 , w7997 , w7998 , w7999 , w8000 , w8001 , w8002 , w8003 , w8004 , w8005 , w8006 , w8007 , w8008 , w8009 , w8010 , w8011 , w8012 , w8013 , w8014 , w8015 , w8016 , w8017 , w8018 , w8019 , w8020 , w8021 , w8022 , w8023 , w8024 , w8025 , w8026 , w8027 , w8028 , w8029 , w8030 , w8031 , w8032 , w8033 , w8034 , w8035 , w8036 , w8037 , w8038 , w8039 , w8040 , w8041 , w8042 , w8043 , w8044 , w8045 , w8046 , w8047 , w8048 , w8049 , w8050 , w8051 , w8052 , w8053 , w8054 , w8055 , w8056 , w8057 , w8058 , w8059 , w8060 , w8061 , w8062 , w8063 , w8064 , w8065 , w8066 , w8067 , w8068 , w8069 , w8070 , w8071 , w8072 , w8073 , w8074 , w8075 , w8076 , w8077 , w8078 , w8079 , w8080 , w8081 , w8082 , w8083 , w8084 , w8085 , w8086 , w8087 , w8088 , w8089 , w8090 , w8091 , w8092 , w8093 , w8094 , w8095 , w8096 , w8097 , w8098 , w8099 , w8100 , w8101 , w8102 , w8103 , w8104 , w8105 , w8106 , w8107 , w8108 , w8109 , w8110 , w8111 , w8112 , w8113 , w8114 , w8115 , w8116 , w8117 , w8118 , w8119 , w8120 , w8121 , w8122 , w8123 , w8124 , w8125 , w8126 , w8127 , w8128 , w8129 , w8130 , w8131 , w8132 , w8133 , w8134 , w8135 , w8136 , w8137 , w8138 , w8139 , w8140 , w8141 , w8142 , w8143 , w8144 , w8145 , w8146 , w8147 , w8148 , w8149 , w8150 , w8151 , w8152 , w8153 , w8154 , w8155 , w8156 , w8157 , w8158 , w8159 , w8160 , w8161 , w8162 , w8163 , w8164 , w8165 , w8166 , w8167 , w8168 , w8169 , w8170 , w8171 , w8172 , w8173 , w8174 , w8175 , w8176 , w8177 , w8178 , w8179 , w8180 , w8181 , w8182 , w8183 , w8184 , w8185 , w8186 , w8187 , w8188 , w8189 , w8190 , w8191 , w8192 , w8193 , w8194 , w8195 , w8196 , w8197 , w8198 , w8199 , w8200 , w8201 , w8202 , w8203 , w8204 , w8205 , w8206 , w8207 , w8208 , w8209 , w8210 , w8211 , w8212 , w8213 , w8214 , w8215 , w8216 , w8217 , w8218 , w8219 , w8220 , w8221 , w8222 , w8223 , w8224 , w8225 , w8226 , w8227 , w8228 , w8229 , w8230 , w8231 , w8232 , w8233 , w8234 , w8235 , w8236 , w8237 , w8238 , w8239 , w8240 , w8241 , w8242 , w8243 , w8244 , w8245 , w8246 , w8247 , w8248 , w8249 , w8250 , w8251 , w8252 , w8253 , w8254 , w8255 , w8256 , w8257 , w8258 , w8259 , w8260 , w8261 , w8262 , w8263 , w8264 , w8265 , w8266 , w8267 , w8268 , w8269 , w8270 , w8271 , w8272 , w8273 , w8274 , w8275 , w8276 , w8277 , w8278 , w8279 , w8280 , w8281 , w8282 , w8283 , w8284 , w8285 , w8286 , w8287 , w8288 , w8289 , w8290 , w8291 , w8292 , w8293 , w8294 , w8295 , w8296 , w8297 , w8298 , w8299 , w8300 , w8301 , w8302 , w8303 , w8304 , w8305 , w8306 , w8307 , w8308 , w8309 , w8310 , w8311 , w8312 , w8313 , w8314 , w8315 , w8316 , w8317 , w8318 , w8319 , w8320 , w8321 , w8322 , w8323 , w8324 , w8325 , w8326 , w8327 , w8328 , w8329 , w8330 , w8331 , w8332 , w8333 , w8334 , w8335 , w8336 , w8337 , w8338 , w8339 , w8340 , w8341 , w8342 , w8343 , w8344 , w8345 , w8346 , w8347 , w8348 , w8349 , w8350 , w8351 , w8352 , w8353 , w8354 , w8355 , w8356 , w8357 , w8358 , w8359 , w8360 , w8361 , w8362 , w8363 , w8364 , w8365 , w8366 , w8367 , w8368 , w8369 , w8370 , w8371 , w8372 , w8373 , w8374 , w8375 , w8376 , w8377 , w8378 , w8379 , w8380 , w8381 , w8382 , w8383 , w8384 , w8385 , w8386 , w8387 , w8388 , w8389 , w8390 , w8391 , w8392 , w8393 , w8394 , w8395 , w8396 , w8397 , w8398 , w8399 , w8400 , w8401 , w8402 , w8403 , w8404 , w8405 , w8406 , w8407 , w8408 , w8409 , w8410 , w8411 , w8412 , w8413 , w8414 , w8415 , w8416 , w8417 , w8418 , w8419 , w8420 , w8421 , w8422 , w8423 , w8424 , w8425 , w8426 , w8427 , w8428 , w8429 , w8430 , w8431 , w8432 , w8433 , w8434 , w8435 , w8436 , w8437 , w8438 , w8439 , w8440 , w8441 , w8442 , w8443 , w8444 , w8445 , w8446 , w8447 , w8448 , w8449 , w8450 , w8451 , w8452 , w8453 , w8454 , w8455 , w8456 , w8457 , w8458 , w8459 , w8460 , w8461 , w8462 , w8463 , w8464 , w8465 , w8466 , w8467 , w8468 , w8469 , w8470 , w8471 , w8472 , w8473 , w8474 , w8475 , w8476 , w8477 , w8478 , w8479 , w8480 , w8481 , w8482 , w8483 , w8484 , w8485 , w8486 , w8487 , w8488 , w8489 , w8490 , w8491 , w8492 , w8493 , w8494 , w8495 , w8496 , w8497 , w8498 , w8499 , w8500 , w8501 , w8502 , w8503 , w8504 , w8505 , w8506 , w8507 , w8508 , w8509 , w8510 , w8511 , w8512 , w8513 , w8514 , w8515 , w8516 , w8517 , w8518 , w8519 , w8520 , w8521 , w8522 , w8523 , w8524 , w8525 , w8526 , w8527 , w8528 , w8529 , w8530 , w8531 , w8532 , w8533 , w8534 , w8535 , w8536 , w8537 , w8538 , w8539 , w8540 , w8541 , w8542 , w8543 , w8544 , w8545 , w8546 , w8547 , w8548 , w8549 , w8550 , w8551 , w8552 , w8553 , w8554 , w8555 , w8556 , w8557 , w8558 , w8559 , w8560 , w8561 , w8562 , w8563 , w8564 , w8565 , w8566 , w8567 , w8568 , w8569 , w8570 , w8571 , w8572 , w8573 , w8574 , w8575 , w8576 , w8577 , w8578 , w8579 , w8580 , w8581 , w8582 , w8583 , w8584 , w8585 , w8586 , w8587 , w8588 , w8589 , w8590 , w8591 ;
  assign zero = 0;
  assign w65 = ~\pi00 & \pi01 ;
  assign w66 = \pi01 ^ \pi02 ;
  assign w67 = \pi00 & w66 ;
  assign w68 = \pi00 | \pi01 ;
  assign w69 = \pi00 & \pi03 ;
  assign w70 = \pi02 ^ w69 ;
  assign w71 = ( \pi00 & ~w68 ) | ( \pi00 & w70 ) | ( ~w68 & w70 ) ;
  assign w72 = \pi02 & \pi03 ;
  assign w73 = ( \pi01 & \pi02 ) | ( \pi01 & \pi03 ) | ( \pi02 & \pi03 ) ;
  assign w74 = \pi00 ^ \pi04 ;
  assign w75 = ( \pi04 & w72 ) | ( \pi04 & ~w74 ) | ( w72 & ~w74 ) ;
  assign w76 = w73 ^ w75 ;
  assign w77 = \pi00 & \pi01 ;
  assign w78 = ( \pi03 & \pi05 ) | ( \pi03 & w77 ) | ( \pi05 & w77 ) ;
  assign w79 = ( \pi04 & ~w77 ) | ( \pi04 & w78 ) | ( ~w77 & w78 ) ;
  assign w80 = w77 & w79 ;
  assign w81 = ( \pi01 & ~\pi04 ) | ( \pi01 & w73 ) | ( ~\pi04 & w73 ) ;
  assign w82 = ( \pi01 & \pi03 ) | ( \pi01 & ~w81 ) | ( \pi03 & ~w81 ) ;
  assign w83 = \pi04 & w73 ;
  assign w84 = \pi00 ^ \pi05 ;
  assign w85 = ( \pi05 & w83 ) | ( \pi05 & ~w84 ) | ( w83 & ~w84 ) ;
  assign w86 = w82 ^ w85 ;
  assign w87 = ( \pi02 & ~\pi05 ) | ( \pi02 & w69 ) | ( ~\pi05 & w69 ) ;
  assign w88 = \pi00 & w87 ;
  assign w89 = \pi03 ^ w88 ;
  assign w90 = ( \pi01 & ~\pi04 ) | ( \pi01 & w89 ) | ( ~\pi04 & w89 ) ;
  assign w91 = \pi05 & w69 ;
  assign w92 = ( \pi04 & w90 ) | ( \pi04 & w91 ) | ( w90 & w91 ) ;
  assign w93 = \pi01 & \pi05 ;
  assign w94 = \pi02 & \pi04 ;
  assign w95 = w93 ^ w94 ;
  assign w96 = w72 ^ w80 ;
  assign w97 = w92 ^ w96 ;
  assign w98 = w95 ^ w97 ;
  assign w99 = \pi00 & \pi06 ;
  assign w100 = w98 ^ w99 ;
  assign w101 = \pi03 & \pi04 ;
  assign w102 = \pi02 & \pi05 ;
  assign w103 = \pi00 & \pi07 ;
  assign w104 = ( w101 & w102 ) | ( w101 & w103 ) | ( w102 & w103 ) ;
  assign w105 = w101 ^ w103 ;
  assign w106 = w102 ^ w105 ;
  assign w107 = ( w72 & w95 ) | ( w72 & w99 ) | ( w95 & w99 ) ;
  assign w108 = ( \pi01 & ~\pi04 ) | ( \pi01 & \pi06 ) | ( ~\pi04 & \pi06 ) ;
  assign w109 = \pi04 & w108 ;
  assign w110 = ~\pi01 & \pi02 ;
  assign w111 = ( ~\pi02 & \pi05 ) | ( ~\pi02 & w110 ) | ( \pi05 & w110 ) ;
  assign w112 = ( \pi04 & ~\pi05 ) | ( \pi04 & w111 ) | ( ~\pi05 & w111 ) ;
  assign w113 = w107 ^ w112 ;
  assign w114 = \pi01 & \pi06 ;
  assign w115 = w113 ^ w114 ;
  assign w116 = w72 ^ w95 ;
  assign w117 = w99 ^ w116 ;
  assign w118 = ( w80 & w92 ) | ( w80 & w117 ) | ( w92 & w117 ) ;
  assign w119 = w115 ^ w118 ;
  assign w120 = w106 ^ w119 ;
  assign w121 = ( ~\pi06 & w102 ) | ( ~\pi06 & w107 ) | ( w102 & w107 ) ;
  assign w122 = \pi04 & w121 ;
  assign w123 = ( \pi01 & \pi04 ) | ( \pi01 & ~\pi06 ) | ( \pi04 & ~\pi06 ) ;
  assign w124 = ( \pi01 & \pi04 ) | ( \pi01 & w107 ) | ( \pi04 & w107 ) ;
  assign w125 = ( w122 & ~w123 ) | ( w122 & w124 ) | ( ~w123 & w124 ) ;
  assign w126 = \pi01 & \pi07 ;
  assign w127 = \pi06 & \pi08 ;
  assign w128 = \pi02 & \pi06 ;
  assign w129 = \pi00 & \pi08 ;
  assign w130 = ( w109 & w128 ) | ( w109 & w129 ) | ( w128 & w129 ) ;
  assign w131 = w109 ^ w129 ;
  assign w132 = w128 ^ w131 ;
  assign w133 = \pi03 & \pi05 ;
  assign w134 = w104 ^ w126 ;
  assign w135 = w132 ^ w134 ;
  assign w136 = w133 ^ w135 ;
  assign w137 = ( w106 & w115 ) | ( w106 & w118 ) | ( w115 & w118 ) ;
  assign w138 = w125 ^ w137 ;
  assign w139 = w136 ^ w138 ;
  assign w140 = w126 ^ w133 ;
  assign w141 = ( w104 & w132 ) | ( w104 & w140 ) | ( w132 & w140 ) ;
  assign w142 = \pi04 & \pi05 ;
  assign w143 = \pi03 & \pi06 ;
  assign w144 = \pi02 & \pi07 ;
  assign w145 = ( w142 & w143 ) | ( w142 & w144 ) | ( w143 & w144 ) ;
  assign w146 = w142 ^ w144 ;
  assign w147 = w143 ^ w146 ;
  assign w148 = \pi00 & \pi09 ;
  assign w149 = \pi03 & w126 ;
  assign w150 = \pi05 & w149 ;
  assign w151 = w148 ^ w150 ;
  assign w152 = \pi05 & \pi08 ;
  assign w153 = w130 ^ w151 ;
  assign w154 = w147 ^ w153 ;
  assign w155 = \pi05 ^ w154 ;
  assign w156 = \pi01 & \pi08 ;
  assign w157 = w155 ^ w156 ;
  assign w158 = ( w125 & w136 ) | ( w125 & w137 ) | ( w136 & w137 ) ;
  assign w159 = w141 ^ w158 ;
  assign w160 = w157 ^ w159 ;
  assign w161 = ( w141 & w157 ) | ( w141 & w158 ) | ( w157 & w158 ) ;
  assign w162 = \pi05 ^ w151 ;
  assign w163 = w156 ^ w162 ;
  assign w164 = ( w130 & w147 ) | ( w130 & w163 ) | ( w147 & w163 ) ;
  assign w165 = \pi08 & \pi10 ;
  assign w166 = \pi07 & \pi08 ;
  assign w167 = \pi03 & \pi07 ;
  assign w168 = \pi02 & \pi08 ;
  assign w169 = \pi00 & \pi10 ;
  assign w170 = ( w167 & w168 ) | ( w167 & w169 ) | ( w168 & w169 ) ;
  assign w171 = w167 ^ w169 ;
  assign w172 = w168 ^ w171 ;
  assign w173 = ( ~\pi08 & w148 ) | ( ~\pi08 & w167 ) | ( w148 & w167 ) ;
  assign w174 = \pi05 & w173 ;
  assign w175 = ( \pi01 & \pi05 ) | ( \pi01 & ~\pi08 ) | ( \pi05 & ~\pi08 ) ;
  assign w176 = ( \pi01 & \pi05 ) | ( \pi01 & w148 ) | ( \pi05 & w148 ) ;
  assign w177 = ( w174 & ~w175 ) | ( w174 & w176 ) | ( ~w175 & w176 ) ;
  assign w178 = \pi04 & \pi06 ;
  assign w179 = w145 ^ w178 ;
  assign w180 = \pi09 ^ w152 ;
  assign w181 = \pi01 & w180 ;
  assign w182 = w179 ^ w181 ;
  assign w183 = w177 ^ w182 ;
  assign w184 = w172 ^ w183 ;
  assign w185 = w161 ^ w164 ;
  assign w186 = w184 ^ w185 ;
  assign w187 = ( w172 & w177 ) | ( w172 & w182 ) | ( w177 & w182 ) ;
  assign w188 = ( \pi03 & \pi08 ) | ( \pi03 & ~\pi09 ) | ( \pi08 & ~\pi09 ) ;
  assign w189 = ( \pi02 & w109 ) | ( \pi02 & w188 ) | ( w109 & w188 ) ;
  assign w190 = \pi09 & w189 ;
  assign w191 = \pi03 & \pi08 ;
  assign w192 = \pi02 ^ w109 ;
  assign w193 = \pi09 & w192 ;
  assign w194 = w191 ^ w193 ;
  assign w195 = \pi01 & \pi10 ;
  assign w196 = \pi06 ^ w170 ;
  assign w197 = w194 ^ w196 ;
  assign w198 = w195 ^ w197 ;
  assign w199 = \pi01 & w152 ;
  assign w200 = \pi01 & \pi09 ;
  assign w201 = w178 ^ w200 ;
  assign w202 = ( w145 & w199 ) | ( w145 & w201 ) | ( w199 & w201 ) ;
  assign w203 = \pi05 & \pi06 ;
  assign w204 = \pi04 & \pi07 ;
  assign w205 = \pi00 & \pi11 ;
  assign w206 = ( w203 & w204 ) | ( w203 & w205 ) | ( w204 & w205 ) ;
  assign w207 = w203 ^ w205 ;
  assign w208 = w204 ^ w207 ;
  assign w209 = w198 ^ w202 ;
  assign w210 = w208 ^ w209 ;
  assign w211 = ( w161 & w164 ) | ( w161 & w184 ) | ( w164 & w184 ) ;
  assign w212 = w210 ^ w211 ;
  assign w213 = w187 ^ w212 ;
  assign w214 = ( w187 & w210 ) | ( w187 & w211 ) | ( w210 & w211 ) ;
  assign w215 = ( w198 & w202 ) | ( w198 & w208 ) | ( w202 & w208 ) ;
  assign w216 = \pi10 & \pi12 ;
  assign w217 = \pi09 & \pi10 ;
  assign w218 = \pi03 & \pi09 ;
  assign w219 = \pi02 & \pi10 ;
  assign w220 = \pi00 & \pi12 ;
  assign w221 = ( w218 & w219 ) | ( w218 & w220 ) | ( w219 & w220 ) ;
  assign w222 = w218 ^ w220 ;
  assign w223 = w219 ^ w222 ;
  assign w224 = w190 ^ w206 ;
  assign w225 = w223 ^ w224 ;
  assign w226 = \pi06 ^ w195 ;
  assign w227 = ( w170 & w194 ) | ( w170 & w226 ) | ( w194 & w226 ) ;
  assign w228 = \pi05 & \pi11 ;
  assign w229 = \pi01 & \pi11 ;
  assign w230 = \pi05 & \pi07 ;
  assign w231 = w229 ^ w230 ;
  assign w232 = ( \pi01 & ~\pi06 ) | ( \pi01 & \pi10 ) | ( ~\pi06 & \pi10 ) ;
  assign w233 = \pi06 & w232 ;
  assign w234 = \pi04 & \pi08 ;
  assign w235 = ( w231 & w233 ) | ( w231 & w234 ) | ( w233 & w234 ) ;
  assign w236 = w231 ^ w233 ;
  assign w237 = w234 ^ w236 ;
  assign w238 = w225 ^ w227 ;
  assign w239 = w237 ^ w238 ;
  assign w240 = w214 ^ w215 ;
  assign w241 = w239 ^ w240 ;
  assign w242 = \pi04 & \pi09 ;
  assign w243 = \pi03 & \pi10 ;
  assign w244 = \pi00 & \pi13 ;
  assign w245 = ( w242 & w243 ) | ( w242 & w244 ) | ( w243 & w244 ) ;
  assign w246 = w242 ^ w244 ;
  assign w247 = w243 ^ w246 ;
  assign w248 = \pi06 & \pi07 ;
  assign w249 = \pi02 & \pi11 ;
  assign w250 = ( w152 & w248 ) | ( w152 & w249 ) | ( w248 & w249 ) ;
  assign w251 = w248 ^ w249 ;
  assign w252 = w152 ^ w251 ;
  assign w253 = w235 ^ w247 ;
  assign w254 = w252 ^ w253 ;
  assign w255 = ( w190 & w206 ) | ( w190 & w223 ) | ( w206 & w223 ) ;
  assign w256 = ( ~\pi01 & \pi07 ) | ( ~\pi01 & w228 ) | ( \pi07 & w228 ) ;
  assign w257 = \pi12 ^ w256 ;
  assign w258 = \pi01 & w257 ;
  assign w259 = \pi07 ^ w221 ;
  assign w260 = w258 ^ w259 ;
  assign w261 = ( w225 & w227 ) | ( w225 & w237 ) | ( w227 & w237 ) ;
  assign w262 = w255 ^ w261 ;
  assign w263 = w260 ^ w262 ;
  assign w264 = ( w214 & w215 ) | ( w214 & w239 ) | ( w215 & w239 ) ;
  assign w265 = w263 ^ w264 ;
  assign w266 = w254 ^ w265 ;
  assign w267 = ( w254 & w263 ) | ( w254 & w264 ) | ( w263 & w264 ) ;
  assign w268 = ( w255 & w260 ) | ( w255 & w261 ) | ( w260 & w261 ) ;
  assign w269 = ( ~\pi01 & \pi13 ) | ( ~\pi01 & w127 ) | ( \pi13 & w127 ) ;
  assign w270 = \pi01 & w269 ;
  assign w271 = \pi01 & \pi13 ;
  assign w272 = w245 ^ w250 ;
  assign w273 = w127 ^ w272 ;
  assign w274 = w271 ^ w273 ;
  assign w275 = ( w235 & w247 ) | ( w235 & w252 ) | ( w247 & w252 ) ;
  assign w276 = \pi03 & \pi11 ;
  assign w277 = \pi02 & \pi12 ;
  assign w278 = \pi00 & \pi14 ;
  assign w279 = ( w276 & w277 ) | ( w276 & w278 ) | ( w277 & w278 ) ;
  assign w280 = w276 ^ w278 ;
  assign w281 = w277 ^ w280 ;
  assign w282 = \pi05 & \pi09 ;
  assign w283 = \pi04 & \pi10 ;
  assign w284 = \pi12 & w126 ;
  assign w285 = ( w282 & w283 ) | ( w282 & w284 ) | ( w283 & w284 ) ;
  assign w286 = w282 ^ w284 ;
  assign w287 = w283 ^ w286 ;
  assign w288 = ( \pi01 & ~\pi07 ) | ( \pi01 & w228 ) | ( ~\pi07 & w228 ) ;
  assign w289 = \pi01 & \pi12 ;
  assign w290 = ( w221 & w288 ) | ( w221 & ~w289 ) | ( w288 & ~w289 ) ;
  assign w291 = ( \pi07 & w289 ) | ( \pi07 & w290 ) | ( w289 & w290 ) ;
  assign w292 = w290 & w291 ;
  assign w293 = w287 ^ w292 ;
  assign w294 = w281 ^ w293 ;
  assign w295 = w275 ^ w294 ;
  assign w296 = w274 ^ w295 ;
  assign w297 = w267 ^ w268 ;
  assign w298 = w296 ^ w297 ;
  assign w299 = ( w267 & w268 ) | ( w267 & w296 ) | ( w268 & w296 ) ;
  assign w300 = ( w274 & w275 ) | ( w274 & w294 ) | ( w275 & w294 ) ;
  assign w301 = \pi01 & \pi14 ;
  assign w302 = \pi08 ^ w301 ;
  assign w303 = \pi04 & \pi11 ;
  assign w304 = ( w270 & w302 ) | ( w270 & w303 ) | ( w302 & w303 ) ;
  assign w305 = w270 ^ w303 ;
  assign w306 = \pi08 ^ w305 ;
  assign w307 = w301 ^ w306 ;
  assign w308 = \pi06 & \pi09 ;
  assign w309 = \pi02 & \pi13 ;
  assign w310 = ( w166 & w308 ) | ( w166 & w309 ) | ( w308 & w309 ) ;
  assign w311 = w166 ^ w309 ;
  assign w312 = w308 ^ w311 ;
  assign w313 = w127 ^ w271 ;
  assign w314 = ( w245 & w250 ) | ( w245 & w313 ) | ( w250 & w313 ) ;
  assign w315 = w307 ^ w312 ;
  assign w316 = w314 ^ w315 ;
  assign w317 = \pi10 & \pi15 ;
  assign w318 = \pi05 & \pi10 ;
  assign w319 = \pi03 & \pi12 ;
  assign w320 = \pi00 & \pi15 ;
  assign w321 = ( w318 & w319 ) | ( w318 & w320 ) | ( w319 & w320 ) ;
  assign w322 = w318 ^ w320 ;
  assign w323 = w319 ^ w322 ;
  assign w324 = w279 ^ w285 ;
  assign w325 = w323 ^ w324 ;
  assign w326 = ( w281 & w287 ) | ( w281 & w292 ) | ( w287 & w292 ) ;
  assign w327 = w316 ^ w325 ;
  assign w328 = w326 ^ w327 ;
  assign w329 = w299 ^ w328 ;
  assign w330 = w300 ^ w329 ;
  assign w331 = ( w316 & w325 ) | ( w316 & w326 ) | ( w325 & w326 ) ;
  assign w332 = \pi06 & \pi16 ;
  assign w333 = \pi06 & \pi10 ;
  assign w334 = \pi00 & \pi16 ;
  assign w335 = ( w228 & w333 ) | ( w228 & w334 ) | ( w333 & w334 ) ;
  assign w336 = w333 ^ w334 ;
  assign w337 = w228 ^ w336 ;
  assign w338 = w304 ^ w321 ;
  assign w339 = w337 ^ w338 ;
  assign w340 = ( w307 & w312 ) | ( w307 & w314 ) | ( w312 & w314 ) ;
  assign w341 = ( w279 & w285 ) | ( w279 & w323 ) | ( w285 & w323 ) ;
  assign w342 = \pi12 & \pi13 ;
  assign w343 = \pi04 & \pi12 ;
  assign w344 = \pi03 & \pi13 ;
  assign w345 = \pi02 & \pi14 ;
  assign w346 = ( w343 & w344 ) | ( w343 & w345 ) | ( w344 & w345 ) ;
  assign w347 = w343 ^ w345 ;
  assign w348 = w344 ^ w347 ;
  assign w349 = \pi07 & \pi09 ;
  assign w350 = ( ~\pi01 & \pi15 ) | ( ~\pi01 & w349 ) | ( \pi15 & w349 ) ;
  assign w351 = \pi01 & w350 ;
  assign w352 = ( ~\pi01 & \pi08 ) | ( ~\pi01 & \pi14 ) | ( \pi08 & \pi14 ) ;
  assign w353 = \pi15 ^ w352 ;
  assign w354 = \pi01 & w353 ;
  assign w355 = w310 ^ w349 ;
  assign w356 = w354 ^ w355 ;
  assign w357 = w341 ^ w356 ;
  assign w358 = w348 ^ w357 ;
  assign w359 = w339 ^ w340 ;
  assign w360 = w358 ^ w359 ;
  assign w361 = ( w299 & w300 ) | ( w299 & w328 ) | ( w300 & w328 ) ;
  assign w362 = w331 ^ w361 ;
  assign w363 = w360 ^ w362 ;
  assign w364 = ( w339 & w340 ) | ( w339 & w358 ) | ( w340 & w358 ) ;
  assign w365 = \pi05 & \pi12 ;
  assign w366 = \pi00 & \pi17 ;
  assign w367 = ( w351 & w365 ) | ( w351 & w366 ) | ( w365 & w366 ) ;
  assign w368 = w351 ^ w366 ;
  assign w369 = w365 ^ w368 ;
  assign w370 = \pi08 & \pi09 ;
  assign w371 = \pi07 & \pi10 ;
  assign w372 = \pi03 & \pi14 ;
  assign w373 = ( w370 & w371 ) | ( w370 & w372 ) | ( w371 & w372 ) ;
  assign w374 = w370 ^ w372 ;
  assign w375 = w371 ^ w374 ;
  assign w376 = \pi11 & \pi13 ;
  assign w377 = \pi13 & \pi15 ;
  assign w378 = \pi06 & \pi11 ;
  assign w379 = \pi04 & \pi13 ;
  assign w380 = \pi02 & \pi15 ;
  assign w381 = ( w378 & w379 ) | ( w378 & w380 ) | ( w379 & w380 ) ;
  assign w382 = w378 ^ w380 ;
  assign w383 = w379 ^ w382 ;
  assign w384 = w369 ^ w375 ;
  assign w385 = w383 ^ w384 ;
  assign w386 = ( w341 & w348 ) | ( w341 & w356 ) | ( w348 & w356 ) ;
  assign w387 = \pi14 & w156 ;
  assign w388 = \pi01 & \pi15 ;
  assign w389 = w349 ^ w388 ;
  assign w390 = ( w310 & w387 ) | ( w310 & w389 ) | ( w387 & w389 ) ;
  assign w391 = ( w304 & w321 ) | ( w304 & w337 ) | ( w321 & w337 ) ;
  assign w392 = \pi09 & \pi16 ;
  assign w393 = \pi01 & \pi16 ;
  assign w394 = \pi09 ^ w346 ;
  assign w395 = w335 ^ w394 ;
  assign w396 = w393 ^ w395 ;
  assign w397 = w390 ^ w391 ;
  assign w398 = w396 ^ w397 ;
  assign w399 = w385 ^ w398 ;
  assign w400 = w386 ^ w399 ;
  assign w401 = ( w331 & w360 ) | ( w331 & w361 ) | ( w360 & w361 ) ;
  assign w402 = w400 ^ w401 ;
  assign w403 = w364 ^ w402 ;
  assign w404 = ( w364 & w400 ) | ( w364 & w401 ) | ( w400 & w401 ) ;
  assign w405 = ( w385 & w386 ) | ( w385 & w398 ) | ( w386 & w398 ) ;
  assign w406 = \pi07 & \pi11 ;
  assign w407 = \pi05 & \pi13 ;
  assign w408 = \pi00 & \pi18 ;
  assign w409 = ( w406 & w407 ) | ( w406 & w408 ) | ( w407 & w408 ) ;
  assign w410 = w406 ^ w408 ;
  assign w411 = w407 ^ w410 ;
  assign w412 = \pi14 & \pi15 ;
  assign w413 = \pi04 & \pi14 ;
  assign w414 = \pi03 & \pi15 ;
  assign w415 = \pi02 & \pi16 ;
  assign w416 = ( w413 & w414 ) | ( w413 & w415 ) | ( w414 & w415 ) ;
  assign w417 = w413 ^ w415 ;
  assign w418 = w414 ^ w417 ;
  assign w419 = \pi01 & w392 ;
  assign w420 = \pi06 & \pi12 ;
  assign w421 = \pi01 & \pi17 ;
  assign w422 = w165 ^ w421 ;
  assign w423 = ( w419 & w420 ) | ( w419 & w422 ) | ( w420 & w422 ) ;
  assign w424 = w165 ^ w420 ;
  assign w425 = \pi17 ^ w392 ;
  assign w426 = \pi01 & w425 ;
  assign w427 = w424 ^ w426 ;
  assign w428 = w411 ^ w427 ;
  assign w429 = w418 ^ w428 ;
  assign w430 = ( w390 & w391 ) | ( w390 & w396 ) | ( w391 & w396 ) ;
  assign w431 = w367 ^ w373 ;
  assign w432 = w381 ^ w431 ;
  assign w433 = \pi09 ^ w393 ;
  assign w434 = ( w335 & w346 ) | ( w335 & w433 ) | ( w346 & w433 ) ;
  assign w435 = ( w369 & w375 ) | ( w369 & w383 ) | ( w375 & w383 ) ;
  assign w436 = w432 ^ w435 ;
  assign w437 = w434 ^ w436 ;
  assign w438 = w430 ^ w437 ;
  assign w439 = w429 ^ w438 ;
  assign w440 = w404 ^ w405 ;
  assign w441 = w439 ^ w440 ;
  assign w442 = \pi08 & \pi11 ;
  assign w443 = \pi03 & \pi16 ;
  assign w444 = ( w217 & w442 ) | ( w217 & w443 ) | ( w442 & w443 ) ;
  assign w445 = w217 ^ w423 ;
  assign w446 = w409 ^ w445 ;
  assign w447 = w442 ^ w446 ;
  assign w448 = w443 ^ w447 ;
  assign w449 = ( w411 & w418 ) | ( w411 & w427 ) | ( w418 & w427 ) ;
  assign w450 = ( \pi01 & ~\pi10 ) | ( \pi01 & \pi18 ) | ( ~\pi10 & \pi18 ) ;
  assign w451 = \pi10 & w450 ;
  assign w452 = ~\pi01 & \pi08 ;
  assign w453 = ( ~\pi08 & \pi17 ) | ( ~\pi08 & w452 ) | ( \pi17 & w452 ) ;
  assign w454 = ( \pi10 & ~\pi17 ) | ( \pi10 & w453 ) | ( ~\pi17 & w453 ) ;
  assign w455 = w416 ^ w454 ;
  assign w456 = \pi01 & \pi18 ;
  assign w457 = w455 ^ w456 ;
  assign w458 = w448 ^ w449 ;
  assign w459 = w457 ^ w458 ;
  assign w460 = \pi15 & \pi17 ;
  assign w461 = \pi04 & \pi15 ;
  assign w462 = \pi02 & \pi17 ;
  assign w463 = \pi00 & \pi19 ;
  assign w464 = ( w461 & w462 ) | ( w461 & w463 ) | ( w462 & w463 ) ;
  assign w465 = w461 ^ w463 ;
  assign w466 = w462 ^ w465 ;
  assign w467 = \pi07 & \pi12 ;
  assign w468 = \pi06 & \pi13 ;
  assign w469 = \pi05 & \pi14 ;
  assign w470 = ( w467 & w468 ) | ( w467 & w469 ) | ( w468 & w469 ) ;
  assign w471 = w467 ^ w469 ;
  assign w472 = w468 ^ w471 ;
  assign w473 = ( w367 & w373 ) | ( w367 & w381 ) | ( w373 & w381 ) ;
  assign w474 = w466 ^ w473 ;
  assign w475 = w472 ^ w474 ;
  assign w476 = ( w432 & w434 ) | ( w432 & w435 ) | ( w434 & w435 ) ;
  assign w477 = w475 ^ w476 ;
  assign w478 = w459 ^ w477 ;
  assign w479 = ( w429 & w430 ) | ( w429 & w437 ) | ( w430 & w437 ) ;
  assign w480 = ( w404 & w405 ) | ( w404 & w439 ) | ( w405 & w439 ) ;
  assign w481 = w478 ^ w480 ;
  assign w482 = w479 ^ w481 ;
  assign w483 = ( w478 & w479 ) | ( w478 & w480 ) | ( w479 & w480 ) ;
  assign w484 = ( w459 & w475 ) | ( w459 & w476 ) | ( w475 & w476 ) ;
  assign w485 = \pi08 & \pi17 ;
  assign w486 = ( ~\pi18 & w416 ) | ( ~\pi18 & w485 ) | ( w416 & w485 ) ;
  assign w487 = \pi10 & w486 ;
  assign w488 = ( \pi01 & \pi10 ) | ( \pi01 & ~\pi18 ) | ( \pi10 & ~\pi18 ) ;
  assign w489 = ( \pi01 & \pi10 ) | ( \pi01 & w416 ) | ( \pi10 & w416 ) ;
  assign w490 = ( w487 & ~w488 ) | ( w487 & w489 ) | ( ~w488 & w489 ) ;
  assign w491 = \pi16 & \pi18 ;
  assign w492 = \pi17 & \pi18 ;
  assign w493 = \pi04 & \pi16 ;
  assign w494 = \pi03 & \pi17 ;
  assign w495 = \pi02 & \pi18 ;
  assign w496 = ( w493 & w494 ) | ( w493 & w495 ) | ( w494 & w495 ) ;
  assign w497 = w493 ^ w495 ;
  assign w498 = w494 ^ w497 ;
  assign w499 = w217 ^ w442 ;
  assign w500 = w443 ^ w499 ;
  assign w501 = ( w409 & w423 ) | ( w409 & w500 ) | ( w423 & w500 ) ;
  assign w502 = w490 ^ w501 ;
  assign w503 = w498 ^ w502 ;
  assign w504 = ( w448 & w449 ) | ( w448 & w457 ) | ( w449 & w457 ) ;
  assign w505 = \pi09 & \pi11 ;
  assign w506 = \pi01 & \pi19 ;
  assign w507 = w464 ^ w505 ;
  assign w508 = w444 ^ w507 ;
  assign w509 = w506 ^ w508 ;
  assign w510 = ( w466 & w472 ) | ( w466 & w473 ) | ( w472 & w473 ) ;
  assign w511 = w509 ^ w510 ;
  assign w512 = \pi00 & \pi20 ;
  assign w513 = \pi07 & \pi13 ;
  assign w514 = w512 ^ w513 ;
  assign w515 = \pi08 & \pi12 ;
  assign w516 = \pi06 & \pi14 ;
  assign w517 = \pi05 & \pi15 ;
  assign w518 = ( w515 & w516 ) | ( w515 & w517 ) | ( w516 & w517 ) ;
  assign w519 = w515 ^ w517 ;
  assign w520 = w516 ^ w519 ;
  assign w521 = w514 ^ w520 ;
  assign w522 = w451 ^ w521 ;
  assign w523 = w470 ^ w522 ;
  assign w524 = w504 ^ w523 ;
  assign w525 = w511 ^ w524 ;
  assign w526 = w503 ^ w525 ;
  assign w527 = w483 ^ w526 ;
  assign w528 = w484 ^ w527 ;
  assign w529 = w511 ^ w523 ;
  assign w530 = ( w503 & w504 ) | ( w503 & w529 ) | ( w504 & w529 ) ;
  assign w531 = ( w451 & w512 ) | ( w451 & w513 ) | ( w512 & w513 ) ;
  assign w532 = w496 ^ w531 ;
  assign w533 = w518 ^ w532 ;
  assign w534 = ( w490 & w498 ) | ( w490 & w501 ) | ( w498 & w501 ) ;
  assign w535 = \pi05 & \pi16 ;
  assign w536 = \pi03 & \pi18 ;
  assign w537 = \pi02 & \pi19 ;
  assign w538 = ( w535 & w536 ) | ( w535 & w537 ) | ( w536 & w537 ) ;
  assign w539 = w535 ^ w537 ;
  assign w540 = w536 ^ w539 ;
  assign w541 = \pi08 & \pi13 ;
  assign w542 = \pi07 & \pi14 ;
  assign w543 = \pi06 & \pi15 ;
  assign w544 = ( w541 & w542 ) | ( w541 & w543 ) | ( w542 & w543 ) ;
  assign w545 = w541 ^ w543 ;
  assign w546 = w542 ^ w545 ;
  assign w547 = \pi04 & \pi17 ;
  assign w548 = \pi10 & \pi11 ;
  assign w549 = \pi09 & \pi12 ;
  assign w550 = ( w547 & w548 ) | ( w547 & w549 ) | ( w548 & w549 ) ;
  assign w551 = w547 ^ w549 ;
  assign w552 = w548 ^ w551 ;
  assign w553 = w540 ^ w552 ;
  assign w554 = w546 ^ w553 ;
  assign w555 = w533 ^ w534 ;
  assign w556 = w554 ^ w555 ;
  assign w557 = w505 ^ w506 ;
  assign w558 = ( w444 & w464 ) | ( w444 & w557 ) | ( w464 & w557 ) ;
  assign w559 = \pi00 & \pi21 ;
  assign w560 = \pi01 & w505 ;
  assign w561 = \pi19 & w560 ;
  assign w562 = w559 ^ w561 ;
  assign w563 = w451 ^ w514 ;
  assign w564 = ( w470 & w520 ) | ( w470 & w563 ) | ( w520 & w563 ) ;
  assign w565 = w558 ^ w562 ;
  assign w566 = w564 ^ w565 ;
  assign w567 = \pi11 ^ w566 ;
  assign w568 = \pi01 & \pi20 ;
  assign w569 = w567 ^ w568 ;
  assign w570 = ( w509 & w510 ) | ( w509 & w523 ) | ( w510 & w523 ) ;
  assign w571 = w556 ^ w570 ;
  assign w572 = w569 ^ w571 ;
  assign w573 = ( w483 & w484 ) | ( w483 & w526 ) | ( w484 & w526 ) ;
  assign w574 = w530 ^ w573 ;
  assign w575 = w572 ^ w574 ;
  assign w576 = ( w530 & w572 ) | ( w530 & w573 ) | ( w572 & w573 ) ;
  assign w577 = ( w556 & w569 ) | ( w556 & w570 ) | ( w569 & w570 ) ;
  assign w578 = \pi09 & \pi19 ;
  assign w579 = ( ~\pi20 & w559 ) | ( ~\pi20 & w578 ) | ( w559 & w578 ) ;
  assign w580 = \pi11 & w579 ;
  assign w581 = ( \pi01 & \pi11 ) | ( \pi01 & ~\pi20 ) | ( \pi11 & ~\pi20 ) ;
  assign w582 = ( \pi01 & \pi11 ) | ( \pi01 & w559 ) | ( \pi11 & w559 ) ;
  assign w583 = ( w580 & ~w581 ) | ( w580 & w582 ) | ( ~w581 & w582 ) ;
  assign w584 = w538 ^ w583 ;
  assign w585 = w544 ^ w584 ;
  assign w586 = \pi11 ^ w562 ;
  assign w587 = w568 ^ w586 ;
  assign w588 = ( w558 & w564 ) | ( w558 & w587 ) | ( w564 & w587 ) ;
  assign w589 = \pi08 & \pi14 ;
  assign w590 = \pi07 & \pi15 ;
  assign w591 = \pi00 & \pi22 ;
  assign w592 = ( w589 & w590 ) | ( w589 & w591 ) | ( w590 & w591 ) ;
  assign w593 = w589 ^ w591 ;
  assign w594 = w590 ^ w593 ;
  assign w595 = \pi09 & \pi13 ;
  assign w596 = \pi02 & \pi20 ;
  assign w597 = ( w332 & w595 ) | ( w332 & w596 ) | ( w595 & w596 ) ;
  assign w598 = w332 ^ w596 ;
  assign w599 = w595 ^ w598 ;
  assign w600 = \pi05 & \pi17 ;
  assign w601 = \pi04 & \pi18 ;
  assign w602 = \pi03 & \pi19 ;
  assign w603 = ( w600 & w601 ) | ( w600 & w602 ) | ( w601 & w602 ) ;
  assign w604 = w600 ^ w602 ;
  assign w605 = w601 ^ w604 ;
  assign w606 = w594 ^ w599 ;
  assign w607 = w605 ^ w606 ;
  assign w608 = w585 ^ w588 ;
  assign w609 = w607 ^ w608 ;
  assign w610 = ( w533 & w534 ) | ( w533 & w554 ) | ( w534 & w554 ) ;
  assign w611 = ( w540 & w546 ) | ( w540 & w552 ) | ( w546 & w552 ) ;
  assign w612 = ( w496 & w518 ) | ( w496 & w531 ) | ( w518 & w531 ) ;
  assign w613 = ( ~\pi01 & \pi11 ) | ( ~\pi01 & \pi20 ) | ( \pi11 & \pi20 ) ;
  assign w614 = \pi21 ^ w613 ;
  assign w615 = \pi01 & w614 ;
  assign w616 = w216 ^ w550 ;
  assign w617 = w615 ^ w616 ;
  assign w618 = w611 ^ w612 ;
  assign w619 = w617 ^ w618 ;
  assign w620 = w609 ^ w610 ;
  assign w621 = w619 ^ w620 ;
  assign w622 = w577 & w621 ;
  assign w623 = w577 | w621 ;
  assign w624 = ~w622 & w623 ;
  assign w625 = w576 ^ w624 ;
  assign w626 = ( w609 & w610 ) | ( w609 & w619 ) | ( w610 & w619 ) ;
  assign w627 = ( w611 & w612 ) | ( w611 & w617 ) | ( w612 & w617 ) ;
  assign w628 = \pi06 & \pi17 ;
  assign w629 = \pi05 & \pi18 ;
  assign w630 = \pi03 & \pi20 ;
  assign w631 = ( w628 & w629 ) | ( w628 & w630 ) | ( w629 & w630 ) ;
  assign w632 = w628 ^ w630 ;
  assign w633 = w629 ^ w632 ;
  assign w634 = \pi11 & \pi12 ;
  assign w635 = \pi10 & \pi13 ;
  assign w636 = \pi04 & \pi19 ;
  assign w637 = ( w634 & w635 ) | ( w634 & w636 ) | ( w635 & w636 ) ;
  assign w638 = w634 ^ w636 ;
  assign w639 = w635 ^ w638 ;
  assign w640 = \pi20 & w229 ;
  assign w641 = \pi01 & \pi21 ;
  assign w642 = w216 ^ w641 ;
  assign w643 = ( w550 & w640 ) | ( w550 & w642 ) | ( w640 & w642 ) ;
  assign w644 = w633 ^ w643 ;
  assign w645 = w639 ^ w644 ;
  assign w646 = \pi21 & \pi23 ;
  assign w647 = ( \pi00 & ~\pi21 ) | ( \pi00 & \pi23 ) | ( ~\pi21 & \pi23 ) ;
  assign w648 = ( \pi01 & ~\pi21 ) | ( \pi01 & w216 ) | ( ~\pi21 & w216 ) ;
  assign w649 = ( \pi02 & w647 ) | ( \pi02 & w648 ) | ( w647 & w648 ) ;
  assign w650 = \pi21 & w649 ;
  assign w651 = \pi00 & \pi23 ;
  assign w652 = \pi02 ^ w648 ;
  assign w653 = \pi21 & w652 ;
  assign w654 = w651 ^ w653 ;
  assign w655 = \pi09 & \pi14 ;
  assign w656 = \pi08 & \pi15 ;
  assign w657 = \pi07 & \pi16 ;
  assign w658 = ( w655 & w656 ) | ( w655 & w657 ) | ( w656 & w657 ) ;
  assign w659 = w655 ^ w657 ;
  assign w660 = w656 ^ w659 ;
  assign w661 = w592 ^ w654 ;
  assign w662 = w660 ^ w661 ;
  assign w663 = w627 ^ w645 ;
  assign w664 = w662 ^ w663 ;
  assign w665 = ( w585 & w588 ) | ( w585 & w607 ) | ( w588 & w607 ) ;
  assign w666 = ( w538 & w544 ) | ( w538 & w583 ) | ( w544 & w583 ) ;
  assign w667 = ( w594 & w599 ) | ( w594 & w605 ) | ( w599 & w605 ) ;
  assign w668 = \pi01 & \pi22 ;
  assign w669 = \pi12 ^ w603 ;
  assign w670 = w597 ^ w669 ;
  assign w671 = w668 ^ w670 ;
  assign w672 = w666 ^ w667 ;
  assign w673 = w671 ^ w672 ;
  assign w674 = w664 ^ w665 ;
  assign w675 = w673 ^ w674 ;
  assign w676 = ( w576 & w622 ) | ( w576 & w623 ) | ( w622 & w623 ) ;
  assign w677 = w622 | w676 ;
  assign w678 = w626 ^ w677 ;
  assign w679 = w675 ^ w678 ;
  assign w680 = ( w626 & w675 ) | ( w626 & w677 ) | ( w675 & w677 ) ;
  assign w681 = ( w664 & w665 ) | ( w664 & w673 ) | ( w665 & w673 ) ;
  assign w682 = ( w627 & w645 ) | ( w627 & w662 ) | ( w645 & w662 ) ;
  assign w683 = w631 ^ w637 ;
  assign w684 = w658 ^ w683 ;
  assign w685 = ( w633 & w639 ) | ( w633 & w643 ) | ( w639 & w643 ) ;
  assign w686 = ( w592 & w654 ) | ( w592 & w660 ) | ( w654 & w660 ) ;
  assign w687 = w685 ^ w686 ;
  assign w688 = w684 ^ w687 ;
  assign w689 = \pi00 & \pi24 ;
  assign w690 = ( \pi01 & \pi12 ) | ( \pi01 & ~\pi22 ) | ( \pi12 & ~\pi22 ) ;
  assign w691 = \pi22 & w690 ;
  assign w692 = w689 ^ w691 ;
  assign w693 = ( ~\pi01 & \pi23 ) | ( ~\pi01 & w376 ) | ( \pi23 & w376 ) ;
  assign w694 = \pi01 & w693 ;
  assign w695 = \pi01 & \pi23 ;
  assign w696 = w376 ^ w695 ;
  assign w697 = \pi18 & \pi22 ;
  assign w698 = \pi07 & \pi17 ;
  assign w699 = \pi06 & \pi18 ;
  assign w700 = \pi02 & \pi22 ;
  assign w701 = ( w698 & w699 ) | ( w698 & w700 ) | ( w699 & w700 ) ;
  assign w702 = w698 ^ w700 ;
  assign w703 = w699 ^ w702 ;
  assign w704 = \pi12 ^ w668 ;
  assign w705 = ( w597 & w603 ) | ( w597 & w704 ) | ( w603 & w704 ) ;
  assign w706 = w692 ^ w703 ;
  assign w707 = w705 ^ w706 ;
  assign w708 = w696 ^ w707 ;
  assign w709 = \pi19 & \pi21 ;
  assign w710 = \pi20 & \pi21 ;
  assign w711 = \pi05 & \pi19 ;
  assign w712 = \pi04 & \pi20 ;
  assign w713 = \pi03 & \pi21 ;
  assign w714 = ( w711 & w712 ) | ( w711 & w713 ) | ( w712 & w713 ) ;
  assign w715 = w711 ^ w713 ;
  assign w716 = w712 ^ w715 ;
  assign w717 = \pi10 & \pi14 ;
  assign w718 = \pi09 & \pi15 ;
  assign w719 = \pi08 & \pi16 ;
  assign w720 = ( w717 & w718 ) | ( w717 & w719 ) | ( w718 & w719 ) ;
  assign w721 = w717 ^ w719 ;
  assign w722 = w718 ^ w721 ;
  assign w723 = w650 ^ w716 ;
  assign w724 = w722 ^ w723 ;
  assign w725 = ( w666 & w667 ) | ( w666 & w671 ) | ( w667 & w671 ) ;
  assign w726 = w708 ^ w725 ;
  assign w727 = w724 ^ w726 ;
  assign w728 = w682 ^ w688 ;
  assign w729 = w727 ^ w728 ;
  assign w730 = w681 & w729 ;
  assign w731 = w681 | w729 ;
  assign w732 = ~w730 & w731 ;
  assign w733 = w680 ^ w732 ;
  assign w734 = ( w682 & w688 ) | ( w682 & w727 ) | ( w688 & w727 ) ;
  assign w735 = \pi02 & \pi23 ;
  assign w736 = \pi00 & \pi25 ;
  assign w737 = ( w317 & w735 ) | ( w317 & w736 ) | ( w735 & w736 ) ;
  assign w738 = w317 ^ w736 ;
  assign w739 = w735 ^ w738 ;
  assign w740 = \pi07 & \pi18 ;
  assign w741 = ( w392 & w485 ) | ( w392 & w740 ) | ( w485 & w740 ) ;
  assign w742 = w392 ^ w740 ;
  assign w743 = w485 ^ w742 ;
  assign w744 = \pi06 & \pi19 ;
  assign w745 = \pi04 & \pi21 ;
  assign w746 = \pi03 & \pi22 ;
  assign w747 = ( w744 & w745 ) | ( w744 & w746 ) | ( w745 & w746 ) ;
  assign w748 = w744 ^ w746 ;
  assign w749 = w745 ^ w748 ;
  assign w750 = w739 ^ w743 ;
  assign w751 = w749 ^ w750 ;
  assign w752 = ( w684 & w685 ) | ( w684 & w686 ) | ( w685 & w686 ) ;
  assign w753 = ( \pi01 & ~\pi13 ) | ( \pi01 & \pi24 ) | ( ~\pi13 & \pi24 ) ;
  assign w754 = \pi13 & w753 ;
  assign w755 = \pi01 & \pi24 ;
  assign w756 = \pi13 ^ w714 ;
  assign w757 = w694 ^ w756 ;
  assign w758 = w755 ^ w757 ;
  assign w759 = ( w631 & w637 ) | ( w631 & w658 ) | ( w637 & w658 ) ;
  assign w760 = \pi11 & \pi14 ;
  assign w761 = \pi05 & \pi20 ;
  assign w762 = ( w342 & w760 ) | ( w342 & w761 ) | ( w760 & w761 ) ;
  assign w763 = w342 ^ w761 ;
  assign w764 = w760 ^ w763 ;
  assign w765 = w758 ^ w759 ;
  assign w766 = w764 ^ w765 ;
  assign w767 = w752 ^ w766 ;
  assign w768 = w751 ^ w767 ;
  assign w769 = ( \pi01 & ~\pi12 ) | ( \pi01 & \pi22 ) | ( ~\pi12 & \pi22 ) ;
  assign w770 = \pi12 & w769 ;
  assign w771 = ( w689 & w696 ) | ( w689 & w770 ) | ( w696 & w770 ) ;
  assign w772 = w701 ^ w771 ;
  assign w773 = w720 ^ w772 ;
  assign w774 = ( w650 & w716 ) | ( w650 & w722 ) | ( w716 & w722 ) ;
  assign w775 = w692 ^ w696 ;
  assign w776 = ( w703 & w705 ) | ( w703 & w775 ) | ( w705 & w775 ) ;
  assign w777 = w773 ^ w776 ;
  assign w778 = w774 ^ w777 ;
  assign w779 = ( w708 & w724 ) | ( w708 & w725 ) | ( w724 & w725 ) ;
  assign w780 = w768 ^ w778 ;
  assign w781 = w779 ^ w780 ;
  assign w782 = ( w680 & w730 ) | ( w680 & w731 ) | ( w730 & w731 ) ;
  assign w783 = w730 | w782 ;
  assign w784 = w781 ^ w783 ;
  assign w785 = w734 ^ w784 ;
  assign w786 = ( w768 & w778 ) | ( w768 & w779 ) | ( w778 & w779 ) ;
  assign w787 = \pi07 & \pi19 ;
  assign w788 = \pi03 & \pi23 ;
  assign w789 = \pi02 & \pi24 ;
  assign w790 = ( w787 & w788 ) | ( w787 & w789 ) | ( w788 & w789 ) ;
  assign w791 = w787 ^ w789 ;
  assign w792 = w788 ^ w791 ;
  assign w793 = \pi11 & \pi15 ;
  assign w794 = \pi10 & \pi16 ;
  assign w795 = \pi09 & \pi17 ;
  assign w796 = ( w793 & w794 ) | ( w793 & w795 ) | ( w794 & w795 ) ;
  assign w797 = w793 ^ w795 ;
  assign w798 = w794 ^ w797 ;
  assign w799 = \pi06 & \pi20 ;
  assign w800 = \pi05 & \pi21 ;
  assign w801 = \pi04 & \pi22 ;
  assign w802 = ( w799 & w800 ) | ( w799 & w801 ) | ( w800 & w801 ) ;
  assign w803 = w799 ^ w801 ;
  assign w804 = w800 ^ w803 ;
  assign w805 = w792 ^ w798 ;
  assign w806 = w804 ^ w805 ;
  assign w807 = ( w773 & w774 ) | ( w773 & w776 ) | ( w774 & w776 ) ;
  assign w808 = ( w701 & w720 ) | ( w701 & w771 ) | ( w720 & w771 ) ;
  assign w809 = \pi13 ^ w755 ;
  assign w810 = ( w694 & w714 ) | ( w694 & w809 ) | ( w714 & w809 ) ;
  assign w811 = w808 ^ w810 ;
  assign w812 = \pi08 & \pi18 ;
  assign w813 = \pi00 & \pi26 ;
  assign w814 = ( w754 & w812 ) | ( w754 & w813 ) | ( w812 & w813 ) ;
  assign w815 = w754 ^ w813 ;
  assign w816 = w812 ^ w815 ;
  assign w817 = w737 ^ w816 ;
  assign w818 = w741 ^ w817 ;
  assign w819 = w806 ^ w818 ;
  assign w820 = w807 ^ w819 ;
  assign w821 = w811 ^ w820 ;
  assign w822 = ( w751 & w752 ) | ( w751 & w766 ) | ( w752 & w766 ) ;
  assign w823 = ( w758 & w759 ) | ( w758 & w764 ) | ( w759 & w764 ) ;
  assign w824 = ( w739 & w743 ) | ( w739 & w749 ) | ( w743 & w749 ) ;
  assign w825 = \pi01 & \pi25 ;
  assign w826 = ( ~\pi12 & \pi14 ) | ( ~\pi12 & w825 ) | ( \pi14 & w825 ) ;
  assign w827 = \pi12 & w826 ;
  assign w828 = \pi12 & \pi14 ;
  assign w829 = w747 ^ w825 ;
  assign w830 = w762 ^ w829 ;
  assign w831 = w828 ^ w830 ;
  assign w832 = w823 ^ w824 ;
  assign w833 = w831 ^ w832 ;
  assign w834 = w821 ^ w822 ;
  assign w835 = w833 ^ w834 ;
  assign w836 = ( w734 & w781 ) | ( w734 & w783 ) | ( w781 & w783 ) ;
  assign w837 = w786 ^ w836 ;
  assign w838 = w835 ^ w837 ;
  assign w839 = ( w821 & w822 ) | ( w821 & w833 ) | ( w822 & w833 ) ;
  assign w840 = w811 ^ w818 ;
  assign w841 = ( w806 & w807 ) | ( w806 & w840 ) | ( w807 & w840 ) ;
  assign w842 = \pi06 & \pi21 ;
  assign w843 = \pi04 & \pi23 ;
  assign w844 = \pi03 & \pi24 ;
  assign w845 = ( w842 & w843 ) | ( w842 & w844 ) | ( w843 & w844 ) ;
  assign w846 = w842 ^ w844 ;
  assign w847 = w843 ^ w846 ;
  assign w848 = \pi13 & \pi14 ;
  assign w849 = \pi12 & \pi15 ;
  assign w850 = \pi05 & \pi22 ;
  assign w851 = ( w848 & w849 ) | ( w848 & w850 ) | ( w849 & w850 ) ;
  assign w852 = w848 ^ w850 ;
  assign w853 = w849 ^ w852 ;
  assign w854 = \pi01 & \pi26 ;
  assign w855 = w827 ^ w854 ;
  assign w856 = \pi14 ^ w855 ;
  assign w857 = \pi00 & \pi27 ;
  assign w858 = w856 ^ w857 ;
  assign w859 = w847 ^ w858 ;
  assign w860 = w853 ^ w859 ;
  assign w861 = w790 ^ w796 ;
  assign w862 = w802 ^ w861 ;
  assign w863 = ( w808 & w810 ) | ( w808 & w818 ) | ( w810 & w818 ) ;
  assign w864 = w860 ^ w863 ;
  assign w865 = w862 ^ w864 ;
  assign w866 = \pi02 & \pi25 ;
  assign w867 = \pi11 & \pi16 ;
  assign w868 = w866 ^ w867 ;
  assign w869 = \pi07 & \pi20 ;
  assign w870 = w868 ^ w869 ;
  assign w871 = \pi10 & \pi17 ;
  assign w872 = \pi09 & \pi18 ;
  assign w873 = \pi08 & \pi19 ;
  assign w874 = ( w871 & w872 ) | ( w871 & w873 ) | ( w872 & w873 ) ;
  assign w875 = w871 ^ w873 ;
  assign w876 = w872 ^ w875 ;
  assign w877 = w814 ^ w870 ;
  assign w878 = w876 ^ w877 ;
  assign w879 = ( w823 & w824 ) | ( w823 & w831 ) | ( w824 & w831 ) ;
  assign w880 = w825 ^ w828 ;
  assign w881 = ( w747 & w762 ) | ( w747 & w880 ) | ( w762 & w880 ) ;
  assign w882 = ( w737 & w741 ) | ( w737 & w816 ) | ( w741 & w816 ) ;
  assign w883 = ( w792 & w798 ) | ( w792 & w804 ) | ( w798 & w804 ) ;
  assign w884 = w881 ^ w882 ;
  assign w885 = w883 ^ w884 ;
  assign w886 = w879 ^ w885 ;
  assign w887 = w878 ^ w886 ;
  assign w888 = w841 ^ w865 ;
  assign w889 = w887 ^ w888 ;
  assign w890 = ( w786 & w835 ) | ( w786 & w836 ) | ( w835 & w836 ) ;
  assign w891 = w839 ^ w890 ;
  assign w892 = w889 ^ w891 ;
  assign w893 = ( w860 & w862 ) | ( w860 & w863 ) | ( w862 & w863 ) ;
  assign w894 = \pi24 & \pi25 ;
  assign w895 = \pi08 & \pi20 ;
  assign w896 = \pi04 & \pi24 ;
  assign w897 = \pi03 & \pi25 ;
  assign w898 = ( w895 & w896 ) | ( w895 & w897 ) | ( w896 & w897 ) ;
  assign w899 = w895 ^ w897 ;
  assign w900 = w896 ^ w899 ;
  assign w901 = \pi14 ^ w854 ;
  assign w902 = ( w827 & w857 ) | ( w827 & w901 ) | ( w857 & w901 ) ;
  assign w903 = \pi07 & \pi21 ;
  assign w904 = \pi06 & \pi22 ;
  assign w905 = \pi05 & \pi23 ;
  assign w906 = ( w903 & w904 ) | ( w903 & w905 ) | ( w904 & w905 ) ;
  assign w907 = w903 ^ w905 ;
  assign w908 = w904 ^ w907 ;
  assign w909 = w900 ^ w902 ;
  assign w910 = w908 ^ w909 ;
  assign w911 = ( w847 & w853 ) | ( w847 & w858 ) | ( w853 & w858 ) ;
  assign w912 = ( w814 & w870 ) | ( w814 & w876 ) | ( w870 & w876 ) ;
  assign w913 = ( ~\pi01 & \pi14 ) | ( ~\pi01 & \pi26 ) | ( \pi14 & \pi26 ) ;
  assign w914 = \pi27 ^ w913 ;
  assign w915 = \pi01 & w914 ;
  assign w916 = w377 ^ w851 ;
  assign w917 = w915 ^ w916 ;
  assign w918 = w911 ^ w912 ;
  assign w919 = w917 ^ w918 ;
  assign w920 = w893 ^ w919 ;
  assign w921 = w910 ^ w920 ;
  assign w922 = ( w841 & w865 ) | ( w841 & w887 ) | ( w865 & w887 ) ;
  assign w923 = ( w878 & w879 ) | ( w878 & w885 ) | ( w879 & w885 ) ;
  assign w924 = ( w866 & w867 ) | ( w866 & w869 ) | ( w867 & w869 ) ;
  assign w925 = w845 ^ w874 ;
  assign w926 = w924 ^ w925 ;
  assign w927 = ( w881 & w882 ) | ( w881 & w883 ) | ( w882 & w883 ) ;
  assign w928 = \pi12 & \pi16 ;
  assign w929 = \pi11 & \pi17 ;
  assign w930 = \pi00 & \pi28 ;
  assign w931 = ( w928 & w929 ) | ( w928 & w930 ) | ( w929 & w930 ) ;
  assign w932 = w928 ^ w930 ;
  assign w933 = w929 ^ w932 ;
  assign w934 = \pi10 & \pi18 ;
  assign w935 = \pi02 & \pi26 ;
  assign w936 = ( w578 & w934 ) | ( w578 & w935 ) | ( w934 & w935 ) ;
  assign w937 = w934 ^ w935 ;
  assign w938 = w578 ^ w937 ;
  assign w939 = ( w790 & w796 ) | ( w790 & w802 ) | ( w796 & w802 ) ;
  assign w940 = w933 ^ w939 ;
  assign w941 = w938 ^ w940 ;
  assign w942 = w927 ^ w941 ;
  assign w943 = w926 ^ w942 ;
  assign w944 = w922 ^ w923 ;
  assign w945 = w943 ^ w944 ;
  assign w946 = ( w839 & w889 ) | ( w839 & w890 ) | ( w889 & w890 ) ;
  assign w947 = w945 ^ w946 ;
  assign w948 = w921 ^ w947 ;
  assign w949 = ( w922 & w923 ) | ( w922 & w943 ) | ( w923 & w943 ) ;
  assign w950 = ( w926 & w927 ) | ( w926 & w941 ) | ( w927 & w941 ) ;
  assign w951 = ( w911 & w912 ) | ( w911 & w917 ) | ( w912 & w917 ) ;
  assign w952 = ( w933 & w938 ) | ( w933 & w939 ) | ( w938 & w939 ) ;
  assign w953 = ( w900 & w902 ) | ( w900 & w908 ) | ( w902 & w908 ) ;
  assign w954 = w952 ^ w953 ;
  assign w955 = ( \pi00 & ~\pi27 ) | ( \pi00 & \pi29 ) | ( ~\pi27 & \pi29 ) ;
  assign w956 = ( \pi01 & ~\pi27 ) | ( \pi01 & w377 ) | ( ~\pi27 & w377 ) ;
  assign w957 = ( \pi02 & w955 ) | ( \pi02 & w956 ) | ( w955 & w956 ) ;
  assign w958 = \pi27 & w957 ;
  assign w959 = \pi00 & \pi29 ;
  assign w960 = \pi02 ^ w956 ;
  assign w961 = \pi27 & w960 ;
  assign w962 = w959 ^ w961 ;
  assign w963 = w931 ^ w962 ;
  assign w964 = w936 ^ w963 ;
  assign w965 = w954 ^ w964 ;
  assign w966 = w950 ^ w965 ;
  assign w967 = w951 ^ w966 ;
  assign w968 = ( w893 & w910 ) | ( w893 & w919 ) | ( w910 & w919 ) ;
  assign w969 = \pi26 & w301 ;
  assign w970 = \pi01 & \pi27 ;
  assign w971 = w377 ^ w970 ;
  assign w972 = ( w851 & w969 ) | ( w851 & w971 ) | ( w969 & w971 ) ;
  assign w973 = \pi13 & \pi16 ;
  assign w974 = \pi06 & \pi23 ;
  assign w975 = ( w412 & w973 ) | ( w412 & w974 ) | ( w973 & w974 ) ;
  assign w976 = w412 ^ w974 ;
  assign w977 = w973 ^ w976 ;
  assign w978 = ( w845 & w874 ) | ( w845 & w924 ) | ( w874 & w924 ) ;
  assign w979 = w972 ^ w977 ;
  assign w980 = w978 ^ w979 ;
  assign w981 = \pi12 & \pi17 ;
  assign w982 = \pi08 & \pi21 ;
  assign w983 = \pi03 & \pi26 ;
  assign w984 = ( w981 & w982 ) | ( w981 & w983 ) | ( w982 & w983 ) ;
  assign w985 = w981 ^ w983 ;
  assign w986 = w982 ^ w985 ;
  assign w987 = \pi11 & \pi18 ;
  assign w988 = \pi10 & \pi19 ;
  assign w989 = \pi09 & \pi20 ;
  assign w990 = ( w987 & w988 ) | ( w987 & w989 ) | ( w988 & w989 ) ;
  assign w991 = w987 ^ w989 ;
  assign w992 = w988 ^ w991 ;
  assign w993 = \pi22 & \pi24 ;
  assign w994 = \pi07 & \pi22 ;
  assign w995 = \pi05 & \pi24 ;
  assign w996 = \pi04 & \pi25 ;
  assign w997 = ( w994 & w995 ) | ( w994 & w996 ) | ( w995 & w996 ) ;
  assign w998 = w994 ^ w996 ;
  assign w999 = w995 ^ w998 ;
  assign w1000 = w986 ^ w992 ;
  assign w1001 = w999 ^ w1000 ;
  assign w1002 = \pi01 & \pi28 ;
  assign w1003 = \pi15 ^ w906 ;
  assign w1004 = w898 ^ w1003 ;
  assign w1005 = w1002 ^ w1004 ;
  assign w1006 = w980 ^ w1001 ;
  assign w1007 = w1005 ^ w1006 ;
  assign w1008 = w967 ^ w968 ;
  assign w1009 = w1007 ^ w1008 ;
  assign w1010 = ( w921 & w945 ) | ( w921 & w946 ) | ( w945 & w946 ) ;
  assign w1011 = w949 ^ w1010 ;
  assign w1012 = w1009 ^ w1011 ;
  assign w1013 = ( w967 & w968 ) | ( w967 & w1007 ) | ( w968 & w1007 ) ;
  assign w1014 = \pi00 & \pi30 ;
  assign w1015 = ( \pi01 & \pi15 ) | ( \pi01 & ~\pi28 ) | ( \pi15 & ~\pi28 ) ;
  assign w1016 = \pi28 & w1015 ;
  assign w1017 = w1014 ^ w1016 ;
  assign w1018 = \pi01 & \pi29 ;
  assign w1019 = \pi14 & \pi16 ;
  assign w1020 = w1018 ^ w1019 ;
  assign w1021 = \pi15 ^ w1002 ;
  assign w1022 = ( w898 & w906 ) | ( w898 & w1021 ) | ( w906 & w1021 ) ;
  assign w1023 = ( w931 & w936 ) | ( w931 & w962 ) | ( w936 & w962 ) ;
  assign w1024 = w1017 ^ w1020 ;
  assign w1025 = w1023 ^ w1024 ;
  assign w1026 = w1022 ^ w1025 ;
  assign w1027 = ( w980 & w1001 ) | ( w980 & w1005 ) | ( w1001 & w1005 ) ;
  assign w1028 = \pi13 & \pi17 ;
  assign w1029 = \pi09 & \pi21 ;
  assign w1030 = \pi02 & \pi28 ;
  assign w1031 = ( w1028 & w1029 ) | ( w1028 & w1030 ) | ( w1029 & w1030 ) ;
  assign w1032 = w1028 ^ w1030 ;
  assign w1033 = w1029 ^ w1032 ;
  assign w1034 = w975 ^ w997 ;
  assign w1035 = w1033 ^ w1034 ;
  assign w1036 = ( w986 & w992 ) | ( w986 & w999 ) | ( w992 & w999 ) ;
  assign w1037 = w958 ^ w984 ;
  assign w1038 = w990 ^ w1037 ;
  assign w1039 = w1035 ^ w1038 ;
  assign w1040 = w1036 ^ w1039 ;
  assign w1041 = w1026 ^ w1027 ;
  assign w1042 = w1040 ^ w1041 ;
  assign w1043 = ( w950 & w951 ) | ( w950 & w965 ) | ( w951 & w965 ) ;
  assign w1044 = \pi08 & \pi22 ;
  assign w1045 = \pi04 & \pi26 ;
  assign w1046 = \pi03 & \pi27 ;
  assign w1047 = ( w1044 & w1045 ) | ( w1044 & w1046 ) | ( w1045 & w1046 ) ;
  assign w1048 = w1044 ^ w1046 ;
  assign w1049 = w1045 ^ w1048 ;
  assign w1050 = \pi07 & \pi23 ;
  assign w1051 = \pi06 & \pi24 ;
  assign w1052 = \pi05 & \pi25 ;
  assign w1053 = ( w1050 & w1051 ) | ( w1050 & w1052 ) | ( w1051 & w1052 ) ;
  assign w1054 = w1050 ^ w1052 ;
  assign w1055 = w1051 ^ w1054 ;
  assign w1056 = \pi12 & \pi18 ;
  assign w1057 = \pi11 & \pi19 ;
  assign w1058 = \pi10 & \pi20 ;
  assign w1059 = ( w1056 & w1057 ) | ( w1056 & w1058 ) | ( w1057 & w1058 ) ;
  assign w1060 = w1056 ^ w1058 ;
  assign w1061 = w1057 ^ w1060 ;
  assign w1062 = w1049 ^ w1055 ;
  assign w1063 = w1061 ^ w1062 ;
  assign w1064 = ( w972 & w977 ) | ( w972 & w978 ) | ( w977 & w978 ) ;
  assign w1065 = ( w952 & w953 ) | ( w952 & w964 ) | ( w953 & w964 ) ;
  assign w1066 = w1064 ^ w1065 ;
  assign w1067 = w1063 ^ w1066 ;
  assign w1068 = w1043 ^ w1067 ;
  assign w1069 = w1042 ^ w1068 ;
  assign w1070 = ( w949 & w1009 ) | ( w949 & w1010 ) | ( w1009 & w1010 ) ;
  assign w1071 = w1013 ^ w1070 ;
  assign w1072 = w1069 ^ w1071 ;
  assign w1073 = ( w1042 & w1043 ) | ( w1042 & w1067 ) | ( w1043 & w1067 ) ;
  assign w1074 = ( w1026 & w1027 ) | ( w1026 & w1040 ) | ( w1027 & w1040 ) ;
  assign w1075 = ( w1035 & w1036 ) | ( w1035 & w1038 ) | ( w1036 & w1038 ) ;
  assign w1076 = \pi08 & \pi23 ;
  assign w1077 = \pi07 & \pi24 ;
  assign w1078 = \pi05 & \pi26 ;
  assign w1079 = ( w1076 & w1077 ) | ( w1076 & w1078 ) | ( w1077 & w1078 ) ;
  assign w1080 = w1076 ^ w1078 ;
  assign w1081 = w1077 ^ w1080 ;
  assign w1082 = \pi15 & \pi16 ;
  assign w1083 = \pi14 & \pi17 ;
  assign w1084 = \pi06 & \pi25 ;
  assign w1085 = ( w1082 & w1083 ) | ( w1082 & w1084 ) | ( w1083 & w1084 ) ;
  assign w1086 = w1082 ^ w1084 ;
  assign w1087 = w1083 ^ w1086 ;
  assign w1088 = \pi27 & \pi28 ;
  assign w1089 = \pi04 & \pi27 ;
  assign w1090 = \pi03 & \pi28 ;
  assign w1091 = \pi02 & \pi29 ;
  assign w1092 = ( w1089 & w1090 ) | ( w1089 & w1091 ) | ( w1090 & w1091 ) ;
  assign w1093 = w1089 ^ w1091 ;
  assign w1094 = w1090 ^ w1093 ;
  assign w1095 = w1081 ^ w1087 ;
  assign w1096 = w1094 ^ w1095 ;
  assign w1097 = \pi10 & \pi21 ;
  assign w1098 = \pi09 & \pi22 ;
  assign w1099 = \pi00 & \pi31 ;
  assign w1100 = ( w1097 & w1098 ) | ( w1097 & w1099 ) | ( w1098 & w1099 ) ;
  assign w1101 = w1097 ^ w1099 ;
  assign w1102 = w1098 ^ w1101 ;
  assign w1103 = ( \pi01 & ~\pi15 ) | ( \pi01 & \pi28 ) | ( ~\pi15 & \pi28 ) ;
  assign w1104 = \pi15 & w1103 ;
  assign w1105 = ( w1014 & w1020 ) | ( w1014 & w1104 ) | ( w1020 & w1104 ) ;
  assign w1106 = \pi13 & \pi18 ;
  assign w1107 = \pi12 & \pi19 ;
  assign w1108 = \pi11 & \pi20 ;
  assign w1109 = ( w1106 & w1107 ) | ( w1106 & w1108 ) | ( w1107 & w1108 ) ;
  assign w1110 = w1106 ^ w1108 ;
  assign w1111 = w1107 ^ w1110 ;
  assign w1112 = w1102 ^ w1105 ;
  assign w1113 = w1111 ^ w1112 ;
  assign w1114 = w1075 ^ w1113 ;
  assign w1115 = w1096 ^ w1114 ;
  assign w1116 = ( w1063 & w1064 ) | ( w1063 & w1065 ) | ( w1064 & w1065 ) ;
  assign w1117 = ( w975 & w997 ) | ( w975 & w1033 ) | ( w997 & w1033 ) ;
  assign w1118 = ( w958 & w984 ) | ( w958 & w990 ) | ( w984 & w990 ) ;
  assign w1119 = ( \pi01 & ~\pi16 ) | ( \pi01 & \pi30 ) | ( ~\pi16 & \pi30 ) ;
  assign w1120 = \pi16 & w1119 ;
  assign w1121 = ~\pi01 & \pi14 ;
  assign w1122 = ( ~\pi14 & \pi29 ) | ( ~\pi14 & w1121 ) | ( \pi29 & w1121 ) ;
  assign w1123 = ( \pi16 & ~\pi29 ) | ( \pi16 & w1122 ) | ( ~\pi29 & w1122 ) ;
  assign w1124 = w1053 ^ w1123 ;
  assign w1125 = \pi01 & \pi30 ;
  assign w1126 = w1124 ^ w1125 ;
  assign w1127 = w1117 ^ w1118 ;
  assign w1128 = w1126 ^ w1127 ;
  assign w1129 = w1031 ^ w1047 ;
  assign w1130 = w1059 ^ w1129 ;
  assign w1131 = ( w1049 & w1055 ) | ( w1049 & w1061 ) | ( w1055 & w1061 ) ;
  assign w1132 = ( w1022 & w1023 ) | ( w1022 & w1024 ) | ( w1023 & w1024 ) ;
  assign w1133 = w1130 ^ w1132 ;
  assign w1134 = w1131 ^ w1133 ;
  assign w1135 = w1116 ^ w1134 ;
  assign w1136 = w1128 ^ w1135 ;
  assign w1137 = w1074 ^ w1136 ;
  assign w1138 = w1115 ^ w1137 ;
  assign w1139 = ( w1013 & w1069 ) | ( w1013 & w1070 ) | ( w1069 & w1070 ) ;
  assign w1140 = w1138 ^ w1139 ;
  assign w1141 = w1073 ^ w1140 ;
  assign w1142 = ( w1073 & w1138 ) | ( w1073 & w1139 ) | ( w1138 & w1139 ) ;
  assign w1143 = ( w1074 & w1115 ) | ( w1074 & w1136 ) | ( w1115 & w1136 ) ;
  assign w1144 = ( w1116 & w1128 ) | ( w1116 & w1134 ) | ( w1128 & w1134 ) ;
  assign w1145 = ( w1130 & w1131 ) | ( w1130 & w1132 ) | ( w1131 & w1132 ) ;
  assign w1146 = \pi09 & \pi23 ;
  assign w1147 = \pi05 & \pi27 ;
  assign w1148 = \pi04 & \pi28 ;
  assign w1149 = ( w1146 & w1147 ) | ( w1146 & w1148 ) | ( w1147 & w1148 ) ;
  assign w1150 = w1146 ^ w1148 ;
  assign w1151 = w1147 ^ w1150 ;
  assign w1152 = \pi08 & \pi24 ;
  assign w1153 = \pi07 & \pi25 ;
  assign w1154 = \pi06 & \pi26 ;
  assign w1155 = ( w1152 & w1153 ) | ( w1152 & w1154 ) | ( w1153 & w1154 ) ;
  assign w1156 = w1152 ^ w1154 ;
  assign w1157 = w1153 ^ w1156 ;
  assign w1158 = \pi14 & \pi29 ;
  assign w1159 = ( ~\pi30 & w1053 ) | ( ~\pi30 & w1158 ) | ( w1053 & w1158 ) ;
  assign w1160 = \pi16 & w1159 ;
  assign w1161 = ( \pi01 & \pi16 ) | ( \pi01 & ~\pi30 ) | ( \pi16 & ~\pi30 ) ;
  assign w1162 = ( \pi01 & \pi16 ) | ( \pi01 & w1053 ) | ( \pi16 & w1053 ) ;
  assign w1163 = ( w1160 & ~w1161 ) | ( w1160 & w1162 ) | ( ~w1161 & w1162 ) ;
  assign w1164 = w1151 ^ w1163 ;
  assign w1165 = w1157 ^ w1164 ;
  assign w1166 = \pi30 & \pi32 ;
  assign w1167 = \pi02 & \pi30 ;
  assign w1168 = \pi00 & \pi32 ;
  assign w1169 = ( w1120 & w1167 ) | ( w1120 & w1168 ) | ( w1167 & w1168 ) ;
  assign w1170 = w1120 ^ w1168 ;
  assign w1171 = w1167 ^ w1170 ;
  assign w1172 = \pi13 & \pi19 ;
  assign w1173 = \pi12 & \pi20 ;
  assign w1174 = \pi11 & \pi21 ;
  assign w1175 = ( w1172 & w1173 ) | ( w1172 & w1174 ) | ( w1173 & w1174 ) ;
  assign w1176 = w1172 ^ w1174 ;
  assign w1177 = w1173 ^ w1176 ;
  assign w1178 = \pi14 & \pi18 ;
  assign w1179 = \pi10 & \pi22 ;
  assign w1180 = \pi03 & \pi29 ;
  assign w1181 = ( w1178 & w1179 ) | ( w1178 & w1180 ) | ( w1179 & w1180 ) ;
  assign w1182 = w1178 ^ w1180 ;
  assign w1183 = w1179 ^ w1182 ;
  assign w1184 = w1171 ^ w1177 ;
  assign w1185 = w1183 ^ w1184 ;
  assign w1186 = w1145 ^ w1165 ;
  assign w1187 = w1185 ^ w1186 ;
  assign w1188 = ( w1117 & w1118 ) | ( w1117 & w1126 ) | ( w1118 & w1126 ) ;
  assign w1189 = w1092 ^ w1100 ;
  assign w1190 = w1109 ^ w1189 ;
  assign w1191 = ( ~\pi01 & \pi31 ) | ( ~\pi01 & w460 ) | ( \pi31 & w460 ) ;
  assign w1192 = \pi01 & w1191 ;
  assign w1193 = \pi01 & \pi31 ;
  assign w1194 = w1079 ^ w1085 ;
  assign w1195 = w460 ^ w1194 ;
  assign w1196 = w1193 ^ w1195 ;
  assign w1197 = w1188 ^ w1190 ;
  assign w1198 = w1196 ^ w1197 ;
  assign w1199 = ( w1102 & w1105 ) | ( w1102 & w1111 ) | ( w1105 & w1111 ) ;
  assign w1200 = ( w1031 & w1047 ) | ( w1031 & w1059 ) | ( w1047 & w1059 ) ;
  assign w1201 = ( w1081 & w1087 ) | ( w1081 & w1094 ) | ( w1087 & w1094 ) ;
  assign w1202 = w1199 ^ w1200 ;
  assign w1203 = w1201 ^ w1202 ;
  assign w1204 = ( w1075 & w1096 ) | ( w1075 & w1113 ) | ( w1096 & w1113 ) ;
  assign w1205 = w1198 ^ w1204 ;
  assign w1206 = w1203 ^ w1205 ;
  assign w1207 = w1144 ^ w1187 ;
  assign w1208 = w1206 ^ w1207 ;
  assign w1209 = w1142 ^ w1143 ;
  assign w1210 = w1208 ^ w1209 ;
  assign w1211 = w1169 ^ w1175 ;
  assign w1212 = w1181 ^ w1211 ;
  assign w1213 = \pi11 & \pi22 ;
  assign w1214 = \pi02 & \pi31 ;
  assign w1215 = \pi00 & \pi33 ;
  assign w1216 = ( w1213 & w1214 ) | ( w1213 & w1215 ) | ( w1214 & w1215 ) ;
  assign w1217 = w1213 ^ w1215 ;
  assign w1218 = w1214 ^ w1217 ;
  assign w1219 = w1149 ^ w1155 ;
  assign w1220 = w1218 ^ w1219 ;
  assign w1221 = \pi29 & \pi30 ;
  assign w1222 = \pi09 & \pi24 ;
  assign w1223 = \pi04 & \pi29 ;
  assign w1224 = \pi03 & \pi30 ;
  assign w1225 = ( w1222 & w1223 ) | ( w1222 & w1224 ) | ( w1223 & w1224 ) ;
  assign w1226 = w1222 ^ w1224 ;
  assign w1227 = w1223 ^ w1226 ;
  assign w1228 = \pi25 & \pi27 ;
  assign w1229 = \pi08 & \pi25 ;
  assign w1230 = \pi06 & \pi27 ;
  assign w1231 = \pi05 & \pi28 ;
  assign w1232 = ( w1229 & w1230 ) | ( w1229 & w1231 ) | ( w1230 & w1231 ) ;
  assign w1233 = w1229 ^ w1231 ;
  assign w1234 = w1230 ^ w1233 ;
  assign w1235 = \pi16 & \pi17 ;
  assign w1236 = \pi15 & \pi18 ;
  assign w1237 = \pi07 & \pi26 ;
  assign w1238 = ( w1235 & w1236 ) | ( w1235 & w1237 ) | ( w1236 & w1237 ) ;
  assign w1239 = w1235 ^ w1237 ;
  assign w1240 = w1236 ^ w1239 ;
  assign w1241 = w1227 ^ w1234 ;
  assign w1242 = w1240 ^ w1241 ;
  assign w1243 = w1212 ^ w1220 ;
  assign w1244 = w1242 ^ w1243 ;
  assign w1245 = ( w1092 & w1100 ) | ( w1092 & w1109 ) | ( w1100 & w1109 ) ;
  assign w1246 = ( w1171 & w1177 ) | ( w1171 & w1183 ) | ( w1177 & w1183 ) ;
  assign w1247 = ( w1151 & w1157 ) | ( w1151 & w1163 ) | ( w1157 & w1163 ) ;
  assign w1248 = w1246 ^ w1247 ;
  assign w1249 = w1245 ^ w1248 ;
  assign w1250 = ( w1145 & w1165 ) | ( w1145 & w1185 ) | ( w1165 & w1185 ) ;
  assign w1251 = w1244 ^ w1250 ;
  assign w1252 = w1249 ^ w1251 ;
  assign w1253 = \pi01 & \pi32 ;
  assign w1254 = \pi17 ^ w1253 ;
  assign w1255 = \pi10 & \pi23 ;
  assign w1256 = ( w1192 & w1254 ) | ( w1192 & w1255 ) | ( w1254 & w1255 ) ;
  assign w1257 = w1192 ^ w1255 ;
  assign w1258 = \pi17 ^ w1257 ;
  assign w1259 = w1253 ^ w1258 ;
  assign w1260 = \pi14 & \pi19 ;
  assign w1261 = \pi13 & \pi20 ;
  assign w1262 = \pi12 & \pi21 ;
  assign w1263 = ( w1260 & w1261 ) | ( w1260 & w1262 ) | ( w1261 & w1262 ) ;
  assign w1264 = w1260 ^ w1262 ;
  assign w1265 = w1261 ^ w1264 ;
  assign w1266 = w460 ^ w1193 ;
  assign w1267 = ( w1079 & w1085 ) | ( w1079 & w1266 ) | ( w1085 & w1266 ) ;
  assign w1268 = w1259 ^ w1267 ;
  assign w1269 = w1265 ^ w1268 ;
  assign w1270 = ( w1199 & w1200 ) | ( w1199 & w1201 ) | ( w1200 & w1201 ) ;
  assign w1271 = ( w1188 & w1190 ) | ( w1188 & w1196 ) | ( w1190 & w1196 ) ;
  assign w1272 = w1269 ^ w1271 ;
  assign w1273 = w1270 ^ w1272 ;
  assign w1274 = ( w1198 & w1203 ) | ( w1198 & w1204 ) | ( w1203 & w1204 ) ;
  assign w1275 = w1252 ^ w1273 ;
  assign w1276 = w1274 ^ w1275 ;
  assign w1277 = ( w1144 & w1187 ) | ( w1144 & w1206 ) | ( w1187 & w1206 ) ;
  assign w1278 = ( w1142 & w1143 ) | ( w1142 & w1208 ) | ( w1143 & w1208 ) ;
  assign w1279 = w1276 ^ w1278 ;
  assign w1280 = w1277 ^ w1279 ;
  assign w1281 = ( w1276 & w1277 ) | ( w1276 & w1278 ) | ( w1277 & w1278 ) ;
  assign w1282 = ( w1252 & w1273 ) | ( w1252 & w1274 ) | ( w1273 & w1274 ) ;
  assign w1283 = \pi12 & \pi22 ;
  assign w1284 = \pi11 & \pi23 ;
  assign w1285 = \pi02 & \pi32 ;
  assign w1286 = ( w1283 & w1284 ) | ( w1283 & w1285 ) | ( w1284 & w1285 ) ;
  assign w1287 = w1283 ^ w1285 ;
  assign w1288 = w1284 ^ w1287 ;
  assign w1289 = w1256 ^ w1263 ;
  assign w1290 = w1288 ^ w1289 ;
  assign w1291 = ( w1259 & w1265 ) | ( w1259 & w1267 ) | ( w1265 & w1267 ) ;
  assign w1292 = w1290 ^ w1291 ;
  assign w1293 = \pi10 & \pi24 ;
  assign w1294 = \pi09 & \pi25 ;
  assign w1295 = \pi05 & \pi29 ;
  assign w1296 = ( w1293 & w1294 ) | ( w1293 & w1295 ) | ( w1294 & w1295 ) ;
  assign w1297 = w1293 ^ w1295 ;
  assign w1298 = w1294 ^ w1297 ;
  assign w1299 = \pi15 & \pi19 ;
  assign w1300 = \pi14 & \pi20 ;
  assign w1301 = \pi13 & \pi21 ;
  assign w1302 = ( w1299 & w1300 ) | ( w1299 & w1301 ) | ( w1300 & w1301 ) ;
  assign w1303 = w1299 ^ w1301 ;
  assign w1304 = w1300 ^ w1303 ;
  assign w1305 = \pi26 & \pi28 ;
  assign w1306 = \pi08 & \pi26 ;
  assign w1307 = \pi07 & \pi27 ;
  assign w1308 = \pi06 & \pi28 ;
  assign w1309 = ( w1306 & w1307 ) | ( w1306 & w1308 ) | ( w1307 & w1308 ) ;
  assign w1310 = w1306 ^ w1308 ;
  assign w1311 = w1307 ^ w1310 ;
  assign w1312 = w1298 ^ w1304 ;
  assign w1313 = w1311 ^ w1312 ;
  assign w1314 = w1216 ^ w1225 ;
  assign w1315 = w1232 ^ w1314 ;
  assign w1316 = ( w1227 & w1234 ) | ( w1227 & w1240 ) | ( w1234 & w1240 ) ;
  assign w1317 = ( ~\pi01 & \pi33 ) | ( ~\pi01 & w491 ) | ( \pi33 & w491 ) ;
  assign w1318 = \pi01 & w1317 ;
  assign w1319 = ( ~\pi01 & \pi17 ) | ( ~\pi01 & \pi32 ) | ( \pi17 & \pi32 ) ;
  assign w1320 = \pi33 ^ w1319 ;
  assign w1321 = \pi01 & w1320 ;
  assign w1322 = w491 ^ w1238 ;
  assign w1323 = w1321 ^ w1322 ;
  assign w1324 = w1315 ^ w1316 ;
  assign w1325 = w1323 ^ w1324 ;
  assign w1326 = ( w1269 & w1270 ) | ( w1269 & w1271 ) | ( w1270 & w1271 ) ;
  assign w1327 = w1313 ^ w1325 ;
  assign w1328 = w1326 ^ w1327 ;
  assign w1329 = w1292 ^ w1328 ;
  assign w1330 = ( w1244 & w1249 ) | ( w1244 & w1250 ) | ( w1249 & w1250 ) ;
  assign w1331 = ( w1212 & w1220 ) | ( w1212 & w1242 ) | ( w1220 & w1242 ) ;
  assign w1332 = ( w1245 & w1246 ) | ( w1245 & w1247 ) | ( w1246 & w1247 ) ;
  assign w1333 = ( w1149 & w1155 ) | ( w1149 & w1218 ) | ( w1155 & w1218 ) ;
  assign w1334 = ( w1169 & w1175 ) | ( w1169 & w1181 ) | ( w1175 & w1181 ) ;
  assign w1335 = \pi30 & \pi31 ;
  assign w1336 = \pi00 & \pi34 ;
  assign w1337 = \pi04 & \pi30 ;
  assign w1338 = w1336 ^ w1337 ;
  assign w1339 = \pi03 & \pi31 ;
  assign w1340 = w1338 ^ w1339 ;
  assign w1341 = w1333 ^ w1334 ;
  assign w1342 = w1340 ^ w1341 ;
  assign w1343 = w1331 ^ w1332 ;
  assign w1344 = w1342 ^ w1343 ;
  assign w1345 = w1329 ^ w1330 ;
  assign w1346 = w1344 ^ w1345 ;
  assign w1347 = w1282 & w1346 ;
  assign w1348 = w1282 | w1346 ;
  assign w1349 = ~w1347 & w1348 ;
  assign w1350 = w1281 ^ w1349 ;
  assign w1351 = ( w1281 & w1347 ) | ( w1281 & w1348 ) | ( w1347 & w1348 ) ;
  assign w1352 = w1347 | w1351 ;
  assign w1353 = ( w1329 & w1330 ) | ( w1329 & w1344 ) | ( w1330 & w1344 ) ;
  assign w1354 = w1292 ^ w1313 ;
  assign w1355 = ( w1325 & w1326 ) | ( w1325 & w1354 ) | ( w1326 & w1354 ) ;
  assign w1356 = ( w1216 & w1225 ) | ( w1216 & w1232 ) | ( w1225 & w1232 ) ;
  assign w1357 = \pi32 & w421 ;
  assign w1358 = \pi01 & \pi33 ;
  assign w1359 = w491 ^ w1358 ;
  assign w1360 = ( w1238 & w1357 ) | ( w1238 & w1359 ) | ( w1357 & w1359 ) ;
  assign w1361 = ( w1256 & w1263 ) | ( w1256 & w1288 ) | ( w1263 & w1288 ) ;
  assign w1362 = w1356 ^ w1361 ;
  assign w1363 = w1360 ^ w1362 ;
  assign w1364 = ( w1315 & w1316 ) | ( w1315 & w1323 ) | ( w1316 & w1323 ) ;
  assign w1365 = ( w1290 & w1291 ) | ( w1290 & w1313 ) | ( w1291 & w1313 ) ;
  assign w1366 = w1363 ^ w1365 ;
  assign w1367 = w1364 ^ w1366 ;
  assign w1368 = \pi08 & \pi27 ;
  assign w1369 = \pi06 & \pi29 ;
  assign w1370 = \pi05 & \pi30 ;
  assign w1371 = ( w1368 & w1369 ) | ( w1368 & w1370 ) | ( w1369 & w1370 ) ;
  assign w1372 = w1368 ^ w1370 ;
  assign w1373 = w1369 ^ w1372 ;
  assign w1374 = \pi16 & \pi19 ;
  assign w1375 = \pi07 & \pi28 ;
  assign w1376 = ( w492 & w1374 ) | ( w492 & w1375 ) | ( w1374 & w1375 ) ;
  assign w1377 = w492 ^ w1375 ;
  assign w1378 = w1374 ^ w1377 ;
  assign w1379 = \pi10 & \pi25 ;
  assign w1380 = \pi09 & \pi26 ;
  assign w1381 = \pi04 & \pi31 ;
  assign w1382 = ( w1379 & w1380 ) | ( w1379 & w1381 ) | ( w1380 & w1381 ) ;
  assign w1383 = w1379 ^ w1381 ;
  assign w1384 = w1380 ^ w1383 ;
  assign w1385 = w1373 ^ w1378 ;
  assign w1386 = w1384 ^ w1385 ;
  assign w1387 = ( w1333 & w1334 ) | ( w1333 & w1340 ) | ( w1334 & w1340 ) ;
  assign w1388 = w1386 ^ w1387 ;
  assign w1389 = \pi33 & \pi35 ;
  assign w1390 = \pi02 & \pi33 ;
  assign w1391 = \pi00 & \pi35 ;
  assign w1392 = ( w1318 & w1390 ) | ( w1318 & w1391 ) | ( w1390 & w1391 ) ;
  assign w1393 = w1318 ^ w1391 ;
  assign w1394 = w1390 ^ w1393 ;
  assign w1395 = \pi12 & \pi23 ;
  assign w1396 = \pi11 & \pi24 ;
  assign w1397 = \pi03 & \pi32 ;
  assign w1398 = ( w1395 & w1396 ) | ( w1395 & w1397 ) | ( w1396 & w1397 ) ;
  assign w1399 = w1395 ^ w1397 ;
  assign w1400 = w1396 ^ w1399 ;
  assign w1401 = \pi15 & \pi20 ;
  assign w1402 = \pi14 & \pi21 ;
  assign w1403 = \pi13 & \pi22 ;
  assign w1404 = ( w1401 & w1402 ) | ( w1401 & w1403 ) | ( w1402 & w1403 ) ;
  assign w1405 = w1401 ^ w1403 ;
  assign w1406 = w1402 ^ w1405 ;
  assign w1407 = w1394 ^ w1400 ;
  assign w1408 = w1406 ^ w1407 ;
  assign w1409 = ( w1331 & w1332 ) | ( w1331 & w1342 ) | ( w1332 & w1342 ) ;
  assign w1410 = ( w1336 & w1337 ) | ( w1336 & w1339 ) | ( w1337 & w1339 ) ;
  assign w1411 = w1286 ^ w1302 ;
  assign w1412 = w1410 ^ w1411 ;
  assign w1413 = ( w1298 & w1304 ) | ( w1298 & w1311 ) | ( w1304 & w1311 ) ;
  assign w1414 = ( \pi01 & ~\pi18 ) | ( \pi01 & \pi34 ) | ( ~\pi18 & \pi34 ) ;
  assign w1415 = \pi18 & w1414 ;
  assign w1416 = \pi01 & \pi34 ;
  assign w1417 = \pi18 ^ w1309 ;
  assign w1418 = w1296 ^ w1417 ;
  assign w1419 = w1416 ^ w1418 ;
  assign w1420 = w1412 ^ w1413 ;
  assign w1421 = w1419 ^ w1420 ;
  assign w1422 = w1408 ^ w1421 ;
  assign w1423 = w1388 ^ w1422 ;
  assign w1424 = w1409 ^ w1423 ;
  assign w1425 = w1355 ^ w1367 ;
  assign w1426 = w1424 ^ w1425 ;
  assign w1427 = w1352 ^ w1353 ;
  assign w1428 = w1426 ^ w1427 ;
  assign w1429 = ( w1355 & w1367 ) | ( w1355 & w1424 ) | ( w1367 & w1424 ) ;
  assign w1430 = w1388 ^ w1408 ;
  assign w1431 = ( w1409 & w1421 ) | ( w1409 & w1430 ) | ( w1421 & w1430 ) ;
  assign w1432 = ( w1286 & w1302 ) | ( w1286 & w1410 ) | ( w1302 & w1410 ) ;
  assign w1433 = \pi18 ^ w1416 ;
  assign w1434 = ( w1296 & w1309 ) | ( w1296 & w1433 ) | ( w1309 & w1433 ) ;
  assign w1435 = ( w1394 & w1400 ) | ( w1394 & w1406 ) | ( w1400 & w1406 ) ;
  assign w1436 = w1432 ^ w1435 ;
  assign w1437 = w1434 ^ w1436 ;
  assign w1438 = ( w1412 & w1413 ) | ( w1412 & w1419 ) | ( w1413 & w1419 ) ;
  assign w1439 = ( w1386 & w1387 ) | ( w1386 & w1408 ) | ( w1387 & w1408 ) ;
  assign w1440 = w1437 ^ w1439 ;
  assign w1441 = w1438 ^ w1440 ;
  assign w1442 = \pi13 & \pi23 ;
  assign w1443 = \pi12 & \pi24 ;
  assign w1444 = \pi02 & \pi34 ;
  assign w1445 = ( w1442 & w1443 ) | ( w1442 & w1444 ) | ( w1443 & w1444 ) ;
  assign w1446 = w1442 ^ w1444 ;
  assign w1447 = w1443 ^ w1446 ;
  assign w1448 = \pi10 & \pi26 ;
  assign w1449 = \pi09 & \pi27 ;
  assign w1450 = \pi05 & \pi31 ;
  assign w1451 = ( w1448 & w1449 ) | ( w1448 & w1450 ) | ( w1449 & w1450 ) ;
  assign w1452 = w1448 ^ w1450 ;
  assign w1453 = w1449 ^ w1452 ;
  assign w1454 = \pi28 & \pi30 ;
  assign w1455 = \pi08 & \pi28 ;
  assign w1456 = \pi07 & \pi29 ;
  assign w1457 = \pi06 & \pi30 ;
  assign w1458 = ( w1455 & w1456 ) | ( w1455 & w1457 ) | ( w1456 & w1457 ) ;
  assign w1459 = w1455 ^ w1457 ;
  assign w1460 = w1456 ^ w1459 ;
  assign w1461 = w1447 ^ w1453 ;
  assign w1462 = w1460 ^ w1461 ;
  assign w1463 = ( w1356 & w1360 ) | ( w1356 & w1361 ) | ( w1360 & w1361 ) ;
  assign w1464 = \pi17 & \pi19 ;
  assign w1465 = \pi01 & \pi35 ;
  assign w1466 = w1415 ^ w1465 ;
  assign w1467 = w1464 ^ w1466 ;
  assign w1468 = \pi00 & \pi36 ;
  assign w1469 = w1467 ^ w1468 ;
  assign w1470 = \pi11 & \pi25 ;
  assign w1471 = \pi04 & \pi32 ;
  assign w1472 = \pi03 & \pi33 ;
  assign w1473 = ( w1470 & w1471 ) | ( w1470 & w1472 ) | ( w1471 & w1472 ) ;
  assign w1474 = w1470 ^ w1472 ;
  assign w1475 = w1471 ^ w1474 ;
  assign w1476 = \pi16 & \pi20 ;
  assign w1477 = \pi15 & \pi21 ;
  assign w1478 = \pi14 & \pi22 ;
  assign w1479 = ( w1476 & w1477 ) | ( w1476 & w1478 ) | ( w1477 & w1478 ) ;
  assign w1480 = w1476 ^ w1478 ;
  assign w1481 = w1477 ^ w1480 ;
  assign w1482 = w1469 ^ w1475 ;
  assign w1483 = w1481 ^ w1482 ;
  assign w1484 = w1463 ^ w1483 ;
  assign w1485 = w1462 ^ w1484 ;
  assign w1486 = ( w1363 & w1364 ) | ( w1363 & w1365 ) | ( w1364 & w1365 ) ;
  assign w1487 = w1371 ^ w1376 ;
  assign w1488 = w1382 ^ w1487 ;
  assign w1489 = w1392 ^ w1398 ;
  assign w1490 = w1404 ^ w1489 ;
  assign w1491 = ( w1373 & w1378 ) | ( w1373 & w1384 ) | ( w1378 & w1384 ) ;
  assign w1492 = w1488 ^ w1490 ;
  assign w1493 = w1491 ^ w1492 ;
  assign w1494 = w1485 ^ w1486 ;
  assign w1495 = w1493 ^ w1494 ;
  assign w1496 = w1431 ^ w1495 ;
  assign w1497 = w1441 ^ w1496 ;
  assign w1498 = ( w1352 & w1353 ) | ( w1352 & w1426 ) | ( w1353 & w1426 ) ;
  assign w1499 = w1429 ^ w1498 ;
  assign w1500 = w1497 ^ w1499 ;
  assign w1501 = ( w1431 & w1441 ) | ( w1431 & w1495 ) | ( w1441 & w1495 ) ;
  assign w1502 = ( w1437 & w1438 ) | ( w1437 & w1439 ) | ( w1438 & w1439 ) ;
  assign w1503 = w1464 ^ w1465 ;
  assign w1504 = ( w1415 & w1468 ) | ( w1415 & w1503 ) | ( w1468 & w1503 ) ;
  assign w1505 = \pi15 & \pi22 ;
  assign w1506 = \pi14 & \pi23 ;
  assign w1507 = \pi13 & \pi24 ;
  assign w1508 = ( w1505 & w1506 ) | ( w1505 & w1507 ) | ( w1506 & w1507 ) ;
  assign w1509 = w1505 ^ w1507 ;
  assign w1510 = w1506 ^ w1509 ;
  assign w1511 = w1451 ^ w1504 ;
  assign w1512 = w1510 ^ w1511 ;
  assign w1513 = w1445 ^ w1473 ;
  assign w1514 = w1479 ^ w1513 ;
  assign w1515 = ( w1469 & w1475 ) | ( w1469 & w1481 ) | ( w1475 & w1481 ) ;
  assign w1516 = w1512 ^ w1515 ;
  assign w1517 = w1514 ^ w1516 ;
  assign w1518 = \pi11 & \pi26 ;
  assign w1519 = \pi10 & \pi27 ;
  assign w1520 = \pi05 & \pi32 ;
  assign w1521 = ( w1518 & w1519 ) | ( w1518 & w1520 ) | ( w1519 & w1520 ) ;
  assign w1522 = w1518 ^ w1520 ;
  assign w1523 = w1519 ^ w1522 ;
  assign w1524 = \pi18 & \pi19 ;
  assign w1525 = \pi17 & \pi20 ;
  assign w1526 = \pi08 & \pi29 ;
  assign w1527 = ( w1524 & w1525 ) | ( w1524 & w1526 ) | ( w1525 & w1526 ) ;
  assign w1528 = w1524 ^ w1526 ;
  assign w1529 = w1525 ^ w1528 ;
  assign w1530 = ( w1392 & w1398 ) | ( w1392 & w1404 ) | ( w1398 & w1404 ) ;
  assign w1531 = w1523 ^ w1530 ;
  assign w1532 = w1529 ^ w1531 ;
  assign w1533 = ( w1432 & w1434 ) | ( w1432 & w1435 ) | ( w1434 & w1435 ) ;
  assign w1534 = \pi12 & \pi25 ;
  assign w1535 = \pi04 & \pi33 ;
  assign w1536 = \pi00 & \pi37 ;
  assign w1537 = ( w1534 & w1535 ) | ( w1534 & w1536 ) | ( w1535 & w1536 ) ;
  assign w1538 = w1534 ^ w1536 ;
  assign w1539 = w1535 ^ w1538 ;
  assign w1540 = \pi34 & \pi35 ;
  assign w1541 = \pi16 & \pi21 ;
  assign w1542 = \pi03 & \pi34 ;
  assign w1543 = \pi02 & \pi35 ;
  assign w1544 = ( w1541 & w1542 ) | ( w1541 & w1543 ) | ( w1542 & w1543 ) ;
  assign w1545 = w1541 ^ w1543 ;
  assign w1546 = w1542 ^ w1545 ;
  assign w1547 = \pi09 & \pi28 ;
  assign w1548 = \pi07 & \pi30 ;
  assign w1549 = \pi06 & \pi31 ;
  assign w1550 = ( w1547 & w1548 ) | ( w1547 & w1549 ) | ( w1548 & w1549 ) ;
  assign w1551 = w1547 ^ w1549 ;
  assign w1552 = w1548 ^ w1551 ;
  assign w1553 = w1539 ^ w1546 ;
  assign w1554 = w1552 ^ w1553 ;
  assign w1555 = w1532 ^ w1533 ;
  assign w1556 = w1554 ^ w1555 ;
  assign w1557 = w1502 ^ w1556 ;
  assign w1558 = w1517 ^ w1557 ;
  assign w1559 = ( w1485 & w1486 ) | ( w1485 & w1493 ) | ( w1486 & w1493 ) ;
  assign w1560 = ( w1462 & w1463 ) | ( w1462 & w1483 ) | ( w1463 & w1483 ) ;
  assign w1561 = ( w1488 & w1490 ) | ( w1488 & w1491 ) | ( w1490 & w1491 ) ;
  assign w1562 = ( w1447 & w1453 ) | ( w1447 & w1460 ) | ( w1453 & w1460 ) ;
  assign w1563 = ( w1371 & w1376 ) | ( w1371 & w1382 ) | ( w1376 & w1382 ) ;
  assign w1564 = ~\pi01 & \pi17 ;
  assign w1565 = ( ~\pi17 & \pi35 ) | ( ~\pi17 & w1564 ) | ( \pi35 & w1564 ) ;
  assign w1566 = ( \pi19 & ~\pi35 ) | ( \pi19 & w1565 ) | ( ~\pi35 & w1565 ) ;
  assign w1567 = w1458 ^ w1566 ;
  assign w1568 = \pi01 & \pi36 ;
  assign w1569 = w1567 ^ w1568 ;
  assign w1570 = w1562 ^ w1563 ;
  assign w1571 = w1569 ^ w1570 ;
  assign w1572 = w1560 ^ w1561 ;
  assign w1573 = w1571 ^ w1572 ;
  assign w1574 = w1558 ^ w1559 ;
  assign w1575 = w1573 ^ w1574 ;
  assign w1576 = ( w1429 & w1497 ) | ( w1429 & w1498 ) | ( w1497 & w1498 ) ;
  assign w1577 = w1501 ^ w1576 ;
  assign w1578 = w1575 ^ w1577 ;
  assign w1579 = ( w1558 & w1559 ) | ( w1558 & w1573 ) | ( w1559 & w1573 ) ;
  assign w1580 = ( w1532 & w1533 ) | ( w1532 & w1554 ) | ( w1533 & w1554 ) ;
  assign w1581 = ( w1512 & w1514 ) | ( w1512 & w1515 ) | ( w1514 & w1515 ) ;
  assign w1582 = w1508 ^ w1537 ;
  assign w1583 = w1544 ^ w1582 ;
  assign w1584 = ( w1523 & w1529 ) | ( w1523 & w1530 ) | ( w1529 & w1530 ) ;
  assign w1585 = w1583 ^ w1584 ;
  assign w1586 = \pi10 & \pi28 ;
  assign w1587 = \pi06 & \pi32 ;
  assign w1588 = \pi05 & \pi33 ;
  assign w1589 = ( w1586 & w1587 ) | ( w1586 & w1588 ) | ( w1587 & w1588 ) ;
  assign w1590 = w1586 ^ w1588 ;
  assign w1591 = w1587 ^ w1590 ;
  assign w1592 = \pi17 & \pi21 ;
  assign w1593 = \pi16 & \pi22 ;
  assign w1594 = \pi15 & \pi23 ;
  assign w1595 = ( w1592 & w1593 ) | ( w1592 & w1594 ) | ( w1593 & w1594 ) ;
  assign w1596 = w1592 ^ w1594 ;
  assign w1597 = w1593 ^ w1596 ;
  assign w1598 = \pi09 & \pi29 ;
  assign w1599 = \pi08 & \pi30 ;
  assign w1600 = \pi07 & \pi31 ;
  assign w1601 = ( w1598 & w1599 ) | ( w1598 & w1600 ) | ( w1599 & w1600 ) ;
  assign w1602 = w1598 ^ w1600 ;
  assign w1603 = w1599 ^ w1602 ;
  assign w1604 = w1591 ^ w1597 ;
  assign w1605 = w1603 ^ w1604 ;
  assign w1606 = w1581 ^ w1605 ;
  assign w1607 = w1580 ^ w1606 ;
  assign w1608 = w1585 ^ w1607 ;
  assign w1609 = ( w1502 & w1517 ) | ( w1502 & w1556 ) | ( w1517 & w1556 ) ;
  assign w1610 = ( w1560 & w1561 ) | ( w1560 & w1571 ) | ( w1561 & w1571 ) ;
  assign w1611 = ( w1451 & w1504 ) | ( w1451 & w1510 ) | ( w1504 & w1510 ) ;
  assign w1612 = ( w1539 & w1546 ) | ( w1539 & w1552 ) | ( w1546 & w1552 ) ;
  assign w1613 = \pi18 & \pi20 ;
  assign w1614 = w1527 ^ w1613 ;
  assign w1615 = w1550 ^ w1614 ;
  assign w1616 = \pi01 & \pi37 ;
  assign w1617 = w1615 ^ w1616 ;
  assign w1618 = w1611 ^ w1612 ;
  assign w1619 = w1617 ^ w1618 ;
  assign w1620 = \pi17 & \pi35 ;
  assign w1621 = ( ~\pi36 & w1458 ) | ( ~\pi36 & w1620 ) | ( w1458 & w1620 ) ;
  assign w1622 = \pi19 & w1621 ;
  assign w1623 = ( \pi01 & \pi19 ) | ( \pi01 & ~\pi36 ) | ( \pi19 & ~\pi36 ) ;
  assign w1624 = ( \pi01 & \pi19 ) | ( \pi01 & w1458 ) | ( \pi19 & w1458 ) ;
  assign w1625 = ( w1622 & ~w1623 ) | ( w1622 & w1624 ) | ( ~w1623 & w1624 ) ;
  assign w1626 = \pi12 & \pi26 ;
  assign w1627 = \pi11 & \pi27 ;
  assign w1628 = \pi04 & \pi34 ;
  assign w1629 = ( w1626 & w1627 ) | ( w1626 & w1628 ) | ( w1627 & w1628 ) ;
  assign w1630 = w1626 ^ w1628 ;
  assign w1631 = w1627 ^ w1630 ;
  assign w1632 = ( w1445 & w1473 ) | ( w1445 & w1479 ) | ( w1473 & w1479 ) ;
  assign w1633 = w1625 ^ w1632 ;
  assign w1634 = w1631 ^ w1633 ;
  assign w1635 = ( w1562 & w1563 ) | ( w1562 & w1569 ) | ( w1563 & w1569 ) ;
  assign w1636 = \pi36 & \pi38 ;
  assign w1637 = ( \pi00 & ~\pi36 ) | ( \pi00 & \pi38 ) | ( ~\pi36 & \pi38 ) ;
  assign w1638 = ( \pi02 & w1623 ) | ( \pi02 & w1637 ) | ( w1623 & w1637 ) ;
  assign w1639 = \pi36 & w1638 ;
  assign w1640 = \pi00 & \pi38 ;
  assign w1641 = \pi02 ^ w1623 ;
  assign w1642 = \pi36 & w1641 ;
  assign w1643 = w1640 ^ w1642 ;
  assign w1644 = \pi14 & \pi24 ;
  assign w1645 = \pi13 & \pi25 ;
  assign w1646 = \pi03 & \pi35 ;
  assign w1647 = ( w1644 & w1645 ) | ( w1644 & w1646 ) | ( w1645 & w1646 ) ;
  assign w1648 = w1644 ^ w1646 ;
  assign w1649 = w1645 ^ w1648 ;
  assign w1650 = w1521 ^ w1643 ;
  assign w1651 = w1649 ^ w1650 ;
  assign w1652 = w1634 ^ w1635 ;
  assign w1653 = w1651 ^ w1652 ;
  assign w1654 = w1610 ^ w1653 ;
  assign w1655 = w1619 ^ w1654 ;
  assign w1656 = w1608 ^ w1655 ;
  assign w1657 = w1609 ^ w1656 ;
  assign w1658 = ( w1501 & w1575 ) | ( w1501 & w1576 ) | ( w1575 & w1576 ) ;
  assign w1659 = w1657 ^ w1658 ;
  assign w1660 = w1579 ^ w1659 ;
  assign w1661 = ( w1608 & w1609 ) | ( w1608 & w1655 ) | ( w1609 & w1655 ) ;
  assign w1662 = ( w1610 & w1619 ) | ( w1610 & w1653 ) | ( w1619 & w1653 ) ;
  assign w1663 = ( w1634 & w1635 ) | ( w1634 & w1651 ) | ( w1635 & w1651 ) ;
  assign w1664 = \pi00 & \pi39 ;
  assign w1665 = ( \pi01 & \pi18 ) | ( \pi01 & ~\pi20 ) | ( \pi18 & ~\pi20 ) ;
  assign w1666 = ( \pi20 & ~\pi37 ) | ( \pi20 & w1665 ) | ( ~\pi37 & w1665 ) ;
  assign w1667 = \pi37 & w1666 ;
  assign w1668 = w1664 ^ w1667 ;
  assign w1669 = w1613 ^ w1616 ;
  assign w1670 = ( w1527 & w1550 ) | ( w1527 & w1669 ) | ( w1550 & w1669 ) ;
  assign w1671 = ( w1508 & w1537 ) | ( w1508 & w1544 ) | ( w1537 & w1544 ) ;
  assign w1672 = w1668 ^ w1670 ;
  assign w1673 = w1671 ^ w1672 ;
  assign w1674 = \pi20 ^ w1673 ;
  assign w1675 = \pi01 & \pi38 ;
  assign w1676 = w1674 ^ w1675 ;
  assign w1677 = w1595 ^ w1639 ;
  assign w1678 = w1647 ^ w1677 ;
  assign w1679 = ( w1591 & w1597 ) | ( w1591 & w1603 ) | ( w1597 & w1603 ) ;
  assign w1680 = ( w1521 & w1643 ) | ( w1521 & w1649 ) | ( w1643 & w1649 ) ;
  assign w1681 = w1678 ^ w1679 ;
  assign w1682 = w1680 ^ w1681 ;
  assign w1683 = w1663 ^ w1682 ;
  assign w1684 = w1676 ^ w1683 ;
  assign w1685 = w1585 ^ w1605 ;
  assign w1686 = ( w1580 & w1581 ) | ( w1580 & w1685 ) | ( w1581 & w1685 ) ;
  assign w1687 = w1589 ^ w1601 ;
  assign w1688 = w1629 ^ w1687 ;
  assign w1689 = ( w1625 & w1631 ) | ( w1625 & w1632 ) | ( w1631 & w1632 ) ;
  assign w1690 = w1688 ^ w1689 ;
  assign w1691 = \pi17 & \pi22 ;
  assign w1692 = \pi12 & \pi27 ;
  assign w1693 = \pi04 & \pi35 ;
  assign w1694 = ( w1691 & w1692 ) | ( w1691 & w1693 ) | ( w1692 & w1693 ) ;
  assign w1695 = w1691 ^ w1693 ;
  assign w1696 = w1692 ^ w1695 ;
  assign w1697 = \pi19 & \pi20 ;
  assign w1698 = \pi18 & \pi21 ;
  assign w1699 = \pi08 & \pi31 ;
  assign w1700 = ( w1697 & w1698 ) | ( w1697 & w1699 ) | ( w1698 & w1699 ) ;
  assign w1701 = w1697 ^ w1699 ;
  assign w1702 = w1698 ^ w1701 ;
  assign w1703 = \pi11 & \pi28 ;
  assign w1704 = \pi10 & \pi29 ;
  assign w1705 = \pi05 & \pi34 ;
  assign w1706 = ( w1703 & w1704 ) | ( w1703 & w1705 ) | ( w1704 & w1705 ) ;
  assign w1707 = w1703 ^ w1705 ;
  assign w1708 = w1704 ^ w1707 ;
  assign w1709 = w1696 ^ w1702 ;
  assign w1710 = w1708 ^ w1709 ;
  assign w1711 = \pi13 & \pi26 ;
  assign w1712 = \pi03 & \pi36 ;
  assign w1713 = \pi02 & \pi37 ;
  assign w1714 = ( w1711 & w1712 ) | ( w1711 & w1713 ) | ( w1712 & w1713 ) ;
  assign w1715 = w1711 ^ w1713 ;
  assign w1716 = w1712 ^ w1715 ;
  assign w1717 = \pi16 & \pi23 ;
  assign w1718 = \pi15 & \pi24 ;
  assign w1719 = \pi14 & \pi25 ;
  assign w1720 = ( w1717 & w1718 ) | ( w1717 & w1719 ) | ( w1718 & w1719 ) ;
  assign w1721 = w1717 ^ w1719 ;
  assign w1722 = w1718 ^ w1721 ;
  assign w1723 = \pi09 & \pi30 ;
  assign w1724 = \pi07 & \pi32 ;
  assign w1725 = \pi06 & \pi33 ;
  assign w1726 = ( w1723 & w1724 ) | ( w1723 & w1725 ) | ( w1724 & w1725 ) ;
  assign w1727 = w1723 ^ w1725 ;
  assign w1728 = w1724 ^ w1727 ;
  assign w1729 = w1716 ^ w1722 ;
  assign w1730 = w1728 ^ w1729 ;
  assign w1731 = ( w1611 & w1612 ) | ( w1611 & w1617 ) | ( w1612 & w1617 ) ;
  assign w1732 = ( w1583 & w1584 ) | ( w1583 & w1605 ) | ( w1584 & w1605 ) ;
  assign w1733 = w1731 ^ w1732 ;
  assign w1734 = w1730 ^ w1733 ;
  assign w1735 = w1690 ^ w1710 ;
  assign w1736 = w1686 ^ w1735 ;
  assign w1737 = w1734 ^ w1736 ;
  assign w1738 = w1662 ^ w1737 ;
  assign w1739 = w1684 ^ w1738 ;
  assign w1740 = ( w1579 & w1657 ) | ( w1579 & w1658 ) | ( w1657 & w1658 ) ;
  assign w1741 = w1661 ^ w1740 ;
  assign w1742 = w1739 ^ w1741 ;
  assign w1743 = ( w1661 & w1739 ) | ( w1661 & w1740 ) | ( w1739 & w1740 ) ;
  assign w1744 = ( w1662 & w1684 ) | ( w1662 & w1737 ) | ( w1684 & w1737 ) ;
  assign w1745 = ( w1686 & w1734 ) | ( w1686 & w1735 ) | ( w1734 & w1735 ) ;
  assign w1746 = ( w1730 & w1731 ) | ( w1730 & w1732 ) | ( w1731 & w1732 ) ;
  assign w1747 = ( w1688 & w1689 ) | ( w1688 & w1710 ) | ( w1689 & w1710 ) ;
  assign w1748 = w1694 ^ w1706 ;
  assign w1749 = w1714 ^ w1748 ;
  assign w1750 = ( w1696 & w1702 ) | ( w1696 & w1708 ) | ( w1702 & w1708 ) ;
  assign w1751 = ( w1716 & w1722 ) | ( w1716 & w1728 ) | ( w1722 & w1728 ) ;
  assign w1752 = w1749 ^ w1750 ;
  assign w1753 = w1751 ^ w1752 ;
  assign w1754 = w1746 ^ w1747 ;
  assign w1755 = w1753 ^ w1754 ;
  assign w1756 = \pi18 & \pi37 ;
  assign w1757 = ( ~\pi38 & w1664 ) | ( ~\pi38 & w1756 ) | ( w1664 & w1756 ) ;
  assign w1758 = \pi20 & w1757 ;
  assign w1759 = ( \pi01 & \pi20 ) | ( \pi01 & ~\pi38 ) | ( \pi20 & ~\pi38 ) ;
  assign w1760 = ( \pi01 & \pi20 ) | ( \pi01 & w1664 ) | ( \pi20 & w1664 ) ;
  assign w1761 = ( w1758 & ~w1759 ) | ( w1758 & w1760 ) | ( ~w1759 & w1760 ) ;
  assign w1762 = w1720 ^ w1761 ;
  assign w1763 = w1726 ^ w1762 ;
  assign w1764 = \pi20 ^ w1668 ;
  assign w1765 = w1675 ^ w1764 ;
  assign w1766 = ( w1670 & w1671 ) | ( w1670 & w1765 ) | ( w1671 & w1765 ) ;
  assign w1767 = \pi02 & \pi38 ;
  assign w1768 = \pi00 & \pi40 ;
  assign w1769 = ( w697 & w1767 ) | ( w697 & w1768 ) | ( w1767 & w1768 ) ;
  assign w1770 = w697 ^ w1768 ;
  assign w1771 = w1767 ^ w1770 ;
  assign w1772 = \pi31 & \pi32 ;
  assign w1773 = \pi09 & \pi31 ;
  assign w1774 = \pi08 & \pi32 ;
  assign w1775 = \pi07 & \pi33 ;
  assign w1776 = ( w1773 & w1774 ) | ( w1773 & w1775 ) | ( w1774 & w1775 ) ;
  assign w1777 = w1773 ^ w1775 ;
  assign w1778 = w1774 ^ w1777 ;
  assign w1779 = \pi35 & \pi36 ;
  assign w1780 = \pi12 & \pi28 ;
  assign w1781 = \pi05 & \pi35 ;
  assign w1782 = \pi04 & \pi36 ;
  assign w1783 = ( w1780 & w1781 ) | ( w1780 & w1782 ) | ( w1781 & w1782 ) ;
  assign w1784 = w1780 ^ w1782 ;
  assign w1785 = w1781 ^ w1784 ;
  assign w1786 = w1771 ^ w1778 ;
  assign w1787 = w1785 ^ w1786 ;
  assign w1788 = w1763 ^ w1766 ;
  assign w1789 = w1787 ^ w1788 ;
  assign w1790 = ( w1663 & w1676 ) | ( w1663 & w1682 ) | ( w1676 & w1682 ) ;
  assign w1791 = \pi14 & \pi26 ;
  assign w1792 = \pi13 & \pi27 ;
  assign w1793 = \pi03 & \pi37 ;
  assign w1794 = ( w1791 & w1792 ) | ( w1791 & w1793 ) | ( w1792 & w1793 ) ;
  assign w1795 = w1791 ^ w1793 ;
  assign w1796 = w1792 ^ w1795 ;
  assign w1797 = \pi17 & \pi23 ;
  assign w1798 = \pi16 & \pi24 ;
  assign w1799 = \pi15 & \pi25 ;
  assign w1800 = ( w1797 & w1798 ) | ( w1797 & w1799 ) | ( w1798 & w1799 ) ;
  assign w1801 = w1797 ^ w1799 ;
  assign w1802 = w1798 ^ w1801 ;
  assign w1803 = \pi11 & \pi29 ;
  assign w1804 = \pi10 & \pi30 ;
  assign w1805 = \pi06 & \pi34 ;
  assign w1806 = ( w1803 & w1804 ) | ( w1803 & w1805 ) | ( w1804 & w1805 ) ;
  assign w1807 = w1803 ^ w1805 ;
  assign w1808 = w1804 ^ w1807 ;
  assign w1809 = w1796 ^ w1802 ;
  assign w1810 = w1808 ^ w1809 ;
  assign w1811 = ( w1678 & w1679 ) | ( w1678 & w1680 ) | ( w1679 & w1680 ) ;
  assign w1812 = ( w1589 & w1601 ) | ( w1589 & w1629 ) | ( w1601 & w1629 ) ;
  assign w1813 = ( w1595 & w1639 ) | ( w1595 & w1647 ) | ( w1639 & w1647 ) ;
  assign w1814 = ( ~\pi01 & \pi20 ) | ( ~\pi01 & \pi38 ) | ( \pi20 & \pi38 ) ;
  assign w1815 = \pi39 ^ w1814 ;
  assign w1816 = \pi01 & w1815 ;
  assign w1817 = w709 ^ w1700 ;
  assign w1818 = w1816 ^ w1817 ;
  assign w1819 = w1812 ^ w1813 ;
  assign w1820 = w1818 ^ w1819 ;
  assign w1821 = w1811 ^ w1820 ;
  assign w1822 = w1810 ^ w1821 ;
  assign w1823 = w1790 ^ w1822 ;
  assign w1824 = w1789 ^ w1823 ;
  assign w1825 = w1745 ^ w1755 ;
  assign w1826 = w1824 ^ w1825 ;
  assign w1827 = w1744 & w1826 ;
  assign w1828 = w1744 | w1826 ;
  assign w1829 = ~w1827 & w1828 ;
  assign w1830 = w1743 ^ w1829 ;
  assign w1831 = ( w1745 & w1755 ) | ( w1745 & w1824 ) | ( w1755 & w1824 ) ;
  assign w1832 = ( w1810 & w1811 ) | ( w1810 & w1820 ) | ( w1811 & w1820 ) ;
  assign w1833 = ( w1763 & w1766 ) | ( w1763 & w1787 ) | ( w1766 & w1787 ) ;
  assign w1834 = w1769 ^ w1794 ;
  assign w1835 = w1800 ^ w1834 ;
  assign w1836 = ( w1771 & w1778 ) | ( w1771 & w1785 ) | ( w1778 & w1785 ) ;
  assign w1837 = \pi01 & \pi40 ;
  assign w1838 = \pi21 ^ w1806 ;
  assign w1839 = w1776 ^ w1838 ;
  assign w1840 = w1837 ^ w1839 ;
  assign w1841 = w1835 ^ w1836 ;
  assign w1842 = w1840 ^ w1841 ;
  assign w1843 = w1832 ^ w1833 ;
  assign w1844 = w1842 ^ w1843 ;
  assign w1845 = ( w1789 & w1790 ) | ( w1789 & w1822 ) | ( w1790 & w1822 ) ;
  assign w1846 = ( w1720 & w1726 ) | ( w1720 & w1761 ) | ( w1726 & w1761 ) ;
  assign w1847 = ( w1694 & w1706 ) | ( w1694 & w1714 ) | ( w1706 & w1714 ) ;
  assign w1848 = ( w1796 & w1802 ) | ( w1796 & w1808 ) | ( w1802 & w1808 ) ;
  assign w1849 = w1846 ^ w1847 ;
  assign w1850 = w1848 ^ w1849 ;
  assign w1851 = \pi39 & \pi41 ;
  assign w1852 = \pi00 & \pi41 ;
  assign w1853 = ( \pi01 & ~\pi39 ) | ( \pi01 & w709 ) | ( ~\pi39 & w709 ) ;
  assign w1854 = \pi02 ^ w1853 ;
  assign w1855 = \pi39 & w1854 ;
  assign w1856 = w1852 ^ w1855 ;
  assign w1857 = \pi15 & \pi26 ;
  assign w1858 = \pi13 & \pi28 ;
  assign w1859 = \pi03 & \pi38 ;
  assign w1860 = ( w1857 & w1858 ) | ( w1857 & w1859 ) | ( w1858 & w1859 ) ;
  assign w1861 = w1857 ^ w1859 ;
  assign w1862 = w1858 ^ w1861 ;
  assign w1863 = w1783 ^ w1856 ;
  assign w1864 = w1862 ^ w1863 ;
  assign w1865 = ( w1749 & w1750 ) | ( w1749 & w1751 ) | ( w1750 & w1751 ) ;
  assign w1866 = w1850 ^ w1864 ;
  assign w1867 = w1865 ^ w1866 ;
  assign w1868 = ( w1746 & w1747 ) | ( w1746 & w1753 ) | ( w1747 & w1753 ) ;
  assign w1869 = \pi11 & \pi30 ;
  assign w1870 = \pi06 & \pi35 ;
  assign w1871 = \pi05 & \pi36 ;
  assign w1872 = ( w1869 & w1870 ) | ( w1869 & w1871 ) | ( w1870 & w1871 ) ;
  assign w1873 = w1869 ^ w1871 ;
  assign w1874 = w1870 ^ w1873 ;
  assign w1875 = \pi19 & \pi22 ;
  assign w1876 = \pi38 & w568 ;
  assign w1877 = \pi01 & \pi39 ;
  assign w1878 = w709 ^ w1877 ;
  assign w1879 = ( w1700 & w1876 ) | ( w1700 & w1878 ) | ( w1876 & w1878 ) ;
  assign w1880 = w710 ^ w1879 ;
  assign w1881 = w1874 ^ w1880 ;
  assign w1882 = w1875 ^ w1881 ;
  assign w1883 = \pi08 & \pi33 ;
  assign w1884 = w1882 ^ w1883 ;
  assign w1885 = ( w1812 & w1813 ) | ( w1812 & w1818 ) | ( w1813 & w1818 ) ;
  assign w1886 = \pi14 & \pi27 ;
  assign w1887 = \pi12 & \pi29 ;
  assign w1888 = \pi04 & \pi37 ;
  assign w1889 = ( w1886 & w1887 ) | ( w1886 & w1888 ) | ( w1887 & w1888 ) ;
  assign w1890 = w1886 ^ w1888 ;
  assign w1891 = w1887 ^ w1890 ;
  assign w1892 = \pi18 & \pi23 ;
  assign w1893 = \pi17 & \pi24 ;
  assign w1894 = \pi16 & \pi25 ;
  assign w1895 = ( w1892 & w1893 ) | ( w1892 & w1894 ) | ( w1893 & w1894 ) ;
  assign w1896 = w1892 ^ w1894 ;
  assign w1897 = w1893 ^ w1896 ;
  assign w1898 = \pi32 & \pi34 ;
  assign w1899 = \pi10 & \pi31 ;
  assign w1900 = \pi09 & \pi32 ;
  assign w1901 = \pi07 & \pi34 ;
  assign w1902 = ( w1899 & w1900 ) | ( w1899 & w1901 ) | ( w1900 & w1901 ) ;
  assign w1903 = w1899 ^ w1901 ;
  assign w1904 = w1900 ^ w1903 ;
  assign w1905 = w1891 ^ w1897 ;
  assign w1906 = w1904 ^ w1905 ;
  assign w1907 = w1884 ^ w1885 ;
  assign w1908 = w1906 ^ w1907 ;
  assign w1909 = w1867 ^ w1868 ;
  assign w1910 = w1908 ^ w1909 ;
  assign w1911 = w1845 ^ w1910 ;
  assign w1912 = w1844 ^ w1911 ;
  assign w1913 = ( w1743 & w1827 ) | ( w1743 & w1828 ) | ( w1827 & w1828 ) ;
  assign w1914 = w1827 | w1913 ;
  assign w1915 = w1912 ^ w1914 ;
  assign w1916 = w1831 ^ w1915 ;
  assign w1917 = ( w1831 & w1912 ) | ( w1831 & w1914 ) | ( w1912 & w1914 ) ;
  assign w1918 = ( w1844 & w1845 ) | ( w1844 & w1910 ) | ( w1845 & w1910 ) ;
  assign w1919 = ( w1832 & w1833 ) | ( w1832 & w1842 ) | ( w1833 & w1842 ) ;
  assign w1920 = ( w1846 & w1847 ) | ( w1846 & w1848 ) | ( w1847 & w1848 ) ;
  assign w1921 = \pi07 & \pi35 ;
  assign w1922 = \pi11 & \pi31 ;
  assign w1923 = \pi06 & \pi36 ;
  assign w1924 = ( w1921 & w1922 ) | ( w1921 & w1923 ) | ( w1922 & w1923 ) ;
  assign w1925 = w1922 ^ w1923 ;
  assign w1926 = w1921 ^ w1925 ;
  assign w1927 = \pi10 & \pi32 ;
  assign w1928 = \pi09 & \pi33 ;
  assign w1929 = \pi08 & \pi34 ;
  assign w1930 = ( w1927 & w1928 ) | ( w1927 & w1929 ) | ( w1928 & w1929 ) ;
  assign w1931 = w1927 ^ w1929 ;
  assign w1932 = w1928 ^ w1931 ;
  assign w1933 = w1902 ^ w1926 ;
  assign w1934 = w1932 ^ w1933 ;
  assign w1935 = w1920 ^ w1934 ;
  assign w1936 = \pi16 & \pi26 ;
  assign w1937 = \pi03 & \pi39 ;
  assign w1938 = \pi02 & \pi40 ;
  assign w1939 = ( w1936 & w1937 ) | ( w1936 & w1938 ) | ( w1937 & w1938 ) ;
  assign w1940 = w1936 ^ w1938 ;
  assign w1941 = w1937 ^ w1940 ;
  assign w1942 = \pi19 & \pi23 ;
  assign w1943 = \pi18 & \pi24 ;
  assign w1944 = \pi17 & \pi25 ;
  assign w1945 = ( w1942 & w1943 ) | ( w1942 & w1944 ) | ( w1943 & w1944 ) ;
  assign w1946 = w1942 ^ w1944 ;
  assign w1947 = w1943 ^ w1946 ;
  assign w1948 = \pi15 & \pi38 ;
  assign w1949 = \pi15 & \pi27 ;
  assign w1950 = \pi14 & \pi28 ;
  assign w1951 = \pi04 & \pi38 ;
  assign w1952 = ( w1949 & w1950 ) | ( w1949 & w1951 ) | ( w1950 & w1951 ) ;
  assign w1953 = w1949 ^ w1951 ;
  assign w1954 = w1950 ^ w1953 ;
  assign w1955 = w1941 ^ w1947 ;
  assign w1956 = w1954 ^ w1955 ;
  assign w1957 = \pi00 & \pi42 ;
  assign w1958 = ( \pi01 & \pi21 ) | ( \pi01 & ~\pi40 ) | ( \pi21 & ~\pi40 ) ;
  assign w1959 = \pi40 & w1958 ;
  assign w1960 = w1957 ^ w1959 ;
  assign w1961 = \pi01 & \pi41 ;
  assign w1962 = \pi20 & \pi22 ;
  assign w1963 = w1961 ^ w1962 ;
  assign w1964 = \pi13 & \pi29 ;
  assign w1965 = \pi12 & \pi30 ;
  assign w1966 = \pi05 & \pi37 ;
  assign w1967 = ( w1964 & w1965 ) | ( w1964 & w1966 ) | ( w1965 & w1966 ) ;
  assign w1968 = w1964 ^ w1966 ;
  assign w1969 = w1965 ^ w1968 ;
  assign w1970 = \pi21 ^ w1837 ;
  assign w1971 = ( w1776 & w1806 ) | ( w1776 & w1970 ) | ( w1806 & w1970 ) ;
  assign w1972 = w1963 ^ w1969 ;
  assign w1973 = w1971 ^ w1972 ;
  assign w1974 = w1960 ^ w1973 ;
  assign w1975 = ( w1835 & w1836 ) | ( w1835 & w1840 ) | ( w1836 & w1840 ) ;
  assign w1976 = ( w710 & w1875 ) | ( w710 & w1883 ) | ( w1875 & w1883 ) ;
  assign w1977 = w1872 ^ w1976 ;
  assign w1978 = w1889 ^ w1977 ;
  assign w1979 = w710 ^ w1875 ;
  assign w1980 = w1883 ^ w1979 ;
  assign w1981 = ( w1874 & w1879 ) | ( w1874 & w1980 ) | ( w1879 & w1980 ) ;
  assign w1982 = ( \pi00 & ~\pi39 ) | ( \pi00 & \pi41 ) | ( ~\pi39 & \pi41 ) ;
  assign w1983 = ( \pi02 & w1853 ) | ( \pi02 & w1982 ) | ( w1853 & w1982 ) ;
  assign w1984 = \pi39 & w1983 ;
  assign w1985 = w1860 ^ w1984 ;
  assign w1986 = w1895 ^ w1985 ;
  assign w1987 = w1981 ^ w1986 ;
  assign w1988 = w1978 ^ w1987 ;
  assign w1989 = w1975 ^ w1988 ;
  assign w1990 = w1974 ^ w1989 ;
  assign w1991 = w1956 ^ w1990 ;
  assign w1992 = w1919 ^ w1991 ;
  assign w1993 = w1935 ^ w1992 ;
  assign w1994 = ( w1867 & w1868 ) | ( w1867 & w1908 ) | ( w1868 & w1908 ) ;
  assign w1995 = ( w1850 & w1864 ) | ( w1850 & w1865 ) | ( w1864 & w1865 ) ;
  assign w1996 = ( w1769 & w1794 ) | ( w1769 & w1800 ) | ( w1794 & w1800 ) ;
  assign w1997 = ( w1783 & w1856 ) | ( w1783 & w1862 ) | ( w1856 & w1862 ) ;
  assign w1998 = ( w1891 & w1897 ) | ( w1891 & w1904 ) | ( w1897 & w1904 ) ;
  assign w1999 = w1996 ^ w1997 ;
  assign w2000 = w1998 ^ w1999 ;
  assign w2001 = ( w1884 & w1885 ) | ( w1884 & w1906 ) | ( w1885 & w1906 ) ;
  assign w2002 = w1995 ^ w2001 ;
  assign w2003 = w2000 ^ w2002 ;
  assign w2004 = w1993 ^ w1994 ;
  assign w2005 = w2003 ^ w2004 ;
  assign w2006 = w1917 ^ w1918 ;
  assign w2007 = w2005 ^ w2006 ;
  assign w2008 = ( w1993 & w1994 ) | ( w1993 & w2003 ) | ( w1994 & w2003 ) ;
  assign w2009 = w1935 ^ w1956 ;
  assign w2010 = ( w1919 & w1990 ) | ( w1919 & w2009 ) | ( w1990 & w2009 ) ;
  assign w2011 = ( w1974 & w1975 ) | ( w1974 & w1988 ) | ( w1975 & w1988 ) ;
  assign w2012 = ( w1920 & w1934 ) | ( w1920 & w1956 ) | ( w1934 & w1956 ) ;
  assign w2013 = ( w1941 & w1947 ) | ( w1941 & w1954 ) | ( w1947 & w1954 ) ;
  assign w2014 = ( w1902 & w1926 ) | ( w1902 & w1932 ) | ( w1926 & w1932 ) ;
  assign w2015 = ~\pi01 & \pi20 ;
  assign w2016 = ( ~\pi20 & \pi41 ) | ( ~\pi20 & w2015 ) | ( \pi41 & w2015 ) ;
  assign w2017 = ( \pi22 & ~\pi41 ) | ( \pi22 & w2016 ) | ( ~\pi41 & w2016 ) ;
  assign w2018 = w1930 ^ w2017 ;
  assign w2019 = \pi01 & \pi42 ;
  assign w2020 = w2018 ^ w2019 ;
  assign w2021 = w2013 ^ w2014 ;
  assign w2022 = w2020 ^ w2021 ;
  assign w2023 = w2011 ^ w2012 ;
  assign w2024 = w2022 ^ w2023 ;
  assign w2025 = ( w1995 & w2000 ) | ( w1995 & w2001 ) | ( w2000 & w2001 ) ;
  assign w2026 = ( w1996 & w1997 ) | ( w1996 & w1998 ) | ( w1997 & w1998 ) ;
  assign w2027 = \pi04 & \pi39 ;
  assign w2028 = \pi03 & \pi40 ;
  assign w2029 = \pi00 & \pi43 ;
  assign w2030 = ( w2027 & w2028 ) | ( w2027 & w2029 ) | ( w2028 & w2029 ) ;
  assign w2031 = w2027 ^ w2029 ;
  assign w2032 = w2028 ^ w2031 ;
  assign w2033 = \pi16 & \pi27 ;
  assign w2034 = \pi15 & \pi28 ;
  assign w2035 = ( w1158 & w2033 ) | ( w1158 & w2034 ) | ( w2033 & w2034 ) ;
  assign w2036 = w1158 ^ w2033 ;
  assign w2037 = w2034 ^ w2036 ;
  assign w2038 = \pi19 & \pi24 ;
  assign w2039 = \pi18 & \pi25 ;
  assign w2040 = \pi17 & \pi26 ;
  assign w2041 = ( w2038 & w2039 ) | ( w2038 & w2040 ) | ( w2039 & w2040 ) ;
  assign w2042 = w2038 ^ w2040 ;
  assign w2043 = w2039 ^ w2042 ;
  assign w2044 = w2032 ^ w2037 ;
  assign w2045 = w2043 ^ w2044 ;
  assign w2046 = \pi10 & \pi33 ;
  assign w2047 = \pi08 & \pi35 ;
  assign w2048 = \pi07 & \pi36 ;
  assign w2049 = ( w2046 & w2047 ) | ( w2046 & w2048 ) | ( w2047 & w2048 ) ;
  assign w2050 = w2046 ^ w2048 ;
  assign w2051 = w2047 ^ w2050 ;
  assign w2052 = \pi21 & \pi22 ;
  assign w2053 = \pi20 & \pi23 ;
  assign w2054 = \pi09 & \pi34 ;
  assign w2055 = ( w2052 & w2053 ) | ( w2052 & w2054 ) | ( w2053 & w2054 ) ;
  assign w2056 = w2052 ^ w2054 ;
  assign w2057 = w2053 ^ w2056 ;
  assign w2058 = \pi13 & \pi30 ;
  assign w2059 = \pi05 & \pi38 ;
  assign w2060 = \pi02 & \pi41 ;
  assign w2061 = ( w2058 & w2059 ) | ( w2058 & w2060 ) | ( w2059 & w2060 ) ;
  assign w2062 = w2058 ^ w2060 ;
  assign w2063 = w2059 ^ w2062 ;
  assign w2064 = w2051 ^ w2057 ;
  assign w2065 = w2063 ^ w2064 ;
  assign w2066 = w2026 ^ w2045 ;
  assign w2067 = w2065 ^ w2066 ;
  assign w2068 = w1960 ^ w1963 ;
  assign w2069 = ( w1969 & w1971 ) | ( w1969 & w2068 ) | ( w1971 & w2068 ) ;
  assign w2070 = w1924 ^ w1945 ;
  assign w2071 = w1952 ^ w2070 ;
  assign w2072 = ( \pi01 & ~\pi21 ) | ( \pi01 & \pi40 ) | ( ~\pi21 & \pi40 ) ;
  assign w2073 = \pi21 & w2072 ;
  assign w2074 = ( w1957 & w1963 ) | ( w1957 & w2073 ) | ( w1963 & w2073 ) ;
  assign w2075 = w1939 ^ w2074 ;
  assign w2076 = w1967 ^ w2075 ;
  assign w2077 = w2069 ^ w2076 ;
  assign w2078 = w2071 ^ w2077 ;
  assign w2079 = ( w1872 & w1889 ) | ( w1872 & w1976 ) | ( w1889 & w1976 ) ;
  assign w2080 = \pi12 & \pi31 ;
  assign w2081 = \pi11 & \pi32 ;
  assign w2082 = \pi06 & \pi37 ;
  assign w2083 = ( w2080 & w2081 ) | ( w2080 & w2082 ) | ( w2081 & w2082 ) ;
  assign w2084 = w2080 ^ w2082 ;
  assign w2085 = w2081 ^ w2084 ;
  assign w2086 = ( w1860 & w1895 ) | ( w1860 & w1984 ) | ( w1895 & w1984 ) ;
  assign w2087 = w2079 ^ w2086 ;
  assign w2088 = w2085 ^ w2087 ;
  assign w2089 = ( w1978 & w1981 ) | ( w1978 & w1986 ) | ( w1981 & w1986 ) ;
  assign w2090 = w2078 ^ w2088 ;
  assign w2091 = w2089 ^ w2090 ;
  assign w2092 = w2025 ^ w2067 ;
  assign w2093 = w2091 ^ w2092 ;
  assign w2094 = w2010 ^ w2093 ;
  assign w2095 = w2024 ^ w2094 ;
  assign w2096 = ( w1917 & w1918 ) | ( w1917 & w2005 ) | ( w1918 & w2005 ) ;
  assign w2097 = w2008 ^ w2096 ;
  assign w2098 = w2095 ^ w2097 ;
  assign w2099 = ( w2010 & w2024 ) | ( w2010 & w2093 ) | ( w2024 & w2093 ) ;
  assign w2100 = ( w2011 & w2012 ) | ( w2011 & w2022 ) | ( w2012 & w2022 ) ;
  assign w2101 = ( w2013 & w2014 ) | ( w2013 & w2020 ) | ( w2014 & w2020 ) ;
  assign w2102 = \pi17 & \pi27 ;
  assign w2103 = \pi15 & \pi29 ;
  assign w2104 = \pi03 & \pi41 ;
  assign w2105 = ( w2102 & w2103 ) | ( w2102 & w2104 ) | ( w2103 & w2104 ) ;
  assign w2106 = w2102 ^ w2104 ;
  assign w2107 = w2103 ^ w2106 ;
  assign w2108 = \pi20 & \pi24 ;
  assign w2109 = \pi19 & \pi25 ;
  assign w2110 = \pi18 & \pi26 ;
  assign w2111 = ( w2108 & w2109 ) | ( w2108 & w2110 ) | ( w2109 & w2110 ) ;
  assign w2112 = w2108 ^ w2110 ;
  assign w2113 = w2109 ^ w2112 ;
  assign w2114 = \pi11 & \pi33 ;
  assign w2115 = \pi07 & \pi37 ;
  assign w2116 = \pi06 & \pi38 ;
  assign w2117 = ( w2114 & w2115 ) | ( w2114 & w2116 ) | ( w2115 & w2116 ) ;
  assign w2118 = w2114 ^ w2116 ;
  assign w2119 = w2115 ^ w2118 ;
  assign w2120 = w2107 ^ w2113 ;
  assign w2121 = w2119 ^ w2120 ;
  assign w2122 = \pi16 & \pi28 ;
  assign w2123 = \pi14 & \pi30 ;
  assign w2124 = \pi04 & \pi40 ;
  assign w2125 = ( w2122 & w2123 ) | ( w2122 & w2124 ) | ( w2123 & w2124 ) ;
  assign w2126 = w2122 ^ w2124 ;
  assign w2127 = w2123 ^ w2126 ;
  assign w2128 = \pi10 & \pi34 ;
  assign w2129 = \pi09 & \pi35 ;
  assign w2130 = \pi08 & \pi36 ;
  assign w2131 = ( w2128 & w2129 ) | ( w2128 & w2130 ) | ( w2129 & w2130 ) ;
  assign w2132 = w2128 ^ w2130 ;
  assign w2133 = w2129 ^ w2132 ;
  assign w2134 = \pi13 & \pi31 ;
  assign w2135 = \pi12 & \pi32 ;
  assign w2136 = \pi05 & \pi39 ;
  assign w2137 = ( w2134 & w2135 ) | ( w2134 & w2136 ) | ( w2135 & w2136 ) ;
  assign w2138 = w2134 ^ w2136 ;
  assign w2139 = w2135 ^ w2138 ;
  assign w2140 = w2127 ^ w2133 ;
  assign w2141 = w2139 ^ w2140 ;
  assign w2142 = w2101 ^ w2121 ;
  assign w2143 = w2141 ^ w2142 ;
  assign w2144 = ( \pi00 & ~\pi42 ) | ( \pi00 & \pi44 ) | ( ~\pi42 & \pi44 ) ;
  assign w2145 = ( \pi01 & \pi22 ) | ( \pi01 & ~\pi42 ) | ( \pi22 & ~\pi42 ) ;
  assign w2146 = ( \pi02 & w2144 ) | ( \pi02 & w2145 ) | ( w2144 & w2145 ) ;
  assign w2147 = \pi42 & w2146 ;
  assign w2148 = \pi00 & \pi44 ;
  assign w2149 = \pi02 ^ w2145 ;
  assign w2150 = \pi42 & w2149 ;
  assign w2151 = w2148 ^ w2150 ;
  assign w2152 = w2035 ^ w2083 ;
  assign w2153 = w2151 ^ w2152 ;
  assign w2154 = ( ~\pi01 & \pi43 ) | ( ~\pi01 & w646 ) | ( \pi43 & w646 ) ;
  assign w2155 = \pi01 & w2154 ;
  assign w2156 = \pi01 & \pi43 ;
  assign w2157 = w2049 ^ w2055 ;
  assign w2158 = w646 ^ w2157 ;
  assign w2159 = w2156 ^ w2158 ;
  assign w2160 = ( w2079 & w2085 ) | ( w2079 & w2086 ) | ( w2085 & w2086 ) ;
  assign w2161 = w2153 ^ w2160 ;
  assign w2162 = w2159 ^ w2161 ;
  assign w2163 = ( w2069 & w2071 ) | ( w2069 & w2076 ) | ( w2071 & w2076 ) ;
  assign w2164 = ( w1939 & w1967 ) | ( w1939 & w2074 ) | ( w1967 & w2074 ) ;
  assign w2165 = \pi20 & \pi41 ;
  assign w2166 = ( ~\pi42 & w1930 ) | ( ~\pi42 & w2165 ) | ( w1930 & w2165 ) ;
  assign w2167 = \pi22 & w2166 ;
  assign w2168 = ( \pi01 & \pi22 ) | ( \pi01 & w1930 ) | ( \pi22 & w1930 ) ;
  assign w2169 = ( ~w2145 & w2167 ) | ( ~w2145 & w2168 ) | ( w2167 & w2168 ) ;
  assign w2170 = ( w1924 & w1945 ) | ( w1924 & w1952 ) | ( w1945 & w1952 ) ;
  assign w2171 = w2164 ^ w2169 ;
  assign w2172 = w2170 ^ w2171 ;
  assign w2173 = w2163 ^ w2172 ;
  assign w2174 = w2143 ^ w2173 ;
  assign w2175 = w2100 ^ w2174 ;
  assign w2176 = w2162 ^ w2175 ;
  assign w2177 = ( w2025 & w2067 ) | ( w2025 & w2091 ) | ( w2067 & w2091 ) ;
  assign w2178 = ( w2078 & w2088 ) | ( w2078 & w2089 ) | ( w2088 & w2089 ) ;
  assign w2179 = ( w2026 & w2045 ) | ( w2026 & w2065 ) | ( w2045 & w2065 ) ;
  assign w2180 = w2030 ^ w2041 ;
  assign w2181 = w2061 ^ w2180 ;
  assign w2182 = ( w2051 & w2057 ) | ( w2051 & w2063 ) | ( w2057 & w2063 ) ;
  assign w2183 = ( w2032 & w2037 ) | ( w2032 & w2043 ) | ( w2037 & w2043 ) ;
  assign w2184 = w2181 ^ w2182 ;
  assign w2185 = w2183 ^ w2184 ;
  assign w2186 = w2178 ^ w2179 ;
  assign w2187 = w2185 ^ w2186 ;
  assign w2188 = w2176 ^ w2177 ;
  assign w2189 = w2187 ^ w2188 ;
  assign w2190 = ( w2008 & w2095 ) | ( w2008 & w2096 ) | ( w2095 & w2096 ) ;
  assign w2191 = w2099 ^ w2190 ;
  assign w2192 = w2189 ^ w2191 ;
  assign w2193 = ( w2101 & w2121 ) | ( w2101 & w2141 ) | ( w2121 & w2141 ) ;
  assign w2194 = ( w2162 & w2163 ) | ( w2162 & w2172 ) | ( w2163 & w2172 ) ;
  assign w2195 = w2105 ^ w2111 ;
  assign w2196 = w2147 ^ w2195 ;
  assign w2197 = ( w2164 & w2169 ) | ( w2164 & w2170 ) | ( w2169 & w2170 ) ;
  assign w2198 = w2196 ^ w2197 ;
  assign w2199 = \pi12 & \pi33 ;
  assign w2200 = \pi11 & \pi34 ;
  assign w2201 = \pi06 & \pi39 ;
  assign w2202 = ( w2199 & w2200 ) | ( w2199 & w2201 ) | ( w2200 & w2201 ) ;
  assign w2203 = w2199 ^ w2201 ;
  assign w2204 = w2200 ^ w2203 ;
  assign w2205 = \pi17 & \pi28 ;
  assign w2206 = \pi16 & \pi29 ;
  assign w2207 = \pi15 & \pi30 ;
  assign w2208 = ( w2205 & w2206 ) | ( w2205 & w2207 ) | ( w2206 & w2207 ) ;
  assign w2209 = w2205 ^ w2207 ;
  assign w2210 = w2206 ^ w2209 ;
  assign w2211 = \pi01 & \pi44 ;
  assign w2212 = \pi23 ^ w2211 ;
  assign w2213 = \pi03 & \pi42 ;
  assign w2214 = ( w2155 & w2212 ) | ( w2155 & w2213 ) | ( w2212 & w2213 ) ;
  assign w2215 = w2155 ^ w2213 ;
  assign w2216 = \pi23 ^ w2215 ;
  assign w2217 = w2211 ^ w2216 ;
  assign w2218 = w2204 ^ w2217 ;
  assign w2219 = w2210 ^ w2218 ;
  assign w2220 = w2193 ^ w2219 ;
  assign w2221 = w2194 ^ w2220 ;
  assign w2222 = w2198 ^ w2221 ;
  assign w2223 = w2162 ^ w2173 ;
  assign w2224 = ( w2100 & w2143 ) | ( w2100 & w2223 ) | ( w2143 & w2223 ) ;
  assign w2225 = \pi04 & \pi41 ;
  assign w2226 = \pi02 & \pi43 ;
  assign w2227 = \pi00 & \pi45 ;
  assign w2228 = ( w2225 & w2226 ) | ( w2225 & w2227 ) | ( w2226 & w2227 ) ;
  assign w2229 = w2225 ^ w2227 ;
  assign w2230 = w2226 ^ w2229 ;
  assign w2231 = \pi09 & \pi36 ;
  assign w2232 = \pi08 & \pi37 ;
  assign w2233 = \pi07 & \pi38 ;
  assign w2234 = ( w2231 & w2232 ) | ( w2231 & w2233 ) | ( w2232 & w2233 ) ;
  assign w2235 = w2231 ^ w2233 ;
  assign w2236 = w2232 ^ w2235 ;
  assign w2237 = \pi22 & \pi23 ;
  assign w2238 = \pi21 & \pi24 ;
  assign w2239 = \pi10 & \pi35 ;
  assign w2240 = ( w2237 & w2238 ) | ( w2237 & w2239 ) | ( w2238 & w2239 ) ;
  assign w2241 = w2237 ^ w2239 ;
  assign w2242 = w2238 ^ w2241 ;
  assign w2243 = w2230 ^ w2236 ;
  assign w2244 = w2242 ^ w2243 ;
  assign w2245 = \pi14 & \pi31 ;
  assign w2246 = \pi13 & \pi32 ;
  assign w2247 = \pi05 & \pi40 ;
  assign w2248 = ( w2245 & w2246 ) | ( w2245 & w2247 ) | ( w2246 & w2247 ) ;
  assign w2249 = w2245 ^ w2247 ;
  assign w2250 = w2246 ^ w2249 ;
  assign w2251 = \pi20 & \pi25 ;
  assign w2252 = \pi19 & \pi26 ;
  assign w2253 = \pi18 & \pi27 ;
  assign w2254 = ( w2251 & w2252 ) | ( w2251 & w2253 ) | ( w2252 & w2253 ) ;
  assign w2255 = w2251 ^ w2253 ;
  assign w2256 = w2252 ^ w2255 ;
  assign w2257 = w2131 ^ w2250 ;
  assign w2258 = w2256 ^ w2257 ;
  assign w2259 = ( w2181 & w2182 ) | ( w2181 & w2183 ) | ( w2182 & w2183 ) ;
  assign w2260 = w2244 ^ w2259 ;
  assign w2261 = w2258 ^ w2260 ;
  assign w2262 = ( w2178 & w2179 ) | ( w2178 & w2185 ) | ( w2179 & w2185 ) ;
  assign w2263 = w2261 ^ w2262 ;
  assign w2264 = ( w2035 & w2083 ) | ( w2035 & w2151 ) | ( w2083 & w2151 ) ;
  assign w2265 = ( w2030 & w2041 ) | ( w2030 & w2061 ) | ( w2041 & w2061 ) ;
  assign w2266 = w646 ^ w2156 ;
  assign w2267 = ( w2049 & w2055 ) | ( w2049 & w2266 ) | ( w2055 & w2266 ) ;
  assign w2268 = w2264 ^ w2265 ;
  assign w2269 = w2267 ^ w2268 ;
  assign w2270 = ( w2153 & w2159 ) | ( w2153 & w2160 ) | ( w2159 & w2160 ) ;
  assign w2271 = w2117 ^ w2125 ;
  assign w2272 = w2137 ^ w2271 ;
  assign w2273 = ( w2127 & w2133 ) | ( w2127 & w2139 ) | ( w2133 & w2139 ) ;
  assign w2274 = ( w2107 & w2113 ) | ( w2107 & w2119 ) | ( w2113 & w2119 ) ;
  assign w2275 = w2272 ^ w2273 ;
  assign w2276 = w2274 ^ w2275 ;
  assign w2277 = w2269 ^ w2270 ;
  assign w2278 = w2276 ^ w2277 ;
  assign w2279 = w2263 ^ w2278 ;
  assign w2280 = w2222 ^ w2279 ;
  assign w2281 = w2224 ^ w2280 ;
  assign w2282 = ( w2176 & w2177 ) | ( w2176 & w2187 ) | ( w2177 & w2187 ) ;
  assign w2283 = ( w2099 & w2189 ) | ( w2099 & w2190 ) | ( w2189 & w2190 ) ;
  assign w2284 = w2281 ^ w2283 ;
  assign w2285 = w2282 ^ w2284 ;
  assign w2286 = ( w2222 & w2224 ) | ( w2222 & w2279 ) | ( w2224 & w2279 ) ;
  assign w2287 = ( w2261 & w2262 ) | ( w2261 & w2278 ) | ( w2262 & w2278 ) ;
  assign w2288 = ( w2269 & w2270 ) | ( w2269 & w2276 ) | ( w2270 & w2276 ) ;
  assign w2289 = ( w2244 & w2258 ) | ( w2244 & w2259 ) | ( w2258 & w2259 ) ;
  assign w2290 = \pi15 & \pi31 ;
  assign w2291 = \pi05 & \pi41 ;
  assign w2292 = \pi02 & \pi44 ;
  assign w2293 = ( w2290 & w2291 ) | ( w2290 & w2292 ) | ( w2291 & w2292 ) ;
  assign w2294 = w2290 ^ w2292 ;
  assign w2295 = w2291 ^ w2294 ;
  assign w2296 = \pi14 & \pi32 ;
  assign w2297 = \pi13 & \pi33 ;
  assign w2298 = \pi06 & \pi40 ;
  assign w2299 = ( w2296 & w2297 ) | ( w2296 & w2298 ) | ( w2297 & w2298 ) ;
  assign w2300 = w2296 ^ w2298 ;
  assign w2301 = w2297 ^ w2300 ;
  assign w2302 = ( w2117 & w2125 ) | ( w2117 & w2137 ) | ( w2125 & w2137 ) ;
  assign w2303 = w2295 ^ w2302 ;
  assign w2304 = w2301 ^ w2303 ;
  assign w2305 = w2202 ^ w2208 ;
  assign w2306 = w2254 ^ w2305 ;
  assign w2307 = ( w2264 & w2265 ) | ( w2264 & w2267 ) | ( w2265 & w2267 ) ;
  assign w2308 = w2304 ^ w2307 ;
  assign w2309 = w2306 ^ w2308 ;
  assign w2310 = w2288 ^ w2289 ;
  assign w2311 = w2309 ^ w2310 ;
  assign w2312 = w2286 ^ w2287 ;
  assign w2313 = w2311 ^ w2312 ;
  assign w2314 = w2198 ^ w2219 ;
  assign w2315 = ( w2193 & w2194 ) | ( w2193 & w2314 ) | ( w2194 & w2314 ) ;
  assign w2316 = ( w2272 & w2273 ) | ( w2272 & w2274 ) | ( w2273 & w2274 ) ;
  assign w2317 = \pi04 & \pi42 ;
  assign w2318 = \pi03 & \pi43 ;
  assign w2319 = \pi00 & \pi46 ;
  assign w2320 = ( w2317 & w2318 ) | ( w2317 & w2319 ) | ( w2318 & w2319 ) ;
  assign w2321 = w2317 ^ w2319 ;
  assign w2322 = w2318 ^ w2321 ;
  assign w2323 = \pi35 & \pi37 ;
  assign w2324 = \pi11 & \pi35 ;
  assign w2325 = \pi10 & \pi36 ;
  assign w2326 = \pi09 & \pi37 ;
  assign w2327 = ( w2324 & w2325 ) | ( w2324 & w2326 ) | ( w2325 & w2326 ) ;
  assign w2328 = w2324 ^ w2326 ;
  assign w2329 = w2325 ^ w2328 ;
  assign w2330 = \pi21 & \pi25 ;
  assign w2331 = \pi20 & \pi26 ;
  assign w2332 = \pi19 & \pi27 ;
  assign w2333 = ( w2330 & w2331 ) | ( w2330 & w2332 ) | ( w2331 & w2332 ) ;
  assign w2334 = w2330 ^ w2332 ;
  assign w2335 = w2331 ^ w2334 ;
  assign w2336 = w2322 ^ w2329 ;
  assign w2337 = w2335 ^ w2336 ;
  assign w2338 = \pi18 & \pi28 ;
  assign w2339 = \pi17 & \pi29 ;
  assign w2340 = \pi16 & \pi30 ;
  assign w2341 = ( w2338 & w2339 ) | ( w2338 & w2340 ) | ( w2339 & w2340 ) ;
  assign w2342 = w2338 ^ w2340 ;
  assign w2343 = w2339 ^ w2342 ;
  assign w2344 = \pi12 & \pi34 ;
  assign w2345 = \pi08 & \pi38 ;
  assign w2346 = \pi07 & \pi39 ;
  assign w2347 = ( w2344 & w2345 ) | ( w2344 & w2346 ) | ( w2345 & w2346 ) ;
  assign w2348 = w2344 ^ w2346 ;
  assign w2349 = w2345 ^ w2348 ;
  assign w2350 = w2214 ^ w2343 ;
  assign w2351 = w2349 ^ w2350 ;
  assign w2352 = w2316 ^ w2351 ;
  assign w2353 = w2337 ^ w2352 ;
  assign w2354 = ( w2131 & w2250 ) | ( w2131 & w2256 ) | ( w2250 & w2256 ) ;
  assign w2355 = ( w2230 & w2236 ) | ( w2230 & w2242 ) | ( w2236 & w2242 ) ;
  assign w2356 = ( w2204 & w2210 ) | ( w2204 & w2217 ) | ( w2210 & w2217 ) ;
  assign w2357 = w2354 ^ w2356 ;
  assign w2358 = w2355 ^ w2357 ;
  assign w2359 = ( w2196 & w2197 ) | ( w2196 & w2219 ) | ( w2197 & w2219 ) ;
  assign w2360 = w2228 ^ w2234 ;
  assign w2361 = w2248 ^ w2360 ;
  assign w2362 = ( w2105 & w2111 ) | ( w2105 & w2147 ) | ( w2111 & w2147 ) ;
  assign w2363 = ( ~\pi01 & \pi45 ) | ( ~\pi01 & w993 ) | ( \pi45 & w993 ) ;
  assign w2364 = \pi01 & w2363 ;
  assign w2365 = ( ~\pi01 & \pi23 ) | ( ~\pi01 & \pi44 ) | ( \pi23 & \pi44 ) ;
  assign w2366 = \pi45 ^ w2365 ;
  assign w2367 = \pi01 & w2366 ;
  assign w2368 = w993 ^ w2240 ;
  assign w2369 = w2367 ^ w2368 ;
  assign w2370 = w2361 ^ w2362 ;
  assign w2371 = w2369 ^ w2370 ;
  assign w2372 = w2358 ^ w2359 ;
  assign w2373 = w2371 ^ w2372 ;
  assign w2374 = w2315 ^ w2373 ;
  assign w2375 = w2353 ^ w2374 ;
  assign w2376 = ( w2281 & w2282 ) | ( w2281 & w2283 ) | ( w2282 & w2283 ) ;
  assign w2377 = w2313 ^ w2376 ;
  assign w2378 = w2375 ^ w2377 ;
  assign w2379 = ( w2286 & w2287 ) | ( w2286 & w2311 ) | ( w2287 & w2311 ) ;
  assign w2380 = ( w2288 & w2289 ) | ( w2288 & w2309 ) | ( w2289 & w2309 ) ;
  assign w2381 = ( w2358 & w2359 ) | ( w2358 & w2371 ) | ( w2359 & w2371 ) ;
  assign w2382 = w2293 ^ w2320 ;
  assign w2383 = w2333 ^ w2382 ;
  assign w2384 = ( w2322 & w2329 ) | ( w2322 & w2335 ) | ( w2329 & w2335 ) ;
  assign w2385 = ( w2295 & w2301 ) | ( w2295 & w2302 ) | ( w2301 & w2302 ) ;
  assign w2386 = w2383 ^ w2385 ;
  assign w2387 = w2384 ^ w2386 ;
  assign w2388 = ( w2316 & w2337 ) | ( w2316 & w2351 ) | ( w2337 & w2351 ) ;
  assign w2389 = ( w2304 & w2306 ) | ( w2304 & w2307 ) | ( w2306 & w2307 ) ;
  assign w2390 = w2388 ^ w2389 ;
  assign w2391 = w2387 ^ w2390 ;
  assign w2392 = w2380 ^ w2391 ;
  assign w2393 = w2381 ^ w2392 ;
  assign w2394 = ( w2315 & w2353 ) | ( w2315 & w2373 ) | ( w2353 & w2373 ) ;
  assign w2395 = \pi44 & w695 ;
  assign w2396 = \pi01 & \pi45 ;
  assign w2397 = w993 ^ w2396 ;
  assign w2398 = ( w2240 & w2395 ) | ( w2240 & w2397 ) | ( w2395 & w2397 ) ;
  assign w2399 = \pi13 & \pi34 ;
  assign w2400 = \pi12 & \pi35 ;
  assign w2401 = \pi07 & \pi40 ;
  assign w2402 = ( w2399 & w2400 ) | ( w2399 & w2401 ) | ( w2400 & w2401 ) ;
  assign w2403 = w2399 ^ w2401 ;
  assign w2404 = w2400 ^ w2403 ;
  assign w2405 = ( w2202 & w2208 ) | ( w2202 & w2254 ) | ( w2208 & w2254 ) ;
  assign w2406 = w2398 ^ w2405 ;
  assign w2407 = w2404 ^ w2406 ;
  assign w2408 = ( w2361 & w2362 ) | ( w2361 & w2369 ) | ( w2362 & w2369 ) ;
  assign w2409 = ( w2354 & w2355 ) | ( w2354 & w2356 ) | ( w2355 & w2356 ) ;
  assign w2410 = w2407 ^ w2409 ;
  assign w2411 = w2408 ^ w2410 ;
  assign w2412 = ( w2214 & w2343 ) | ( w2214 & w2349 ) | ( w2343 & w2349 ) ;
  assign w2413 = ( w2228 & w2234 ) | ( w2228 & w2248 ) | ( w2234 & w2248 ) ;
  assign w2414 = \pi01 & \pi46 ;
  assign w2415 = \pi24 ^ w2347 ;
  assign w2416 = w2327 ^ w2415 ;
  assign w2417 = w2414 ^ w2416 ;
  assign w2418 = w2412 ^ w2413 ;
  assign w2419 = w2417 ^ w2418 ;
  assign w2420 = \pi02 & \pi45 ;
  assign w2421 = \pi00 & \pi47 ;
  assign w2422 = ( w2364 & w2420 ) | ( w2364 & w2421 ) | ( w2420 & w2421 ) ;
  assign w2423 = w2364 ^ w2421 ;
  assign w2424 = w2420 ^ w2423 ;
  assign w2425 = \pi18 & \pi29 ;
  assign w2426 = \pi17 & \pi30 ;
  assign w2427 = \pi16 & \pi31 ;
  assign w2428 = ( w2425 & w2426 ) | ( w2425 & w2427 ) | ( w2426 & w2427 ) ;
  assign w2429 = w2425 ^ w2427 ;
  assign w2430 = w2426 ^ w2429 ;
  assign w2431 = \pi21 & \pi26 ;
  assign w2432 = \pi20 & \pi27 ;
  assign w2433 = \pi19 & \pi28 ;
  assign w2434 = ( w2431 & w2432 ) | ( w2431 & w2433 ) | ( w2432 & w2433 ) ;
  assign w2435 = w2431 ^ w2433 ;
  assign w2436 = w2432 ^ w2435 ;
  assign w2437 = w2424 ^ w2430 ;
  assign w2438 = w2436 ^ w2437 ;
  assign w2439 = \pi15 & \pi32 ;
  assign w2440 = \pi04 & \pi43 ;
  assign w2441 = \pi03 & \pi44 ;
  assign w2442 = ( w2439 & w2440 ) | ( w2439 & w2441 ) | ( w2440 & w2441 ) ;
  assign w2443 = w2439 ^ w2441 ;
  assign w2444 = w2440 ^ w2443 ;
  assign w2445 = w2299 ^ w2341 ;
  assign w2446 = w2444 ^ w2445 ;
  assign w2447 = \pi11 & \pi36 ;
  assign w2448 = \pi09 & \pi38 ;
  assign w2449 = \pi08 & \pi39 ;
  assign w2450 = ( w2447 & w2448 ) | ( w2447 & w2449 ) | ( w2448 & w2449 ) ;
  assign w2451 = w2447 ^ w2449 ;
  assign w2452 = w2448 ^ w2451 ;
  assign w2453 = \pi23 & \pi24 ;
  assign w2454 = \pi22 & \pi25 ;
  assign w2455 = \pi10 & \pi37 ;
  assign w2456 = ( w2453 & w2454 ) | ( w2453 & w2455 ) | ( w2454 & w2455 ) ;
  assign w2457 = w2453 ^ w2455 ;
  assign w2458 = w2454 ^ w2457 ;
  assign w2459 = \pi33 & \pi41 ;
  assign w2460 = \pi14 & \pi33 ;
  assign w2461 = \pi06 & \pi41 ;
  assign w2462 = \pi05 & \pi42 ;
  assign w2463 = ( w2460 & w2461 ) | ( w2460 & w2462 ) | ( w2461 & w2462 ) ;
  assign w2464 = w2460 ^ w2462 ;
  assign w2465 = w2461 ^ w2464 ;
  assign w2466 = w2452 ^ w2458 ;
  assign w2467 = w2465 ^ w2466 ;
  assign w2468 = w2438 ^ w2446 ;
  assign w2469 = w2467 ^ w2468 ;
  assign w2470 = w2411 ^ w2419 ;
  assign w2471 = w2469 ^ w2470 ;
  assign w2472 = w2393 ^ w2394 ;
  assign w2473 = w2471 ^ w2472 ;
  assign w2474 = ( w2313 & w2375 ) | ( w2313 & w2376 ) | ( w2375 & w2376 ) ;
  assign w2475 = w2379 ^ w2474 ;
  assign w2476 = w2473 ^ w2475 ;
  assign w2477 = ( w2379 & w2473 ) | ( w2379 & w2474 ) | ( w2473 & w2474 ) ;
  assign w2478 = ( w2393 & w2394 ) | ( w2393 & w2471 ) | ( w2394 & w2471 ) ;
  assign w2479 = ( w2380 & w2381 ) | ( w2380 & w2391 ) | ( w2381 & w2391 ) ;
  assign w2480 = ( w2387 & w2388 ) | ( w2387 & w2389 ) | ( w2388 & w2389 ) ;
  assign w2481 = ( w2407 & w2408 ) | ( w2407 & w2409 ) | ( w2408 & w2409 ) ;
  assign w2482 = \pi14 & \pi34 ;
  assign w2483 = \pi13 & \pi35 ;
  assign w2484 = \pi06 & \pi42 ;
  assign w2485 = ( w2482 & w2483 ) | ( w2482 & w2484 ) | ( w2483 & w2484 ) ;
  assign w2486 = w2482 ^ w2484 ;
  assign w2487 = w2483 ^ w2486 ;
  assign w2488 = \pi12 & \pi36 ;
  assign w2489 = \pi08 & \pi40 ;
  assign w2490 = \pi07 & \pi41 ;
  assign w2491 = ( w2488 & w2489 ) | ( w2488 & w2490 ) | ( w2489 & w2490 ) ;
  assign w2492 = w2488 ^ w2490 ;
  assign w2493 = w2489 ^ w2492 ;
  assign w2494 = \pi37 & \pi39 ;
  assign w2495 = \pi11 & \pi37 ;
  assign w2496 = \pi10 & \pi38 ;
  assign w2497 = \pi09 & \pi39 ;
  assign w2498 = ( w2495 & w2496 ) | ( w2495 & w2497 ) | ( w2496 & w2497 ) ;
  assign w2499 = w2495 ^ w2497 ;
  assign w2500 = w2496 ^ w2499 ;
  assign w2501 = w2487 ^ w2493 ;
  assign w2502 = w2500 ^ w2501 ;
  assign w2503 = ( w2398 & w2404 ) | ( w2398 & w2405 ) | ( w2404 & w2405 ) ;
  assign w2504 = \pi33 & \pi43 ;
  assign w2505 = \pi15 & \pi33 ;
  assign w2506 = \pi05 & \pi43 ;
  assign w2507 = \pi04 & \pi44 ;
  assign w2508 = ( w2505 & w2506 ) | ( w2505 & w2507 ) | ( w2506 & w2507 ) ;
  assign w2509 = w2505 ^ w2507 ;
  assign w2510 = w2506 ^ w2509 ;
  assign w2511 = \pi22 & \pi26 ;
  assign w2512 = \pi21 & \pi27 ;
  assign w2513 = \pi20 & \pi28 ;
  assign w2514 = ( w2511 & w2512 ) | ( w2511 & w2513 ) | ( w2512 & w2513 ) ;
  assign w2515 = w2511 ^ w2513 ;
  assign w2516 = w2512 ^ w2515 ;
  assign w2517 = \pi19 & \pi29 ;
  assign w2518 = \pi18 & \pi30 ;
  assign w2519 = \pi17 & \pi31 ;
  assign w2520 = ( w2517 & w2518 ) | ( w2517 & w2519 ) | ( w2518 & w2519 ) ;
  assign w2521 = w2517 ^ w2519 ;
  assign w2522 = w2518 ^ w2521 ;
  assign w2523 = w2510 ^ w2516 ;
  assign w2524 = w2522 ^ w2523 ;
  assign w2525 = w2502 ^ w2503 ;
  assign w2526 = w2524 ^ w2525 ;
  assign w2527 = w2480 ^ w2481 ;
  assign w2528 = w2526 ^ w2527 ;
  assign w2529 = ( w2411 & w2419 ) | ( w2411 & w2469 ) | ( w2419 & w2469 ) ;
  assign w2530 = ( w2383 & w2384 ) | ( w2383 & w2385 ) | ( w2384 & w2385 ) ;
  assign w2531 = ( w2412 & w2413 ) | ( w2412 & w2417 ) | ( w2413 & w2417 ) ;
  assign w2532 = \pi00 & \pi48 ;
  assign w2533 = ( \pi01 & \pi24 ) | ( \pi01 & ~\pi46 ) | ( \pi24 & ~\pi46 ) ;
  assign w2534 = \pi46 & w2533 ;
  assign w2535 = w2532 ^ w2534 ;
  assign w2536 = \pi01 & \pi47 ;
  assign w2537 = \pi23 & \pi25 ;
  assign w2538 = w2536 ^ w2537 ;
  assign w2539 = ( w2293 & w2320 ) | ( w2293 & w2333 ) | ( w2320 & w2333 ) ;
  assign w2540 = ( w2299 & w2341 ) | ( w2299 & w2444 ) | ( w2341 & w2444 ) ;
  assign w2541 = w2535 ^ w2538 ;
  assign w2542 = w2539 ^ w2541 ;
  assign w2543 = w2540 ^ w2542 ;
  assign w2544 = w2530 ^ w2531 ;
  assign w2545 = w2543 ^ w2544 ;
  assign w2546 = w2434 ^ w2450 ;
  assign w2547 = w2463 ^ w2546 ;
  assign w2548 = ( w2452 & w2458 ) | ( w2452 & w2465 ) | ( w2458 & w2465 ) ;
  assign w2549 = \pi16 & \pi32 ;
  assign w2550 = \pi03 & \pi45 ;
  assign w2551 = \pi02 & \pi46 ;
  assign w2552 = ( w2549 & w2550 ) | ( w2549 & w2551 ) | ( w2550 & w2551 ) ;
  assign w2553 = w2549 ^ w2551 ;
  assign w2554 = w2550 ^ w2553 ;
  assign w2555 = w2402 ^ w2456 ;
  assign w2556 = w2554 ^ w2555 ;
  assign w2557 = w2547 ^ w2548 ;
  assign w2558 = w2556 ^ w2557 ;
  assign w2559 = ( w2438 & w2446 ) | ( w2438 & w2467 ) | ( w2446 & w2467 ) ;
  assign w2560 = w2422 ^ w2428 ;
  assign w2561 = w2442 ^ w2560 ;
  assign w2562 = \pi24 ^ w2414 ;
  assign w2563 = ( w2327 & w2347 ) | ( w2327 & w2562 ) | ( w2347 & w2562 ) ;
  assign w2564 = ( w2424 & w2430 ) | ( w2424 & w2436 ) | ( w2430 & w2436 ) ;
  assign w2565 = w2561 ^ w2564 ;
  assign w2566 = w2563 ^ w2565 ;
  assign w2567 = w2559 ^ w2566 ;
  assign w2568 = w2558 ^ w2567 ;
  assign w2569 = w2529 ^ w2545 ;
  assign w2570 = w2568 ^ w2569 ;
  assign w2571 = w2479 ^ w2570 ;
  assign w2572 = w2528 ^ w2571 ;
  assign w2573 = w2478 | w2572 ;
  assign w2574 = w2478 & w2572 ;
  assign w2575 = w2573 & ~w2574 ;
  assign w2576 = w2477 ^ w2575 ;
  assign w2577 = ( w2529 & w2545 ) | ( w2529 & w2568 ) | ( w2545 & w2568 ) ;
  assign w2578 = ( w2558 & w2559 ) | ( w2558 & w2566 ) | ( w2559 & w2566 ) ;
  assign w2579 = ( w2530 & w2531 ) | ( w2530 & w2543 ) | ( w2531 & w2543 ) ;
  assign w2580 = \pi13 & \pi36 ;
  assign w2581 = \pi08 & \pi41 ;
  assign w2582 = \pi07 & \pi42 ;
  assign w2583 = ( w2580 & w2581 ) | ( w2580 & w2582 ) | ( w2581 & w2582 ) ;
  assign w2584 = w2580 ^ w2582 ;
  assign w2585 = w2581 ^ w2584 ;
  assign w2586 = \pi23 & \pi26 ;
  assign w2587 = \pi11 & \pi38 ;
  assign w2588 = ( w894 & w2586 ) | ( w894 & w2587 ) | ( w2586 & w2587 ) ;
  assign w2589 = w894 ^ w2587 ;
  assign w2590 = w2586 ^ w2589 ;
  assign w2591 = \pi15 & \pi34 ;
  assign w2592 = \pi14 & \pi35 ;
  assign w2593 = \pi06 & \pi43 ;
  assign w2594 = ( w2591 & w2592 ) | ( w2591 & w2593 ) | ( w2592 & w2593 ) ;
  assign w2595 = w2591 ^ w2593 ;
  assign w2596 = w2592 ^ w2595 ;
  assign w2597 = w2585 ^ w2590 ;
  assign w2598 = w2596 ^ w2597 ;
  assign w2599 = \pi22 & \pi27 ;
  assign w2600 = \pi03 & \pi46 ;
  assign w2601 = \pi02 & \pi47 ;
  assign w2602 = ( w2599 & w2600 ) | ( w2599 & w2601 ) | ( w2600 & w2601 ) ;
  assign w2603 = w2599 ^ w2601 ;
  assign w2604 = w2600 ^ w2603 ;
  assign w2605 = \pi21 & \pi28 ;
  assign w2606 = \pi20 & \pi29 ;
  assign w2607 = \pi19 & \pi30 ;
  assign w2608 = ( w2605 & w2606 ) | ( w2605 & w2607 ) | ( w2606 & w2607 ) ;
  assign w2609 = w2605 ^ w2607 ;
  assign w2610 = w2606 ^ w2609 ;
  assign w2611 = \pi12 & \pi37 ;
  assign w2612 = \pi10 & \pi39 ;
  assign w2613 = \pi09 & \pi40 ;
  assign w2614 = ( w2611 & w2612 ) | ( w2611 & w2613 ) | ( w2612 & w2613 ) ;
  assign w2615 = w2611 ^ w2613 ;
  assign w2616 = w2612 ^ w2615 ;
  assign w2617 = w2604 ^ w2610 ;
  assign w2618 = w2616 ^ w2617 ;
  assign w2619 = \pi05 & \pi44 ;
  assign w2620 = \pi04 & \pi45 ;
  assign w2621 = \pi00 & \pi49 ;
  assign w2622 = ( w2619 & w2620 ) | ( w2619 & w2621 ) | ( w2620 & w2621 ) ;
  assign w2623 = w2619 ^ w2621 ;
  assign w2624 = w2620 ^ w2623 ;
  assign w2625 = ( \pi01 & ~\pi24 ) | ( \pi01 & \pi46 ) | ( ~\pi24 & \pi46 ) ;
  assign w2626 = \pi24 & w2625 ;
  assign w2627 = ( w2532 & w2538 ) | ( w2532 & w2626 ) | ( w2538 & w2626 ) ;
  assign w2628 = \pi18 & \pi31 ;
  assign w2629 = \pi17 & \pi32 ;
  assign w2630 = \pi16 & \pi33 ;
  assign w2631 = ( w2628 & w2629 ) | ( w2628 & w2630 ) | ( w2629 & w2630 ) ;
  assign w2632 = w2628 ^ w2630 ;
  assign w2633 = w2629 ^ w2632 ;
  assign w2634 = w2624 ^ w2627 ;
  assign w2635 = w2633 ^ w2634 ;
  assign w2636 = w2598 ^ w2635 ;
  assign w2637 = w2618 ^ w2636 ;
  assign w2638 = w2578 ^ w2579 ;
  assign w2639 = w2637 ^ w2638 ;
  assign w2640 = ( w2480 & w2481 ) | ( w2480 & w2526 ) | ( w2481 & w2526 ) ;
  assign w2641 = ( w2434 & w2450 ) | ( w2434 & w2463 ) | ( w2450 & w2463 ) ;
  assign w2642 = ( w2402 & w2456 ) | ( w2402 & w2554 ) | ( w2456 & w2554 ) ;
  assign w2643 = ( w2422 & w2428 ) | ( w2422 & w2442 ) | ( w2428 & w2442 ) ;
  assign w2644 = w2641 ^ w2643 ;
  assign w2645 = w2642 ^ w2644 ;
  assign w2646 = ( w2547 & w2548 ) | ( w2547 & w2556 ) | ( w2548 & w2556 ) ;
  assign w2647 = ( w2561 & w2563 ) | ( w2561 & w2564 ) | ( w2563 & w2564 ) ;
  assign w2648 = w2645 ^ w2647 ;
  assign w2649 = w2646 ^ w2648 ;
  assign w2650 = w2485 ^ w2491 ;
  assign w2651 = w2520 ^ w2650 ;
  assign w2652 = ( w2510 & w2516 ) | ( w2510 & w2522 ) | ( w2516 & w2522 ) ;
  assign w2653 = ( w2539 & w2540 ) | ( w2539 & w2541 ) | ( w2540 & w2541 ) ;
  assign w2654 = w2651 ^ w2653 ;
  assign w2655 = w2652 ^ w2654 ;
  assign w2656 = ( w2502 & w2503 ) | ( w2502 & w2524 ) | ( w2503 & w2524 ) ;
  assign w2657 = w2508 ^ w2514 ;
  assign w2658 = w2552 ^ w2657 ;
  assign w2659 = ( w2487 & w2493 ) | ( w2487 & w2500 ) | ( w2493 & w2500 ) ;
  assign w2660 = ~\pi01 & \pi23 ;
  assign w2661 = ( ~\pi23 & \pi47 ) | ( ~\pi23 & w2660 ) | ( \pi47 & w2660 ) ;
  assign w2662 = ( \pi25 & ~\pi47 ) | ( \pi25 & w2661 ) | ( ~\pi47 & w2661 ) ;
  assign w2663 = w2498 ^ w2662 ;
  assign w2664 = \pi01 & \pi48 ;
  assign w2665 = w2663 ^ w2664 ;
  assign w2666 = w2658 ^ w2659 ;
  assign w2667 = w2665 ^ w2666 ;
  assign w2668 = w2655 ^ w2656 ;
  assign w2669 = w2667 ^ w2668 ;
  assign w2670 = w2640 ^ w2649 ;
  assign w2671 = w2669 ^ w2670 ;
  assign w2672 = w2577 ^ w2671 ;
  assign w2673 = w2639 ^ w2672 ;
  assign w2674 = ( w2479 & w2528 ) | ( w2479 & w2570 ) | ( w2528 & w2570 ) ;
  assign w2675 = ( w2477 & w2573 ) | ( w2477 & w2574 ) | ( w2573 & w2574 ) ;
  assign w2676 = w2574 | w2675 ;
  assign w2677 = w2673 ^ w2676 ;
  assign w2678 = w2674 ^ w2677 ;
  assign w2679 = ( w2673 & w2674 ) | ( w2673 & w2676 ) | ( w2674 & w2676 ) ;
  assign w2680 = ( w2577 & w2639 ) | ( w2577 & w2671 ) | ( w2639 & w2671 ) ;
  assign w2681 = ( w2640 & w2649 ) | ( w2640 & w2669 ) | ( w2649 & w2669 ) ;
  assign w2682 = ( w2655 & w2656 ) | ( w2655 & w2667 ) | ( w2656 & w2667 ) ;
  assign w2683 = ( w2645 & w2646 ) | ( w2645 & w2647 ) | ( w2646 & w2647 ) ;
  assign w2684 = \pi16 & \pi34 ;
  assign w2685 = \pi15 & \pi35 ;
  assign w2686 = \pi05 & \pi45 ;
  assign w2687 = ( w2684 & w2685 ) | ( w2684 & w2686 ) | ( w2685 & w2686 ) ;
  assign w2688 = w2684 ^ w2686 ;
  assign w2689 = w2685 ^ w2688 ;
  assign w2690 = \pi23 & \pi27 ;
  assign w2691 = \pi22 & \pi28 ;
  assign w2692 = \pi18 & \pi32 ;
  assign w2693 = ( w2690 & w2691 ) | ( w2690 & w2692 ) | ( w2691 & w2692 ) ;
  assign w2694 = w2690 ^ w2692 ;
  assign w2695 = w2691 ^ w2694 ;
  assign w2696 = \pi23 & \pi47 ;
  assign w2697 = ( ~\pi48 & w2498 ) | ( ~\pi48 & w2696 ) | ( w2498 & w2696 ) ;
  assign w2698 = \pi25 & w2697 ;
  assign w2699 = ( \pi01 & \pi25 ) | ( \pi01 & ~\pi48 ) | ( \pi25 & ~\pi48 ) ;
  assign w2700 = ( \pi01 & \pi25 ) | ( \pi01 & w2498 ) | ( \pi25 & w2498 ) ;
  assign w2701 = ( w2698 & ~w2699 ) | ( w2698 & w2700 ) | ( ~w2699 & w2700 ) ;
  assign w2702 = w2689 ^ w2701 ;
  assign w2703 = w2695 ^ w2702 ;
  assign w2704 = ( \pi00 & ~\pi48 ) | ( \pi00 & \pi50 ) | ( ~\pi48 & \pi50 ) ;
  assign w2705 = ( \pi02 & w825 ) | ( \pi02 & w2704 ) | ( w825 & w2704 ) ;
  assign w2706 = \pi48 & w2705 ;
  assign w2707 = \pi00 & \pi50 ;
  assign w2708 = \pi02 ^ w825 ;
  assign w2709 = \pi48 & w2708 ;
  assign w2710 = w2707 ^ w2709 ;
  assign w2711 = \pi17 & \pi33 ;
  assign w2712 = \pi04 & \pi46 ;
  assign w2713 = \pi03 & \pi47 ;
  assign w2714 = ( w2711 & w2712 ) | ( w2711 & w2713 ) | ( w2712 & w2713 ) ;
  assign w2715 = w2711 ^ w2713 ;
  assign w2716 = w2712 ^ w2715 ;
  assign w2717 = \pi21 & \pi29 ;
  assign w2718 = \pi20 & \pi30 ;
  assign w2719 = \pi19 & \pi31 ;
  assign w2720 = ( w2717 & w2718 ) | ( w2717 & w2719 ) | ( w2718 & w2719 ) ;
  assign w2721 = w2717 ^ w2719 ;
  assign w2722 = w2718 ^ w2721 ;
  assign w2723 = w2710 ^ w2716 ;
  assign w2724 = w2722 ^ w2723 ;
  assign w2725 = \pi14 & \pi36 ;
  assign w2726 = \pi07 & \pi43 ;
  assign w2727 = \pi06 & \pi44 ;
  assign w2728 = ( w2725 & w2726 ) | ( w2725 & w2727 ) | ( w2726 & w2727 ) ;
  assign w2729 = w2725 ^ w2727 ;
  assign w2730 = w2726 ^ w2729 ;
  assign w2731 = \pi13 & \pi37 ;
  assign w2732 = \pi09 & \pi41 ;
  assign w2733 = \pi08 & \pi42 ;
  assign w2734 = ( w2731 & w2732 ) | ( w2731 & w2733 ) | ( w2732 & w2733 ) ;
  assign w2735 = w2731 ^ w2733 ;
  assign w2736 = w2732 ^ w2735 ;
  assign w2737 = \pi12 & \pi38 ;
  assign w2738 = \pi11 & \pi39 ;
  assign w2739 = \pi10 & \pi40 ;
  assign w2740 = ( w2737 & w2738 ) | ( w2737 & w2739 ) | ( w2738 & w2739 ) ;
  assign w2741 = w2737 ^ w2739 ;
  assign w2742 = w2738 ^ w2741 ;
  assign w2743 = w2730 ^ w2736 ;
  assign w2744 = w2742 ^ w2743 ;
  assign w2745 = w2703 ^ w2724 ;
  assign w2746 = w2744 ^ w2745 ;
  assign w2747 = w2682 ^ w2683 ;
  assign w2748 = w2746 ^ w2747 ;
  assign w2749 = ( w2578 & w2579 ) | ( w2578 & w2637 ) | ( w2579 & w2637 ) ;
  assign w2750 = ( w2651 & w2652 ) | ( w2651 & w2653 ) | ( w2652 & w2653 ) ;
  assign w2751 = ( w2658 & w2659 ) | ( w2658 & w2665 ) | ( w2659 & w2665 ) ;
  assign w2752 = ( w2485 & w2491 ) | ( w2485 & w2520 ) | ( w2491 & w2520 ) ;
  assign w2753 = ( w2508 & w2514 ) | ( w2508 & w2552 ) | ( w2514 & w2552 ) ;
  assign w2754 = w2594 ^ w2602 ;
  assign w2755 = w2622 ^ w2754 ;
  assign w2756 = w2752 ^ w2753 ;
  assign w2757 = w2755 ^ w2756 ;
  assign w2758 = w2750 ^ w2751 ;
  assign w2759 = w2757 ^ w2758 ;
  assign w2760 = ( w2604 & w2610 ) | ( w2604 & w2616 ) | ( w2610 & w2616 ) ;
  assign w2761 = ( w2624 & w2627 ) | ( w2624 & w2633 ) | ( w2627 & w2633 ) ;
  assign w2762 = \pi24 & \pi26 ;
  assign w2763 = w2588 ^ w2762 ;
  assign w2764 = w2614 ^ w2763 ;
  assign w2765 = \pi01 & \pi49 ;
  assign w2766 = w2764 ^ w2765 ;
  assign w2767 = w2761 ^ w2766 ;
  assign w2768 = w2760 ^ w2767 ;
  assign w2769 = w2583 ^ w2608 ;
  assign w2770 = w2631 ^ w2769 ;
  assign w2771 = ( w2585 & w2590 ) | ( w2585 & w2596 ) | ( w2590 & w2596 ) ;
  assign w2772 = ( w2641 & w2642 ) | ( w2641 & w2643 ) | ( w2642 & w2643 ) ;
  assign w2773 = w2771 ^ w2772 ;
  assign w2774 = w2770 ^ w2773 ;
  assign w2775 = ( w2598 & w2618 ) | ( w2598 & w2635 ) | ( w2618 & w2635 ) ;
  assign w2776 = w2768 ^ w2774 ;
  assign w2777 = w2775 ^ w2776 ;
  assign w2778 = w2749 ^ w2777 ;
  assign w2779 = w2759 ^ w2778 ;
  assign w2780 = w2681 ^ w2779 ;
  assign w2781 = w2748 ^ w2780 ;
  assign w2782 = w2680 | w2781 ;
  assign w2783 = w2680 & w2781 ;
  assign w2784 = w2782 & ~w2783 ;
  assign w2785 = w2679 ^ w2784 ;
  assign w2786 = ( w2679 & w2782 ) | ( w2679 & w2783 ) | ( w2782 & w2783 ) ;
  assign w2787 = w2783 | w2786 ;
  assign w2788 = ( w2681 & w2748 ) | ( w2681 & w2779 ) | ( w2748 & w2779 ) ;
  assign w2789 = ( w2749 & w2759 ) | ( w2749 & w2777 ) | ( w2759 & w2777 ) ;
  assign w2790 = ( w2768 & w2774 ) | ( w2768 & w2775 ) | ( w2774 & w2775 ) ;
  assign w2791 = ( w2750 & w2751 ) | ( w2750 & w2757 ) | ( w2751 & w2757 ) ;
  assign w2792 = \pi00 & \pi51 ;
  assign w2793 = ( \pi01 & \pi24 ) | ( \pi01 & ~\pi26 ) | ( \pi24 & ~\pi26 ) ;
  assign w2794 = ( \pi26 & ~\pi49 ) | ( \pi26 & w2793 ) | ( ~\pi49 & w2793 ) ;
  assign w2795 = \pi49 & w2794 ;
  assign w2796 = w2792 ^ w2795 ;
  assign w2797 = \pi20 & \pi31 ;
  assign w2798 = \pi19 & \pi32 ;
  assign w2799 = \pi17 & \pi34 ;
  assign w2800 = ( w2797 & w2798 ) | ( w2797 & w2799 ) | ( w2798 & w2799 ) ;
  assign w2801 = w2797 ^ w2799 ;
  assign w2802 = w2798 ^ w2801 ;
  assign w2803 = ( w2583 & w2608 ) | ( w2583 & w2631 ) | ( w2608 & w2631 ) ;
  assign w2804 = w2796 ^ w2803 ;
  assign w2805 = w2802 ^ w2804 ;
  assign w2806 = \pi26 ^ w2805 ;
  assign w2807 = \pi01 & \pi50 ;
  assign w2808 = w2806 ^ w2807 ;
  assign w2809 = \pi18 & \pi33 ;
  assign w2810 = \pi16 & \pi35 ;
  assign w2811 = \pi05 & \pi46 ;
  assign w2812 = ( w2809 & w2810 ) | ( w2809 & w2811 ) | ( w2810 & w2811 ) ;
  assign w2813 = w2809 ^ w2811 ;
  assign w2814 = w2810 ^ w2813 ;
  assign w2815 = \pi23 & \pi28 ;
  assign w2816 = \pi22 & \pi29 ;
  assign w2817 = \pi21 & \pi30 ;
  assign w2818 = ( w2815 & w2816 ) | ( w2815 & w2817 ) | ( w2816 & w2817 ) ;
  assign w2819 = w2815 ^ w2817 ;
  assign w2820 = w2816 ^ w2819 ;
  assign w2821 = \pi15 & \pi36 ;
  assign w2822 = \pi14 & \pi37 ;
  assign w2823 = \pi06 & \pi45 ;
  assign w2824 = ( w2821 & w2822 ) | ( w2821 & w2823 ) | ( w2822 & w2823 ) ;
  assign w2825 = w2821 ^ w2823 ;
  assign w2826 = w2822 ^ w2825 ;
  assign w2827 = w2814 ^ w2820 ;
  assign w2828 = w2826 ^ w2827 ;
  assign w2829 = \pi13 & \pi38 ;
  assign w2830 = \pi08 & \pi43 ;
  assign w2831 = \pi07 & \pi44 ;
  assign w2832 = ( w2829 & w2830 ) | ( w2829 & w2831 ) | ( w2830 & w2831 ) ;
  assign w2833 = w2829 ^ w2831 ;
  assign w2834 = w2830 ^ w2833 ;
  assign w2835 = \pi12 & \pi39 ;
  assign w2836 = \pi10 & \pi41 ;
  assign w2837 = \pi09 & \pi42 ;
  assign w2838 = ( w2835 & w2836 ) | ( w2835 & w2837 ) | ( w2836 & w2837 ) ;
  assign w2839 = w2835 ^ w2837 ;
  assign w2840 = w2836 ^ w2839 ;
  assign w2841 = \pi25 & \pi26 ;
  assign w2842 = \pi24 & \pi27 ;
  assign w2843 = \pi11 & \pi40 ;
  assign w2844 = ( w2841 & w2842 ) | ( w2841 & w2843 ) | ( w2842 & w2843 ) ;
  assign w2845 = w2841 ^ w2843 ;
  assign w2846 = w2842 ^ w2845 ;
  assign w2847 = w2834 ^ w2840 ;
  assign w2848 = w2846 ^ w2847 ;
  assign w2849 = w2808 ^ w2828 ;
  assign w2850 = w2848 ^ w2849 ;
  assign w2851 = w2790 ^ w2791 ;
  assign w2852 = w2850 ^ w2851 ;
  assign w2853 = ( w2682 & w2683 ) | ( w2682 & w2746 ) | ( w2683 & w2746 ) ;
  assign w2854 = ( w2770 & w2771 ) | ( w2770 & w2772 ) | ( w2771 & w2772 ) ;
  assign w2855 = ( w2760 & w2761 ) | ( w2760 & w2766 ) | ( w2761 & w2766 ) ;
  assign w2856 = ( w2594 & w2602 ) | ( w2594 & w2622 ) | ( w2602 & w2622 ) ;
  assign w2857 = w2762 ^ w2765 ;
  assign w2858 = ( w2588 & w2614 ) | ( w2588 & w2857 ) | ( w2614 & w2857 ) ;
  assign w2859 = ( w2710 & w2716 ) | ( w2710 & w2722 ) | ( w2716 & w2722 ) ;
  assign w2860 = w2858 ^ w2859 ;
  assign w2861 = w2856 ^ w2860 ;
  assign w2862 = w2854 ^ w2855 ;
  assign w2863 = w2861 ^ w2862 ;
  assign w2864 = ( w2703 & w2724 ) | ( w2703 & w2744 ) | ( w2724 & w2744 ) ;
  assign w2865 = \pi04 & \pi47 ;
  assign w2866 = \pi03 & \pi48 ;
  assign w2867 = \pi02 & \pi49 ;
  assign w2868 = ( w2865 & w2866 ) | ( w2865 & w2867 ) | ( w2866 & w2867 ) ;
  assign w2869 = w2865 ^ w2867 ;
  assign w2870 = w2866 ^ w2869 ;
  assign w2871 = w2687 ^ w2740 ;
  assign w2872 = w2870 ^ w2871 ;
  assign w2873 = ( w2689 & w2695 ) | ( w2689 & w2701 ) | ( w2695 & w2701 ) ;
  assign w2874 = ( w2752 & w2753 ) | ( w2752 & w2755 ) | ( w2753 & w2755 ) ;
  assign w2875 = w2873 ^ w2874 ;
  assign w2876 = w2872 ^ w2875 ;
  assign w2877 = w2693 ^ w2728 ;
  assign w2878 = w2734 ^ w2877 ;
  assign w2879 = ( w2730 & w2736 ) | ( w2730 & w2742 ) | ( w2736 & w2742 ) ;
  assign w2880 = w2706 ^ w2714 ;
  assign w2881 = w2720 ^ w2880 ;
  assign w2882 = w2878 ^ w2881 ;
  assign w2883 = w2879 ^ w2882 ;
  assign w2884 = w2864 ^ w2876 ;
  assign w2885 = w2883 ^ w2884 ;
  assign w2886 = w2853 ^ w2863 ;
  assign w2887 = w2885 ^ w2886 ;
  assign w2888 = w2789 ^ w2852 ;
  assign w2889 = w2887 ^ w2888 ;
  assign w2890 = w2787 ^ w2788 ;
  assign w2891 = w2889 ^ w2890 ;
  assign w2892 = ( w2787 & w2788 ) | ( w2787 & w2889 ) | ( w2788 & w2889 ) ;
  assign w2893 = ( w2789 & w2852 ) | ( w2789 & w2887 ) | ( w2852 & w2887 ) ;
  assign w2894 = ( w2790 & w2791 ) | ( w2790 & w2850 ) | ( w2791 & w2850 ) ;
  assign w2895 = ( w2706 & w2714 ) | ( w2706 & w2720 ) | ( w2714 & w2720 ) ;
  assign w2896 = \pi19 & \pi33 ;
  assign w2897 = \pi03 & \pi49 ;
  assign w2898 = \pi02 & \pi50 ;
  assign w2899 = ( w2896 & w2897 ) | ( w2896 & w2898 ) | ( w2897 & w2898 ) ;
  assign w2900 = w2896 ^ w2898 ;
  assign w2901 = w2897 ^ w2900 ;
  assign w2902 = ( w2693 & w2728 ) | ( w2693 & w2734 ) | ( w2728 & w2734 ) ;
  assign w2903 = w2895 ^ w2902 ;
  assign w2904 = w2901 ^ w2903 ;
  assign w2905 = ( w2872 & w2873 ) | ( w2872 & w2874 ) | ( w2873 & w2874 ) ;
  assign w2906 = ( w2834 & w2840 ) | ( w2834 & w2846 ) | ( w2840 & w2846 ) ;
  assign w2907 = ( w2687 & w2740 ) | ( w2687 & w2870 ) | ( w2740 & w2870 ) ;
  assign w2908 = ( ~\pi01 & \pi51 ) | ( ~\pi01 & w1228 ) | ( \pi51 & w1228 ) ;
  assign w2909 = \pi01 & w2908 ;
  assign w2910 = ( ~\pi01 & \pi26 ) | ( ~\pi01 & \pi50 ) | ( \pi26 & \pi50 ) ;
  assign w2911 = \pi51 ^ w2910 ;
  assign w2912 = \pi01 & w2911 ;
  assign w2913 = w1228 ^ w2844 ;
  assign w2914 = w2912 ^ w2913 ;
  assign w2915 = w2906 ^ w2907 ;
  assign w2916 = w2914 ^ w2915 ;
  assign w2917 = w2904 ^ w2905 ;
  assign w2918 = w2916 ^ w2917 ;
  assign w2919 = \pi24 & \pi49 ;
  assign w2920 = ( ~\pi50 & w2792 ) | ( ~\pi50 & w2919 ) | ( w2792 & w2919 ) ;
  assign w2921 = \pi26 & w2920 ;
  assign w2922 = ( \pi01 & \pi26 ) | ( \pi01 & ~\pi50 ) | ( \pi26 & ~\pi50 ) ;
  assign w2923 = ( \pi01 & \pi26 ) | ( \pi01 & w2792 ) | ( \pi26 & w2792 ) ;
  assign w2924 = ( w2921 & ~w2922 ) | ( w2921 & w2923 ) | ( ~w2922 & w2923 ) ;
  assign w2925 = \pi04 & \pi48 ;
  assign w2926 = \pi00 & \pi52 ;
  assign w2927 = ( w1620 & w2925 ) | ( w1620 & w2926 ) | ( w2925 & w2926 ) ;
  assign w2928 = w1620 ^ w2926 ;
  assign w2929 = w2925 ^ w2928 ;
  assign w2930 = w2838 ^ w2924 ;
  assign w2931 = w2929 ^ w2930 ;
  assign w2932 = \pi26 ^ w2796 ;
  assign w2933 = w2807 ^ w2932 ;
  assign w2934 = ( w2802 & w2803 ) | ( w2802 & w2933 ) | ( w2803 & w2933 ) ;
  assign w2935 = ( w2856 & w2858 ) | ( w2856 & w2859 ) | ( w2858 & w2859 ) ;
  assign w2936 = w2931 ^ w2935 ;
  assign w2937 = w2934 ^ w2936 ;
  assign w2938 = ( w2808 & w2828 ) | ( w2808 & w2848 ) | ( w2828 & w2848 ) ;
  assign w2939 = w2812 ^ w2818 ;
  assign w2940 = w2832 ^ w2939 ;
  assign w2941 = w2800 ^ w2824 ;
  assign w2942 = w2868 ^ w2941 ;
  assign w2943 = ( w2814 & w2820 ) | ( w2814 & w2826 ) | ( w2820 & w2826 ) ;
  assign w2944 = w2940 ^ w2942 ;
  assign w2945 = w2943 ^ w2944 ;
  assign w2946 = w2937 ^ w2938 ;
  assign w2947 = w2945 ^ w2946 ;
  assign w2948 = w2894 ^ w2947 ;
  assign w2949 = w2918 ^ w2948 ;
  assign w2950 = ( w2864 & w2876 ) | ( w2864 & w2883 ) | ( w2876 & w2883 ) ;
  assign w2951 = ( w2854 & w2855 ) | ( w2854 & w2861 ) | ( w2855 & w2861 ) ;
  assign w2952 = ( w2878 & w2879 ) | ( w2878 & w2881 ) | ( w2879 & w2881 ) ;
  assign w2953 = \pi16 & \pi36 ;
  assign w2954 = \pi06 & \pi46 ;
  assign w2955 = \pi05 & \pi47 ;
  assign w2956 = ( w2953 & w2954 ) | ( w2953 & w2955 ) | ( w2954 & w2955 ) ;
  assign w2957 = w2953 ^ w2955 ;
  assign w2958 = w2954 ^ w2957 ;
  assign w2959 = \pi40 & \pi42 ;
  assign w2960 = \pi12 & \pi40 ;
  assign w2961 = \pi11 & \pi41 ;
  assign w2962 = \pi10 & \pi42 ;
  assign w2963 = ( w2960 & w2961 ) | ( w2960 & w2962 ) | ( w2961 & w2962 ) ;
  assign w2964 = w2960 ^ w2962 ;
  assign w2965 = w2961 ^ w2964 ;
  assign w2966 = \pi15 & \pi37 ;
  assign w2967 = \pi08 & \pi44 ;
  assign w2968 = \pi07 & \pi45 ;
  assign w2969 = ( w2966 & w2967 ) | ( w2966 & w2968 ) | ( w2967 & w2968 ) ;
  assign w2970 = w2966 ^ w2968 ;
  assign w2971 = w2967 ^ w2970 ;
  assign w2972 = w2958 ^ w2965 ;
  assign w2973 = w2971 ^ w2972 ;
  assign w2974 = \pi21 & \pi31 ;
  assign w2975 = \pi20 & \pi32 ;
  assign w2976 = \pi18 & \pi34 ;
  assign w2977 = ( w2974 & w2975 ) | ( w2974 & w2976 ) | ( w2975 & w2976 ) ;
  assign w2978 = w2974 ^ w2976 ;
  assign w2979 = w2975 ^ w2978 ;
  assign w2980 = \pi24 & \pi28 ;
  assign w2981 = \pi23 & \pi29 ;
  assign w2982 = \pi22 & \pi30 ;
  assign w2983 = ( w2980 & w2981 ) | ( w2980 & w2982 ) | ( w2981 & w2982 ) ;
  assign w2984 = w2980 ^ w2982 ;
  assign w2985 = w2981 ^ w2984 ;
  assign w2986 = \pi14 & \pi38 ;
  assign w2987 = \pi13 & \pi39 ;
  assign w2988 = \pi09 & \pi43 ;
  assign w2989 = ( w2986 & w2987 ) | ( w2986 & w2988 ) | ( w2987 & w2988 ) ;
  assign w2990 = w2986 ^ w2988 ;
  assign w2991 = w2987 ^ w2990 ;
  assign w2992 = w2979 ^ w2985 ;
  assign w2993 = w2991 ^ w2992 ;
  assign w2994 = w2952 ^ w2973 ;
  assign w2995 = w2993 ^ w2994 ;
  assign w2996 = w2950 ^ w2951 ;
  assign w2997 = w2995 ^ w2996 ;
  assign w2998 = ( w2853 & w2863 ) | ( w2853 & w2885 ) | ( w2863 & w2885 ) ;
  assign w2999 = w2949 ^ w2997 ;
  assign w3000 = w2998 ^ w2999 ;
  assign w3001 = w2893 | w3000 ;
  assign w3002 = w2893 & w3000 ;
  assign w3003 = w3001 & ~w3002 ;
  assign w3004 = w2892 ^ w3003 ;
  assign w3005 = ( w2892 & w3001 ) | ( w2892 & w3002 ) | ( w3001 & w3002 ) ;
  assign w3006 = w3002 | w3005 ;
  assign w3007 = ( w2949 & w2997 ) | ( w2949 & w2998 ) | ( w2997 & w2998 ) ;
  assign w3008 = ( w2894 & w2918 ) | ( w2894 & w2947 ) | ( w2918 & w2947 ) ;
  assign w3009 = ( w2937 & w2938 ) | ( w2937 & w2945 ) | ( w2938 & w2945 ) ;
  assign w3010 = \pi03 & \pi50 ;
  assign w3011 = \pi02 & \pi51 ;
  assign w3012 = ( w2909 & w3010 ) | ( w2909 & w3011 ) | ( w3010 & w3011 ) ;
  assign w3013 = w2909 ^ w3011 ;
  assign w3014 = w3010 ^ w3013 ;
  assign w3015 = \pi18 & \pi35 ;
  assign w3016 = \pi17 & \pi36 ;
  assign w3017 = \pi04 & \pi49 ;
  assign w3018 = ( w3015 & w3016 ) | ( w3015 & w3017 ) | ( w3016 & w3017 ) ;
  assign w3019 = w3015 ^ w3017 ;
  assign w3020 = w3016 ^ w3019 ;
  assign w3021 = \pi21 & \pi32 ;
  assign w3022 = \pi20 & \pi33 ;
  assign w3023 = \pi19 & \pi34 ;
  assign w3024 = ( w3021 & w3022 ) | ( w3021 & w3023 ) | ( w3022 & w3023 ) ;
  assign w3025 = w3021 ^ w3023 ;
  assign w3026 = w3022 ^ w3025 ;
  assign w3027 = w3014 ^ w3020 ;
  assign w3028 = w3026 ^ w3027 ;
  assign w3029 = ( w2895 & w2901 ) | ( w2895 & w2902 ) | ( w2901 & w2902 ) ;
  assign w3030 = \pi07 & \pi46 ;
  assign w3031 = \pi06 & \pi47 ;
  assign w3032 = ( w1948 & w3030 ) | ( w1948 & w3031 ) | ( w3030 & w3031 ) ;
  assign w3033 = w1948 ^ w3031 ;
  assign w3034 = w3030 ^ w3033 ;
  assign w3035 = \pi14 & \pi39 ;
  assign w3036 = \pi09 & \pi44 ;
  assign w3037 = \pi08 & \pi45 ;
  assign w3038 = ( w3035 & w3036 ) | ( w3035 & w3037 ) | ( w3036 & w3037 ) ;
  assign w3039 = w3035 ^ w3037 ;
  assign w3040 = w3036 ^ w3039 ;
  assign w3041 = \pi16 & \pi37 ;
  assign w3042 = \pi05 & \pi48 ;
  assign w3043 = \pi00 & \pi53 ;
  assign w3044 = ( w3041 & w3042 ) | ( w3041 & w3043 ) | ( w3042 & w3043 ) ;
  assign w3045 = w3041 ^ w3043 ;
  assign w3046 = w3042 ^ w3045 ;
  assign w3047 = w3034 ^ w3040 ;
  assign w3048 = w3046 ^ w3047 ;
  assign w3049 = w3028 ^ w3029 ;
  assign w3050 = w3048 ^ w3049 ;
  assign w3051 = \pi13 & \pi40 ;
  assign w3052 = \pi12 & \pi41 ;
  assign w3053 = \pi10 & \pi43 ;
  assign w3054 = ( w3051 & w3052 ) | ( w3051 & w3053 ) | ( w3052 & w3053 ) ;
  assign w3055 = w3051 ^ w3053 ;
  assign w3056 = w3052 ^ w3055 ;
  assign w3057 = \pi24 & \pi29 ;
  assign w3058 = \pi23 & \pi30 ;
  assign w3059 = \pi22 & \pi31 ;
  assign w3060 = ( w3057 & w3058 ) | ( w3057 & w3059 ) | ( w3058 & w3059 ) ;
  assign w3061 = w3057 ^ w3059 ;
  assign w3062 = w3058 ^ w3061 ;
  assign w3063 = \pi26 & \pi27 ;
  assign w3064 = \pi25 & \pi28 ;
  assign w3065 = \pi11 & \pi42 ;
  assign w3066 = ( w3063 & w3064 ) | ( w3063 & w3065 ) | ( w3064 & w3065 ) ;
  assign w3067 = w3063 ^ w3065 ;
  assign w3068 = w3064 ^ w3067 ;
  assign w3069 = w3056 ^ w3062 ;
  assign w3070 = w3068 ^ w3069 ;
  assign w3071 = ( w2906 & w2907 ) | ( w2906 & w2914 ) | ( w2907 & w2914 ) ;
  assign w3072 = ( w2940 & w2942 ) | ( w2940 & w2943 ) | ( w2942 & w2943 ) ;
  assign w3073 = w3071 ^ w3072 ;
  assign w3074 = w3070 ^ w3073 ;
  assign w3075 = w3009 ^ w3050 ;
  assign w3076 = w3074 ^ w3075 ;
  assign w3077 = w2956 ^ w2969 ;
  assign w3078 = w2977 ^ w3077 ;
  assign w3079 = ( w2958 & w2965 ) | ( w2958 & w2971 ) | ( w2965 & w2971 ) ;
  assign w3080 = ( \pi01 & ~\pi27 ) | ( \pi01 & \pi52 ) | ( ~\pi27 & \pi52 ) ;
  assign w3081 = \pi27 & w3080 ;
  assign w3082 = \pi01 & \pi52 ;
  assign w3083 = \pi27 ^ w2989 ;
  assign w3084 = w2963 ^ w3083 ;
  assign w3085 = w3082 ^ w3084 ;
  assign w3086 = w3078 ^ w3079 ;
  assign w3087 = w3085 ^ w3086 ;
  assign w3088 = w2899 ^ w2927 ;
  assign w3089 = w2983 ^ w3088 ;
  assign w3090 = ( w2979 & w2985 ) | ( w2979 & w2991 ) | ( w2985 & w2991 ) ;
  assign w3091 = ( w2838 & w2924 ) | ( w2838 & w2929 ) | ( w2924 & w2929 ) ;
  assign w3092 = w3089 ^ w3091 ;
  assign w3093 = w3090 ^ w3092 ;
  assign w3094 = ( w2904 & w2905 ) | ( w2904 & w2916 ) | ( w2905 & w2916 ) ;
  assign w3095 = w3093 ^ w3094 ;
  assign w3096 = w3087 ^ w3095 ;
  assign w3097 = ( w2952 & w2973 ) | ( w2952 & w2993 ) | ( w2973 & w2993 ) ;
  assign w3098 = ( w2812 & w2818 ) | ( w2812 & w2832 ) | ( w2818 & w2832 ) ;
  assign w3099 = \pi50 & w854 ;
  assign w3100 = \pi01 & \pi51 ;
  assign w3101 = w1228 ^ w3100 ;
  assign w3102 = ( w2844 & w3099 ) | ( w2844 & w3101 ) | ( w3099 & w3101 ) ;
  assign w3103 = ( w2800 & w2824 ) | ( w2800 & w2868 ) | ( w2824 & w2868 ) ;
  assign w3104 = w3098 ^ w3102 ;
  assign w3105 = w3103 ^ w3104 ;
  assign w3106 = ( w2931 & w2934 ) | ( w2931 & w2935 ) | ( w2934 & w2935 ) ;
  assign w3107 = w3097 ^ w3106 ;
  assign w3108 = w3105 ^ w3107 ;
  assign w3109 = ( w2950 & w2951 ) | ( w2950 & w2995 ) | ( w2951 & w2995 ) ;
  assign w3110 = w3096 ^ w3109 ;
  assign w3111 = w3108 ^ w3110 ;
  assign w3112 = w3008 ^ w3111 ;
  assign w3113 = w3076 ^ w3112 ;
  assign w3114 = w3006 ^ w3007 ;
  assign w3115 = w3113 ^ w3114 ;
  assign w3116 = ( w3008 & w3076 ) | ( w3008 & w3111 ) | ( w3076 & w3111 ) ;
  assign w3117 = ( w3087 & w3093 ) | ( w3087 & w3094 ) | ( w3093 & w3094 ) ;
  assign w3118 = ( w3097 & w3105 ) | ( w3097 & w3106 ) | ( w3105 & w3106 ) ;
  assign w3119 = ( w3078 & w3079 ) | ( w3078 & w3085 ) | ( w3079 & w3085 ) ;
  assign w3120 = ( w3089 & w3090 ) | ( w3089 & w3091 ) | ( w3090 & w3091 ) ;
  assign w3121 = ( ~\pi01 & \pi53 ) | ( ~\pi01 & w1305 ) | ( \pi53 & w1305 ) ;
  assign w3122 = \pi01 & w3121 ;
  assign w3123 = \pi01 & \pi53 ;
  assign w3124 = w1305 ^ w3123 ;
  assign w3125 = w3081 ^ w3124 ;
  assign w3126 = \pi00 & \pi54 ;
  assign w3127 = w3125 ^ w3126 ;
  assign w3128 = \pi22 & \pi32 ;
  assign w3129 = \pi21 & \pi33 ;
  assign w3130 = \pi19 & \pi35 ;
  assign w3131 = ( w3128 & w3129 ) | ( w3128 & w3130 ) | ( w3129 & w3130 ) ;
  assign w3132 = w3128 ^ w3130 ;
  assign w3133 = w3129 ^ w3132 ;
  assign w3134 = \pi25 & \pi29 ;
  assign w3135 = \pi24 & \pi30 ;
  assign w3136 = \pi23 & \pi31 ;
  assign w3137 = ( w3134 & w3135 ) | ( w3134 & w3136 ) | ( w3135 & w3136 ) ;
  assign w3138 = w3134 ^ w3136 ;
  assign w3139 = w3135 ^ w3138 ;
  assign w3140 = w3127 ^ w3133 ;
  assign w3141 = w3139 ^ w3140 ;
  assign w3142 = w3119 ^ w3120 ;
  assign w3143 = w3141 ^ w3142 ;
  assign w3144 = w3117 ^ w3118 ;
  assign w3145 = w3143 ^ w3144 ;
  assign w3146 = ( w3096 & w3108 ) | ( w3096 & w3109 ) | ( w3108 & w3109 ) ;
  assign w3147 = ( w3009 & w3050 ) | ( w3009 & w3074 ) | ( w3050 & w3074 ) ;
  assign w3148 = ( w2956 & w2969 ) | ( w2956 & w2977 ) | ( w2969 & w2977 ) ;
  assign w3149 = ( w2899 & w2927 ) | ( w2899 & w2983 ) | ( w2927 & w2983 ) ;
  assign w3150 = \pi27 ^ w3082 ;
  assign w3151 = ( w2963 & w2989 ) | ( w2963 & w3150 ) | ( w2989 & w3150 ) ;
  assign w3152 = w3148 ^ w3149 ;
  assign w3153 = w3151 ^ w3152 ;
  assign w3154 = ( w3028 & w3029 ) | ( w3028 & w3048 ) | ( w3029 & w3048 ) ;
  assign w3155 = w3032 ^ w3044 ;
  assign w3156 = w3066 ^ w3155 ;
  assign w3157 = w3018 ^ w3024 ;
  assign w3158 = w3060 ^ w3157 ;
  assign w3159 = ( w3034 & w3040 ) | ( w3034 & w3046 ) | ( w3040 & w3046 ) ;
  assign w3160 = w3156 ^ w3159 ;
  assign w3161 = w3158 ^ w3160 ;
  assign w3162 = w3154 ^ w3161 ;
  assign w3163 = w3153 ^ w3162 ;
  assign w3164 = \pi20 & \pi34 ;
  assign w3165 = \pi18 & \pi36 ;
  assign w3166 = \pi05 & \pi49 ;
  assign w3167 = ( w3164 & w3165 ) | ( w3164 & w3166 ) | ( w3165 & w3166 ) ;
  assign w3168 = w3164 ^ w3166 ;
  assign w3169 = w3165 ^ w3168 ;
  assign w3170 = \pi13 & \pi41 ;
  assign w3171 = \pi12 & \pi42 ;
  assign w3172 = \pi11 & \pi43 ;
  assign w3173 = ( w3170 & w3171 ) | ( w3170 & w3172 ) | ( w3171 & w3172 ) ;
  assign w3174 = w3170 ^ w3172 ;
  assign w3175 = w3171 ^ w3174 ;
  assign w3176 = \pi38 & \pi48 ;
  assign w3177 = \pi17 & \pi37 ;
  assign w3178 = \pi16 & \pi38 ;
  assign w3179 = \pi06 & \pi48 ;
  assign w3180 = ( w3177 & w3178 ) | ( w3177 & w3179 ) | ( w3178 & w3179 ) ;
  assign w3181 = w3177 ^ w3179 ;
  assign w3182 = w3178 ^ w3181 ;
  assign w3183 = w3169 ^ w3175 ;
  assign w3184 = w3182 ^ w3183 ;
  assign w3185 = ( w3098 & w3102 ) | ( w3098 & w3103 ) | ( w3102 & w3103 ) ;
  assign w3186 = \pi04 & \pi50 ;
  assign w3187 = \pi03 & \pi51 ;
  assign w3188 = \pi02 & \pi52 ;
  assign w3189 = ( w3186 & w3187 ) | ( w3186 & w3188 ) | ( w3187 & w3188 ) ;
  assign w3190 = w3186 ^ w3188 ;
  assign w3191 = w3187 ^ w3190 ;
  assign w3192 = \pi15 & \pi39 ;
  assign w3193 = \pi08 & \pi46 ;
  assign w3194 = \pi07 & \pi47 ;
  assign w3195 = ( w3192 & w3193 ) | ( w3192 & w3194 ) | ( w3193 & w3194 ) ;
  assign w3196 = w3192 ^ w3194 ;
  assign w3197 = w3193 ^ w3196 ;
  assign w3198 = \pi14 & \pi40 ;
  assign w3199 = \pi10 & \pi44 ;
  assign w3200 = \pi09 & \pi45 ;
  assign w3201 = ( w3198 & w3199 ) | ( w3198 & w3200 ) | ( w3199 & w3200 ) ;
  assign w3202 = w3198 ^ w3200 ;
  assign w3203 = w3199 ^ w3202 ;
  assign w3204 = w3191 ^ w3197 ;
  assign w3205 = w3203 ^ w3204 ;
  assign w3206 = w3185 ^ w3205 ;
  assign w3207 = w3184 ^ w3206 ;
  assign w3208 = ( w3070 & w3071 ) | ( w3070 & w3072 ) | ( w3071 & w3072 ) ;
  assign w3209 = w3012 ^ w3038 ;
  assign w3210 = w3054 ^ w3209 ;
  assign w3211 = ( w3056 & w3062 ) | ( w3056 & w3068 ) | ( w3062 & w3068 ) ;
  assign w3212 = ( w3014 & w3020 ) | ( w3014 & w3026 ) | ( w3020 & w3026 ) ;
  assign w3213 = w3210 ^ w3212 ;
  assign w3214 = w3211 ^ w3213 ;
  assign w3215 = w3207 ^ w3214 ;
  assign w3216 = w3208 ^ w3215 ;
  assign w3217 = w3147 ^ w3163 ;
  assign w3218 = w3216 ^ w3217 ;
  assign w3219 = w3146 ^ w3218 ;
  assign w3220 = w3145 ^ w3219 ;
  assign w3221 = ( w3006 & w3007 ) | ( w3006 & w3113 ) | ( w3007 & w3113 ) ;
  assign w3222 = w3116 ^ w3221 ;
  assign w3223 = w3220 ^ w3222 ;
  assign w3224 = ( w3145 & w3146 ) | ( w3145 & w3218 ) | ( w3146 & w3218 ) ;
  assign w3225 = ( w3147 & w3163 ) | ( w3147 & w3216 ) | ( w3163 & w3216 ) ;
  assign w3226 = ( w3207 & w3208 ) | ( w3207 & w3214 ) | ( w3208 & w3214 ) ;
  assign w3227 = ( w3153 & w3154 ) | ( w3153 & w3161 ) | ( w3154 & w3161 ) ;
  assign w3228 = ( w3156 & w3158 ) | ( w3156 & w3159 ) | ( w3158 & w3159 ) ;
  assign w3229 = \pi17 & \pi38 ;
  assign w3230 = \pi06 & \pi49 ;
  assign w3231 = \pi03 & \pi52 ;
  assign w3232 = ( w3229 & w3230 ) | ( w3229 & w3231 ) | ( w3230 & w3231 ) ;
  assign w3233 = w3229 ^ w3231 ;
  assign w3234 = w3230 ^ w3233 ;
  assign w3235 = \pi15 & \pi40 ;
  assign w3236 = \pi14 & \pi41 ;
  assign w3237 = \pi09 & \pi46 ;
  assign w3238 = ( w3235 & w3236 ) | ( w3235 & w3237 ) | ( w3236 & w3237 ) ;
  assign w3239 = w3235 ^ w3237 ;
  assign w3240 = w3236 ^ w3239 ;
  assign w3241 = ( w3018 & w3024 ) | ( w3018 & w3060 ) | ( w3024 & w3060 ) ;
  assign w3242 = w3234 ^ w3241 ;
  assign w3243 = w3240 ^ w3242 ;
  assign w3244 = ( w3210 & w3211 ) | ( w3210 & w3212 ) | ( w3211 & w3212 ) ;
  assign w3245 = w3228 ^ w3244 ;
  assign w3246 = w3243 ^ w3245 ;
  assign w3247 = w3226 ^ w3227 ;
  assign w3248 = w3246 ^ w3247 ;
  assign w3249 = ( w3032 & w3044 ) | ( w3032 & w3066 ) | ( w3044 & w3066 ) ;
  assign w3250 = ( w3012 & w3038 ) | ( w3012 & w3054 ) | ( w3038 & w3054 ) ;
  assign w3251 = \pi01 & \pi54 ;
  assign w3252 = \pi28 ^ w3173 ;
  assign w3253 = w3122 ^ w3252 ;
  assign w3254 = w3251 ^ w3253 ;
  assign w3255 = w3249 ^ w3250 ;
  assign w3256 = w3254 ^ w3255 ;
  assign w3257 = ( w3184 & w3185 ) | ( w3184 & w3205 ) | ( w3185 & w3205 ) ;
  assign w3258 = ( w3081 & w3124 ) | ( w3081 & w3126 ) | ( w3124 & w3126 ) ;
  assign w3259 = \pi19 & \pi36 ;
  assign w3260 = \pi05 & \pi50 ;
  assign w3261 = ( w1756 & w3259 ) | ( w1756 & w3260 ) | ( w3259 & w3260 ) ;
  assign w3262 = w3259 ^ w3260 ;
  assign w3263 = w1756 ^ w3262 ;
  assign w3264 = w3195 ^ w3258 ;
  assign w3265 = w3263 ^ w3264 ;
  assign w3266 = w3167 ^ w3189 ;
  assign w3267 = w3201 ^ w3266 ;
  assign w3268 = ( w3127 & w3133 ) | ( w3127 & w3139 ) | ( w3133 & w3139 ) ;
  assign w3269 = w3265 ^ w3268 ;
  assign w3270 = w3267 ^ w3269 ;
  assign w3271 = w3256 ^ w3257 ;
  assign w3272 = w3270 ^ w3271 ;
  assign w3273 = ( w3117 & w3118 ) | ( w3117 & w3143 ) | ( w3118 & w3143 ) ;
  assign w3274 = \pi13 & \pi42 ;
  assign w3275 = \pi11 & \pi44 ;
  assign w3276 = \pi10 & \pi45 ;
  assign w3277 = ( w3274 & w3275 ) | ( w3274 & w3276 ) | ( w3275 & w3276 ) ;
  assign w3278 = w3274 ^ w3276 ;
  assign w3279 = w3275 ^ w3278 ;
  assign w3280 = \pi26 & \pi29 ;
  assign w3281 = \pi12 & \pi43 ;
  assign w3282 = ( w1088 & w3280 ) | ( w1088 & w3281 ) | ( w3280 & w3281 ) ;
  assign w3283 = w1088 ^ w3281 ;
  assign w3284 = w3280 ^ w3283 ;
  assign w3285 = \pi16 & \pi39 ;
  assign w3286 = \pi08 & \pi47 ;
  assign w3287 = \pi07 & \pi48 ;
  assign w3288 = ( w3285 & w3286 ) | ( w3285 & w3287 ) | ( w3286 & w3287 ) ;
  assign w3289 = w3285 ^ w3287 ;
  assign w3290 = w3286 ^ w3289 ;
  assign w3291 = w3279 ^ w3284 ;
  assign w3292 = w3290 ^ w3291 ;
  assign w3293 = ( w3148 & w3149 ) | ( w3148 & w3151 ) | ( w3149 & w3151 ) ;
  assign w3294 = w3292 ^ w3293 ;
  assign w3295 = \pi04 & \pi51 ;
  assign w3296 = \pi02 & \pi53 ;
  assign w3297 = \pi00 & \pi55 ;
  assign w3298 = ( w3295 & w3296 ) | ( w3295 & w3297 ) | ( w3296 & w3297 ) ;
  assign w3299 = w3295 ^ w3297 ;
  assign w3300 = w3296 ^ w3299 ;
  assign w3301 = \pi22 & \pi33 ;
  assign w3302 = \pi21 & \pi34 ;
  assign w3303 = \pi20 & \pi35 ;
  assign w3304 = ( w3301 & w3302 ) | ( w3301 & w3303 ) | ( w3302 & w3303 ) ;
  assign w3305 = w3301 ^ w3303 ;
  assign w3306 = w3302 ^ w3305 ;
  assign w3307 = \pi25 & \pi30 ;
  assign w3308 = \pi24 & \pi31 ;
  assign w3309 = \pi23 & \pi32 ;
  assign w3310 = ( w3307 & w3308 ) | ( w3307 & w3309 ) | ( w3308 & w3309 ) ;
  assign w3311 = w3307 ^ w3309 ;
  assign w3312 = w3308 ^ w3311 ;
  assign w3313 = w3300 ^ w3306 ;
  assign w3314 = w3312 ^ w3313 ;
  assign w3315 = ( w3119 & w3120 ) | ( w3119 & w3141 ) | ( w3120 & w3141 ) ;
  assign w3316 = w3131 ^ w3137 ;
  assign w3317 = w3180 ^ w3316 ;
  assign w3318 = ( w3169 & w3175 ) | ( w3169 & w3182 ) | ( w3175 & w3182 ) ;
  assign w3319 = ( w3191 & w3197 ) | ( w3191 & w3203 ) | ( w3197 & w3203 ) ;
  assign w3320 = w3317 ^ w3319 ;
  assign w3321 = w3318 ^ w3320 ;
  assign w3322 = w3314 ^ w3321 ;
  assign w3323 = w3315 ^ w3322 ;
  assign w3324 = w3294 ^ w3323 ;
  assign w3325 = w3272 ^ w3273 ;
  assign w3326 = w3324 ^ w3325 ;
  assign w3327 = w3225 ^ w3326 ;
  assign w3328 = w3248 ^ w3327 ;
  assign w3329 = ( w3116 & w3220 ) | ( w3116 & w3221 ) | ( w3220 & w3221 ) ;
  assign w3330 = w3224 ^ w3329 ;
  assign w3331 = w3328 ^ w3330 ;
  assign w3332 = ( w3225 & w3248 ) | ( w3225 & w3326 ) | ( w3248 & w3326 ) ;
  assign w3333 = \pi17 & \pi39 ;
  assign w3334 = \pi07 & \pi49 ;
  assign w3335 = \pi06 & \pi50 ;
  assign w3336 = ( w3333 & w3334 ) | ( w3333 & w3335 ) | ( w3334 & w3335 ) ;
  assign w3337 = w3333 ^ w3335 ;
  assign w3338 = w3334 ^ w3337 ;
  assign w3339 = \pi13 & \pi43 ;
  assign w3340 = \pi12 & \pi44 ;
  assign w3341 = \pi11 & \pi45 ;
  assign w3342 = ( w3339 & w3340 ) | ( w3339 & w3341 ) | ( w3340 & w3341 ) ;
  assign w3343 = w3339 ^ w3341 ;
  assign w3344 = w3340 ^ w3343 ;
  assign w3345 = \pi16 & \pi40 ;
  assign w3346 = \pi15 & \pi41 ;
  assign w3347 = \pi08 & \pi48 ;
  assign w3348 = ( w3345 & w3346 ) | ( w3345 & w3347 ) | ( w3346 & w3347 ) ;
  assign w3349 = w3345 ^ w3347 ;
  assign w3350 = w3346 ^ w3349 ;
  assign w3351 = w3338 ^ w3344 ;
  assign w3352 = w3350 ^ w3351 ;
  assign w3353 = \pi23 & \pi33 ;
  assign w3354 = \pi22 & \pi34 ;
  assign w3355 = \pi20 & \pi36 ;
  assign w3356 = ( w3353 & w3354 ) | ( w3353 & w3355 ) | ( w3354 & w3355 ) ;
  assign w3357 = w3353 ^ w3355 ;
  assign w3358 = w3354 ^ w3357 ;
  assign w3359 = \pi26 & \pi30 ;
  assign w3360 = \pi25 & \pi31 ;
  assign w3361 = \pi24 & \pi32 ;
  assign w3362 = ( w3359 & w3360 ) | ( w3359 & w3361 ) | ( w3360 & w3361 ) ;
  assign w3363 = w3359 ^ w3361 ;
  assign w3364 = w3360 ^ w3363 ;
  assign w3365 = \pi14 & \pi42 ;
  assign w3366 = \pi10 & \pi46 ;
  assign w3367 = \pi09 & \pi47 ;
  assign w3368 = ( w3365 & w3366 ) | ( w3365 & w3367 ) | ( w3366 & w3367 ) ;
  assign w3369 = w3365 ^ w3367 ;
  assign w3370 = w3366 ^ w3369 ;
  assign w3371 = w3358 ^ w3364 ;
  assign w3372 = w3370 ^ w3371 ;
  assign w3373 = \pi00 & \pi56 ;
  assign w3374 = ( \pi01 & \pi28 ) | ( \pi01 & ~\pi54 ) | ( \pi28 & ~\pi54 ) ;
  assign w3375 = \pi02 ^ w3374 ;
  assign w3376 = \pi54 & w3375 ;
  assign w3377 = w3373 ^ w3376 ;
  assign w3378 = \pi19 & \pi37 ;
  assign w3379 = \pi04 & \pi52 ;
  assign w3380 = \pi03 & \pi53 ;
  assign w3381 = ( w3378 & w3379 ) | ( w3378 & w3380 ) | ( w3379 & w3380 ) ;
  assign w3382 = w3378 ^ w3380 ;
  assign w3383 = w3379 ^ w3382 ;
  assign w3384 = w3288 ^ w3377 ;
  assign w3385 = w3383 ^ w3384 ;
  assign w3386 = w3352 ^ w3372 ;
  assign w3387 = w3385 ^ w3386 ;
  assign w3388 = ( w3228 & w3243 ) | ( w3228 & w3244 ) | ( w3243 & w3244 ) ;
  assign w3389 = w3232 ^ w3304 ;
  assign w3390 = w3310 ^ w3389 ;
  assign w3391 = ( w3279 & w3284 ) | ( w3279 & w3290 ) | ( w3284 & w3290 ) ;
  assign w3392 = \pi27 & \pi29 ;
  assign w3393 = w3282 ^ w3392 ;
  assign w3394 = w3277 ^ w3393 ;
  assign w3395 = \pi01 & \pi55 ;
  assign w3396 = w3394 ^ w3395 ;
  assign w3397 = w3391 ^ w3396 ;
  assign w3398 = w3390 ^ w3397 ;
  assign w3399 = w3388 ^ w3398 ;
  assign w3400 = w3387 ^ w3399 ;
  assign w3401 = ( w3226 & w3227 ) | ( w3226 & w3246 ) | ( w3227 & w3246 ) ;
  assign w3402 = w3238 ^ w3261 ;
  assign w3403 = w3298 ^ w3402 ;
  assign w3404 = ( w3234 & w3240 ) | ( w3234 & w3241 ) | ( w3240 & w3241 ) ;
  assign w3405 = ( w3249 & w3250 ) | ( w3249 & w3254 ) | ( w3250 & w3254 ) ;
  assign w3406 = w3404 ^ w3405 ;
  assign w3407 = w3403 ^ w3406 ;
  assign w3408 = ( w3131 & w3137 ) | ( w3131 & w3180 ) | ( w3137 & w3180 ) ;
  assign w3409 = ( w3195 & w3258 ) | ( w3195 & w3263 ) | ( w3258 & w3263 ) ;
  assign w3410 = ( w3300 & w3306 ) | ( w3300 & w3312 ) | ( w3306 & w3312 ) ;
  assign w3411 = w3408 ^ w3409 ;
  assign w3412 = w3410 ^ w3411 ;
  assign w3413 = ( w3292 & w3293 ) | ( w3292 & w3314 ) | ( w3293 & w3314 ) ;
  assign w3414 = w3407 ^ w3412 ;
  assign w3415 = w3413 ^ w3414 ;
  assign w3416 = w3400 ^ w3401 ;
  assign w3417 = w3415 ^ w3416 ;
  assign w3418 = ( w3265 & w3267 ) | ( w3265 & w3268 ) | ( w3267 & w3268 ) ;
  assign w3419 = \pi28 ^ w3251 ;
  assign w3420 = ( w3122 & w3173 ) | ( w3122 & w3419 ) | ( w3173 & w3419 ) ;
  assign w3421 = \pi21 & \pi35 ;
  assign w3422 = \pi18 & \pi38 ;
  assign w3423 = \pi05 & \pi51 ;
  assign w3424 = ( w3421 & w3422 ) | ( w3421 & w3423 ) | ( w3422 & w3423 ) ;
  assign w3425 = w3421 ^ w3423 ;
  assign w3426 = w3422 ^ w3425 ;
  assign w3427 = ( w3167 & w3189 ) | ( w3167 & w3201 ) | ( w3189 & w3201 ) ;
  assign w3428 = w3420 ^ w3427 ;
  assign w3429 = w3426 ^ w3428 ;
  assign w3430 = ( w3317 & w3318 ) | ( w3317 & w3319 ) | ( w3318 & w3319 ) ;
  assign w3431 = w3418 ^ w3429 ;
  assign w3432 = w3430 ^ w3431 ;
  assign w3433 = ( w3256 & w3257 ) | ( w3256 & w3270 ) | ( w3257 & w3270 ) ;
  assign w3434 = w3294 ^ w3314 ;
  assign w3435 = ( w3315 & w3321 ) | ( w3315 & w3434 ) | ( w3321 & w3434 ) ;
  assign w3436 = w3433 ^ w3435 ;
  assign w3437 = w3432 ^ w3436 ;
  assign w3438 = ( w3272 & w3273 ) | ( w3272 & w3324 ) | ( w3273 & w3324 ) ;
  assign w3439 = w3417 ^ w3438 ;
  assign w3440 = w3437 ^ w3439 ;
  assign w3441 = ( w3224 & w3328 ) | ( w3224 & w3329 ) | ( w3328 & w3329 ) ;
  assign w3442 = w3332 ^ w3441 ;
  assign w3443 = w3440 ^ w3442 ;
  assign w3444 = ( w3417 & w3437 ) | ( w3417 & w3438 ) | ( w3437 & w3438 ) ;
  assign w3445 = ( w3432 & w3433 ) | ( w3432 & w3435 ) | ( w3433 & w3435 ) ;
  assign w3446 = w3392 ^ w3395 ;
  assign w3447 = ( w3277 & w3282 ) | ( w3277 & w3446 ) | ( w3282 & w3446 ) ;
  assign w3448 = ( w3288 & w3377 ) | ( w3288 & w3383 ) | ( w3377 & w3383 ) ;
  assign w3449 = ( w3358 & w3364 ) | ( w3358 & w3370 ) | ( w3364 & w3370 ) ;
  assign w3450 = w3447 ^ w3448 ;
  assign w3451 = w3449 ^ w3450 ;
  assign w3452 = ( w3352 & w3372 ) | ( w3352 & w3385 ) | ( w3372 & w3385 ) ;
  assign w3453 = ( w3338 & w3344 ) | ( w3338 & w3350 ) | ( w3344 & w3350 ) ;
  assign w3454 = w3336 ^ w3348 ;
  assign w3455 = w3362 ^ w3454 ;
  assign w3456 = ( \pi00 & ~\pi54 ) | ( \pi00 & \pi56 ) | ( ~\pi54 & \pi56 ) ;
  assign w3457 = ( \pi02 & w3374 ) | ( \pi02 & w3456 ) | ( w3374 & w3456 ) ;
  assign w3458 = \pi54 & w3457 ;
  assign w3459 = w3356 ^ w3381 ;
  assign w3460 = w3458 ^ w3459 ;
  assign w3461 = w3453 ^ w3455 ;
  assign w3462 = w3460 ^ w3461 ;
  assign w3463 = w3451 ^ w3452 ;
  assign w3464 = w3462 ^ w3463 ;
  assign w3465 = ( w3418 & w3429 ) | ( w3418 & w3430 ) | ( w3429 & w3430 ) ;
  assign w3466 = w3342 ^ w3368 ;
  assign w3467 = w3424 ^ w3466 ;
  assign w3468 = ( w3420 & w3426 ) | ( w3420 & w3427 ) | ( w3426 & w3427 ) ;
  assign w3469 = w3467 ^ w3468 ;
  assign w3470 = \pi16 & \pi41 ;
  assign w3471 = \pi08 & \pi49 ;
  assign w3472 = \pi07 & \pi50 ;
  assign w3473 = ( w3470 & w3471 ) | ( w3470 & w3472 ) | ( w3471 & w3472 ) ;
  assign w3474 = w3470 ^ w3472 ;
  assign w3475 = w3471 ^ w3474 ;
  assign w3476 = \pi23 & \pi34 ;
  assign w3477 = \pi22 & \pi35 ;
  assign w3478 = \pi21 & \pi36 ;
  assign w3479 = ( w3476 & w3477 ) | ( w3476 & w3478 ) | ( w3477 & w3478 ) ;
  assign w3480 = w3476 ^ w3478 ;
  assign w3481 = w3477 ^ w3480 ;
  assign w3482 = \pi26 & \pi31 ;
  assign w3483 = \pi25 & \pi32 ;
  assign w3484 = \pi24 & \pi33 ;
  assign w3485 = ( w3482 & w3483 ) | ( w3482 & w3484 ) | ( w3483 & w3484 ) ;
  assign w3486 = w3482 ^ w3484 ;
  assign w3487 = w3483 ^ w3486 ;
  assign w3488 = w3475 ^ w3481 ;
  assign w3489 = w3487 ^ w3488 ;
  assign w3490 = ( w3408 & w3409 ) | ( w3408 & w3410 ) | ( w3409 & w3410 ) ;
  assign w3491 = \pi53 & \pi54 ;
  assign w3492 = \pi04 & \pi53 ;
  assign w3493 = \pi03 & \pi54 ;
  assign w3494 = \pi02 & \pi55 ;
  assign w3495 = ( w3492 & w3493 ) | ( w3492 & w3494 ) | ( w3493 & w3494 ) ;
  assign w3496 = w3492 ^ w3494 ;
  assign w3497 = w3493 ^ w3496 ;
  assign w3498 = \pi20 & \pi37 ;
  assign w3499 = \pi19 & \pi38 ;
  assign w3500 = \pi05 & \pi52 ;
  assign w3501 = ( w3498 & w3499 ) | ( w3498 & w3500 ) | ( w3499 & w3500 ) ;
  assign w3502 = w3498 ^ w3500 ;
  assign w3503 = w3499 ^ w3502 ;
  assign w3504 = \pi15 & \pi42 ;
  assign w3505 = \pi10 & \pi47 ;
  assign w3506 = \pi09 & \pi48 ;
  assign w3507 = ( w3504 & w3505 ) | ( w3504 & w3506 ) | ( w3505 & w3506 ) ;
  assign w3508 = w3504 ^ w3506 ;
  assign w3509 = w3505 ^ w3508 ;
  assign w3510 = w3497 ^ w3503 ;
  assign w3511 = w3509 ^ w3510 ;
  assign w3512 = \pi14 & \pi43 ;
  assign w3513 = \pi13 & \pi44 ;
  assign w3514 = \pi11 & \pi46 ;
  assign w3515 = ( w3512 & w3513 ) | ( w3512 & w3514 ) | ( w3513 & w3514 ) ;
  assign w3516 = w3512 ^ w3514 ;
  assign w3517 = w3513 ^ w3516 ;
  assign w3518 = \pi28 & \pi29 ;
  assign w3519 = \pi27 & \pi30 ;
  assign w3520 = \pi12 & \pi45 ;
  assign w3521 = ( w3518 & w3519 ) | ( w3518 & w3520 ) | ( w3519 & w3520 ) ;
  assign w3522 = w3518 ^ w3520 ;
  assign w3523 = w3519 ^ w3522 ;
  assign w3524 = \pi17 & \pi51 ;
  assign w3525 = \pi18 & \pi39 ;
  assign w3526 = \pi17 & \pi40 ;
  assign w3527 = \pi06 & \pi51 ;
  assign w3528 = ( w3525 & w3526 ) | ( w3525 & w3527 ) | ( w3526 & w3527 ) ;
  assign w3529 = w3525 ^ w3527 ;
  assign w3530 = w3526 ^ w3529 ;
  assign w3531 = w3517 ^ w3523 ;
  assign w3532 = w3530 ^ w3531 ;
  assign w3533 = w3490 ^ w3511 ;
  assign w3534 = w3532 ^ w3533 ;
  assign w3535 = w3489 ^ w3534 ;
  assign w3536 = w3465 ^ w3535 ;
  assign w3537 = w3469 ^ w3536 ;
  assign w3538 = w3445 ^ w3537 ;
  assign w3539 = w3464 ^ w3538 ;
  assign w3540 = ( w3400 & w3401 ) | ( w3400 & w3415 ) | ( w3401 & w3415 ) ;
  assign w3541 = ( w3387 & w3388 ) | ( w3387 & w3398 ) | ( w3388 & w3398 ) ;
  assign w3542 = ( w3407 & w3412 ) | ( w3407 & w3413 ) | ( w3412 & w3413 ) ;
  assign w3543 = ( w3403 & w3404 ) | ( w3403 & w3405 ) | ( w3404 & w3405 ) ;
  assign w3544 = ( w3390 & w3391 ) | ( w3390 & w3396 ) | ( w3391 & w3396 ) ;
  assign w3545 = \pi00 & \pi57 ;
  assign w3546 = ( \pi01 & \pi27 ) | ( \pi01 & ~\pi29 ) | ( \pi27 & ~\pi29 ) ;
  assign w3547 = ( \pi29 & ~\pi55 ) | ( \pi29 & w3546 ) | ( ~\pi55 & w3546 ) ;
  assign w3548 = \pi55 & w3547 ;
  assign w3549 = w3545 ^ w3548 ;
  assign w3550 = ( w3232 & w3304 ) | ( w3232 & w3310 ) | ( w3304 & w3310 ) ;
  assign w3551 = ( w3238 & w3261 ) | ( w3238 & w3298 ) | ( w3261 & w3298 ) ;
  assign w3552 = w3549 ^ w3550 ;
  assign w3553 = w3551 ^ w3552 ;
  assign w3554 = \pi29 ^ w3553 ;
  assign w3555 = \pi01 & \pi56 ;
  assign w3556 = w3554 ^ w3555 ;
  assign w3557 = w3543 ^ w3544 ;
  assign w3558 = w3556 ^ w3557 ;
  assign w3559 = w3541 ^ w3542 ;
  assign w3560 = w3558 ^ w3559 ;
  assign w3561 = w3539 ^ w3540 ;
  assign w3562 = w3560 ^ w3561 ;
  assign w3563 = ( w3332 & w3440 ) | ( w3332 & w3441 ) | ( w3440 & w3441 ) ;
  assign w3564 = w3444 ^ w3563 ;
  assign w3565 = w3562 ^ w3564 ;
  assign w3566 = ( w3444 & w3562 ) | ( w3444 & w3563 ) | ( w3562 & w3563 ) ;
  assign w3567 = ( w3539 & w3540 ) | ( w3539 & w3560 ) | ( w3540 & w3560 ) ;
  assign w3568 = ( w3445 & w3464 ) | ( w3445 & w3537 ) | ( w3464 & w3537 ) ;
  assign w3569 = ( w3451 & w3452 ) | ( w3451 & w3462 ) | ( w3452 & w3462 ) ;
  assign w3570 = ( w3467 & w3468 ) | ( w3467 & w3489 ) | ( w3468 & w3489 ) ;
  assign w3571 = ( w3342 & w3368 ) | ( w3342 & w3424 ) | ( w3368 & w3424 ) ;
  assign w3572 = ( w3356 & w3381 ) | ( w3356 & w3458 ) | ( w3381 & w3458 ) ;
  assign w3573 = ( w3336 & w3348 ) | ( w3336 & w3362 ) | ( w3348 & w3362 ) ;
  assign w3574 = w3571 ^ w3572 ;
  assign w3575 = w3573 ^ w3574 ;
  assign w3576 = ( w3453 & w3455 ) | ( w3453 & w3460 ) | ( w3455 & w3460 ) ;
  assign w3577 = w3570 ^ w3575 ;
  assign w3578 = w3576 ^ w3577 ;
  assign w3579 = w3469 ^ w3489 ;
  assign w3580 = ( w3465 & w3534 ) | ( w3465 & w3579 ) | ( w3534 & w3579 ) ;
  assign w3581 = w3578 ^ w3580 ;
  assign w3582 = w3569 ^ w3581 ;
  assign w3583 = ( w3541 & w3542 ) | ( w3541 & w3558 ) | ( w3542 & w3558 ) ;
  assign w3584 = ( w3490 & w3511 ) | ( w3490 & w3532 ) | ( w3511 & w3532 ) ;
  assign w3585 = ( w3517 & w3523 ) | ( w3517 & w3530 ) | ( w3523 & w3530 ) ;
  assign w3586 = ( w3497 & w3503 ) | ( w3497 & w3509 ) | ( w3503 & w3509 ) ;
  assign w3587 = ( ~\pi01 & \pi29 ) | ( ~\pi01 & \pi56 ) | ( \pi29 & \pi56 ) ;
  assign w3588 = \pi57 ^ w3587 ;
  assign w3589 = \pi01 & w3588 ;
  assign w3590 = w1454 ^ w3521 ;
  assign w3591 = w3589 ^ w3590 ;
  assign w3592 = w3585 ^ w3586 ;
  assign w3593 = w3591 ^ w3592 ;
  assign w3594 = ( w3475 & w3481 ) | ( w3475 & w3487 ) | ( w3481 & w3487 ) ;
  assign w3595 = w3479 ^ w3485 ;
  assign w3596 = w3507 ^ w3595 ;
  assign w3597 = w3495 ^ w3501 ;
  assign w3598 = w3515 ^ w3597 ;
  assign w3599 = w3594 ^ w3596 ;
  assign w3600 = w3598 ^ w3599 ;
  assign w3601 = w3584 ^ w3593 ;
  assign w3602 = w3600 ^ w3601 ;
  assign w3603 = \pi04 & \pi54 ;
  assign w3604 = \pi02 & \pi56 ;
  assign w3605 = \pi00 & \pi58 ;
  assign w3606 = ( w3603 & w3604 ) | ( w3603 & w3605 ) | ( w3604 & w3605 ) ;
  assign w3607 = w3603 ^ w3605 ;
  assign w3608 = w3604 ^ w3607 ;
  assign w3609 = \pi21 & \pi37 ;
  assign w3610 = \pi20 & \pi38 ;
  assign w3611 = \pi05 & \pi53 ;
  assign w3612 = ( w3609 & w3610 ) | ( w3609 & w3611 ) | ( w3610 & w3611 ) ;
  assign w3613 = w3609 ^ w3611 ;
  assign w3614 = w3610 ^ w3613 ;
  assign w3615 = \pi42 & \pi49 ;
  assign w3616 = \pi17 & \pi41 ;
  assign w3617 = \pi16 & \pi42 ;
  assign w3618 = \pi09 & \pi49 ;
  assign w3619 = ( w3616 & w3617 ) | ( w3616 & w3618 ) | ( w3617 & w3618 ) ;
  assign w3620 = w3616 ^ w3618 ;
  assign w3621 = w3617 ^ w3620 ;
  assign w3622 = w3608 ^ w3614 ;
  assign w3623 = w3621 ^ w3622 ;
  assign w3624 = \pi18 & \pi40 ;
  assign w3625 = \pi08 & \pi50 ;
  assign w3626 = \pi07 & \pi51 ;
  assign w3627 = ( w3624 & w3625 ) | ( w3624 & w3626 ) | ( w3625 & w3626 ) ;
  assign w3628 = w3624 ^ w3626 ;
  assign w3629 = w3625 ^ w3628 ;
  assign w3630 = \pi24 & \pi34 ;
  assign w3631 = \pi23 & \pi35 ;
  assign w3632 = \pi22 & \pi36 ;
  assign w3633 = ( w3630 & w3631 ) | ( w3630 & w3632 ) | ( w3631 & w3632 ) ;
  assign w3634 = w3630 ^ w3632 ;
  assign w3635 = w3631 ^ w3634 ;
  assign w3636 = \pi27 & \pi31 ;
  assign w3637 = \pi26 & \pi32 ;
  assign w3638 = \pi25 & \pi33 ;
  assign w3639 = ( w3636 & w3637 ) | ( w3636 & w3638 ) | ( w3637 & w3638 ) ;
  assign w3640 = w3636 ^ w3638 ;
  assign w3641 = w3637 ^ w3640 ;
  assign w3642 = w3629 ^ w3635 ;
  assign w3643 = w3641 ^ w3642 ;
  assign w3644 = ( w3447 & w3448 ) | ( w3447 & w3449 ) | ( w3448 & w3449 ) ;
  assign w3645 = w3623 ^ w3644 ;
  assign w3646 = w3643 ^ w3645 ;
  assign w3647 = ( w3543 & w3544 ) | ( w3543 & w3556 ) | ( w3544 & w3556 ) ;
  assign w3648 = \pi27 & \pi55 ;
  assign w3649 = ( ~\pi56 & w3545 ) | ( ~\pi56 & w3648 ) | ( w3545 & w3648 ) ;
  assign w3650 = \pi29 & w3649 ;
  assign w3651 = ( \pi01 & \pi29 ) | ( \pi01 & ~\pi56 ) | ( \pi29 & ~\pi56 ) ;
  assign w3652 = ( \pi01 & \pi29 ) | ( \pi01 & w3545 ) | ( \pi29 & w3545 ) ;
  assign w3653 = ( w3650 & ~w3651 ) | ( w3650 & w3652 ) | ( ~w3651 & w3652 ) ;
  assign w3654 = w3473 ^ w3653 ;
  assign w3655 = w3528 ^ w3654 ;
  assign w3656 = \pi29 ^ w3549 ;
  assign w3657 = w3555 ^ w3656 ;
  assign w3658 = ( w3550 & w3551 ) | ( w3550 & w3657 ) | ( w3551 & w3657 ) ;
  assign w3659 = \pi15 & \pi43 ;
  assign w3660 = \pi11 & \pi47 ;
  assign w3661 = \pi10 & \pi48 ;
  assign w3662 = ( w3659 & w3660 ) | ( w3659 & w3661 ) | ( w3660 & w3661 ) ;
  assign w3663 = w3659 ^ w3661 ;
  assign w3664 = w3660 ^ w3663 ;
  assign w3665 = \pi14 & \pi44 ;
  assign w3666 = \pi13 & \pi45 ;
  assign w3667 = \pi12 & \pi46 ;
  assign w3668 = ( w3665 & w3666 ) | ( w3665 & w3667 ) | ( w3666 & w3667 ) ;
  assign w3669 = w3665 ^ w3667 ;
  assign w3670 = w3666 ^ w3669 ;
  assign w3671 = \pi19 & \pi39 ;
  assign w3672 = \pi06 & \pi52 ;
  assign w3673 = \pi03 & \pi55 ;
  assign w3674 = ( w3671 & w3672 ) | ( w3671 & w3673 ) | ( w3672 & w3673 ) ;
  assign w3675 = w3671 ^ w3673 ;
  assign w3676 = w3672 ^ w3675 ;
  assign w3677 = w3664 ^ w3670 ;
  assign w3678 = w3676 ^ w3677 ;
  assign w3679 = w3655 ^ w3658 ;
  assign w3680 = w3678 ^ w3679 ;
  assign w3681 = w3646 ^ w3647 ;
  assign w3682 = w3680 ^ w3681 ;
  assign w3683 = w3583 ^ w3682 ;
  assign w3684 = w3602 ^ w3683 ;
  assign w3685 = w3568 ^ w3684 ;
  assign w3686 = w3582 ^ w3685 ;
  assign w3687 = w3567 & w3686 ;
  assign w3688 = w3567 | w3686 ;
  assign w3689 = ~w3687 & w3688 ;
  assign w3690 = w3566 ^ w3689 ;
  assign w3691 = ( w3583 & w3602 ) | ( w3583 & w3682 ) | ( w3602 & w3682 ) ;
  assign w3692 = ( w3646 & w3647 ) | ( w3646 & w3680 ) | ( w3647 & w3680 ) ;
  assign w3693 = ( w3584 & w3593 ) | ( w3584 & w3600 ) | ( w3593 & w3600 ) ;
  assign w3694 = ( w3655 & w3658 ) | ( w3655 & w3678 ) | ( w3658 & w3678 ) ;
  assign w3695 = ( w3473 & w3528 ) | ( w3473 & w3653 ) | ( w3528 & w3653 ) ;
  assign w3696 = ( w3495 & w3501 ) | ( w3495 & w3515 ) | ( w3501 & w3515 ) ;
  assign w3697 = ( w3479 & w3485 ) | ( w3479 & w3507 ) | ( w3485 & w3507 ) ;
  assign w3698 = w3695 ^ w3696 ;
  assign w3699 = w3697 ^ w3698 ;
  assign w3700 = ( w3594 & w3596 ) | ( w3594 & w3598 ) | ( w3596 & w3598 ) ;
  assign w3701 = w3694 ^ w3699 ;
  assign w3702 = w3700 ^ w3701 ;
  assign w3703 = w3692 ^ w3693 ;
  assign w3704 = w3702 ^ w3703 ;
  assign w3705 = ( w3570 & w3575 ) | ( w3570 & w3576 ) | ( w3575 & w3576 ) ;
  assign w3706 = ( w3585 & w3586 ) | ( w3585 & w3591 ) | ( w3586 & w3591 ) ;
  assign w3707 = \pi14 & \pi45 ;
  assign w3708 = \pi12 & \pi47 ;
  assign w3709 = \pi11 & \pi48 ;
  assign w3710 = ( w3707 & w3708 ) | ( w3707 & w3709 ) | ( w3708 & w3709 ) ;
  assign w3711 = w3707 ^ w3709 ;
  assign w3712 = w3708 ^ w3711 ;
  assign w3713 = \pi28 & \pi31 ;
  assign w3714 = \pi13 & \pi46 ;
  assign w3715 = ( w1221 & w3713 ) | ( w1221 & w3714 ) | ( w3713 & w3714 ) ;
  assign w3716 = w1221 ^ w3714 ;
  assign w3717 = w3713 ^ w3716 ;
  assign w3718 = \pi17 & \pi42 ;
  assign w3719 = \pi16 & \pi43 ;
  assign w3720 = \pi08 & \pi51 ;
  assign w3721 = ( w3718 & w3719 ) | ( w3718 & w3720 ) | ( w3719 & w3720 ) ;
  assign w3722 = w3718 ^ w3720 ;
  assign w3723 = w3719 ^ w3722 ;
  assign w3724 = w3712 ^ w3717 ;
  assign w3725 = w3723 ^ w3724 ;
  assign w3726 = ( \pi01 & ~\pi57 ) | ( \pi01 & w1454 ) | ( ~\pi57 & w1454 ) ;
  assign w3727 = ( \pi03 & \pi56 ) | ( \pi03 & ~\pi57 ) | ( \pi56 & ~\pi57 ) ;
  assign w3728 = ( \pi02 & w3726 ) | ( \pi02 & w3727 ) | ( w3726 & w3727 ) ;
  assign w3729 = \pi57 & w3728 ;
  assign w3730 = \pi03 & \pi56 ;
  assign w3731 = \pi02 ^ w3726 ;
  assign w3732 = \pi57 & w3731 ;
  assign w3733 = w3730 ^ w3732 ;
  assign w3734 = \pi19 & \pi40 ;
  assign w3735 = \pi05 & \pi54 ;
  assign w3736 = \pi04 & \pi55 ;
  assign w3737 = ( w3734 & w3735 ) | ( w3734 & w3736 ) | ( w3735 & w3736 ) ;
  assign w3738 = w3734 ^ w3736 ;
  assign w3739 = w3735 ^ w3738 ;
  assign w3740 = w3639 ^ w3733 ;
  assign w3741 = w3739 ^ w3740 ;
  assign w3742 = w3706 ^ w3725 ;
  assign w3743 = w3741 ^ w3742 ;
  assign w3744 = \pi18 & \pi41 ;
  assign w3745 = \pi07 & \pi52 ;
  assign w3746 = \pi06 & \pi53 ;
  assign w3747 = ( w3744 & w3745 ) | ( w3744 & w3746 ) | ( w3745 & w3746 ) ;
  assign w3748 = w3744 ^ w3746 ;
  assign w3749 = w3745 ^ w3748 ;
  assign w3750 = \pi15 & \pi44 ;
  assign w3751 = \pi10 & \pi49 ;
  assign w3752 = \pi09 & \pi50 ;
  assign w3753 = ( w3750 & w3751 ) | ( w3750 & w3752 ) | ( w3751 & w3752 ) ;
  assign w3754 = w3750 ^ w3752 ;
  assign w3755 = w3751 ^ w3754 ;
  assign w3756 = \pi56 & w1018 ;
  assign w3757 = \pi01 & \pi57 ;
  assign w3758 = w1454 ^ w3757 ;
  assign w3759 = ( w3521 & w3756 ) | ( w3521 & w3758 ) | ( w3756 & w3758 ) ;
  assign w3760 = w3749 ^ w3759 ;
  assign w3761 = w3755 ^ w3760 ;
  assign w3762 = ( w3571 & w3572 ) | ( w3571 & w3573 ) | ( w3572 & w3573 ) ;
  assign w3763 = w3761 ^ w3762 ;
  assign w3764 = \pi22 & \pi37 ;
  assign w3765 = \pi21 & \pi38 ;
  assign w3766 = \pi20 & \pi39 ;
  assign w3767 = ( w3764 & w3765 ) | ( w3764 & w3766 ) | ( w3765 & w3766 ) ;
  assign w3768 = w3764 ^ w3766 ;
  assign w3769 = w3765 ^ w3768 ;
  assign w3770 = \pi25 & \pi34 ;
  assign w3771 = \pi24 & \pi35 ;
  assign w3772 = \pi23 & \pi36 ;
  assign w3773 = ( w3770 & w3771 ) | ( w3770 & w3772 ) | ( w3771 & w3772 ) ;
  assign w3774 = w3770 ^ w3772 ;
  assign w3775 = w3771 ^ w3774 ;
  assign w3776 = \pi27 & \pi32 ;
  assign w3777 = \pi26 & \pi33 ;
  assign w3778 = \pi00 & \pi59 ;
  assign w3779 = ( w3776 & w3777 ) | ( w3776 & w3778 ) | ( w3777 & w3778 ) ;
  assign w3780 = w3776 ^ w3778 ;
  assign w3781 = w3777 ^ w3780 ;
  assign w3782 = w3769 ^ w3775 ;
  assign w3783 = w3781 ^ w3782 ;
  assign w3784 = w3763 ^ w3783 ;
  assign w3785 = w3705 ^ w3784 ;
  assign w3786 = w3743 ^ w3785 ;
  assign w3787 = ( w3569 & w3578 ) | ( w3569 & w3580 ) | ( w3578 & w3580 ) ;
  assign w3788 = ( w3664 & w3670 ) | ( w3664 & w3676 ) | ( w3670 & w3676 ) ;
  assign w3789 = ( w3629 & w3635 ) | ( w3629 & w3641 ) | ( w3635 & w3641 ) ;
  assign w3790 = ( w3608 & w3614 ) | ( w3608 & w3621 ) | ( w3614 & w3621 ) ;
  assign w3791 = w3788 ^ w3789 ;
  assign w3792 = w3790 ^ w3791 ;
  assign w3793 = ( w3623 & w3643 ) | ( w3623 & w3644 ) | ( w3643 & w3644 ) ;
  assign w3794 = w3606 ^ w3619 ;
  assign w3795 = w3674 ^ w3794 ;
  assign w3796 = w3612 ^ w3627 ;
  assign w3797 = w3633 ^ w3796 ;
  assign w3798 = \pi01 & \pi58 ;
  assign w3799 = \pi30 ^ w3668 ;
  assign w3800 = w3662 ^ w3799 ;
  assign w3801 = w3798 ^ w3800 ;
  assign w3802 = w3795 ^ w3797 ;
  assign w3803 = w3801 ^ w3802 ;
  assign w3804 = w3792 ^ w3793 ;
  assign w3805 = w3803 ^ w3804 ;
  assign w3806 = w3786 ^ w3787 ;
  assign w3807 = w3805 ^ w3806 ;
  assign w3808 = w3691 ^ w3704 ;
  assign w3809 = w3807 ^ w3808 ;
  assign w3810 = ( w3568 & w3582 ) | ( w3568 & w3684 ) | ( w3582 & w3684 ) ;
  assign w3811 = ( w3566 & w3687 ) | ( w3566 & w3688 ) | ( w3687 & w3688 ) ;
  assign w3812 = w3687 | w3811 ;
  assign w3813 = w3809 ^ w3812 ;
  assign w3814 = w3810 ^ w3813 ;
  assign w3815 = ( w3691 & w3704 ) | ( w3691 & w3807 ) | ( w3704 & w3807 ) ;
  assign w3816 = ( w3786 & w3787 ) | ( w3786 & w3805 ) | ( w3787 & w3805 ) ;
  assign w3817 = ( w3705 & w3743 ) | ( w3705 & w3784 ) | ( w3743 & w3784 ) ;
  assign w3818 = ( w3792 & w3793 ) | ( w3792 & w3803 ) | ( w3793 & w3803 ) ;
  assign w3819 = ( w3612 & w3627 ) | ( w3612 & w3633 ) | ( w3627 & w3633 ) ;
  assign w3820 = ( w3606 & w3619 ) | ( w3606 & w3674 ) | ( w3619 & w3674 ) ;
  assign w3821 = ( w3639 & w3733 ) | ( w3639 & w3739 ) | ( w3733 & w3739 ) ;
  assign w3822 = w3819 ^ w3821 ;
  assign w3823 = w3820 ^ w3822 ;
  assign w3824 = ( w3788 & w3789 ) | ( w3788 & w3790 ) | ( w3789 & w3790 ) ;
  assign w3825 = ( w3761 & w3762 ) | ( w3761 & w3783 ) | ( w3762 & w3783 ) ;
  assign w3826 = w3823 ^ w3825 ;
  assign w3827 = w3824 ^ w3826 ;
  assign w3828 = w3817 ^ w3818 ;
  assign w3829 = w3827 ^ w3828 ;
  assign w3830 = ( w3694 & w3699 ) | ( w3694 & w3700 ) | ( w3699 & w3700 ) ;
  assign w3831 = \pi04 & \pi56 ;
  assign w3832 = \pi03 & \pi57 ;
  assign w3833 = \pi02 & \pi58 ;
  assign w3834 = ( w3831 & w3832 ) | ( w3831 & w3833 ) | ( w3832 & w3833 ) ;
  assign w3835 = w3831 ^ w3833 ;
  assign w3836 = w3832 ^ w3835 ;
  assign w3837 = \pi22 & \pi38 ;
  assign w3838 = \pi21 & \pi39 ;
  assign w3839 = \pi20 & \pi40 ;
  assign w3840 = ( w3837 & w3838 ) | ( w3837 & w3839 ) | ( w3838 & w3839 ) ;
  assign w3841 = w3837 ^ w3839 ;
  assign w3842 = w3838 ^ w3841 ;
  assign w3843 = \pi26 & \pi34 ;
  assign w3844 = \pi25 & \pi35 ;
  assign w3845 = \pi24 & \pi36 ;
  assign w3846 = ( w3843 & w3844 ) | ( w3843 & w3845 ) | ( w3844 & w3845 ) ;
  assign w3847 = w3843 ^ w3845 ;
  assign w3848 = w3844 ^ w3847 ;
  assign w3849 = w3836 ^ w3842 ;
  assign w3850 = w3848 ^ w3849 ;
  assign w3851 = ( w3695 & w3696 ) | ( w3695 & w3697 ) | ( w3696 & w3697 ) ;
  assign w3852 = \pi17 & \pi43 ;
  assign w3853 = \pi16 & \pi44 ;
  assign w3854 = \pi09 & \pi51 ;
  assign w3855 = ( w3852 & w3853 ) | ( w3852 & w3854 ) | ( w3853 & w3854 ) ;
  assign w3856 = w3852 ^ w3854 ;
  assign w3857 = w3853 ^ w3856 ;
  assign w3858 = \pi15 & \pi45 ;
  assign w3859 = \pi11 & \pi49 ;
  assign w3860 = \pi10 & \pi50 ;
  assign w3861 = ( w3858 & w3859 ) | ( w3858 & w3860 ) | ( w3859 & w3860 ) ;
  assign w3862 = w3858 ^ w3860 ;
  assign w3863 = w3859 ^ w3862 ;
  assign w3864 = w3710 ^ w3857 ;
  assign w3865 = w3863 ^ w3864 ;
  assign w3866 = w3850 ^ w3851 ;
  assign w3867 = w3865 ^ w3866 ;
  assign w3868 = ( w3795 & w3797 ) | ( w3795 & w3801 ) | ( w3797 & w3801 ) ;
  assign w3869 = \pi00 & \pi60 ;
  assign w3870 = ( \pi01 & \pi30 ) | ( \pi01 & ~\pi58 ) | ( \pi30 & ~\pi58 ) ;
  assign w3871 = \pi58 & w3870 ;
  assign w3872 = w3869 ^ w3871 ;
  assign w3873 = \pi01 & \pi59 ;
  assign w3874 = \pi29 & \pi31 ;
  assign w3875 = w3873 ^ w3874 ;
  assign w3876 = \pi28 & \pi32 ;
  assign w3877 = \pi27 & \pi33 ;
  assign w3878 = \pi23 & \pi37 ;
  assign w3879 = ( w3876 & w3877 ) | ( w3876 & w3878 ) | ( w3877 & w3878 ) ;
  assign w3880 = w3876 ^ w3878 ;
  assign w3881 = w3877 ^ w3880 ;
  assign w3882 = \pi30 ^ w3798 ;
  assign w3883 = ( w3662 & w3668 ) | ( w3662 & w3882 ) | ( w3668 & w3882 ) ;
  assign w3884 = w3875 ^ w3881 ;
  assign w3885 = w3883 ^ w3884 ;
  assign w3886 = w3872 ^ w3885 ;
  assign w3887 = \pi18 & \pi42 ;
  assign w3888 = \pi08 & \pi52 ;
  assign w3889 = \pi07 & \pi53 ;
  assign w3890 = ( w3887 & w3888 ) | ( w3887 & w3889 ) | ( w3888 & w3889 ) ;
  assign w3891 = w3887 ^ w3889 ;
  assign w3892 = w3888 ^ w3891 ;
  assign w3893 = \pi14 & \pi46 ;
  assign w3894 = \pi13 & \pi47 ;
  assign w3895 = \pi12 & \pi48 ;
  assign w3896 = ( w3893 & w3894 ) | ( w3893 & w3895 ) | ( w3894 & w3895 ) ;
  assign w3897 = w3893 ^ w3895 ;
  assign w3898 = w3894 ^ w3897 ;
  assign w3899 = \pi19 & \pi41 ;
  assign w3900 = \pi06 & \pi54 ;
  assign w3901 = \pi05 & \pi55 ;
  assign w3902 = ( w3899 & w3900 ) | ( w3899 & w3901 ) | ( w3900 & w3901 ) ;
  assign w3903 = w3899 ^ w3901 ;
  assign w3904 = w3900 ^ w3903 ;
  assign w3905 = w3892 ^ w3898 ;
  assign w3906 = w3904 ^ w3905 ;
  assign w3907 = w3868 ^ w3886 ;
  assign w3908 = w3906 ^ w3907 ;
  assign w3909 = w3830 ^ w3867 ;
  assign w3910 = w3908 ^ w3909 ;
  assign w3911 = ( w3692 & w3693 ) | ( w3692 & w3702 ) | ( w3693 & w3702 ) ;
  assign w3912 = w3715 ^ w3721 ;
  assign w3913 = w3747 ^ w3912 ;
  assign w3914 = ( w3769 & w3775 ) | ( w3769 & w3781 ) | ( w3775 & w3781 ) ;
  assign w3915 = ( w3712 & w3717 ) | ( w3712 & w3723 ) | ( w3717 & w3723 ) ;
  assign w3916 = w3913 ^ w3915 ;
  assign w3917 = w3914 ^ w3916 ;
  assign w3918 = ( w3706 & w3725 ) | ( w3706 & w3741 ) | ( w3725 & w3741 ) ;
  assign w3919 = ( w3749 & w3755 ) | ( w3749 & w3759 ) | ( w3755 & w3759 ) ;
  assign w3920 = w3737 ^ w3767 ;
  assign w3921 = w3773 ^ w3920 ;
  assign w3922 = w3729 ^ w3753 ;
  assign w3923 = w3779 ^ w3922 ;
  assign w3924 = w3919 ^ w3923 ;
  assign w3925 = w3921 ^ w3924 ;
  assign w3926 = w3917 ^ w3918 ;
  assign w3927 = w3925 ^ w3926 ;
  assign w3928 = w3910 ^ w3911 ;
  assign w3929 = w3927 ^ w3928 ;
  assign w3930 = w3816 ^ w3929 ;
  assign w3931 = w3829 ^ w3930 ;
  assign w3932 = ( w3809 & w3810 ) | ( w3809 & w3812 ) | ( w3810 & w3812 ) ;
  assign w3933 = w3931 ^ w3932 ;
  assign w3934 = w3815 ^ w3933 ;
  assign w3935 = ( w3816 & w3829 ) | ( w3816 & w3929 ) | ( w3829 & w3929 ) ;
  assign w3936 = ( w3910 & w3911 ) | ( w3910 & w3927 ) | ( w3911 & w3927 ) ;
  assign w3937 = ( w3830 & w3867 ) | ( w3830 & w3908 ) | ( w3867 & w3908 ) ;
  assign w3938 = ( w3913 & w3914 ) | ( w3913 & w3915 ) | ( w3914 & w3915 ) ;
  assign w3939 = \pi19 & \pi42 ;
  assign w3940 = \pi08 & \pi53 ;
  assign w3941 = \pi07 & \pi54 ;
  assign w3942 = ( w3939 & w3940 ) | ( w3939 & w3941 ) | ( w3940 & w3941 ) ;
  assign w3943 = w3939 ^ w3941 ;
  assign w3944 = w3940 ^ w3943 ;
  assign w3945 = \pi44 & \pi52 ;
  assign w3946 = \pi18 & \pi43 ;
  assign w3947 = \pi17 & \pi44 ;
  assign w3948 = \pi09 & \pi52 ;
  assign w3949 = ( w3946 & w3947 ) | ( w3946 & w3948 ) | ( w3947 & w3948 ) ;
  assign w3950 = w3946 ^ w3948 ;
  assign w3951 = w3947 ^ w3950 ;
  assign w3952 = \pi28 & \pi33 ;
  assign w3953 = \pi27 & \pi34 ;
  assign w3954 = \pi26 & \pi35 ;
  assign w3955 = ( w3952 & w3953 ) | ( w3952 & w3954 ) | ( w3953 & w3954 ) ;
  assign w3956 = w3952 ^ w3954 ;
  assign w3957 = w3953 ^ w3956 ;
  assign w3958 = w3944 ^ w3951 ;
  assign w3959 = w3957 ^ w3958 ;
  assign w3960 = ( w3919 & w3921 ) | ( w3919 & w3923 ) | ( w3921 & w3923 ) ;
  assign w3961 = w3938 ^ w3960 ;
  assign w3962 = w3959 ^ w3961 ;
  assign w3963 = ( w3850 & w3851 ) | ( w3850 & w3865 ) | ( w3851 & w3865 ) ;
  assign w3964 = ( w3729 & w3753 ) | ( w3729 & w3779 ) | ( w3753 & w3779 ) ;
  assign w3965 = ( w3715 & w3721 ) | ( w3715 & w3747 ) | ( w3721 & w3747 ) ;
  assign w3966 = \pi23 & \pi38 ;
  assign w3967 = \pi04 & \pi57 ;
  assign w3968 = \pi03 & \pi58 ;
  assign w3969 = ( w3966 & w3967 ) | ( w3966 & w3968 ) | ( w3967 & w3968 ) ;
  assign w3970 = w3966 ^ w3968 ;
  assign w3971 = w3967 ^ w3970 ;
  assign w3972 = w3964 ^ w3965 ;
  assign w3973 = w3971 ^ w3972 ;
  assign w3974 = ( w3710 & w3857 ) | ( w3710 & w3863 ) | ( w3857 & w3863 ) ;
  assign w3975 = ( w3737 & w3767 ) | ( w3737 & w3773 ) | ( w3767 & w3773 ) ;
  assign w3976 = ( \pi01 & ~\pi31 ) | ( \pi01 & \pi60 ) | ( ~\pi31 & \pi60 ) ;
  assign w3977 = \pi31 & w3976 ;
  assign w3978 = ~\pi01 & \pi29 ;
  assign w3979 = ( ~\pi29 & \pi59 ) | ( ~\pi29 & w3978 ) | ( \pi59 & w3978 ) ;
  assign w3980 = ( \pi31 & ~\pi59 ) | ( \pi31 & w3979 ) | ( ~\pi59 & w3979 ) ;
  assign w3981 = w3896 ^ w3980 ;
  assign w3982 = \pi01 & \pi60 ;
  assign w3983 = w3981 ^ w3982 ;
  assign w3984 = w3974 ^ w3975 ;
  assign w3985 = w3983 ^ w3984 ;
  assign w3986 = w3963 ^ w3973 ;
  assign w3987 = w3985 ^ w3986 ;
  assign w3988 = w3937 ^ w3987 ;
  assign w3989 = w3962 ^ w3988 ;
  assign w3990 = ( w3868 & w3886 ) | ( w3868 & w3906 ) | ( w3886 & w3906 ) ;
  assign w3991 = ( \pi01 & ~\pi30 ) | ( \pi01 & \pi58 ) | ( ~\pi30 & \pi58 ) ;
  assign w3992 = \pi30 & w3991 ;
  assign w3993 = ( w3869 & w3875 ) | ( w3869 & w3992 ) | ( w3875 & w3992 ) ;
  assign w3994 = w3855 ^ w3993 ;
  assign w3995 = w3890 ^ w3994 ;
  assign w3996 = ( w3892 & w3898 ) | ( w3892 & w3904 ) | ( w3898 & w3904 ) ;
  assign w3997 = w3872 ^ w3875 ;
  assign w3998 = ( w3881 & w3883 ) | ( w3881 & w3997 ) | ( w3883 & w3997 ) ;
  assign w3999 = w3995 ^ w3998 ;
  assign w4000 = w3996 ^ w3999 ;
  assign w4001 = ( w3836 & w3842 ) | ( w3836 & w3848 ) | ( w3842 & w3848 ) ;
  assign w4002 = w3840 ^ w3846 ;
  assign w4003 = w3879 ^ w4002 ;
  assign w4004 = w3834 ^ w3861 ;
  assign w4005 = w3902 ^ w4004 ;
  assign w4006 = w4001 ^ w4003 ;
  assign w4007 = w4005 ^ w4006 ;
  assign w4008 = ( w3990 & w4000 ) | ( w3990 & w4007 ) | ( w4000 & w4007 ) ;
  assign w4009 = w3990 ^ w4000 ;
  assign w4010 = w4007 ^ w4009 ;
  assign w4011 = ( w3817 & w3818 ) | ( w3817 & w3827 ) | ( w3818 & w3827 ) ;
  assign w4012 = ( w3917 & w3918 ) | ( w3917 & w3925 ) | ( w3918 & w3925 ) ;
  assign w4013 = ( w3823 & w3824 ) | ( w3823 & w3825 ) | ( w3824 & w3825 ) ;
  assign w4014 = \pi16 & \pi45 ;
  assign w4015 = \pi15 & \pi46 ;
  assign w4016 = \pi10 & \pi51 ;
  assign w4017 = ( w4014 & w4015 ) | ( w4014 & w4016 ) | ( w4015 & w4016 ) ;
  assign w4018 = w4014 ^ w4016 ;
  assign w4019 = w4015 ^ w4018 ;
  assign w4020 = \pi14 & \pi50 ;
  assign w4021 = \pi14 & \pi47 ;
  assign w4022 = \pi12 & \pi49 ;
  assign w4023 = \pi11 & \pi50 ;
  assign w4024 = ( w4021 & w4022 ) | ( w4021 & w4023 ) | ( w4022 & w4023 ) ;
  assign w4025 = w4021 ^ w4023 ;
  assign w4026 = w4022 ^ w4025 ;
  assign w4027 = \pi29 & \pi32 ;
  assign w4028 = \pi13 & \pi48 ;
  assign w4029 = ( w1335 & w4027 ) | ( w1335 & w4028 ) | ( w4027 & w4028 ) ;
  assign w4030 = w1335 ^ w4028 ;
  assign w4031 = w4027 ^ w4030 ;
  assign w4032 = w4019 ^ w4026 ;
  assign w4033 = w4031 ^ w4032 ;
  assign w4034 = ( w3819 & w3820 ) | ( w3819 & w3821 ) | ( w3820 & w3821 ) ;
  assign w4035 = \pi05 & \pi56 ;
  assign w4036 = \pi02 & \pi59 ;
  assign w4037 = \pi00 & \pi61 ;
  assign w4038 = ( w4035 & w4036 ) | ( w4035 & w4037 ) | ( w4036 & w4037 ) ;
  assign w4039 = w4035 ^ w4037 ;
  assign w4040 = w4036 ^ w4039 ;
  assign w4041 = \pi21 & \pi40 ;
  assign w4042 = \pi06 & \pi55 ;
  assign w4043 = ( w2165 & w4041 ) | ( w2165 & w4042 ) | ( w4041 & w4042 ) ;
  assign w4044 = w4041 ^ w4042 ;
  assign w4045 = w2165 ^ w4044 ;
  assign w4046 = \pi25 & \pi36 ;
  assign w4047 = \pi24 & \pi37 ;
  assign w4048 = \pi22 & \pi39 ;
  assign w4049 = ( w4046 & w4047 ) | ( w4046 & w4048 ) | ( w4047 & w4048 ) ;
  assign w4050 = w4046 ^ w4048 ;
  assign w4051 = w4047 ^ w4050 ;
  assign w4052 = w4040 ^ w4045 ;
  assign w4053 = w4051 ^ w4052 ;
  assign w4054 = w4033 ^ w4034 ;
  assign w4055 = w4053 ^ w4054 ;
  assign w4056 = w4012 ^ w4013 ;
  assign w4057 = w4055 ^ w4056 ;
  assign w4058 = w4011 ^ w4057 ;
  assign w4059 = w4010 ^ w4058 ;
  assign w4060 = w3936 ^ w4059 ;
  assign w4061 = w3989 ^ w4060 ;
  assign w4062 = ( w3815 & w3931 ) | ( w3815 & w3932 ) | ( w3931 & w3932 ) ;
  assign w4063 = w3935 ^ w4062 ;
  assign w4064 = w4061 ^ w4063 ;
  assign w4065 = ( w3935 & w4061 ) | ( w3935 & w4062 ) | ( w4061 & w4062 ) ;
  assign w4066 = ( w3936 & w3989 ) | ( w3936 & w4059 ) | ( w3989 & w4059 ) ;
  assign w4067 = ( w3937 & w3962 ) | ( w3937 & w3987 ) | ( w3962 & w3987 ) ;
  assign w4068 = \pi58 & \pi59 ;
  assign w4069 = \pi05 & \pi57 ;
  assign w4070 = \pi04 & \pi58 ;
  assign w4071 = \pi03 & \pi59 ;
  assign w4072 = ( w4069 & w4070 ) | ( w4069 & w4071 ) | ( w4070 & w4071 ) ;
  assign w4073 = w4069 ^ w4071 ;
  assign w4074 = w4070 ^ w4073 ;
  assign w4075 = w3949 ^ w4017 ;
  assign w4076 = w4074 ^ w4075 ;
  assign w4077 = ( w3944 & w3951 ) | ( w3944 & w3957 ) | ( w3951 & w3957 ) ;
  assign w4078 = ( w3964 & w3965 ) | ( w3964 & w3971 ) | ( w3965 & w3971 ) ;
  assign w4079 = w4076 ^ w4078 ;
  assign w4080 = w4077 ^ w4079 ;
  assign w4081 = ( w3855 & w3890 ) | ( w3855 & w3993 ) | ( w3890 & w3993 ) ;
  assign w4082 = \pi29 & \pi59 ;
  assign w4083 = ( ~\pi60 & w3896 ) | ( ~\pi60 & w4082 ) | ( w3896 & w4082 ) ;
  assign w4084 = \pi31 & w4083 ;
  assign w4085 = ( \pi01 & \pi31 ) | ( \pi01 & ~\pi60 ) | ( \pi31 & ~\pi60 ) ;
  assign w4086 = ( \pi01 & \pi31 ) | ( \pi01 & w3896 ) | ( \pi31 & w3896 ) ;
  assign w4087 = ( w4084 & ~w4085 ) | ( w4084 & w4086 ) | ( ~w4085 & w4086 ) ;
  assign w4088 = ( w3840 & w3846 ) | ( w3840 & w3879 ) | ( w3846 & w3879 ) ;
  assign w4089 = w4081 ^ w4087 ;
  assign w4090 = w4088 ^ w4089 ;
  assign w4091 = ( w4033 & w4034 ) | ( w4033 & w4053 ) | ( w4034 & w4053 ) ;
  assign w4092 = w4080 ^ w4091 ;
  assign w4093 = w4090 ^ w4092 ;
  assign w4094 = ( w3963 & w3973 ) | ( w3963 & w3985 ) | ( w3973 & w3985 ) ;
  assign w4095 = \pi19 & \pi43 ;
  assign w4096 = \pi18 & \pi44 ;
  assign w4097 = \pi08 & \pi54 ;
  assign w4098 = ( w4095 & w4096 ) | ( w4095 & w4097 ) | ( w4096 & w4097 ) ;
  assign w4099 = w4095 ^ w4097 ;
  assign w4100 = w4096 ^ w4099 ;
  assign w4101 = \pi29 & \pi33 ;
  assign w4102 = \pi28 & \pi34 ;
  assign w4103 = \pi27 & \pi35 ;
  assign w4104 = ( w4101 & w4102 ) | ( w4101 & w4103 ) | ( w4102 & w4103 ) ;
  assign w4105 = w4101 ^ w4103 ;
  assign w4106 = w4102 ^ w4105 ;
  assign w4107 = \pi24 & \pi38 ;
  assign w4108 = \pi23 & \pi39 ;
  assign w4109 = \pi22 & \pi40 ;
  assign w4110 = ( w4107 & w4108 ) | ( w4107 & w4109 ) | ( w4108 & w4109 ) ;
  assign w4111 = w4107 ^ w4109 ;
  assign w4112 = w4108 ^ w4111 ;
  assign w4113 = w4100 ^ w4106 ;
  assign w4114 = w4112 ^ w4113 ;
  assign w4115 = \pi02 & \pi60 ;
  assign w4116 = \pi00 & \pi62 ;
  assign w4117 = ( w3977 & w4115 ) | ( w3977 & w4116 ) | ( w4115 & w4116 ) ;
  assign w4118 = w3977 ^ w4116 ;
  assign w4119 = w4115 ^ w4118 ;
  assign w4120 = \pi26 & \pi36 ;
  assign w4121 = \pi25 & \pi37 ;
  assign w4122 = \pi21 & \pi41 ;
  assign w4123 = ( w4120 & w4121 ) | ( w4120 & w4122 ) | ( w4121 & w4122 ) ;
  assign w4124 = w4120 ^ w4122 ;
  assign w4125 = w4121 ^ w4124 ;
  assign w4126 = \pi17 & \pi45 ;
  assign w4127 = \pi10 & \pi52 ;
  assign w4128 = \pi09 & \pi53 ;
  assign w4129 = ( w4126 & w4127 ) | ( w4126 & w4128 ) | ( w4127 & w4128 ) ;
  assign w4130 = w4126 ^ w4128 ;
  assign w4131 = w4127 ^ w4130 ;
  assign w4132 = w4119 ^ w4125 ;
  assign w4133 = w4131 ^ w4132 ;
  assign w4134 = \pi16 & \pi46 ;
  assign w4135 = \pi15 & \pi47 ;
  assign w4136 = \pi11 & \pi51 ;
  assign w4137 = ( w4134 & w4135 ) | ( w4134 & w4136 ) | ( w4135 & w4136 ) ;
  assign w4138 = w4134 ^ w4136 ;
  assign w4139 = w4135 ^ w4138 ;
  assign w4140 = \pi14 & \pi48 ;
  assign w4141 = \pi13 & \pi49 ;
  assign w4142 = \pi12 & \pi50 ;
  assign w4143 = ( w4140 & w4141 ) | ( w4140 & w4142 ) | ( w4141 & w4142 ) ;
  assign w4144 = w4140 ^ w4142 ;
  assign w4145 = w4141 ^ w4144 ;
  assign w4146 = \pi20 & \pi42 ;
  assign w4147 = \pi07 & \pi55 ;
  assign w4148 = \pi06 & \pi56 ;
  assign w4149 = ( w4146 & w4147 ) | ( w4146 & w4148 ) | ( w4147 & w4148 ) ;
  assign w4150 = w4146 ^ w4148 ;
  assign w4151 = w4147 ^ w4150 ;
  assign w4152 = w4139 ^ w4145 ;
  assign w4153 = w4151 ^ w4152 ;
  assign w4154 = w4114 ^ w4133 ;
  assign w4155 = w4153 ^ w4154 ;
  assign w4156 = w4008 ^ w4094 ;
  assign w4157 = w4155 ^ w4156 ;
  assign w4158 = w4067 ^ w4157 ;
  assign w4159 = w4093 ^ w4158 ;
  assign w4160 = ( w4010 & w4011 ) | ( w4010 & w4057 ) | ( w4011 & w4057 ) ;
  assign w4161 = ( w3834 & w3861 ) | ( w3834 & w3902 ) | ( w3861 & w3902 ) ;
  assign w4162 = ( w4040 & w4045 ) | ( w4040 & w4051 ) | ( w4045 & w4051 ) ;
  assign w4163 = ( w4019 & w4026 ) | ( w4019 & w4031 ) | ( w4026 & w4031 ) ;
  assign w4164 = w4161 ^ w4162 ;
  assign w4165 = w4163 ^ w4164 ;
  assign w4166 = w3942 ^ w4038 ;
  assign w4167 = w4043 ^ w4166 ;
  assign w4168 = w3955 ^ w3969 ;
  assign w4169 = w4049 ^ w4168 ;
  assign w4170 = ( ~\pi01 & \pi61 ) | ( ~\pi01 & w1166 ) | ( \pi61 & w1166 ) ;
  assign w4171 = \pi01 & w4170 ;
  assign w4172 = \pi01 & \pi61 ;
  assign w4173 = w4024 ^ w4029 ;
  assign w4174 = w1166 ^ w4173 ;
  assign w4175 = w4172 ^ w4174 ;
  assign w4176 = w4167 ^ w4169 ;
  assign w4177 = w4175 ^ w4176 ;
  assign w4178 = ( w3938 & w3959 ) | ( w3938 & w3960 ) | ( w3959 & w3960 ) ;
  assign w4179 = w4165 ^ w4178 ;
  assign w4180 = w4177 ^ w4179 ;
  assign w4181 = ( w4001 & w4003 ) | ( w4001 & w4005 ) | ( w4003 & w4005 ) ;
  assign w4182 = ( w3974 & w3975 ) | ( w3974 & w3983 ) | ( w3975 & w3983 ) ;
  assign w4183 = ( w3995 & w3996 ) | ( w3995 & w3998 ) | ( w3996 & w3998 ) ;
  assign w4184 = w4181 ^ w4183 ;
  assign w4185 = w4182 ^ w4184 ;
  assign w4186 = ( w4012 & w4013 ) | ( w4012 & w4055 ) | ( w4013 & w4055 ) ;
  assign w4187 = w4180 ^ w4186 ;
  assign w4188 = w4185 ^ w4187 ;
  assign w4189 = w4159 ^ w4160 ;
  assign w4190 = w4188 ^ w4189 ;
  assign w4191 = w4066 & w4190 ;
  assign w4192 = w4066 | w4190 ;
  assign w4193 = ~w4191 & w4192 ;
  assign w4194 = w4065 ^ w4193 ;
  assign w4195 = ( w4065 & w4191 ) | ( w4065 & w4192 ) | ( w4191 & w4192 ) ;
  assign w4196 = w4191 | w4195 ;
  assign w4197 = ( w4159 & w4160 ) | ( w4159 & w4188 ) | ( w4160 & w4188 ) ;
  assign w4198 = ( w4008 & w4094 ) | ( w4008 & w4155 ) | ( w4094 & w4155 ) ;
  assign w4199 = ( w4167 & w4169 ) | ( w4167 & w4175 ) | ( w4169 & w4175 ) ;
  assign w4200 = ( w4161 & w4162 ) | ( w4161 & w4163 ) | ( w4162 & w4163 ) ;
  assign w4201 = ( w4076 & w4077 ) | ( w4076 & w4078 ) | ( w4077 & w4078 ) ;
  assign w4202 = w4199 ^ w4201 ;
  assign w4203 = w4200 ^ w4202 ;
  assign w4204 = ( w3949 & w4017 ) | ( w3949 & w4074 ) | ( w4017 & w4074 ) ;
  assign w4205 = ( w3955 & w3969 ) | ( w3955 & w4049 ) | ( w3969 & w4049 ) ;
  assign w4206 = w1166 ^ w4172 ;
  assign w4207 = ( w4024 & w4029 ) | ( w4024 & w4206 ) | ( w4029 & w4206 ) ;
  assign w4208 = w4204 ^ w4205 ;
  assign w4209 = w4207 ^ w4208 ;
  assign w4210 = ( w4114 & w4133 ) | ( w4114 & w4153 ) | ( w4133 & w4153 ) ;
  assign w4211 = w4110 ^ w4143 ;
  assign w4212 = w4149 ^ w4211 ;
  assign w4213 = w4072 ^ w4117 ;
  assign w4214 = w4123 ^ w4213 ;
  assign w4215 = ( w3942 & w4038 ) | ( w3942 & w4043 ) | ( w4038 & w4043 ) ;
  assign w4216 = w4212 ^ w4214 ;
  assign w4217 = w4215 ^ w4216 ;
  assign w4218 = w4210 ^ w4217 ;
  assign w4219 = w4209 ^ w4218 ;
  assign w4220 = ( w4198 & w4203 ) | ( w4198 & w4219 ) | ( w4203 & w4219 ) ;
  assign w4221 = w4198 ^ w4203 ;
  assign w4222 = w4219 ^ w4221 ;
  assign w4223 = ( w4067 & w4093 ) | ( w4067 & w4157 ) | ( w4093 & w4157 ) ;
  assign w4224 = ( w4180 & w4185 ) | ( w4180 & w4186 ) | ( w4185 & w4186 ) ;
  assign w4225 = ( w4181 & w4182 ) | ( w4181 & w4183 ) | ( w4182 & w4183 ) ;
  assign w4226 = w4098 ^ w4104 ;
  assign w4227 = w4129 ^ w4226 ;
  assign w4228 = ( w4100 & w4106 ) | ( w4100 & w4112 ) | ( w4106 & w4112 ) ;
  assign w4229 = ( w4139 & w4145 ) | ( w4139 & w4151 ) | ( w4145 & w4151 ) ;
  assign w4230 = w4227 ^ w4228 ;
  assign w4231 = w4229 ^ w4230 ;
  assign w4232 = ( w4081 & w4087 ) | ( w4081 & w4088 ) | ( w4087 & w4088 ) ;
  assign w4233 = ( w4119 & w4125 ) | ( w4119 & w4131 ) | ( w4125 & w4131 ) ;
  assign w4234 = \pi01 & \pi62 ;
  assign w4235 = w4171 ^ w4234 ;
  assign w4236 = \pi32 ^ w4235 ;
  assign w4237 = \pi00 & \pi63 ;
  assign w4238 = w4236 ^ w4237 ;
  assign w4239 = \pi26 & \pi37 ;
  assign w4240 = \pi25 & \pi38 ;
  assign w4241 = \pi24 & \pi39 ;
  assign w4242 = ( w4239 & w4240 ) | ( w4239 & w4241 ) | ( w4240 & w4241 ) ;
  assign w4243 = w4239 ^ w4241 ;
  assign w4244 = w4240 ^ w4243 ;
  assign w4245 = \pi29 & \pi34 ;
  assign w4246 = \pi28 & \pi35 ;
  assign w4247 = \pi27 & \pi36 ;
  assign w4248 = ( w4245 & w4246 ) | ( w4245 & w4247 ) | ( w4246 & w4247 ) ;
  assign w4249 = w4245 ^ w4247 ;
  assign w4250 = w4246 ^ w4249 ;
  assign w4251 = w4238 ^ w4244 ;
  assign w4252 = w4250 ^ w4251 ;
  assign w4253 = w4232 ^ w4252 ;
  assign w4254 = w4233 ^ w4253 ;
  assign w4255 = w4225 ^ w4254 ;
  assign w4256 = w4231 ^ w4255 ;
  assign w4257 = ( w4165 & w4177 ) | ( w4165 & w4178 ) | ( w4177 & w4178 ) ;
  assign w4258 = ( w4080 & w4090 ) | ( w4080 & w4091 ) | ( w4090 & w4091 ) ;
  assign w4259 = \pi46 & \pi54 ;
  assign w4260 = \pi18 & \pi45 ;
  assign w4261 = \pi17 & \pi46 ;
  assign w4262 = \pi09 & \pi54 ;
  assign w4263 = ( w4260 & w4261 ) | ( w4260 & w4262 ) | ( w4261 & w4262 ) ;
  assign w4264 = w4260 ^ w4262 ;
  assign w4265 = w4261 ^ w4264 ;
  assign w4266 = \pi16 & \pi47 ;
  assign w4267 = \pi11 & \pi52 ;
  assign w4268 = \pi10 & \pi53 ;
  assign w4269 = ( w4266 & w4267 ) | ( w4266 & w4268 ) | ( w4267 & w4268 ) ;
  assign w4270 = w4266 ^ w4268 ;
  assign w4271 = w4267 ^ w4270 ;
  assign w4272 = \pi15 & \pi48 ;
  assign w4273 = \pi13 & \pi50 ;
  assign w4274 = \pi12 & \pi51 ;
  assign w4275 = ( w4272 & w4273 ) | ( w4272 & w4274 ) | ( w4273 & w4274 ) ;
  assign w4276 = w4272 ^ w4274 ;
  assign w4277 = w4273 ^ w4276 ;
  assign w4278 = w4265 ^ w4271 ;
  assign w4279 = w4277 ^ w4278 ;
  assign w4280 = \pi23 & \pi40 ;
  assign w4281 = \pi20 & \pi43 ;
  assign w4282 = \pi06 & \pi57 ;
  assign w4283 = ( w4280 & w4281 ) | ( w4280 & w4282 ) | ( w4281 & w4282 ) ;
  assign w4284 = w4280 ^ w4282 ;
  assign w4285 = w4281 ^ w4284 ;
  assign w4286 = \pi30 & \pi33 ;
  assign w4287 = \pi14 & \pi49 ;
  assign w4288 = ( w1772 & w4286 ) | ( w1772 & w4287 ) | ( w4286 & w4287 ) ;
  assign w4289 = w1772 ^ w4287 ;
  assign w4290 = w4286 ^ w4289 ;
  assign w4291 = \pi19 & \pi44 ;
  assign w4292 = \pi08 & \pi55 ;
  assign w4293 = \pi07 & \pi56 ;
  assign w4294 = ( w4291 & w4292 ) | ( w4291 & w4293 ) | ( w4292 & w4293 ) ;
  assign w4295 = w4291 ^ w4293 ;
  assign w4296 = w4292 ^ w4295 ;
  assign w4297 = w4285 ^ w4290 ;
  assign w4298 = w4296 ^ w4297 ;
  assign w4299 = \pi59 & \pi60 ;
  assign w4300 = \pi60 & \pi61 ;
  assign w4301 = \pi04 & \pi59 ;
  assign w4302 = \pi03 & \pi60 ;
  assign w4303 = \pi02 & \pi61 ;
  assign w4304 = ( w4301 & w4302 ) | ( w4301 & w4303 ) | ( w4302 & w4303 ) ;
  assign w4305 = w4301 ^ w4303 ;
  assign w4306 = w4302 ^ w4305 ;
  assign w4307 = \pi22 & \pi41 ;
  assign w4308 = \pi21 & \pi42 ;
  assign w4309 = \pi05 & \pi58 ;
  assign w4310 = ( w4307 & w4308 ) | ( w4307 & w4309 ) | ( w4308 & w4309 ) ;
  assign w4311 = w4307 ^ w4309 ;
  assign w4312 = w4308 ^ w4311 ;
  assign w4313 = w4137 ^ w4306 ;
  assign w4314 = w4312 ^ w4313 ;
  assign w4315 = w4279 ^ w4298 ;
  assign w4316 = w4314 ^ w4315 ;
  assign w4317 = w4257 ^ w4258 ;
  assign w4318 = w4316 ^ w4317 ;
  assign w4319 = w4224 ^ w4318 ;
  assign w4320 = w4256 ^ w4319 ;
  assign w4321 = w4222 ^ w4223 ;
  assign w4322 = w4320 ^ w4321 ;
  assign w4323 = w4196 ^ w4197 ;
  assign w4324 = w4322 ^ w4323 ;
  assign w4325 = ( w4196 & w4197 ) | ( w4196 & w4322 ) | ( w4197 & w4322 ) ;
  assign w4326 = ( w4224 & w4256 ) | ( w4224 & w4318 ) | ( w4256 & w4318 ) ;
  assign w4327 = ( w4257 & w4258 ) | ( w4257 & w4316 ) | ( w4258 & w4316 ) ;
  assign w4328 = ( w4225 & w4231 ) | ( w4225 & w4254 ) | ( w4231 & w4254 ) ;
  assign w4329 = ( w4279 & w4298 ) | ( w4279 & w4314 ) | ( w4298 & w4314 ) ;
  assign w4330 = ( w4232 & w4233 ) | ( w4232 & w4252 ) | ( w4233 & w4252 ) ;
  assign w4331 = ( w4238 & w4244 ) | ( w4238 & w4250 ) | ( w4244 & w4250 ) ;
  assign w4332 = w4248 ^ w4263 ;
  assign w4333 = w4283 ^ w4332 ;
  assign w4334 = w4294 ^ w4304 ;
  assign w4335 = w4310 ^ w4334 ;
  assign w4336 = w4331 ^ w4333 ;
  assign w4337 = w4335 ^ w4336 ;
  assign w4338 = w4330 ^ w4337 ;
  assign w4339 = w4329 ^ w4338 ;
  assign w4340 = w4327 ^ w4328 ;
  assign w4341 = w4339 ^ w4340 ;
  assign w4342 = ( w4209 & w4210 ) | ( w4209 & w4217 ) | ( w4210 & w4217 ) ;
  assign w4343 = \pi17 & \pi47 ;
  assign w4344 = \pi07 & \pi57 ;
  assign w4345 = \pi06 & \pi58 ;
  assign w4346 = ( w4343 & w4344 ) | ( w4343 & w4345 ) | ( w4344 & w4345 ) ;
  assign w4347 = w4343 ^ w4345 ;
  assign w4348 = w4344 ^ w4347 ;
  assign w4349 = \pi22 & \pi42 ;
  assign w4350 = \pi21 & \pi43 ;
  assign w4351 = \pi20 & \pi44 ;
  assign w4352 = ( w4349 & w4350 ) | ( w4349 & w4351 ) | ( w4350 & w4351 ) ;
  assign w4353 = w4349 ^ w4351 ;
  assign w4354 = w4350 ^ w4353 ;
  assign w4355 = \pi25 & \pi39 ;
  assign w4356 = \pi24 & \pi40 ;
  assign w4357 = \pi23 & \pi41 ;
  assign w4358 = ( w4355 & w4356 ) | ( w4355 & w4357 ) | ( w4356 & w4357 ) ;
  assign w4359 = w4355 ^ w4357 ;
  assign w4360 = w4356 ^ w4359 ;
  assign w4361 = w4348 ^ w4354 ;
  assign w4362 = w4360 ^ w4361 ;
  assign w4363 = \pi26 & \pi38 ;
  assign w4364 = \pi16 & \pi48 ;
  assign w4365 = \pi08 & \pi56 ;
  assign w4366 = ( w4363 & w4364 ) | ( w4363 & w4365 ) | ( w4364 & w4365 ) ;
  assign w4367 = w4363 ^ w4365 ;
  assign w4368 = w4364 ^ w4367 ;
  assign w4369 = \pi29 & \pi35 ;
  assign w4370 = \pi28 & \pi36 ;
  assign w4371 = \pi27 & \pi37 ;
  assign w4372 = ( w4369 & w4370 ) | ( w4369 & w4371 ) | ( w4370 & w4371 ) ;
  assign w4373 = w4369 ^ w4371 ;
  assign w4374 = w4370 ^ w4373 ;
  assign w4375 = \pi31 & \pi33 ;
  assign w4376 = \pi30 & \pi34 ;
  assign w4377 = ( w4020 & w4375 ) | ( w4020 & w4376 ) | ( w4375 & w4376 ) ;
  assign w4378 = w4020 ^ w4376 ;
  assign w4379 = w4375 ^ w4378 ;
  assign w4380 = w4368 ^ w4379 ;
  assign w4381 = w4374 ^ w4380 ;
  assign w4382 = \pi19 & \pi45 ;
  assign w4383 = \pi18 & \pi46 ;
  assign w4384 = \pi05 & \pi59 ;
  assign w4385 = ( w4382 & w4383 ) | ( w4382 & w4384 ) | ( w4383 & w4384 ) ;
  assign w4386 = w4382 ^ w4384 ;
  assign w4387 = w4383 ^ w4386 ;
  assign w4388 = \pi32 ^ w4234 ;
  assign w4389 = ( w4171 & w4237 ) | ( w4171 & w4388 ) | ( w4237 & w4388 ) ;
  assign w4390 = \pi61 & \pi62 ;
  assign w4391 = \pi04 & \pi60 ;
  assign w4392 = \pi03 & \pi61 ;
  assign w4393 = \pi02 & \pi62 ;
  assign w4394 = ( w4391 & w4392 ) | ( w4391 & w4393 ) | ( w4392 & w4393 ) ;
  assign w4395 = w4391 ^ w4393 ;
  assign w4396 = w4392 ^ w4395 ;
  assign w4397 = w4387 ^ w4389 ;
  assign w4398 = w4396 ^ w4397 ;
  assign w4399 = w4381 ^ w4398 ;
  assign w4400 = w4362 ^ w4399 ;
  assign w4401 = ( w4110 & w4143 ) | ( w4110 & w4149 ) | ( w4143 & w4149 ) ;
  assign w4402 = ( w4098 & w4104 ) | ( w4098 & w4129 ) | ( w4104 & w4129 ) ;
  assign w4403 = ( w4072 & w4117 ) | ( w4072 & w4123 ) | ( w4117 & w4123 ) ;
  assign w4404 = w4401 ^ w4403 ;
  assign w4405 = w4402 ^ w4404 ;
  assign w4406 = ( w4227 & w4228 ) | ( w4227 & w4229 ) | ( w4228 & w4229 ) ;
  assign w4407 = ( w4212 & w4214 ) | ( w4212 & w4215 ) | ( w4214 & w4215 ) ;
  assign w4408 = w4406 ^ w4407 ;
  assign w4409 = w4405 ^ w4408 ;
  assign w4410 = w4342 ^ w4409 ;
  assign w4411 = w4400 ^ w4410 ;
  assign w4412 = w4242 ^ w4269 ;
  assign w4413 = w4275 ^ w4412 ;
  assign w4414 = ( w4285 & w4290 ) | ( w4285 & w4296 ) | ( w4290 & w4296 ) ;
  assign w4415 = ( w4265 & w4271 ) | ( w4265 & w4277 ) | ( w4271 & w4277 ) ;
  assign w4416 = w4413 ^ w4414 ;
  assign w4417 = w4415 ^ w4416 ;
  assign w4418 = ( w4199 & w4200 ) | ( w4199 & w4201 ) | ( w4200 & w4201 ) ;
  assign w4419 = ( w4204 & w4205 ) | ( w4204 & w4207 ) | ( w4205 & w4207 ) ;
  assign w4420 = ( w4137 & w4306 ) | ( w4137 & w4312 ) | ( w4306 & w4312 ) ;
  assign w4421 = ( ~\pi01 & \pi32 ) | ( ~\pi01 & \pi62 ) | ( \pi32 & \pi62 ) ;
  assign w4422 = \pi63 ^ w4421 ;
  assign w4423 = \pi01 & w4422 ;
  assign w4424 = w4288 ^ w4423 ;
  assign w4425 = \pi15 & \pi49 ;
  assign w4426 = \pi10 & \pi54 ;
  assign w4427 = \pi09 & \pi55 ;
  assign w4428 = ( w4425 & w4426 ) | ( w4425 & w4427 ) | ( w4426 & w4427 ) ;
  assign w4429 = w4425 ^ w4427 ;
  assign w4430 = w4426 ^ w4429 ;
  assign w4431 = \pi13 & \pi51 ;
  assign w4432 = \pi12 & \pi52 ;
  assign w4433 = \pi11 & \pi53 ;
  assign w4434 = ( w4431 & w4432 ) | ( w4431 & w4433 ) | ( w4432 & w4433 ) ;
  assign w4435 = w4431 ^ w4433 ;
  assign w4436 = w4432 ^ w4435 ;
  assign w4437 = w4424 ^ w4430 ;
  assign w4438 = w4436 ^ w4437 ;
  assign w4439 = w4419 ^ w4438 ;
  assign w4440 = w4420 ^ w4439 ;
  assign w4441 = w4418 ^ w4440 ;
  assign w4442 = w4417 ^ w4441 ;
  assign w4443 = w4220 ^ w4442 ;
  assign w4444 = w4411 ^ w4443 ;
  assign w4445 = w4326 ^ w4444 ;
  assign w4446 = w4341 ^ w4445 ;
  assign w4447 = ( w4222 & w4223 ) | ( w4222 & w4320 ) | ( w4223 & w4320 ) ;
  assign w4448 = w4446 | w4447 ;
  assign w4449 = w4446 & w4447 ;
  assign w4450 = w4448 & ~w4449 ;
  assign w4451 = w4325 ^ w4450 ;
  assign w4452 = ( w4325 & w4448 ) | ( w4325 & w4449 ) | ( w4448 & w4449 ) ;
  assign w4453 = w4449 | w4452 ;
  assign w4454 = ( w4326 & w4341 ) | ( w4326 & w4444 ) | ( w4341 & w4444 ) ;
  assign w4455 = ( w4220 & w4411 ) | ( w4220 & w4442 ) | ( w4411 & w4442 ) ;
  assign w4456 = ( w4342 & w4400 ) | ( w4342 & w4409 ) | ( w4400 & w4409 ) ;
  assign w4457 = ( w4417 & w4418 ) | ( w4417 & w4440 ) | ( w4418 & w4440 ) ;
  assign w4458 = ( w4362 & w4381 ) | ( w4362 & w4398 ) | ( w4381 & w4398 ) ;
  assign w4459 = ( w4419 & w4420 ) | ( w4419 & w4438 ) | ( w4420 & w4438 ) ;
  assign w4460 = ( w4424 & w4430 ) | ( w4424 & w4436 ) | ( w4430 & w4436 ) ;
  assign w4461 = w4346 ^ w4358 ;
  assign w4462 = w4428 ^ w4461 ;
  assign w4463 = w4366 ^ w4385 ;
  assign w4464 = w4394 ^ w4463 ;
  assign w4465 = w4460 ^ w4462 ;
  assign w4466 = w4464 ^ w4465 ;
  assign w4467 = w4458 ^ w4459 ;
  assign w4468 = w4466 ^ w4467 ;
  assign w4469 = w4456 ^ w4457 ;
  assign w4470 = w4468 ^ w4469 ;
  assign w4471 = ( w4327 & w4328 ) | ( w4327 & w4339 ) | ( w4328 & w4339 ) ;
  assign w4472 = ( w4401 & w4402 ) | ( w4401 & w4403 ) | ( w4402 & w4403 ) ;
  assign w4473 = ( w4387 & w4389 ) | ( w4387 & w4396 ) | ( w4389 & w4396 ) ;
  assign w4474 = \pi61 & \pi63 ;
  assign w4475 = \pi04 & \pi61 ;
  assign w4476 = ( \pi02 & \pi63 ) | ( \pi02 & ~w4377 ) | ( \pi63 & ~w4377 ) ;
  assign w4477 = w4475 ^ w4476 ;
  assign w4478 = w4377 & w4477 ;
  assign w4479 = \pi02 & \pi63 ;
  assign w4480 = w4377 ^ w4479 ;
  assign w4481 = w4475 ^ w4480 ;
  assign w4482 = \pi18 & \pi47 ;
  assign w4483 = \pi13 & \pi52 ;
  assign w4484 = \pi12 & \pi53 ;
  assign w4485 = ( w4482 & w4483 ) | ( w4482 & w4484 ) | ( w4483 & w4484 ) ;
  assign w4486 = w4482 ^ w4484 ;
  assign w4487 = w4483 ^ w4486 ;
  assign w4488 = \pi16 & \pi49 ;
  assign w4489 = \pi15 & \pi50 ;
  assign w4490 = \pi14 & \pi51 ;
  assign w4491 = ( w4488 & w4489 ) | ( w4488 & w4490 ) | ( w4489 & w4490 ) ;
  assign w4492 = w4488 ^ w4490 ;
  assign w4493 = w4489 ^ w4492 ;
  assign w4494 = w4481 ^ w4487 ;
  assign w4495 = w4493 ^ w4494 ;
  assign w4496 = w4472 ^ w4473 ;
  assign w4497 = w4495 ^ w4496 ;
  assign w4498 = w4352 ^ w4372 ;
  assign w4499 = w4434 ^ w4498 ;
  assign w4500 = ( w4368 & w4374 ) | ( w4368 & w4379 ) | ( w4374 & w4379 ) ;
  assign w4501 = ( w4348 & w4354 ) | ( w4348 & w4360 ) | ( w4354 & w4360 ) ;
  assign w4502 = w4499 ^ w4500 ;
  assign w4503 = w4501 ^ w4502 ;
  assign w4504 = ( w4405 & w4406 ) | ( w4405 & w4407 ) | ( w4406 & w4407 ) ;
  assign w4505 = w4497 ^ w4504 ;
  assign w4506 = w4503 ^ w4505 ;
  assign w4507 = ( w4329 & w4330 ) | ( w4329 & w4337 ) | ( w4330 & w4337 ) ;
  assign w4508 = \pi20 & \pi45 ;
  assign w4509 = \pi10 & \pi55 ;
  assign w4510 = \pi09 & \pi56 ;
  assign w4511 = ( w4508 & w4509 ) | ( w4508 & w4510 ) | ( w4509 & w4510 ) ;
  assign w4512 = w4508 ^ w4510 ;
  assign w4513 = w4509 ^ w4512 ;
  assign w4514 = \pi25 & \pi40 ;
  assign w4515 = \pi24 & \pi41 ;
  assign w4516 = \pi23 & \pi42 ;
  assign w4517 = ( w4514 & w4515 ) | ( w4514 & w4516 ) | ( w4515 & w4516 ) ;
  assign w4518 = w4514 ^ w4516 ;
  assign w4519 = w4515 ^ w4518 ;
  assign w4520 = \pi28 & \pi37 ;
  assign w4521 = \pi27 & \pi38 ;
  assign w4522 = \pi26 & \pi39 ;
  assign w4523 = ( w4520 & w4521 ) | ( w4520 & w4522 ) | ( w4521 & w4522 ) ;
  assign w4524 = w4520 ^ w4522 ;
  assign w4525 = w4521 ^ w4524 ;
  assign w4526 = w4513 ^ w4519 ;
  assign w4527 = w4525 ^ w4526 ;
  assign w4528 = \pi29 & \pi36 ;
  assign w4529 = \pi19 & \pi46 ;
  assign w4530 = \pi11 & \pi54 ;
  assign w4531 = ( w4528 & w4529 ) | ( w4528 & w4530 ) | ( w4529 & w4530 ) ;
  assign w4532 = w4528 ^ w4530 ;
  assign w4533 = w4529 ^ w4532 ;
  assign w4534 = \pi32 & \pi33 ;
  assign w4535 = \pi31 & \pi34 ;
  assign w4536 = \pi30 & \pi35 ;
  assign w4537 = ( w4534 & w4535 ) | ( w4534 & w4536 ) | ( w4535 & w4536 ) ;
  assign w4538 = w4534 ^ w4536 ;
  assign w4539 = w4535 ^ w4538 ;
  assign w4540 = \pi17 & \pi48 ;
  assign w4541 = \pi03 & \pi62 ;
  assign w4542 = ( \pi33 & w4540 ) | ( \pi33 & w4541 ) | ( w4540 & w4541 ) ;
  assign w4543 = \pi33 ^ w4541 ;
  assign w4544 = w4540 ^ w4543 ;
  assign w4545 = w4533 ^ w4539 ;
  assign w4546 = w4544 ^ w4545 ;
  assign w4547 = \pi22 & \pi43 ;
  assign w4548 = \pi21 & \pi44 ;
  assign w4549 = \pi08 & \pi57 ;
  assign w4550 = ( w4547 & w4548 ) | ( w4547 & w4549 ) | ( w4548 & w4549 ) ;
  assign w4551 = w4547 ^ w4549 ;
  assign w4552 = w4548 ^ w4551 ;
  assign w4553 = ( \pi63 & w4288 ) | ( \pi63 & w4421 ) | ( w4288 & w4421 ) ;
  assign w4554 = \pi01 & w4553 ;
  assign w4555 = \pi07 & \pi58 ;
  assign w4556 = \pi06 & \pi59 ;
  assign w4557 = \pi05 & \pi60 ;
  assign w4558 = ( w4555 & w4556 ) | ( w4555 & w4557 ) | ( w4556 & w4557 ) ;
  assign w4559 = w4555 ^ w4557 ;
  assign w4560 = w4556 ^ w4559 ;
  assign w4561 = w4552 ^ w4554 ;
  assign w4562 = w4560 ^ w4561 ;
  assign w4563 = w4527 ^ w4562 ;
  assign w4564 = w4546 ^ w4563 ;
  assign w4565 = ( w4242 & w4269 ) | ( w4242 & w4275 ) | ( w4269 & w4275 ) ;
  assign w4566 = ( w4248 & w4263 ) | ( w4248 & w4283 ) | ( w4263 & w4283 ) ;
  assign w4567 = ( w4294 & w4304 ) | ( w4294 & w4310 ) | ( w4304 & w4310 ) ;
  assign w4568 = w4565 ^ w4566 ;
  assign w4569 = w4567 ^ w4568 ;
  assign w4570 = ( w4331 & w4333 ) | ( w4331 & w4335 ) | ( w4333 & w4335 ) ;
  assign w4571 = ( w4413 & w4414 ) | ( w4413 & w4415 ) | ( w4414 & w4415 ) ;
  assign w4572 = w4570 ^ w4571 ;
  assign w4573 = w4569 ^ w4572 ;
  assign w4574 = w4507 ^ w4573 ;
  assign w4575 = w4564 ^ w4574 ;
  assign w4576 = w4471 ^ w4575 ;
  assign w4577 = w4506 ^ w4576 ;
  assign w4578 = w4455 ^ w4577 ;
  assign w4579 = w4470 ^ w4578 ;
  assign w4580 = w4453 ^ w4454 ;
  assign w4581 = w4579 ^ w4580 ;
  assign w4582 = ( w4453 & w4454 ) | ( w4453 & w4579 ) | ( w4454 & w4579 ) ;
  assign w4583 = ( w4455 & w4470 ) | ( w4455 & w4577 ) | ( w4470 & w4577 ) ;
  assign w4584 = ( w4471 & w4506 ) | ( w4471 & w4575 ) | ( w4506 & w4575 ) ;
  assign w4585 = ( w4497 & w4503 ) | ( w4497 & w4504 ) | ( w4503 & w4504 ) ;
  assign w4586 = w4485 ^ w4511 ;
  assign w4587 = w4517 ^ w4586 ;
  assign w4588 = ( w4552 & w4554 ) | ( w4552 & w4560 ) | ( w4554 & w4560 ) ;
  assign w4589 = ( w4513 & w4519 ) | ( w4513 & w4525 ) | ( w4519 & w4525 ) ;
  assign w4590 = w4587 ^ w4588 ;
  assign w4591 = w4589 ^ w4590 ;
  assign w4592 = ( w4527 & w4546 ) | ( w4527 & w4562 ) | ( w4546 & w4562 ) ;
  assign w4593 = ( w4472 & w4473 ) | ( w4472 & w4495 ) | ( w4473 & w4495 ) ;
  assign w4594 = w4591 ^ w4592 ;
  assign w4595 = w4593 ^ w4594 ;
  assign w4596 = ( w4569 & w4570 ) | ( w4569 & w4571 ) | ( w4570 & w4571 ) ;
  assign w4597 = \pi08 & \pi58 ;
  assign w4598 = \pi07 & \pi59 ;
  assign w4599 = \pi06 & \pi60 ;
  assign w4600 = ( w4597 & w4598 ) | ( w4597 & w4599 ) | ( w4598 & w4599 ) ;
  assign w4601 = w4597 ^ w4599 ;
  assign w4602 = w4598 ^ w4601 ;
  assign w4603 = ~\pi02 & w4474 ;
  assign w4604 = ( w4474 & w4478 ) | ( w4474 & ~w4603 ) | ( w4478 & ~w4603 ) ;
  assign w4605 = ( \pi04 & w4478 ) | ( \pi04 & w4604 ) | ( w4478 & w4604 ) ;
  assign w4606 = w4523 ^ w4602 ;
  assign w4607 = w4605 ^ w4606 ;
  assign w4608 = ( w4481 & w4487 ) | ( w4481 & w4493 ) | ( w4487 & w4493 ) ;
  assign w4609 = ( w4565 & w4566 ) | ( w4565 & w4567 ) | ( w4566 & w4567 ) ;
  assign w4610 = w4607 ^ w4608 ;
  assign w4611 = w4609 ^ w4610 ;
  assign w4612 = w4491 ^ w4537 ;
  assign w4613 = w4542 ^ w4612 ;
  assign w4614 = w4531 ^ w4550 ;
  assign w4615 = w4558 ^ w4614 ;
  assign w4616 = ( w4533 & w4539 ) | ( w4533 & w4544 ) | ( w4539 & w4544 ) ;
  assign w4617 = w4613 ^ w4615 ;
  assign w4618 = w4616 ^ w4617 ;
  assign w4619 = w4596 ^ w4611 ;
  assign w4620 = w4618 ^ w4619 ;
  assign w4621 = w4585 ^ w4620 ;
  assign w4622 = w4595 ^ w4621 ;
  assign w4623 = ( w4456 & w4457 ) | ( w4456 & w4468 ) | ( w4457 & w4468 ) ;
  assign w4624 = ( w4507 & w4564 ) | ( w4507 & w4573 ) | ( w4564 & w4573 ) ;
  assign w4625 = w4623 ^ w4624 ;
  assign w4626 = ( w4458 & w4459 ) | ( w4458 & w4466 ) | ( w4459 & w4466 ) ;
  assign w4627 = \pi05 & \pi61 ;
  assign w4628 = \pi04 & \pi62 ;
  assign w4629 = \pi03 & \pi63 ;
  assign w4630 = ( w4627 & w4628 ) | ( w4627 & w4629 ) | ( w4628 & w4629 ) ;
  assign w4631 = w4627 ^ w4629 ;
  assign w4632 = w4628 ^ w4631 ;
  assign w4633 = \pi29 & \pi37 ;
  assign w4634 = \pi28 & \pi38 ;
  assign w4635 = \pi27 & \pi39 ;
  assign w4636 = ( w4633 & w4634 ) | ( w4633 & w4635 ) | ( w4634 & w4635 ) ;
  assign w4637 = w4633 ^ w4635 ;
  assign w4638 = w4634 ^ w4637 ;
  assign w4639 = \pi19 & \pi47 ;
  assign w4640 = \pi12 & \pi54 ;
  assign w4641 = \pi11 & \pi55 ;
  assign w4642 = ( w4639 & w4640 ) | ( w4639 & w4641 ) | ( w4640 & w4641 ) ;
  assign w4643 = w4639 ^ w4641 ;
  assign w4644 = w4640 ^ w4643 ;
  assign w4645 = w4632 ^ w4638 ;
  assign w4646 = w4644 ^ w4645 ;
  assign w4647 = \pi24 & \pi42 ;
  assign w4648 = \pi23 & \pi43 ;
  assign w4649 = \pi09 & \pi57 ;
  assign w4650 = ( w4647 & w4648 ) | ( w4647 & w4649 ) | ( w4648 & w4649 ) ;
  assign w4651 = w4647 ^ w4649 ;
  assign w4652 = w4648 ^ w4651 ;
  assign w4653 = \pi22 & \pi44 ;
  assign w4654 = \pi21 & \pi45 ;
  assign w4655 = \pi20 & \pi46 ;
  assign w4656 = ( w4653 & w4654 ) | ( w4653 & w4655 ) | ( w4654 & w4655 ) ;
  assign w4657 = w4653 ^ w4655 ;
  assign w4658 = w4654 ^ w4657 ;
  assign w4659 = \pi26 & \pi40 ;
  assign w4660 = \pi25 & \pi41 ;
  assign w4661 = \pi10 & \pi56 ;
  assign w4662 = ( w4659 & w4660 ) | ( w4659 & w4661 ) | ( w4660 & w4661 ) ;
  assign w4663 = w4659 ^ w4661 ;
  assign w4664 = w4660 ^ w4663 ;
  assign w4665 = w4652 ^ w4658 ;
  assign w4666 = w4664 ^ w4665 ;
  assign w4667 = \pi18 & \pi48 ;
  assign w4668 = \pi15 & \pi51 ;
  assign w4669 = \pi13 & \pi53 ;
  assign w4670 = ( w4667 & w4668 ) | ( w4667 & w4669 ) | ( w4668 & w4669 ) ;
  assign w4671 = w4667 ^ w4669 ;
  assign w4672 = w4668 ^ w4671 ;
  assign w4673 = \pi31 & \pi35 ;
  assign w4674 = \pi30 & \pi36 ;
  assign w4675 = \pi14 & \pi52 ;
  assign w4676 = ( w4673 & w4674 ) | ( w4673 & w4675 ) | ( w4674 & w4675 ) ;
  assign w4677 = w4673 ^ w4675 ;
  assign w4678 = w4674 ^ w4677 ;
  assign w4679 = \pi17 & \pi49 ;
  assign w4680 = \pi16 & \pi50 ;
  assign w4681 = ( w1898 & w4679 ) | ( w1898 & w4680 ) | ( w4679 & w4680 ) ;
  assign w4682 = w1898 ^ w4680 ;
  assign w4683 = w4679 ^ w4682 ;
  assign w4684 = w4672 ^ w4683 ;
  assign w4685 = w4678 ^ w4684 ;
  assign w4686 = w4646 ^ w4685 ;
  assign w4687 = w4666 ^ w4686 ;
  assign w4688 = ( w4346 & w4358 ) | ( w4346 & w4428 ) | ( w4358 & w4428 ) ;
  assign w4689 = ( w4366 & w4385 ) | ( w4366 & w4394 ) | ( w4385 & w4394 ) ;
  assign w4690 = ( w4352 & w4372 ) | ( w4352 & w4434 ) | ( w4372 & w4434 ) ;
  assign w4691 = w4688 ^ w4689 ;
  assign w4692 = w4690 ^ w4691 ;
  assign w4693 = ( w4460 & w4462 ) | ( w4460 & w4464 ) | ( w4462 & w4464 ) ;
  assign w4694 = ( w4499 & w4500 ) | ( w4499 & w4501 ) | ( w4500 & w4501 ) ;
  assign w4695 = w4693 ^ w4694 ;
  assign w4696 = w4692 ^ w4695 ;
  assign w4697 = w4626 ^ w4696 ;
  assign w4698 = w4687 ^ w4697 ;
  assign w4699 = w4622 ^ w4698 ;
  assign w4700 = w4584 ^ w4699 ;
  assign w4701 = w4625 ^ w4700 ;
  assign w4702 = w4582 ^ w4583 ;
  assign w4703 = w4701 ^ w4702 ;
  assign w4704 = w4625 ^ w4698 ;
  assign w4705 = ( w4584 & w4622 ) | ( w4584 & w4704 ) | ( w4622 & w4704 ) ;
  assign w4706 = ( w4585 & w4595 ) | ( w4585 & w4620 ) | ( w4595 & w4620 ) ;
  assign w4707 = ( w4626 & w4687 ) | ( w4626 & w4696 ) | ( w4687 & w4696 ) ;
  assign w4708 = w4706 ^ w4707 ;
  assign w4709 = ( w4591 & w4592 ) | ( w4591 & w4593 ) | ( w4592 & w4593 ) ;
  assign w4710 = \pi19 & \pi48 ;
  assign w4711 = \pi17 & \pi50 ;
  assign w4712 = \pi14 & \pi53 ;
  assign w4713 = ( w4710 & w4711 ) | ( w4710 & w4712 ) | ( w4711 & w4712 ) ;
  assign w4714 = w4710 ^ w4712 ;
  assign w4715 = w4711 ^ w4714 ;
  assign w4716 = \pi26 & \pi41 ;
  assign w4717 = \pi25 & \pi42 ;
  assign w4718 = \pi21 & \pi46 ;
  assign w4719 = ( w4716 & w4717 ) | ( w4716 & w4718 ) | ( w4717 & w4718 ) ;
  assign w4720 = w4716 ^ w4718 ;
  assign w4721 = w4717 ^ w4720 ;
  assign w4722 = \pi28 & \pi39 ;
  assign w4723 = \pi27 & \pi40 ;
  assign w4724 = \pi04 & \pi63 ;
  assign w4725 = ( w4722 & w4723 ) | ( w4722 & w4724 ) | ( w4723 & w4724 ) ;
  assign w4726 = w4722 ^ w4724 ;
  assign w4727 = w4723 ^ w4726 ;
  assign w4728 = w4715 ^ w4721 ;
  assign w4729 = w4727 ^ w4728 ;
  assign w4730 = \pi18 & \pi49 ;
  assign w4731 = \pi05 & \pi62 ;
  assign w4732 = ( \pi34 & w4730 ) | ( \pi34 & w4731 ) | ( w4730 & w4731 ) ;
  assign w4733 = \pi34 ^ w4731 ;
  assign w4734 = w4730 ^ w4733 ;
  assign w4735 = \pi33 & \pi34 ;
  assign w4736 = \pi32 & \pi35 ;
  assign w4737 = \pi31 & \pi36 ;
  assign w4738 = ( w4735 & w4736 ) | ( w4735 & w4737 ) | ( w4736 & w4737 ) ;
  assign w4739 = w4735 ^ w4737 ;
  assign w4740 = w4736 ^ w4739 ;
  assign w4741 = \pi29 & \pi38 ;
  assign w4742 = \pi13 & \pi54 ;
  assign w4743 = \pi12 & \pi55 ;
  assign w4744 = ( w4741 & w4742 ) | ( w4741 & w4743 ) | ( w4742 & w4743 ) ;
  assign w4745 = w4741 ^ w4743 ;
  assign w4746 = w4742 ^ w4745 ;
  assign w4747 = w4734 ^ w4740 ;
  assign w4748 = w4746 ^ w4747 ;
  assign w4749 = \pi09 & \pi58 ;
  assign w4750 = \pi08 & \pi59 ;
  assign w4751 = \pi07 & \pi60 ;
  assign w4752 = ( w4749 & w4750 ) | ( w4749 & w4751 ) | ( w4750 & w4751 ) ;
  assign w4753 = w4749 ^ w4751 ;
  assign w4754 = w4750 ^ w4753 ;
  assign w4755 = \pi24 & \pi43 ;
  assign w4756 = \pi23 & \pi44 ;
  assign w4757 = \pi22 & \pi45 ;
  assign w4758 = ( w4755 & w4756 ) | ( w4755 & w4757 ) | ( w4756 & w4757 ) ;
  assign w4759 = w4755 ^ w4757 ;
  assign w4760 = w4756 ^ w4759 ;
  assign w4761 = \pi30 & \pi37 ;
  assign w4762 = \pi16 & \pi51 ;
  assign w4763 = \pi15 & \pi52 ;
  assign w4764 = ( w4761 & w4762 ) | ( w4761 & w4763 ) | ( w4762 & w4763 ) ;
  assign w4765 = w4761 ^ w4763 ;
  assign w4766 = w4762 ^ w4765 ;
  assign w4767 = w4754 ^ w4760 ;
  assign w4768 = w4766 ^ w4767 ;
  assign w4769 = w4729 ^ w4748 ;
  assign w4770 = w4768 ^ w4769 ;
  assign w4771 = ( w4531 & w4550 ) | ( w4531 & w4558 ) | ( w4550 & w4558 ) ;
  assign w4772 = ( w4485 & w4511 ) | ( w4485 & w4517 ) | ( w4511 & w4517 ) ;
  assign w4773 = ( w4491 & w4537 ) | ( w4491 & w4542 ) | ( w4537 & w4542 ) ;
  assign w4774 = w4771 ^ w4772 ;
  assign w4775 = w4773 ^ w4774 ;
  assign w4776 = ( w4613 & w4615 ) | ( w4613 & w4616 ) | ( w4615 & w4616 ) ;
  assign w4777 = ( w4587 & w4588 ) | ( w4587 & w4589 ) | ( w4588 & w4589 ) ;
  assign w4778 = w4775 ^ w4777 ;
  assign w4779 = w4776 ^ w4778 ;
  assign w4780 = w4709 ^ w4779 ;
  assign w4781 = w4770 ^ w4780 ;
  assign w4782 = ( w4623 & w4624 ) | ( w4623 & w4698 ) | ( w4624 & w4698 ) ;
  assign w4783 = ( w4596 & w4611 ) | ( w4596 & w4618 ) | ( w4611 & w4618 ) ;
  assign w4784 = ( w4692 & w4693 ) | ( w4692 & w4694 ) | ( w4693 & w4694 ) ;
  assign w4785 = ( w4652 & w4658 ) | ( w4652 & w4664 ) | ( w4658 & w4664 ) ;
  assign w4786 = \pi02 | w4478 ;
  assign w4787 = ( \pi04 & w4478 ) | ( \pi04 & w4786 ) | ( w4478 & w4786 ) ;
  assign w4788 = ( w4474 & w4478 ) | ( w4474 & w4787 ) | ( w4478 & w4787 ) ;
  assign w4789 = ( w4523 & w4602 ) | ( w4523 & w4788 ) | ( w4602 & w4788 ) ;
  assign w4790 = ( w4632 & w4638 ) | ( w4632 & w4644 ) | ( w4638 & w4644 ) ;
  assign w4791 = w4785 ^ w4789 ;
  assign w4792 = w4790 ^ w4791 ;
  assign w4793 = w4600 ^ w4630 ;
  assign w4794 = w4636 ^ w4793 ;
  assign w4795 = w4650 ^ w4656 ;
  assign w4796 = w4662 ^ w4795 ;
  assign w4797 = w4681 ^ w4794 ;
  assign w4798 = w4796 ^ w4797 ;
  assign w4799 = w4676 ^ w4798 ;
  assign w4800 = \pi06 & \pi61 ;
  assign w4801 = w4799 ^ w4800 ;
  assign w4802 = w4784 ^ w4792 ;
  assign w4803 = w4801 ^ w4802 ;
  assign w4804 = \pi20 & \pi47 ;
  assign w4805 = \pi11 & \pi56 ;
  assign w4806 = \pi10 & \pi57 ;
  assign w4807 = ( w4804 & w4805 ) | ( w4804 & w4806 ) | ( w4805 & w4806 ) ;
  assign w4808 = w4804 ^ w4806 ;
  assign w4809 = w4805 ^ w4808 ;
  assign w4810 = w4642 ^ w4670 ;
  assign w4811 = w4809 ^ w4810 ;
  assign w4812 = ( w4672 & w4678 ) | ( w4672 & w4683 ) | ( w4678 & w4683 ) ;
  assign w4813 = ( w4688 & w4689 ) | ( w4688 & w4690 ) | ( w4689 & w4690 ) ;
  assign w4814 = w4812 ^ w4813 ;
  assign w4815 = w4811 ^ w4814 ;
  assign w4816 = ( w4646 & w4666 ) | ( w4646 & w4685 ) | ( w4666 & w4685 ) ;
  assign w4817 = ( w4607 & w4608 ) | ( w4607 & w4609 ) | ( w4608 & w4609 ) ;
  assign w4818 = w4815 ^ w4817 ;
  assign w4819 = w4816 ^ w4818 ;
  assign w4820 = w4783 ^ w4803 ;
  assign w4821 = w4819 ^ w4820 ;
  assign w4822 = w4781 ^ w4821 ;
  assign w4823 = w4708 ^ w4822 ;
  assign w4824 = w4782 ^ w4823 ;
  assign w4825 = ( w4582 & w4583 ) | ( w4582 & w4701 ) | ( w4583 & w4701 ) ;
  assign w4826 = w4705 ^ w4825 ;
  assign w4827 = w4824 ^ w4826 ;
  assign w4828 = ( w4706 & w4707 ) | ( w4706 & w4781 ) | ( w4707 & w4781 ) ;
  assign w4829 = ( w4784 & w4792 ) | ( w4784 & w4801 ) | ( w4792 & w4801 ) ;
  assign w4830 = ( w4729 & w4748 ) | ( w4729 & w4768 ) | ( w4748 & w4768 ) ;
  assign w4831 = ( w4642 & w4670 ) | ( w4642 & w4809 ) | ( w4670 & w4809 ) ;
  assign w4832 = ( w4650 & w4656 ) | ( w4650 & w4662 ) | ( w4656 & w4662 ) ;
  assign w4833 = ( w4754 & w4760 ) | ( w4754 & w4766 ) | ( w4760 & w4766 ) ;
  assign w4834 = w4831 ^ w4832 ;
  assign w4835 = w4833 ^ w4834 ;
  assign w4836 = \pi08 & \pi60 ;
  assign w4837 = \pi07 & \pi61 ;
  assign w4838 = w4732 ^ w4837 ;
  assign w4839 = w4836 ^ w4838 ;
  assign w4840 = ( w4600 & w4630 ) | ( w4600 & w4636 ) | ( w4630 & w4636 ) ;
  assign w4841 = ( w4676 & w4681 ) | ( w4676 & w4800 ) | ( w4681 & w4800 ) ;
  assign w4842 = w4839 ^ w4841 ;
  assign w4843 = w4840 ^ w4842 ;
  assign w4844 = w4830 ^ w4835 ;
  assign w4845 = w4843 ^ w4844 ;
  assign w4846 = ( w4775 & w4776 ) | ( w4775 & w4777 ) | ( w4776 & w4777 ) ;
  assign w4847 = w4713 ^ w4719 ;
  assign w4848 = w4744 ^ w4847 ;
  assign w4849 = ( w4715 & w4721 ) | ( w4715 & w4727 ) | ( w4721 & w4727 ) ;
  assign w4850 = ( w4734 & w4740 ) | ( w4734 & w4746 ) | ( w4740 & w4746 ) ;
  assign w4851 = w4848 ^ w4849 ;
  assign w4852 = w4850 ^ w4851 ;
  assign w4853 = ( w4771 & w4772 ) | ( w4771 & w4773 ) | ( w4772 & w4773 ) ;
  assign w4854 = w4752 ^ w4758 ;
  assign w4855 = w4807 ^ w4854 ;
  assign w4856 = w4725 ^ w4738 ;
  assign w4857 = w4764 ^ w4856 ;
  assign w4858 = w4853 ^ w4855 ;
  assign w4859 = w4857 ^ w4858 ;
  assign w4860 = w4846 ^ w4859 ;
  assign w4861 = w4852 ^ w4860 ;
  assign w4862 = w4829 ^ w4861 ;
  assign w4863 = w4845 ^ w4862 ;
  assign w4864 = ( w4783 & w4803 ) | ( w4783 & w4819 ) | ( w4803 & w4819 ) ;
  assign w4865 = ( w4709 & w4770 ) | ( w4709 & w4779 ) | ( w4770 & w4779 ) ;
  assign w4866 = ( w4815 & w4816 ) | ( w4815 & w4817 ) | ( w4816 & w4817 ) ;
  assign w4867 = w4676 ^ w4681 ;
  assign w4868 = w4800 ^ w4867 ;
  assign w4869 = ( w4794 & w4796 ) | ( w4794 & w4868 ) | ( w4796 & w4868 ) ;
  assign w4870 = ( w4785 & w4789 ) | ( w4785 & w4790 ) | ( w4789 & w4790 ) ;
  assign w4871 = ( w4811 & w4812 ) | ( w4811 & w4813 ) | ( w4812 & w4813 ) ;
  assign w4872 = w4870 ^ w4871 ;
  assign w4873 = w4869 ^ w4872 ;
  assign w4874 = \pi11 & \pi57 ;
  assign w4875 = \pi10 & \pi58 ;
  assign w4876 = \pi09 & \pi59 ;
  assign w4877 = ( w4874 & w4875 ) | ( w4874 & w4876 ) | ( w4875 & w4876 ) ;
  assign w4878 = w4874 ^ w4876 ;
  assign w4879 = w4875 ^ w4878 ;
  assign w4880 = \pi29 & \pi39 ;
  assign w4881 = \pi28 & \pi40 ;
  assign w4882 = \pi27 & \pi41 ;
  assign w4883 = ( w4880 & w4881 ) | ( w4880 & w4882 ) | ( w4881 & w4882 ) ;
  assign w4884 = w4880 ^ w4882 ;
  assign w4885 = w4881 ^ w4884 ;
  assign w4886 = \pi21 & \pi47 ;
  assign w4887 = \pi06 & \pi62 ;
  assign w4888 = \pi05 & \pi63 ;
  assign w4889 = ( w4886 & w4887 ) | ( w4886 & w4888 ) | ( w4887 & w4888 ) ;
  assign w4890 = w4886 ^ w4888 ;
  assign w4891 = w4887 ^ w4890 ;
  assign w4892 = w4879 ^ w4885 ;
  assign w4893 = w4891 ^ w4892 ;
  assign w4894 = \pi19 & \pi49 ;
  assign w4895 = \pi18 & \pi50 ;
  assign w4896 = ( w1389 & w4894 ) | ( w1389 & w4895 ) | ( w4894 & w4895 ) ;
  assign w4897 = w1389 ^ w4895 ;
  assign w4898 = w4894 ^ w4897 ;
  assign w4899 = \pi32 & \pi36 ;
  assign w4900 = \pi31 & \pi37 ;
  assign w4901 = \pi30 & \pi38 ;
  assign w4902 = ( w4899 & w4900 ) | ( w4899 & w4901 ) | ( w4900 & w4901 ) ;
  assign w4903 = w4899 ^ w4901 ;
  assign w4904 = w4900 ^ w4903 ;
  assign w4905 = \pi13 & \pi55 ;
  assign w4906 = \pi12 & \pi56 ;
  assign w4907 = ( w3524 & w4905 ) | ( w3524 & w4906 ) | ( w4905 & w4906 ) ;
  assign w4908 = w3524 ^ w4906 ;
  assign w4909 = w4905 ^ w4908 ;
  assign w4910 = w4898 ^ w4909 ;
  assign w4911 = w4904 ^ w4910 ;
  assign w4912 = \pi16 & \pi52 ;
  assign w4913 = \pi15 & \pi53 ;
  assign w4914 = \pi14 & \pi54 ;
  assign w4915 = ( w4912 & w4913 ) | ( w4912 & w4914 ) | ( w4913 & w4914 ) ;
  assign w4916 = w4912 ^ w4914 ;
  assign w4917 = w4913 ^ w4916 ;
  assign w4918 = \pi23 & \pi45 ;
  assign w4919 = \pi22 & \pi46 ;
  assign w4920 = \pi20 & \pi48 ;
  assign w4921 = ( w4918 & w4919 ) | ( w4918 & w4920 ) | ( w4919 & w4920 ) ;
  assign w4922 = w4918 ^ w4920 ;
  assign w4923 = w4919 ^ w4922 ;
  assign w4924 = \pi26 & \pi42 ;
  assign w4925 = \pi25 & \pi43 ;
  assign w4926 = \pi24 & \pi44 ;
  assign w4927 = ( w4924 & w4925 ) | ( w4924 & w4926 ) | ( w4925 & w4926 ) ;
  assign w4928 = w4924 ^ w4926 ;
  assign w4929 = w4925 ^ w4928 ;
  assign w4930 = w4917 ^ w4923 ;
  assign w4931 = w4929 ^ w4930 ;
  assign w4932 = w4893 ^ w4911 ;
  assign w4933 = w4931 ^ w4932 ;
  assign w4934 = w4866 ^ w4873 ;
  assign w4935 = w4933 ^ w4934 ;
  assign w4936 = w4864 ^ w4865 ;
  assign w4937 = w4935 ^ w4936 ;
  assign w4938 = w4828 ^ w4937 ;
  assign w4939 = w4863 ^ w4938 ;
  assign w4940 = w4708 ^ w4781 ;
  assign w4941 = ( w4782 & w4821 ) | ( w4782 & w4940 ) | ( w4821 & w4940 ) ;
  assign w4942 = ( w4705 & w4824 ) | ( w4705 & w4825 ) | ( w4824 & w4825 ) ;
  assign w4943 = w4939 ^ w4942 ;
  assign w4944 = w4941 ^ w4943 ;
  assign w4945 = ( w4829 & w4845 ) | ( w4829 & w4861 ) | ( w4845 & w4861 ) ;
  assign w4946 = ( w4866 & w4873 ) | ( w4866 & w4933 ) | ( w4873 & w4933 ) ;
  assign w4947 = w4945 ^ w4946 ;
  assign w4948 = ( w4848 & w4849 ) | ( w4848 & w4850 ) | ( w4849 & w4850 ) ;
  assign w4949 = \pi19 & \pi50 ;
  assign w4950 = \pi18 & \pi51 ;
  assign w4951 = \pi17 & \pi52 ;
  assign w4952 = ( w4949 & w4950 ) | ( w4949 & w4951 ) | ( w4950 & w4951 ) ;
  assign w4953 = w4949 ^ w4951 ;
  assign w4954 = w4950 ^ w4953 ;
  assign w4955 = \pi30 & \pi39 ;
  assign w4956 = \pi29 & \pi40 ;
  assign w4957 = \pi28 & \pi41 ;
  assign w4958 = ( w4955 & w4956 ) | ( w4955 & w4957 ) | ( w4956 & w4957 ) ;
  assign w4959 = w4955 ^ w4957 ;
  assign w4960 = w4956 ^ w4959 ;
  assign w4961 = ( w4752 & w4758 ) | ( w4752 & w4807 ) | ( w4758 & w4807 ) ;
  assign w4962 = w4954 ^ w4961 ;
  assign w4963 = w4960 ^ w4962 ;
  assign w4964 = \pi33 & \pi36 ;
  assign w4965 = \pi32 & \pi37 ;
  assign w4966 = \pi31 & \pi38 ;
  assign w4967 = ( w4964 & w4965 ) | ( w4964 & w4966 ) | ( w4965 & w4966 ) ;
  assign w4968 = w4964 ^ w4966 ;
  assign w4969 = w4965 ^ w4968 ;
  assign w4970 = \pi20 & \pi54 ;
  assign w4971 = \pi20 & \pi49 ;
  assign w4972 = \pi16 & \pi53 ;
  assign w4973 = \pi15 & \pi54 ;
  assign w4974 = ( w4971 & w4972 ) | ( w4971 & w4973 ) | ( w4972 & w4973 ) ;
  assign w4975 = w4971 ^ w4973 ;
  assign w4976 = w4972 ^ w4975 ;
  assign w4977 = ~\pi34 & \pi35 ;
  assign w4978 = w4969 ^ w4977 ;
  assign w4979 = w4976 ^ w4978 ;
  assign w4980 = \pi07 & \pi62 ;
  assign w4981 = w4979 ^ w4980 ;
  assign w4982 = ( w4948 & w4963 ) | ( w4948 & w4981 ) | ( w4963 & w4981 ) ;
  assign w4983 = w4948 ^ w4963 ;
  assign w4984 = w4981 ^ w4983 ;
  assign w4985 = ( w4830 & w4835 ) | ( w4830 & w4843 ) | ( w4835 & w4843 ) ;
  assign w4986 = \pi10 & \pi59 ;
  assign w4987 = \pi09 & \pi60 ;
  assign w4988 = \pi08 & \pi61 ;
  assign w4989 = ( w4986 & w4987 ) | ( w4986 & w4988 ) | ( w4987 & w4988 ) ;
  assign w4990 = w4986 ^ w4988 ;
  assign w4991 = w4987 ^ w4990 ;
  assign w4992 = \pi25 & \pi44 ;
  assign w4993 = \pi24 & \pi45 ;
  assign w4994 = \pi23 & \pi46 ;
  assign w4995 = ( w4992 & w4993 ) | ( w4992 & w4994 ) | ( w4993 & w4994 ) ;
  assign w4996 = w4992 ^ w4994 ;
  assign w4997 = w4993 ^ w4996 ;
  assign w4998 = \pi27 & \pi42 ;
  assign w4999 = \pi26 & \pi43 ;
  assign w5000 = \pi06 & \pi63 ;
  assign w5001 = ( w4998 & w4999 ) | ( w4998 & w5000 ) | ( w4999 & w5000 ) ;
  assign w5002 = w4998 ^ w5000 ;
  assign w5003 = w4999 ^ w5002 ;
  assign w5004 = w4991 ^ w4997 ;
  assign w5005 = w5003 ^ w5004 ;
  assign w5006 = ( w4831 & w4832 ) | ( w4831 & w4833 ) | ( w4832 & w4833 ) ;
  assign w5007 = w5005 ^ w5006 ;
  assign w5008 = \pi13 & \pi56 ;
  assign w5009 = \pi12 & \pi57 ;
  assign w5010 = \pi11 & \pi58 ;
  assign w5011 = ( w5008 & w5009 ) | ( w5008 & w5010 ) | ( w5009 & w5010 ) ;
  assign w5012 = w5008 ^ w5010 ;
  assign w5013 = w5009 ^ w5012 ;
  assign w5014 = ( w4732 & w4836 ) | ( w4732 & w4837 ) | ( w4836 & w4837 ) ;
  assign w5015 = \pi22 & \pi47 ;
  assign w5016 = \pi21 & \pi48 ;
  assign w5017 = \pi14 & \pi55 ;
  assign w5018 = ( w5015 & w5016 ) | ( w5015 & w5017 ) | ( w5016 & w5017 ) ;
  assign w5019 = w5015 ^ w5017 ;
  assign w5020 = w5016 ^ w5019 ;
  assign w5021 = w5013 ^ w5014 ;
  assign w5022 = w5020 ^ w5021 ;
  assign w5023 = w5007 ^ w5022 ;
  assign w5024 = w4984 ^ w5023 ;
  assign w5025 = w4985 ^ w5024 ;
  assign w5026 = ( w4864 & w4865 ) | ( w4864 & w4935 ) | ( w4865 & w4935 ) ;
  assign w5027 = ( w4846 & w4852 ) | ( w4846 & w4859 ) | ( w4852 & w4859 ) ;
  assign w5028 = ( w4893 & w4911 ) | ( w4893 & w4931 ) | ( w4911 & w4931 ) ;
  assign w5029 = ( w4853 & w4855 ) | ( w4853 & w4857 ) | ( w4855 & w4857 ) ;
  assign w5030 = w4883 ^ w4907 ;
  assign w5031 = w4927 ^ w5030 ;
  assign w5032 = ( w4725 & w4738 ) | ( w4725 & w4764 ) | ( w4738 & w4764 ) ;
  assign w5033 = ( w4713 & w4719 ) | ( w4713 & w4744 ) | ( w4719 & w4744 ) ;
  assign w5034 = w5031 ^ w5032 ;
  assign w5035 = w5033 ^ w5034 ;
  assign w5036 = w5028 ^ w5029 ;
  assign w5037 = w5035 ^ w5036 ;
  assign w5038 = ( w4869 & w4870 ) | ( w4869 & w4871 ) | ( w4870 & w4871 ) ;
  assign w5039 = ( w4898 & w4904 ) | ( w4898 & w4909 ) | ( w4904 & w4909 ) ;
  assign w5040 = ( w4917 & w4923 ) | ( w4917 & w4929 ) | ( w4923 & w4929 ) ;
  assign w5041 = ( w4839 & w4840 ) | ( w4839 & w4841 ) | ( w4840 & w4841 ) ;
  assign w5042 = w5039 ^ w5041 ;
  assign w5043 = w5040 ^ w5042 ;
  assign w5044 = w4877 ^ w4889 ;
  assign w5045 = w4921 ^ w5044 ;
  assign w5046 = w4896 ^ w4902 ;
  assign w5047 = w4915 ^ w5046 ;
  assign w5048 = ( w4879 & w4885 ) | ( w4879 & w4891 ) | ( w4885 & w4891 ) ;
  assign w5049 = w5045 ^ w5047 ;
  assign w5050 = w5048 ^ w5049 ;
  assign w5051 = w5038 ^ w5043 ;
  assign w5052 = w5050 ^ w5051 ;
  assign w5053 = w5027 ^ w5052 ;
  assign w5054 = w5037 ^ w5053 ;
  assign w5055 = w5025 ^ w5054 ;
  assign w5056 = w4947 ^ w5055 ;
  assign w5057 = w5026 ^ w5056 ;
  assign w5058 = ( w4828 & w4863 ) | ( w4828 & w4937 ) | ( w4863 & w4937 ) ;
  assign w5059 = ( w4939 & w4941 ) | ( w4939 & w4942 ) | ( w4941 & w4942 ) ;
  assign w5060 = w5057 ^ w5059 ;
  assign w5061 = w5058 ^ w5060 ;
  assign w5062 = ( w5057 & w5058 ) | ( w5057 & w5059 ) | ( w5058 & w5059 ) ;
  assign w5063 = w4947 ^ w5025 ;
  assign w5064 = ( w5026 & w5054 ) | ( w5026 & w5063 ) | ( w5054 & w5063 ) ;
  assign w5065 = ( w5027 & w5037 ) | ( w5027 & w5052 ) | ( w5037 & w5052 ) ;
  assign w5066 = w4958 ^ w4995 ;
  assign w5067 = w5001 ^ w5066 ;
  assign w5068 = \pi08 & \pi62 ;
  assign w5069 = ~\pi62 & w1921 ;
  assign w5070 = ( w1540 & w1921 ) | ( w1540 & ~w5069 ) | ( w1921 & ~w5069 ) ;
  assign w5071 = ( w4967 & w5068 ) | ( w4967 & w5070 ) | ( w5068 & w5070 ) ;
  assign w5072 = ( \pi62 & w1540 ) | ( \pi62 & ~w1921 ) | ( w1540 & ~w1921 ) ;
  assign w5073 = \pi08 ^ w5072 ;
  assign w5074 = \pi62 & ~w5073 ;
  assign w5075 = w1540 ^ w4967 ;
  assign w5076 = w5074 ^ w5075 ;
  assign w5077 = ( w4954 & w4960 ) | ( w4954 & w4961 ) | ( w4960 & w4961 ) ;
  assign w5078 = w5067 ^ w5077 ;
  assign w5079 = w5076 ^ w5078 ;
  assign w5080 = ( w4991 & w4997 ) | ( w4991 & w5003 ) | ( w4997 & w5003 ) ;
  assign w5081 = ( w5013 & w5014 ) | ( w5013 & w5020 ) | ( w5014 & w5020 ) ;
  assign w5082 = w4977 ^ w4980 ;
  assign w5083 = ( w4969 & w4976 ) | ( w4969 & w5082 ) | ( w4976 & w5082 ) ;
  assign w5084 = w5080 ^ w5081 ;
  assign w5085 = w5083 ^ w5084 ;
  assign w5086 = w4982 ^ w5085 ;
  assign w5087 = ( w5045 & w5047 ) | ( w5045 & w5048 ) | ( w5047 & w5048 ) ;
  assign w5088 = \pi28 & \pi42 ;
  assign w5089 = \pi07 & \pi63 ;
  assign w5090 = ( w2696 & w5088 ) | ( w2696 & w5089 ) | ( w5088 & w5089 ) ;
  assign w5091 = w5088 ^ w5089 ;
  assign w5092 = w2696 ^ w5091 ;
  assign w5093 = \pi31 & \pi39 ;
  assign w5094 = \pi30 & \pi40 ;
  assign w5095 = \pi29 & \pi41 ;
  assign w5096 = ( w5093 & w5094 ) | ( w5093 & w5095 ) | ( w5094 & w5095 ) ;
  assign w5097 = w5093 ^ w5095 ;
  assign w5098 = w5094 ^ w5097 ;
  assign w5099 = ( w4896 & w4902 ) | ( w4896 & w4915 ) | ( w4902 & w4915 ) ;
  assign w5100 = w5092 ^ w5099 ;
  assign w5101 = w5098 ^ w5100 ;
  assign w5102 = \pi22 & \pi48 ;
  assign w5103 = \pi15 & \pi55 ;
  assign w5104 = \pi14 & \pi56 ;
  assign w5105 = ( w5102 & w5103 ) | ( w5102 & w5104 ) | ( w5103 & w5104 ) ;
  assign w5106 = w5102 ^ w5104 ;
  assign w5107 = w5103 ^ w5106 ;
  assign w5108 = \pi27 & \pi43 ;
  assign w5109 = \pi26 & \pi44 ;
  assign w5110 = \pi25 & \pi45 ;
  assign w5111 = ( w5108 & w5109 ) | ( w5108 & w5110 ) | ( w5109 & w5110 ) ;
  assign w5112 = w5108 ^ w5110 ;
  assign w5113 = w5109 ^ w5112 ;
  assign w5114 = \pi21 & \pi49 ;
  assign w5115 = \pi20 & \pi50 ;
  assign w5116 = \pi19 & \pi51 ;
  assign w5117 = ( w5114 & w5115 ) | ( w5114 & w5116 ) | ( w5115 & w5116 ) ;
  assign w5118 = w5114 ^ w5116 ;
  assign w5119 = w5115 ^ w5118 ;
  assign w5120 = w5107 ^ w5113 ;
  assign w5121 = w5119 ^ w5120 ;
  assign w5122 = ( w5087 & w5101 ) | ( w5087 & w5121 ) | ( w5101 & w5121 ) ;
  assign w5123 = w5087 ^ w5101 ;
  assign w5124 = w5121 ^ w5123 ;
  assign w5125 = ( w5028 & w5029 ) | ( w5028 & w5035 ) | ( w5029 & w5035 ) ;
  assign w5126 = \pi11 & \pi59 ;
  assign w5127 = \pi10 & \pi60 ;
  assign w5128 = \pi09 & \pi61 ;
  assign w5129 = ( w5126 & w5127 ) | ( w5126 & w5128 ) | ( w5127 & w5128 ) ;
  assign w5130 = w5126 ^ w5128 ;
  assign w5131 = w5127 ^ w5130 ;
  assign w5132 = \pi18 & \pi52 ;
  assign w5133 = \pi17 & \pi53 ;
  assign w5134 = \pi16 & \pi54 ;
  assign w5135 = ( w5132 & w5133 ) | ( w5132 & w5134 ) | ( w5133 & w5134 ) ;
  assign w5136 = w5132 ^ w5134 ;
  assign w5137 = w5133 ^ w5136 ;
  assign w5138 = \pi24 & \pi46 ;
  assign w5139 = \pi13 & \pi57 ;
  assign w5140 = \pi12 & \pi58 ;
  assign w5141 = ( w5138 & w5139 ) | ( w5138 & w5140 ) | ( w5139 & w5140 ) ;
  assign w5142 = w5138 ^ w5140 ;
  assign w5143 = w5139 ^ w5142 ;
  assign w5144 = w5131 ^ w5137 ;
  assign w5145 = w5143 ^ w5144 ;
  assign w5146 = \pi34 & \pi36 ;
  assign w5147 = \pi33 & \pi37 ;
  assign w5148 = \pi32 & \pi38 ;
  assign w5149 = ( w5146 & w5147 ) | ( w5146 & w5148 ) | ( w5147 & w5148 ) ;
  assign w5150 = w5146 ^ w5148 ;
  assign w5151 = w5147 ^ w5150 ;
  assign w5152 = w4952 ^ w4974 ;
  assign w5153 = w5151 ^ w5152 ;
  assign w5154 = ( w5031 & w5032 ) | ( w5031 & w5033 ) | ( w5032 & w5033 ) ;
  assign w5155 = w5145 ^ w5154 ;
  assign w5156 = w5153 ^ w5155 ;
  assign w5157 = w5124 ^ w5125 ;
  assign w5158 = w5156 ^ w5157 ;
  assign w5159 = w5079 ^ w5086 ;
  assign w5160 = w5065 ^ w5159 ;
  assign w5161 = w5158 ^ w5160 ;
  assign w5162 = ( w5038 & w5043 ) | ( w5038 & w5050 ) | ( w5043 & w5050 ) ;
  assign w5163 = ( w5005 & w5006 ) | ( w5005 & w5022 ) | ( w5006 & w5022 ) ;
  assign w5164 = ( w5039 & w5040 ) | ( w5039 & w5041 ) | ( w5040 & w5041 ) ;
  assign w5165 = w4989 ^ w5011 ;
  assign w5166 = w5018 ^ w5165 ;
  assign w5167 = ( w4877 & w4889 ) | ( w4877 & w4921 ) | ( w4889 & w4921 ) ;
  assign w5168 = ( w4883 & w4907 ) | ( w4883 & w4927 ) | ( w4907 & w4927 ) ;
  assign w5169 = w5166 ^ w5168 ;
  assign w5170 = w5167 ^ w5169 ;
  assign w5171 = w5163 ^ w5164 ;
  assign w5172 = w5170 ^ w5171 ;
  assign w5173 = ( w4984 & w4985 ) | ( w4984 & w5023 ) | ( w4985 & w5023 ) ;
  assign w5174 = w5162 ^ w5172 ;
  assign w5175 = w5173 ^ w5174 ;
  assign w5176 = ( w4945 & w4946 ) | ( w4945 & w5025 ) | ( w4946 & w5025 ) ;
  assign w5177 = w5161 ^ w5176 ;
  assign w5178 = w5175 ^ w5177 ;
  assign w5179 = w5064 | w5178 ;
  assign w5180 = w5064 & w5178 ;
  assign w5181 = w5179 & ~w5180 ;
  assign w5182 = w5062 ^ w5181 ;
  assign w5183 = ( w5062 & w5179 ) | ( w5062 & w5180 ) | ( w5179 & w5180 ) ;
  assign w5184 = w5180 | w5183 ;
  assign w5185 = ( w5161 & w5175 ) | ( w5161 & w5176 ) | ( w5175 & w5176 ) ;
  assign w5186 = ( w5124 & w5125 ) | ( w5124 & w5156 ) | ( w5125 & w5156 ) ;
  assign w5187 = ( w4952 & w4974 ) | ( w4952 & w5151 ) | ( w4974 & w5151 ) ;
  assign w5188 = ( w4958 & w4995 ) | ( w4958 & w5001 ) | ( w4995 & w5001 ) ;
  assign w5189 = w5071 ^ w5187 ;
  assign w5190 = w5188 ^ w5189 ;
  assign w5191 = ( w5067 & w5076 ) | ( w5067 & w5077 ) | ( w5076 & w5077 ) ;
  assign w5192 = ( w5145 & w5153 ) | ( w5145 & w5154 ) | ( w5153 & w5154 ) ;
  assign w5193 = w5191 ^ w5192 ;
  assign w5194 = w5190 ^ w5193 ;
  assign w5195 = ( w4982 & w5079 ) | ( w4982 & w5085 ) | ( w5079 & w5085 ) ;
  assign w5196 = w5186 ^ w5194 ;
  assign w5197 = w5195 ^ w5196 ;
  assign w5198 = ( w5065 & w5158 ) | ( w5065 & w5159 ) | ( w5158 & w5159 ) ;
  assign w5199 = ( w5162 & w5172 ) | ( w5162 & w5173 ) | ( w5172 & w5173 ) ;
  assign w5200 = ( w5131 & w5137 ) | ( w5131 & w5143 ) | ( w5137 & w5143 ) ;
  assign w5201 = ( w4989 & w5011 ) | ( w4989 & w5018 ) | ( w5011 & w5018 ) ;
  assign w5202 = ( w5107 & w5113 ) | ( w5107 & w5119 ) | ( w5113 & w5119 ) ;
  assign w5203 = w5200 ^ w5201 ;
  assign w5204 = w5202 ^ w5203 ;
  assign w5205 = ( w5092 & w5098 ) | ( w5092 & w5099 ) | ( w5098 & w5099 ) ;
  assign w5206 = w5111 ^ w5129 ;
  assign w5207 = w5141 ^ w5206 ;
  assign w5208 = w5090 ^ w5096 ;
  assign w5209 = w5105 ^ w5208 ;
  assign w5210 = w5205 ^ w5207 ;
  assign w5211 = w5209 ^ w5210 ;
  assign w5212 = w5122 ^ w5211 ;
  assign w5213 = w5204 ^ w5212 ;
  assign w5214 = ( w5163 & w5164 ) | ( w5163 & w5170 ) | ( w5164 & w5170 ) ;
  assign w5215 = \pi22 & \pi49 ;
  assign w5216 = \pi09 & \pi62 ;
  assign w5217 = ( \pi36 & w5215 ) | ( \pi36 & w5216 ) | ( w5215 & w5216 ) ;
  assign w5218 = \pi36 ^ w5216 ;
  assign w5219 = w5215 ^ w5218 ;
  assign w5220 = \pi21 & \pi50 ;
  assign w5221 = \pi20 & \pi51 ;
  assign w5222 = \pi19 & \pi52 ;
  assign w5223 = ( w5220 & w5221 ) | ( w5220 & w5222 ) | ( w5221 & w5222 ) ;
  assign w5224 = w5220 ^ w5222 ;
  assign w5225 = w5221 ^ w5224 ;
  assign w5226 = \pi34 & \pi37 ;
  assign w5227 = \pi33 & \pi38 ;
  assign w5228 = ( w1779 & w5226 ) | ( w1779 & w5227 ) | ( w5226 & w5227 ) ;
  assign w5229 = w1779 ^ w5227 ;
  assign w5230 = w5226 ^ w5229 ;
  assign w5231 = w5219 ^ w5230 ;
  assign w5232 = w5225 ^ w5231 ;
  assign w5233 = \pi11 & \pi60 ;
  assign w5234 = \pi10 & \pi61 ;
  assign w5235 = \pi08 & \pi63 ;
  assign w5236 = ( w5233 & w5234 ) | ( w5233 & w5235 ) | ( w5234 & w5235 ) ;
  assign w5237 = w5233 ^ w5235 ;
  assign w5238 = w5234 ^ w5237 ;
  assign w5239 = w5135 ^ w5149 ;
  assign w5240 = w5238 ^ w5239 ;
  assign w5241 = ( w5166 & w5167 ) | ( w5166 & w5168 ) | ( w5167 & w5168 ) ;
  assign w5242 = w5232 ^ w5241 ;
  assign w5243 = w5240 ^ w5242 ;
  assign w5244 = ( w5080 & w5081 ) | ( w5080 & w5083 ) | ( w5081 & w5083 ) ;
  assign w5245 = \pi29 & \pi42 ;
  assign w5246 = \pi28 & \pi43 ;
  assign w5247 = \pi27 & \pi44 ;
  assign w5248 = ( w5245 & w5246 ) | ( w5245 & w5247 ) | ( w5246 & w5247 ) ;
  assign w5249 = w5245 ^ w5247 ;
  assign w5250 = w5246 ^ w5249 ;
  assign w5251 = \pi32 & \pi39 ;
  assign w5252 = \pi31 & \pi40 ;
  assign w5253 = \pi30 & \pi41 ;
  assign w5254 = ( w5251 & w5252 ) | ( w5251 & w5253 ) | ( w5252 & w5253 ) ;
  assign w5255 = w5251 ^ w5253 ;
  assign w5256 = w5252 ^ w5255 ;
  assign w5257 = \pi23 & \pi48 ;
  assign w5258 = \pi18 & \pi53 ;
  assign w5259 = \pi17 & \pi54 ;
  assign w5260 = ( w5257 & w5258 ) | ( w5257 & w5259 ) | ( w5258 & w5259 ) ;
  assign w5261 = w5257 ^ w5259 ;
  assign w5262 = w5258 ^ w5261 ;
  assign w5263 = w5250 ^ w5256 ;
  assign w5264 = w5262 ^ w5263 ;
  assign w5265 = \pi13 & \pi58 ;
  assign w5266 = ( \pi12 & \pi59 ) | ( \pi12 & ~w5117 ) | ( \pi59 & ~w5117 ) ;
  assign w5267 = w5265 ^ w5266 ;
  assign w5268 = w5117 & w5267 ;
  assign w5269 = \pi12 & \pi59 ;
  assign w5270 = w5117 ^ w5269 ;
  assign w5271 = w5265 ^ w5270 ;
  assign w5272 = \pi16 & \pi55 ;
  assign w5273 = \pi15 & \pi56 ;
  assign w5274 = \pi14 & \pi57 ;
  assign w5275 = ( w5272 & w5273 ) | ( w5272 & w5274 ) | ( w5273 & w5274 ) ;
  assign w5276 = w5272 ^ w5274 ;
  assign w5277 = w5273 ^ w5276 ;
  assign w5278 = \pi26 & \pi45 ;
  assign w5279 = \pi25 & \pi46 ;
  assign w5280 = \pi24 & \pi47 ;
  assign w5281 = ( w5278 & w5279 ) | ( w5278 & w5280 ) | ( w5279 & w5280 ) ;
  assign w5282 = w5278 ^ w5280 ;
  assign w5283 = w5279 ^ w5282 ;
  assign w5284 = w5271 ^ w5277 ;
  assign w5285 = w5283 ^ w5284 ;
  assign w5286 = w5244 ^ w5285 ;
  assign w5287 = w5264 ^ w5286 ;
  assign w5288 = w5214 ^ w5243 ;
  assign w5289 = w5287 ^ w5288 ;
  assign w5290 = w5199 ^ w5213 ;
  assign w5291 = w5289 ^ w5290 ;
  assign w5292 = w5198 ^ w5291 ;
  assign w5293 = w5197 ^ w5292 ;
  assign w5294 = w5184 ^ w5185 ;
  assign w5295 = w5293 ^ w5294 ;
  assign w5296 = ( w5184 & w5185 ) | ( w5184 & w5293 ) | ( w5185 & w5293 ) ;
  assign w5297 = ( w5214 & w5243 ) | ( w5214 & w5287 ) | ( w5243 & w5287 ) ;
  assign w5298 = ( w5205 & w5207 ) | ( w5205 & w5209 ) | ( w5207 & w5209 ) ;
  assign w5299 = ( w5135 & w5149 ) | ( w5135 & w5238 ) | ( w5149 & w5238 ) ;
  assign w5300 = \pi31 & \pi41 ;
  assign w5301 = \pi30 & \pi42 ;
  assign w5302 = \pi29 & \pi43 ;
  assign w5303 = ( w5300 & w5301 ) | ( w5300 & w5302 ) | ( w5301 & w5302 ) ;
  assign w5304 = w5300 ^ w5302 ;
  assign w5305 = w5301 ^ w5304 ;
  assign w5306 = ( w5090 & w5096 ) | ( w5090 & w5105 ) | ( w5096 & w5105 ) ;
  assign w5307 = w5299 ^ w5306 ;
  assign w5308 = w5305 ^ w5307 ;
  assign w5309 = ( w5232 & w5240 ) | ( w5232 & w5241 ) | ( w5240 & w5241 ) ;
  assign w5310 = w5298 ^ w5309 ;
  assign w5311 = w5308 ^ w5310 ;
  assign w5312 = ( w5122 & w5204 ) | ( w5122 & w5211 ) | ( w5204 & w5211 ) ;
  assign w5313 = w5297 ^ w5311 ;
  assign w5314 = w5312 ^ w5313 ;
  assign w5315 = ( w5199 & w5213 ) | ( w5199 & w5289 ) | ( w5213 & w5289 ) ;
  assign w5316 = ( w5186 & w5194 ) | ( w5186 & w5195 ) | ( w5194 & w5195 ) ;
  assign w5317 = ( w5250 & w5256 ) | ( w5250 & w5262 ) | ( w5256 & w5262 ) ;
  assign w5318 = ( w5111 & w5129 ) | ( w5111 & w5141 ) | ( w5129 & w5141 ) ;
  assign w5319 = ( w5219 & w5225 ) | ( w5219 & w5230 ) | ( w5225 & w5230 ) ;
  assign w5320 = w5317 ^ w5319 ;
  assign w5321 = w5318 ^ w5320 ;
  assign w5322 = ( w5244 & w5264 ) | ( w5244 & w5285 ) | ( w5264 & w5285 ) ;
  assign w5323 = ( w5271 & w5277 ) | ( w5271 & w5283 ) | ( w5277 & w5283 ) ;
  assign w5324 = w5248 ^ w5254 ;
  assign w5325 = w5260 ^ w5324 ;
  assign w5326 = w5217 ^ w5228 ;
  assign w5327 = w5223 ^ w5326 ;
  assign w5328 = w5323 ^ w5327 ;
  assign w5329 = w5325 ^ w5328 ;
  assign w5330 = w5321 ^ w5322 ;
  assign w5331 = w5329 ^ w5330 ;
  assign w5332 = ( w5200 & w5201 ) | ( w5200 & w5202 ) | ( w5201 & w5202 ) ;
  assign w5333 = \pi32 & \pi40 ;
  assign w5334 = \pi23 & \pi49 ;
  assign w5335 = \pi16 & \pi56 ;
  assign w5336 = ( w5333 & w5334 ) | ( w5333 & w5335 ) | ( w5334 & w5335 ) ;
  assign w5337 = w5333 ^ w5335 ;
  assign w5338 = w5334 ^ w5337 ;
  assign w5339 = \pi22 & \pi50 ;
  assign w5340 = \pi21 & \pi51 ;
  assign w5341 = ( w2323 & w5339 ) | ( w2323 & w5340 ) | ( w5339 & w5340 ) ;
  assign w5342 = w2323 ^ w5340 ;
  assign w5343 = w5339 ^ w5342 ;
  assign w5344 = \pi20 & \pi52 ;
  assign w5345 = \pi18 & \pi54 ;
  assign w5346 = \pi17 & \pi55 ;
  assign w5347 = ( w5344 & w5345 ) | ( w5344 & w5346 ) | ( w5345 & w5346 ) ;
  assign w5348 = w5344 ^ w5346 ;
  assign w5349 = w5345 ^ w5348 ;
  assign w5350 = w5338 ^ w5343 ;
  assign w5351 = w5349 ^ w5350 ;
  assign w5352 = \pi11 & \pi61 ;
  assign w5353 = \pi10 & \pi62 ;
  assign w5354 = \pi09 & \pi63 ;
  assign w5355 = ( w5352 & w5353 ) | ( w5352 & w5354 ) | ( w5353 & w5354 ) ;
  assign w5356 = w5352 ^ w5354 ;
  assign w5357 = w5353 ^ w5356 ;
  assign w5358 = \pi25 & \pi47 ;
  assign w5359 = \pi24 & \pi48 ;
  assign w5360 = \pi12 & \pi60 ;
  assign w5361 = ( w5358 & w5359 ) | ( w5358 & w5360 ) | ( w5359 & w5360 ) ;
  assign w5362 = w5358 ^ w5360 ;
  assign w5363 = w5359 ^ w5362 ;
  assign w5364 = w5357 ^ w5363 ;
  assign w5365 = w4068 | w5268 ;
  assign w5366 = ( w342 & w5268 ) | ( w342 & w5365 ) | ( w5268 & w5365 ) ;
  assign w5367 = w5364 ^ w5366 ;
  assign w5368 = w5332 ^ w5351 ;
  assign w5369 = w5367 ^ w5368 ;
  assign w5370 = ( w5190 & w5191 ) | ( w5190 & w5192 ) | ( w5191 & w5192 ) ;
  assign w5371 = w5236 ^ w5275 ;
  assign w5372 = w5281 ^ w5371 ;
  assign w5373 = ( w5071 & w5187 ) | ( w5071 & w5188 ) | ( w5187 & w5188 ) ;
  assign w5374 = \pi15 & \pi57 ;
  assign w5375 = \pi14 & \pi58 ;
  assign w5376 = \pi13 & \pi59 ;
  assign w5377 = ( w5374 & w5375 ) | ( w5374 & w5376 ) | ( w5375 & w5376 ) ;
  assign w5378 = w5374 ^ w5376 ;
  assign w5379 = w5375 ^ w5378 ;
  assign w5380 = \pi28 & \pi44 ;
  assign w5381 = \pi27 & \pi45 ;
  assign w5382 = \pi26 & \pi46 ;
  assign w5383 = ( w5380 & w5381 ) | ( w5380 & w5382 ) | ( w5381 & w5382 ) ;
  assign w5384 = w5380 ^ w5382 ;
  assign w5385 = w5381 ^ w5384 ;
  assign w5386 = \pi34 & \pi38 ;
  assign w5387 = \pi33 & \pi39 ;
  assign w5388 = \pi19 & \pi53 ;
  assign w5389 = ( w5386 & w5387 ) | ( w5386 & w5388 ) | ( w5387 & w5388 ) ;
  assign w5390 = w5386 ^ w5388 ;
  assign w5391 = w5387 ^ w5390 ;
  assign w5392 = w5379 ^ w5385 ;
  assign w5393 = w5391 ^ w5392 ;
  assign w5394 = w5372 ^ w5373 ;
  assign w5395 = w5393 ^ w5394 ;
  assign w5396 = w5369 ^ w5370 ;
  assign w5397 = w5395 ^ w5396 ;
  assign w5398 = w5316 ^ w5397 ;
  assign w5399 = w5331 ^ w5398 ;
  assign w5400 = w5315 ^ w5399 ;
  assign w5401 = w5314 ^ w5400 ;
  assign w5402 = ( w5197 & w5198 ) | ( w5197 & w5291 ) | ( w5198 & w5291 ) ;
  assign w5403 = w5401 | w5402 ;
  assign w5404 = w5401 & w5402 ;
  assign w5405 = w5403 & ~w5404 ;
  assign w5406 = w5296 ^ w5405 ;
  assign w5407 = ( w5296 & w5403 ) | ( w5296 & w5404 ) | ( w5403 & w5404 ) ;
  assign w5408 = w5404 | w5407 ;
  assign w5409 = ( w5314 & w5315 ) | ( w5314 & w5399 ) | ( w5315 & w5399 ) ;
  assign w5410 = ( w5316 & w5331 ) | ( w5316 & w5397 ) | ( w5331 & w5397 ) ;
  assign w5411 = ( w5369 & w5370 ) | ( w5369 & w5395 ) | ( w5370 & w5395 ) ;
  assign w5412 = ( w5321 & w5322 ) | ( w5321 & w5329 ) | ( w5322 & w5329 ) ;
  assign w5413 = ( w5372 & w5373 ) | ( w5372 & w5393 ) | ( w5373 & w5393 ) ;
  assign w5414 = ( w5236 & w5275 ) | ( w5236 & w5281 ) | ( w5275 & w5281 ) ;
  assign w5415 = \pi33 & \pi40 ;
  assign w5416 = \pi32 & \pi41 ;
  assign w5417 = \pi31 & \pi42 ;
  assign w5418 = ( w5415 & w5416 ) | ( w5415 & w5417 ) | ( w5416 & w5417 ) ;
  assign w5419 = w5415 ^ w5417 ;
  assign w5420 = w5416 ^ w5419 ;
  assign w5421 = ( w5248 & w5254 ) | ( w5248 & w5260 ) | ( w5254 & w5260 ) ;
  assign w5422 = w5414 ^ w5421 ;
  assign w5423 = w5420 ^ w5422 ;
  assign w5424 = ( w5323 & w5325 ) | ( w5323 & w5327 ) | ( w5325 & w5327 ) ;
  assign w5425 = w5413 ^ w5424 ;
  assign w5426 = w5423 ^ w5425 ;
  assign w5427 = w5411 ^ w5412 ;
  assign w5428 = w5426 ^ w5427 ;
  assign w5429 = ( w5297 & w5311 ) | ( w5297 & w5312 ) | ( w5311 & w5312 ) ;
  assign w5430 = w342 & w4068 ;
  assign w5431 = w5268 | w5430 ;
  assign w5432 = ( w5357 & w5363 ) | ( w5357 & w5431 ) | ( w5363 & w5431 ) ;
  assign w5433 = ( w5217 & w5223 ) | ( w5217 & w5228 ) | ( w5223 & w5228 ) ;
  assign w5434 = ( w5379 & w5385 ) | ( w5379 & w5391 ) | ( w5385 & w5391 ) ;
  assign w5435 = w5432 ^ w5433 ;
  assign w5436 = w5434 ^ w5435 ;
  assign w5437 = ( w5332 & w5351 ) | ( w5332 & w5367 ) | ( w5351 & w5367 ) ;
  assign w5438 = ( w5338 & w5343 ) | ( w5338 & w5349 ) | ( w5343 & w5349 ) ;
  assign w5439 = w5347 ^ w5355 ;
  assign w5440 = w5361 ^ w5439 ;
  assign w5441 = w5341 ^ w5438 ;
  assign w5442 = w5440 ^ w5441 ;
  assign w5443 = w5389 ^ w5442 ;
  assign w5444 = \pi13 & \pi60 ;
  assign w5445 = w5443 ^ w5444 ;
  assign w5446 = w5436 ^ w5437 ;
  assign w5447 = w5445 ^ w5446 ;
  assign w5448 = \pi23 & \pi50 ;
  assign w5449 = \pi11 & \pi62 ;
  assign w5450 = ( \pi37 & w5448 ) | ( \pi37 & w5449 ) | ( w5448 & w5449 ) ;
  assign w5451 = \pi37 ^ w5449 ;
  assign w5452 = w5448 ^ w5451 ;
  assign w5453 = \pi19 & \pi54 ;
  assign w5454 = \pi18 & \pi55 ;
  assign w5455 = ( w2919 & w5453 ) | ( w2919 & w5454 ) | ( w5453 & w5454 ) ;
  assign w5456 = w2919 ^ w5454 ;
  assign w5457 = w5453 ^ w5456 ;
  assign w5458 = \pi22 & \pi51 ;
  assign w5459 = \pi21 & \pi52 ;
  assign w5460 = \pi20 & \pi53 ;
  assign w5461 = ( w5458 & w5459 ) | ( w5458 & w5460 ) | ( w5459 & w5460 ) ;
  assign w5462 = w5458 ^ w5460 ;
  assign w5463 = w5459 ^ w5462 ;
  assign w5464 = w5452 ^ w5457 ;
  assign w5465 = w5463 ^ w5464 ;
  assign w5466 = \pi16 & \pi57 ;
  assign w5467 = \pi15 & \pi58 ;
  assign w5468 = \pi14 & \pi59 ;
  assign w5469 = ( w5466 & w5467 ) | ( w5466 & w5468 ) | ( w5467 & w5468 ) ;
  assign w5470 = w5466 ^ w5468 ;
  assign w5471 = w5467 ^ w5470 ;
  assign w5472 = \pi27 & \pi46 ;
  assign w5473 = \pi26 & \pi47 ;
  assign w5474 = \pi17 & \pi56 ;
  assign w5475 = ( w5472 & w5473 ) | ( w5472 & w5474 ) | ( w5473 & w5474 ) ;
  assign w5476 = w5472 ^ w5474 ;
  assign w5477 = w5473 ^ w5476 ;
  assign w5478 = w5336 ^ w5471 ;
  assign w5479 = w5477 ^ w5478 ;
  assign w5480 = ( w5317 & w5318 ) | ( w5317 & w5319 ) | ( w5318 & w5319 ) ;
  assign w5481 = w5465 ^ w5480 ;
  assign w5482 = w5479 ^ w5481 ;
  assign w5483 = ( w5298 & w5308 ) | ( w5298 & w5309 ) | ( w5308 & w5309 ) ;
  assign w5484 = w5303 ^ w5377 ;
  assign w5485 = w5383 ^ w5484 ;
  assign w5486 = ( w5299 & w5305 ) | ( w5299 & w5306 ) | ( w5305 & w5306 ) ;
  assign w5487 = \pi25 & \pi48 ;
  assign w5488 = \pi12 & \pi61 ;
  assign w5489 = \pi10 & \pi63 ;
  assign w5490 = ( w5487 & w5488 ) | ( w5487 & w5489 ) | ( w5488 & w5489 ) ;
  assign w5491 = w5487 ^ w5489 ;
  assign w5492 = w5488 ^ w5491 ;
  assign w5493 = \pi30 & \pi43 ;
  assign w5494 = \pi29 & \pi44 ;
  assign w5495 = \pi28 & \pi45 ;
  assign w5496 = ( w5493 & w5494 ) | ( w5493 & w5495 ) | ( w5494 & w5495 ) ;
  assign w5497 = w5493 ^ w5495 ;
  assign w5498 = w5494 ^ w5497 ;
  assign w5499 = \pi36 & \pi37 ;
  assign w5500 = \pi35 & \pi38 ;
  assign w5501 = \pi34 & \pi39 ;
  assign w5502 = ( w5499 & w5500 ) | ( w5499 & w5501 ) | ( w5500 & w5501 ) ;
  assign w5503 = w5499 ^ w5501 ;
  assign w5504 = w5500 ^ w5503 ;
  assign w5505 = w5492 ^ w5498 ;
  assign w5506 = w5504 ^ w5505 ;
  assign w5507 = w5485 ^ w5486 ;
  assign w5508 = w5506 ^ w5507 ;
  assign w5509 = w5482 ^ w5483 ;
  assign w5510 = w5508 ^ w5509 ;
  assign w5511 = w5429 ^ w5510 ;
  assign w5512 = w5447 ^ w5511 ;
  assign w5513 = w5410 ^ w5428 ;
  assign w5514 = w5512 ^ w5513 ;
  assign w5515 = w5408 ^ w5409 ;
  assign w5516 = w5514 ^ w5515 ;
  assign w5517 = ( w5410 & w5428 ) | ( w5410 & w5512 ) | ( w5428 & w5512 ) ;
  assign w5518 = ( w5411 & w5412 ) | ( w5411 & w5426 ) | ( w5412 & w5426 ) ;
  assign w5519 = \pi16 & \pi58 ;
  assign w5520 = \pi15 & \pi59 ;
  assign w5521 = \pi14 & \pi60 ;
  assign w5522 = ( w5519 & w5520 ) | ( w5519 & w5521 ) | ( w5520 & w5521 ) ;
  assign w5523 = w5519 ^ w5521 ;
  assign w5524 = w5520 ^ w5523 ;
  assign w5525 = w5418 ^ w5502 ;
  assign w5526 = w5524 ^ w5525 ;
  assign w5527 = ( w5452 & w5457 ) | ( w5452 & w5463 ) | ( w5457 & w5463 ) ;
  assign w5528 = ( w5414 & w5420 ) | ( w5414 & w5421 ) | ( w5420 & w5421 ) ;
  assign w5529 = w5526 ^ w5528 ;
  assign w5530 = w5527 ^ w5529 ;
  assign w5531 = ( w5465 & w5479 ) | ( w5465 & w5480 ) | ( w5479 & w5480 ) ;
  assign w5532 = ( w5485 & w5486 ) | ( w5485 & w5506 ) | ( w5486 & w5506 ) ;
  assign w5533 = w5531 ^ w5532 ;
  assign w5534 = w5530 & w5533 ;
  assign w5535 = w5530 | w5533 ;
  assign w5536 = \pi13 & \pi61 ;
  assign w5537 = ( \pi12 & \pi62 ) | ( \pi12 & ~w5450 ) | ( \pi62 & ~w5450 ) ;
  assign w5538 = w5536 ^ w5537 ;
  assign w5539 = w5450 & w5538 ;
  assign w5540 = \pi12 & \pi62 ;
  assign w5541 = w5450 ^ w5540 ;
  assign w5542 = w5536 ^ w5541 ;
  assign w5543 = \pi30 & \pi44 ;
  assign w5544 = \pi29 & \pi45 ;
  assign w5545 = \pi17 & \pi57 ;
  assign w5546 = ( w5543 & w5544 ) | ( w5543 & w5545 ) | ( w5544 & w5545 ) ;
  assign w5547 = w5543 ^ w5545 ;
  assign w5548 = w5544 ^ w5547 ;
  assign w5549 = ( w5303 & w5377 ) | ( w5303 & w5383 ) | ( w5377 & w5383 ) ;
  assign w5550 = w5542 ^ w5549 ;
  assign w5551 = w5548 ^ w5550 ;
  assign w5552 = \pi32 & \pi42 ;
  assign w5553 = \pi31 & \pi43 ;
  assign w5554 = \pi11 & \pi63 ;
  assign w5555 = ( w5552 & w5553 ) | ( w5552 & w5554 ) | ( w5553 & w5554 ) ;
  assign w5556 = w5552 ^ w5554 ;
  assign w5557 = w5553 ^ w5556 ;
  assign w5558 = \pi25 & \pi49 ;
  assign w5559 = \pi18 & \pi56 ;
  assign w5560 = ( w2459 & w5558 ) | ( w2459 & w5559 ) | ( w5558 & w5559 ) ;
  assign w5561 = w2459 ^ w5559 ;
  assign w5562 = w5558 ^ w5561 ;
  assign w5563 = \pi28 & \pi46 ;
  assign w5564 = \pi27 & \pi47 ;
  assign w5565 = \pi26 & \pi48 ;
  assign w5566 = ( w5563 & w5564 ) | ( w5563 & w5565 ) | ( w5564 & w5565 ) ;
  assign w5567 = w5563 ^ w5565 ;
  assign w5568 = w5564 ^ w5567 ;
  assign w5569 = w5557 ^ w5562 ;
  assign w5570 = w5568 ^ w5569 ;
  assign w5571 = \pi22 & \pi52 ;
  assign w5572 = \pi21 & \pi53 ;
  assign w5573 = \pi19 & \pi55 ;
  assign w5574 = ( w5571 & w5572 ) | ( w5571 & w5573 ) | ( w5572 & w5573 ) ;
  assign w5575 = w5571 ^ w5573 ;
  assign w5576 = w5572 ^ w5575 ;
  assign w5577 = \pi35 & \pi39 ;
  assign w5578 = \pi34 & \pi40 ;
  assign w5579 = ( w4970 & w5577 ) | ( w4970 & w5578 ) | ( w5577 & w5578 ) ;
  assign w5580 = w4970 ^ w5578 ;
  assign w5581 = w5577 ^ w5580 ;
  assign w5582 = \pi24 & \pi50 ;
  assign w5583 = \pi23 & \pi51 ;
  assign w5584 = ( w1636 & w5582 ) | ( w1636 & w5583 ) | ( w5582 & w5583 ) ;
  assign w5585 = w1636 ^ w5583 ;
  assign w5586 = w5582 ^ w5585 ;
  assign w5587 = w5581 ^ w5586 ;
  assign w5588 = w5576 ^ w5587 ;
  assign w5589 = w5551 ^ w5570 ;
  assign w5590 = w5588 ^ w5589 ;
  assign w5591 = ( w5413 & w5423 ) | ( w5413 & w5424 ) | ( w5423 & w5424 ) ;
  assign w5592 = w5469 ^ w5475 ;
  assign w5593 = w5496 ^ w5592 ;
  assign w5594 = w5455 ^ w5461 ;
  assign w5595 = w5490 ^ w5594 ;
  assign w5596 = ( w5492 & w5498 ) | ( w5492 & w5504 ) | ( w5498 & w5504 ) ;
  assign w5597 = w5593 ^ w5595 ;
  assign w5598 = w5596 ^ w5597 ;
  assign w5599 = w5590 ^ w5591 ;
  assign w5600 = w5598 ^ w5599 ;
  assign w5601 = ~w5534 & w5535 ;
  assign w5602 = w5600 ^ w5601 ;
  assign w5603 = w5518 ^ w5602 ;
  assign w5604 = ( w5429 & w5447 ) | ( w5429 & w5510 ) | ( w5447 & w5510 ) ;
  assign w5605 = ( w5482 & w5483 ) | ( w5482 & w5508 ) | ( w5483 & w5508 ) ;
  assign w5606 = ( w5436 & w5437 ) | ( w5436 & w5445 ) | ( w5437 & w5445 ) ;
  assign w5607 = ( w5347 & w5355 ) | ( w5347 & w5361 ) | ( w5355 & w5361 ) ;
  assign w5608 = ( w5336 & w5471 ) | ( w5336 & w5477 ) | ( w5471 & w5477 ) ;
  assign w5609 = ( w5341 & w5389 ) | ( w5341 & w5444 ) | ( w5389 & w5444 ) ;
  assign w5610 = w5607 ^ w5609 ;
  assign w5611 = w5608 ^ w5610 ;
  assign w5612 = w5341 ^ w5389 ;
  assign w5613 = w5444 ^ w5612 ;
  assign w5614 = ( w5438 & w5440 ) | ( w5438 & w5613 ) | ( w5440 & w5613 ) ;
  assign w5615 = ( w5432 & w5433 ) | ( w5432 & w5434 ) | ( w5433 & w5434 ) ;
  assign w5616 = w5614 ^ w5615 ;
  assign w5617 = w5611 ^ w5616 ;
  assign w5618 = w5605 ^ w5606 ;
  assign w5619 = w5617 ^ w5618 ;
  assign w5620 = w5603 ^ w5604 ;
  assign w5621 = w5619 ^ w5620 ;
  assign w5622 = ( w5408 & w5409 ) | ( w5408 & w5514 ) | ( w5409 & w5514 ) ;
  assign w5623 = w5621 ^ w5622 ;
  assign w5624 = w5517 ^ w5623 ;
  assign w5625 = ( w5603 & w5604 ) | ( w5603 & w5619 ) | ( w5604 & w5619 ) ;
  assign w5626 = ( w5605 & w5606 ) | ( w5605 & w5617 ) | ( w5606 & w5617 ) ;
  assign w5627 = ( w5418 & w5502 ) | ( w5418 & w5524 ) | ( w5502 & w5524 ) ;
  assign w5628 = ( w5455 & w5461 ) | ( w5455 & w5490 ) | ( w5461 & w5490 ) ;
  assign w5629 = ( w5469 & w5475 ) | ( w5469 & w5496 ) | ( w5475 & w5496 ) ;
  assign w5630 = w5627 ^ w5628 ;
  assign w5631 = w5629 ^ w5630 ;
  assign w5632 = ( w5551 & w5570 ) | ( w5551 & w5588 ) | ( w5570 & w5588 ) ;
  assign w5633 = ( w5542 & w5548 ) | ( w5542 & w5549 ) | ( w5548 & w5549 ) ;
  assign w5634 = w5579 ^ w5584 ;
  assign w5635 = w5574 ^ w5634 ;
  assign w5636 = w5555 ^ w5560 ;
  assign w5637 = w342 | w5539 ;
  assign w5638 = ( w4390 & w5539 ) | ( w4390 & w5637 ) | ( w5539 & w5637 ) ;
  assign w5639 = w5636 ^ w5638 ;
  assign w5640 = w5633 ^ w5635 ;
  assign w5641 = w5639 ^ w5640 ;
  assign w5642 = w5632 ^ w5641 ;
  assign w5643 = w5631 ^ w5642 ;
  assign w5644 = \pi30 & \pi45 ;
  assign w5645 = \pi19 & \pi56 ;
  assign w5646 = \pi12 & \pi63 ;
  assign w5647 = ( w5644 & w5645 ) | ( w5644 & w5646 ) | ( w5645 & w5646 ) ;
  assign w5648 = w5644 ^ w5646 ;
  assign w5649 = w5645 ^ w5648 ;
  assign w5650 = \pi36 & \pi39 ;
  assign w5651 = \pi35 & \pi40 ;
  assign w5652 = \pi23 & \pi52 ;
  assign w5653 = ( w5650 & w5651 ) | ( w5650 & w5652 ) | ( w5651 & w5652 ) ;
  assign w5654 = w5650 ^ w5652 ;
  assign w5655 = w5651 ^ w5654 ;
  assign w5656 = w5649 ^ w5655 ;
  assign w5657 = ~\pi37 & \pi38 ;
  assign w5658 = \pi13 & \pi62 ;
  assign w5659 = w5656 ^ w5658 ;
  assign w5660 = w5657 ^ w5659 ;
  assign w5661 = ( w5607 & w5608 ) | ( w5607 & w5609 ) | ( w5608 & w5609 ) ;
  assign w5662 = w5660 ^ w5661 ;
  assign w5663 = \pi16 & \pi59 ;
  assign w5664 = \pi15 & \pi60 ;
  assign w5665 = \pi14 & \pi61 ;
  assign w5666 = ( w5663 & w5664 ) | ( w5663 & w5665 ) | ( w5664 & w5665 ) ;
  assign w5667 = w5663 ^ w5665 ;
  assign w5668 = w5664 ^ w5667 ;
  assign w5669 = \pi26 & \pi49 ;
  assign w5670 = \pi18 & \pi57 ;
  assign w5671 = \pi17 & \pi58 ;
  assign w5672 = ( w5669 & w5670 ) | ( w5669 & w5671 ) | ( w5670 & w5671 ) ;
  assign w5673 = w5669 ^ w5671 ;
  assign w5674 = w5670 ^ w5673 ;
  assign w5675 = \pi29 & \pi46 ;
  assign w5676 = \pi28 & \pi47 ;
  assign w5677 = \pi27 & \pi48 ;
  assign w5678 = ( w5675 & w5676 ) | ( w5675 & w5677 ) | ( w5676 & w5677 ) ;
  assign w5679 = w5675 ^ w5677 ;
  assign w5680 = w5676 ^ w5679 ;
  assign w5681 = w5668 ^ w5674 ;
  assign w5682 = w5680 ^ w5681 ;
  assign w5683 = ( w5611 & w5614 ) | ( w5611 & w5615 ) | ( w5614 & w5615 ) ;
  assign w5684 = w5522 ^ w5546 ;
  assign w5685 = w5566 ^ w5684 ;
  assign w5686 = ( w5576 & w5581 ) | ( w5576 & w5586 ) | ( w5581 & w5586 ) ;
  assign w5687 = ( w5557 & w5562 ) | ( w5557 & w5568 ) | ( w5562 & w5568 ) ;
  assign w5688 = w5686 ^ w5687 ;
  assign w5689 = w5685 ^ w5688 ;
  assign w5690 = w5682 ^ w5689 ;
  assign w5691 = w5683 ^ w5690 ;
  assign w5692 = w5662 ^ w5691 ;
  assign w5693 = w5626 ^ w5692 ;
  assign w5694 = w5643 ^ w5693 ;
  assign w5695 = ( w5526 & w5527 ) | ( w5526 & w5528 ) | ( w5527 & w5528 ) ;
  assign w5696 = \pi34 & \pi41 ;
  assign w5697 = \pi25 & \pi50 ;
  assign w5698 = \pi20 & \pi55 ;
  assign w5699 = ( w5696 & w5697 ) | ( w5696 & w5698 ) | ( w5697 & w5698 ) ;
  assign w5700 = w5696 ^ w5698 ;
  assign w5701 = w5697 ^ w5700 ;
  assign w5702 = \pi33 & \pi42 ;
  assign w5703 = \pi32 & \pi43 ;
  assign w5704 = \pi31 & \pi44 ;
  assign w5705 = ( w5702 & w5703 ) | ( w5702 & w5704 ) | ( w5703 & w5704 ) ;
  assign w5706 = w5702 ^ w5704 ;
  assign w5707 = w5703 ^ w5706 ;
  assign w5708 = \pi24 & \pi51 ;
  assign w5709 = \pi22 & \pi53 ;
  assign w5710 = \pi21 & \pi54 ;
  assign w5711 = ( w5708 & w5709 ) | ( w5708 & w5710 ) | ( w5709 & w5710 ) ;
  assign w5712 = w5708 ^ w5710 ;
  assign w5713 = w5709 ^ w5712 ;
  assign w5714 = w5701 ^ w5707 ;
  assign w5715 = w5713 ^ w5714 ;
  assign w5716 = ( w5593 & w5595 ) | ( w5593 & w5596 ) | ( w5595 & w5596 ) ;
  assign w5717 = w5695 ^ w5716 ;
  assign w5718 = w5715 ^ w5717 ;
  assign w5719 = ( w5530 & w5531 ) | ( w5530 & w5532 ) | ( w5531 & w5532 ) ;
  assign w5720 = ( w5590 & w5591 ) | ( w5590 & w5598 ) | ( w5591 & w5598 ) ;
  assign w5721 = w5719 ^ w5720 ;
  assign w5722 = w5718 ^ w5721 ;
  assign w5723 = ( w5518 & w5600 ) | ( w5518 & w5601 ) | ( w5600 & w5601 ) ;
  assign w5724 = w5694 ^ w5723 ;
  assign w5725 = w5722 ^ w5724 ;
  assign w5726 = ( w5517 & w5621 ) | ( w5517 & w5622 ) | ( w5621 & w5622 ) ;
  assign w5727 = w5625 ^ w5726 ;
  assign w5728 = w5725 ^ w5727 ;
  assign w5729 = ( w5625 & w5725 ) | ( w5625 & w5726 ) | ( w5725 & w5726 ) ;
  assign w5730 = ( w5694 & w5722 ) | ( w5694 & w5723 ) | ( w5722 & w5723 ) ;
  assign w5731 = w342 & w4390 ;
  assign w5732 = w5539 | w5731 ;
  assign w5733 = ( w5555 & w5560 ) | ( w5555 & w5732 ) | ( w5560 & w5732 ) ;
  assign w5734 = ( w5522 & w5546 ) | ( w5522 & w5566 ) | ( w5546 & w5566 ) ;
  assign w5735 = ( w5574 & w5579 ) | ( w5574 & w5584 ) | ( w5579 & w5584 ) ;
  assign w5736 = w5733 ^ w5735 ;
  assign w5737 = w5734 ^ w5736 ;
  assign w5738 = ( w5660 & w5661 ) | ( w5660 & w5682 ) | ( w5661 & w5682 ) ;
  assign w5739 = w5647 ^ w5678 ;
  assign w5740 = w5699 ^ w5739 ;
  assign w5741 = ( w5701 & w5707 ) | ( w5701 & w5713 ) | ( w5707 & w5713 ) ;
  assign w5742 = \pi37 & \pi38 ;
  assign w5743 = w5653 & w5742 ;
  assign w5744 = ( \pi13 & \pi38 ) | ( \pi13 & w5742 ) | ( \pi38 & w5742 ) ;
  assign w5745 = ( \pi14 & w5653 ) | ( \pi14 & w5744 ) | ( w5653 & w5744 ) ;
  assign w5746 = ( \pi62 & w5743 ) | ( \pi62 & w5745 ) | ( w5743 & w5745 ) ;
  assign w5747 = \pi14 & \pi62 ;
  assign w5748 = w5653 ^ w5747 ;
  assign w5749 = \pi13 & ~\pi37 ;
  assign w5750 = \pi62 & w5749 ;
  assign w5751 = ( \pi37 & \pi38 ) | ( \pi37 & w5750 ) | ( \pi38 & w5750 ) ;
  assign w5752 = w5748 ^ w5751 ;
  assign w5753 = w5740 ^ w5741 ;
  assign w5754 = w5752 ^ w5753 ;
  assign w5755 = w5737 ^ w5738 ;
  assign w5756 = w5754 ^ w5755 ;
  assign w5757 = ( w5718 & w5719 ) | ( w5718 & w5720 ) | ( w5719 & w5720 ) ;
  assign w5758 = w5756 ^ w5757 ;
  assign w5759 = ( w5695 & w5715 ) | ( w5695 & w5716 ) | ( w5715 & w5716 ) ;
  assign w5760 = w5666 ^ w5672 ;
  assign w5761 = w5705 ^ w5760 ;
  assign w5762 = ( w5668 & w5674 ) | ( w5668 & w5680 ) | ( w5674 & w5680 ) ;
  assign w5763 = w5657 ^ w5658 ;
  assign w5764 = ( w5649 & w5655 ) | ( w5649 & w5763 ) | ( w5655 & w5763 ) ;
  assign w5765 = w5761 ^ w5762 ;
  assign w5766 = w5764 ^ w5765 ;
  assign w5767 = \pi30 & \pi46 ;
  assign w5768 = \pi29 & \pi47 ;
  assign w5769 = \pi28 & \pi48 ;
  assign w5770 = ( w5767 & w5768 ) | ( w5767 & w5769 ) | ( w5768 & w5769 ) ;
  assign w5771 = w5767 ^ w5769 ;
  assign w5772 = w5768 ^ w5771 ;
  assign w5773 = \pi36 & \pi40 ;
  assign w5774 = \pi35 & \pi41 ;
  assign w5775 = \pi34 & \pi42 ;
  assign w5776 = ( w5773 & w5774 ) | ( w5773 & w5775 ) | ( w5774 & w5775 ) ;
  assign w5777 = w5773 ^ w5775 ;
  assign w5778 = w5774 ^ w5777 ;
  assign w5779 = \pi25 & \pi51 ;
  assign w5780 = \pi24 & \pi52 ;
  assign w5781 = ( w2494 & w5779 ) | ( w2494 & w5780 ) | ( w5779 & w5780 ) ;
  assign w5782 = w2494 ^ w5780 ;
  assign w5783 = w5779 ^ w5782 ;
  assign w5784 = w5772 ^ w5783 ;
  assign w5785 = w5778 ^ w5784 ;
  assign w5786 = ( w5627 & w5628 ) | ( w5627 & w5629 ) | ( w5628 & w5629 ) ;
  assign w5787 = w5785 ^ w5786 ;
  assign w5788 = \pi17 & \pi59 ;
  assign w5789 = \pi16 & \pi60 ;
  assign w5790 = \pi15 & \pi61 ;
  assign w5791 = ( w5788 & w5789 ) | ( w5788 & w5790 ) | ( w5789 & w5790 ) ;
  assign w5792 = w5788 ^ w5790 ;
  assign w5793 = w5789 ^ w5792 ;
  assign w5794 = \pi27 & \pi49 ;
  assign w5795 = \pi26 & \pi50 ;
  assign w5796 = \pi18 & \pi58 ;
  assign w5797 = ( w5794 & w5795 ) | ( w5794 & w5796 ) | ( w5795 & w5796 ) ;
  assign w5798 = w5794 ^ w5796 ;
  assign w5799 = w5795 ^ w5798 ;
  assign w5800 = w5711 ^ w5793 ;
  assign w5801 = w5799 ^ w5800 ;
  assign w5802 = w5766 ^ w5801 ;
  assign w5803 = w5759 ^ w5802 ;
  assign w5804 = w5787 ^ w5803 ;
  assign w5805 = ( w5626 & w5643 ) | ( w5626 & w5692 ) | ( w5643 & w5692 ) ;
  assign w5806 = w5662 ^ w5682 ;
  assign w5807 = ( w5683 & w5689 ) | ( w5683 & w5806 ) | ( w5689 & w5806 ) ;
  assign w5808 = ( w5631 & w5632 ) | ( w5631 & w5641 ) | ( w5632 & w5641 ) ;
  assign w5809 = ( w5633 & w5635 ) | ( w5633 & w5639 ) | ( w5635 & w5639 ) ;
  assign w5810 = \pi32 & \pi44 ;
  assign w5811 = \pi31 & \pi45 ;
  assign w5812 = \pi13 & \pi63 ;
  assign w5813 = ( w5810 & w5811 ) | ( w5810 & w5812 ) | ( w5811 & w5812 ) ;
  assign w5814 = w5810 ^ w5812 ;
  assign w5815 = w5811 ^ w5814 ;
  assign w5816 = \pi23 & \pi53 ;
  assign w5817 = \pi19 & \pi57 ;
  assign w5818 = ( w2504 & w5816 ) | ( w2504 & w5817 ) | ( w5816 & w5817 ) ;
  assign w5819 = w2504 ^ w5817 ;
  assign w5820 = w5816 ^ w5819 ;
  assign w5821 = \pi22 & \pi54 ;
  assign w5822 = \pi21 & \pi55 ;
  assign w5823 = \pi20 & \pi56 ;
  assign w5824 = ( w5821 & w5822 ) | ( w5821 & w5823 ) | ( w5822 & w5823 ) ;
  assign w5825 = w5821 ^ w5823 ;
  assign w5826 = w5822 ^ w5825 ;
  assign w5827 = w5815 ^ w5820 ;
  assign w5828 = w5826 ^ w5827 ;
  assign w5829 = ( w5685 & w5686 ) | ( w5685 & w5687 ) | ( w5686 & w5687 ) ;
  assign w5830 = w5809 ^ w5829 ;
  assign w5831 = w5828 ^ w5830 ;
  assign w5832 = w5807 ^ w5808 ;
  assign w5833 = w5831 ^ w5832 ;
  assign w5834 = w5804 ^ w5833 ;
  assign w5835 = w5805 ^ w5834 ;
  assign w5836 = w5758 ^ w5835 ;
  assign w5837 = w5729 ^ w5730 ;
  assign w5838 = w5836 ^ w5837 ;
  assign w5839 = w5758 ^ w5804 ;
  assign w5840 = ( w5805 & w5833 ) | ( w5805 & w5839 ) | ( w5833 & w5839 ) ;
  assign w5841 = ( w5807 & w5808 ) | ( w5807 & w5831 ) | ( w5808 & w5831 ) ;
  assign w5842 = \pi18 & \pi59 ;
  assign w5843 = ( \pi17 & \pi60 ) | ( \pi17 & ~w5781 ) | ( \pi60 & ~w5781 ) ;
  assign w5844 = w5842 ^ w5843 ;
  assign w5845 = w5781 & w5844 ;
  assign w5846 = \pi17 & \pi60 ;
  assign w5847 = w5781 ^ w5846 ;
  assign w5848 = w5842 ^ w5847 ;
  assign w5849 = ( w5666 & w5672 ) | ( w5666 & w5705 ) | ( w5672 & w5705 ) ;
  assign w5850 = ( w5647 & w5678 ) | ( w5647 & w5699 ) | ( w5678 & w5699 ) ;
  assign w5851 = w5848 ^ w5849 ;
  assign w5852 = w5850 ^ w5851 ;
  assign w5853 = ( w5785 & w5786 ) | ( w5785 & w5801 ) | ( w5786 & w5801 ) ;
  assign w5854 = w5770 ^ w5813 ;
  assign w5855 = w5824 ^ w5854 ;
  assign w5856 = w5791 ^ w5818 ;
  assign w5857 = w5797 ^ w5856 ;
  assign w5858 = ( w5815 & w5820 ) | ( w5815 & w5826 ) | ( w5820 & w5826 ) ;
  assign w5859 = w5857 ^ w5858 ;
  assign w5860 = w5855 ^ w5859 ;
  assign w5861 = w5852 ^ w5853 ;
  assign w5862 = w5860 ^ w5861 ;
  assign w5863 = w5841 ^ w5862 ;
  assign w5864 = ( w5711 & w5793 ) | ( w5711 & w5799 ) | ( w5793 & w5799 ) ;
  assign w5865 = ( w5772 & w5778 ) | ( w5772 & w5783 ) | ( w5778 & w5783 ) ;
  assign w5866 = w5746 ^ w5865 ;
  assign w5867 = w5864 ^ w5866 ;
  assign w5868 = ( w5809 & w5828 ) | ( w5809 & w5829 ) | ( w5828 & w5829 ) ;
  assign w5869 = \pi31 & \pi46 ;
  assign w5870 = \pi30 & \pi47 ;
  assign w5871 = \pi14 & \pi63 ;
  assign w5872 = ( w5869 & w5870 ) | ( w5869 & w5871 ) | ( w5870 & w5871 ) ;
  assign w5873 = w5869 ^ w5871 ;
  assign w5874 = w5870 ^ w5873 ;
  assign w5875 = \pi37 & \pi40 ;
  assign w5876 = \pi36 & \pi41 ;
  assign w5877 = \pi35 & \pi42 ;
  assign w5878 = ( w5875 & w5876 ) | ( w5875 & w5877 ) | ( w5876 & w5877 ) ;
  assign w5879 = w5875 ^ w5877 ;
  assign w5880 = w5876 ^ w5879 ;
  assign w5881 = ~\pi38 & \pi39 ;
  assign w5882 = w5874 ^ w5881 ;
  assign w5883 = w5880 ^ w5882 ;
  assign w5884 = \pi15 & \pi62 ;
  assign w5885 = w5883 ^ w5884 ;
  assign w5886 = ( w5733 & w5734 ) | ( w5733 & w5735 ) | ( w5734 & w5735 ) ;
  assign w5887 = w5885 ^ w5886 ;
  assign w5888 = \pi21 & \pi56 ;
  assign w5889 = \pi20 & \pi57 ;
  assign w5890 = \pi19 & \pi58 ;
  assign w5891 = ( w5888 & w5889 ) | ( w5888 & w5890 ) | ( w5889 & w5890 ) ;
  assign w5892 = w5888 ^ w5890 ;
  assign w5893 = w5889 ^ w5892 ;
  assign w5894 = \pi29 & \pi48 ;
  assign w5895 = \pi28 & \pi49 ;
  assign w5896 = \pi27 & \pi50 ;
  assign w5897 = ( w5894 & w5895 ) | ( w5894 & w5896 ) | ( w5895 & w5896 ) ;
  assign w5898 = w5894 ^ w5896 ;
  assign w5899 = w5895 ^ w5898 ;
  assign w5900 = w5776 ^ w5893 ;
  assign w5901 = w5899 ^ w5900 ;
  assign w5902 = w5867 ^ w5901 ;
  assign w5903 = w5868 ^ w5902 ;
  assign w5904 = w5887 ^ w5903 ;
  assign w5905 = ( w5756 & w5757 ) | ( w5756 & w5804 ) | ( w5757 & w5804 ) ;
  assign w5906 = w5787 ^ w5801 ;
  assign w5907 = ( w5759 & w5766 ) | ( w5759 & w5906 ) | ( w5766 & w5906 ) ;
  assign w5908 = ( w5737 & w5738 ) | ( w5737 & w5754 ) | ( w5738 & w5754 ) ;
  assign w5909 = ( w5740 & w5741 ) | ( w5740 & w5752 ) | ( w5741 & w5752 ) ;
  assign w5910 = \pi34 & \pi43 ;
  assign w5911 = \pi26 & \pi51 ;
  assign w5912 = \pi22 & \pi55 ;
  assign w5913 = ( w5910 & w5911 ) | ( w5910 & w5912 ) | ( w5911 & w5912 ) ;
  assign w5914 = w5910 ^ w5912 ;
  assign w5915 = w5911 ^ w5914 ;
  assign w5916 = \pi25 & \pi52 ;
  assign w5917 = \pi24 & \pi53 ;
  assign w5918 = \pi23 & \pi54 ;
  assign w5919 = ( w5916 & w5917 ) | ( w5916 & w5918 ) | ( w5917 & w5918 ) ;
  assign w5920 = w5916 ^ w5918 ;
  assign w5921 = w5917 ^ w5920 ;
  assign w5922 = \pi33 & \pi44 ;
  assign w5923 = \pi32 & \pi45 ;
  assign w5924 = \pi16 & \pi61 ;
  assign w5925 = ( w5922 & w5923 ) | ( w5922 & w5924 ) | ( w5923 & w5924 ) ;
  assign w5926 = w5922 ^ w5924 ;
  assign w5927 = w5923 ^ w5926 ;
  assign w5928 = w5915 ^ w5921 ;
  assign w5929 = w5927 ^ w5928 ;
  assign w5930 = ( w5761 & w5762 ) | ( w5761 & w5764 ) | ( w5762 & w5764 ) ;
  assign w5931 = w5909 ^ w5930 ;
  assign w5932 = w5929 ^ w5931 ;
  assign w5933 = w5907 ^ w5908 ;
  assign w5934 = w5932 ^ w5933 ;
  assign w5935 = w5904 ^ w5934 ;
  assign w5936 = w5863 ^ w5935 ;
  assign w5937 = w5905 ^ w5936 ;
  assign w5938 = ( w5729 & w5730 ) | ( w5729 & w5836 ) | ( w5730 & w5836 ) ;
  assign w5939 = w5840 ^ w5938 ;
  assign w5940 = w5937 ^ w5939 ;
  assign w5941 = ( w5840 & w5937 ) | ( w5840 & w5938 ) | ( w5937 & w5938 ) ;
  assign w5942 = w5863 ^ w5904 ;
  assign w5943 = ( w5905 & w5934 ) | ( w5905 & w5942 ) | ( w5934 & w5942 ) ;
  assign w5944 = w5887 ^ w5901 ;
  assign w5945 = ( w5867 & w5868 ) | ( w5867 & w5944 ) | ( w5868 & w5944 ) ;
  assign w5946 = ( w5852 & w5853 ) | ( w5852 & w5860 ) | ( w5853 & w5860 ) ;
  assign w5947 = ( w5746 & w5864 ) | ( w5746 & w5865 ) | ( w5864 & w5865 ) ;
  assign w5948 = \pi21 & \pi57 ;
  assign w5949 = \pi19 & \pi59 ;
  assign w5950 = \pi18 & \pi60 ;
  assign w5951 = ( w5948 & w5949 ) | ( w5948 & w5950 ) | ( w5949 & w5950 ) ;
  assign w5952 = w5948 ^ w5950 ;
  assign w5953 = w5949 ^ w5952 ;
  assign w5954 = \pi29 & \pi49 ;
  assign w5955 = \pi28 & \pi50 ;
  assign w5956 = \pi27 & \pi51 ;
  assign w5957 = ( w5954 & w5955 ) | ( w5954 & w5956 ) | ( w5955 & w5956 ) ;
  assign w5958 = w5954 ^ w5956 ;
  assign w5959 = w5955 ^ w5958 ;
  assign w5960 = \pi17 & \pi61 ;
  assign w5961 = \pi16 & \pi62 ;
  assign w5962 = \pi15 & \pi63 ;
  assign w5963 = ( w5960 & w5961 ) | ( w5960 & w5962 ) | ( w5961 & w5962 ) ;
  assign w5964 = w5960 ^ w5962 ;
  assign w5965 = w5961 ^ w5964 ;
  assign w5966 = w5953 ^ w5959 ;
  assign w5967 = w5965 ^ w5966 ;
  assign w5968 = \pi31 & \pi47 ;
  assign w5969 = \pi30 & \pi48 ;
  assign w5970 = \pi20 & \pi58 ;
  assign w5971 = ( w5968 & w5969 ) | ( w5968 & w5970 ) | ( w5969 & w5970 ) ;
  assign w5972 = w5968 ^ w5970 ;
  assign w5973 = w5969 ^ w5972 ;
  assign w5974 = \pi34 & \pi44 ;
  assign w5975 = \pi33 & \pi45 ;
  assign w5976 = \pi32 & \pi46 ;
  assign w5977 = ( w5974 & w5975 ) | ( w5974 & w5976 ) | ( w5975 & w5976 ) ;
  assign w5978 = w5974 ^ w5976 ;
  assign w5979 = w5975 ^ w5978 ;
  assign w5980 = \pi25 & \pi53 ;
  assign w5981 = \pi24 & \pi54 ;
  assign w5982 = \pi22 & \pi56 ;
  assign w5983 = ( w5980 & w5981 ) | ( w5980 & w5982 ) | ( w5981 & w5982 ) ;
  assign w5984 = w5980 ^ w5982 ;
  assign w5985 = w5981 ^ w5984 ;
  assign w5986 = w5973 ^ w5979 ;
  assign w5987 = w5985 ^ w5986 ;
  assign w5988 = w5947 ^ w5967 ;
  assign w5989 = w5987 ^ w5988 ;
  assign w5990 = w5945 ^ w5946 ;
  assign w5991 = w5989 ^ w5990 ;
  assign w5992 = ( w5841 & w5862 ) | ( w5841 & w5904 ) | ( w5862 & w5904 ) ;
  assign w5993 = ( w5907 & w5908 ) | ( w5907 & w5932 ) | ( w5908 & w5932 ) ;
  assign w5994 = ( w5776 & w5893 ) | ( w5776 & w5899 ) | ( w5893 & w5899 ) ;
  assign w5995 = w5881 ^ w5884 ;
  assign w5996 = ( w5874 & w5880 ) | ( w5874 & w5995 ) | ( w5880 & w5995 ) ;
  assign w5997 = ( w5915 & w5921 ) | ( w5915 & w5927 ) | ( w5921 & w5927 ) ;
  assign w5998 = w5994 ^ w5996 ;
  assign w5999 = w5997 ^ w5998 ;
  assign w6000 = ( w5855 & w5857 ) | ( w5855 & w5858 ) | ( w5857 & w5858 ) ;
  assign w6001 = w5878 ^ w5919 ;
  assign w6002 = ( \pi15 & \pi38 ) | ( \pi15 & \pi62 ) | ( \pi38 & \pi62 ) ;
  assign w6003 = ~\pi38 & w6002 ;
  assign w6004 = ( \pi38 & \pi39 ) | ( \pi38 & w6003 ) | ( \pi39 & w6003 ) ;
  assign w6005 = w6001 ^ w6004 ;
  assign w6006 = w5872 ^ w5897 ;
  assign w6007 = w5925 ^ w6006 ;
  assign w6008 = ( w5791 & w5797 ) | ( w5791 & w5818 ) | ( w5797 & w5818 ) ;
  assign w6009 = w6005 ^ w6008 ;
  assign w6010 = w6007 ^ w6009 ;
  assign w6011 = w6000 ^ w6010 ;
  assign w6012 = w5999 ^ w6011 ;
  assign w6013 = w5993 ^ w6012 ;
  assign w6014 = ( w5909 & w5929 ) | ( w5909 & w5930 ) | ( w5929 & w5930 ) ;
  assign w6015 = ( w5885 & w5886 ) | ( w5885 & w5901 ) | ( w5886 & w5901 ) ;
  assign w6016 = \pi36 & \pi42 ;
  assign w6017 = \pi35 & \pi43 ;
  assign w6018 = \pi23 & \pi55 ;
  assign w6019 = ( w6016 & w6017 ) | ( w6016 & w6018 ) | ( w6017 & w6018 ) ;
  assign w6020 = w6016 ^ w6018 ;
  assign w6021 = w6017 ^ w6020 ;
  assign w6022 = \pi38 & \pi40 ;
  assign w6023 = \pi37 & \pi41 ;
  assign w6024 = \pi26 & \pi52 ;
  assign w6025 = ( w6022 & w6023 ) | ( w6022 & w6024 ) | ( w6023 & w6024 ) ;
  assign w6026 = w6022 ^ w6024 ;
  assign w6027 = w6023 ^ w6026 ;
  assign w6028 = ( w5770 & w5813 ) | ( w5770 & w5824 ) | ( w5813 & w5824 ) ;
  assign w6029 = w6021 ^ w6028 ;
  assign w6030 = w6027 ^ w6029 ;
  assign w6031 = w5891 ^ w5913 ;
  assign w6032 = w4299 | w5845 ;
  assign w6033 = ( w492 & w5845 ) | ( w492 & w6032 ) | ( w5845 & w6032 ) ;
  assign w6034 = w6031 ^ w6033 ;
  assign w6035 = ( w5848 & w5849 ) | ( w5848 & w5850 ) | ( w5849 & w5850 ) ;
  assign w6036 = w6034 ^ w6035 ;
  assign w6037 = w6030 ^ w6036 ;
  assign w6038 = w6015 ^ w6037 ;
  assign w6039 = w6014 ^ w6038 ;
  assign w6040 = w5991 ^ w6039 ;
  assign w6041 = w5992 ^ w6040 ;
  assign w6042 = w6013 ^ w6041 ;
  assign w6043 = w5941 ^ w5943 ;
  assign w6044 = w6042 ^ w6043 ;
  assign w6045 = w6013 ^ w6039 ;
  assign w6046 = ( w5991 & w5992 ) | ( w5991 & w6045 ) | ( w5992 & w6045 ) ;
  assign w6047 = ( w6014 & w6015 ) | ( w6014 & w6037 ) | ( w6015 & w6037 ) ;
  assign w6048 = ( w5947 & w5967 ) | ( w5947 & w5987 ) | ( w5967 & w5987 ) ;
  assign w6049 = w5951 ^ w5957 ;
  assign w6050 = w5983 ^ w6049 ;
  assign w6051 = ( w6021 & w6027 ) | ( w6021 & w6028 ) | ( w6027 & w6028 ) ;
  assign w6052 = \pi35 & \pi44 ;
  assign w6053 = \pi34 & \pi45 ;
  assign w6054 = \pi16 & \pi63 ;
  assign w6055 = ( w6052 & w6053 ) | ( w6052 & w6054 ) | ( w6053 & w6054 ) ;
  assign w6056 = w6052 ^ w6054 ;
  assign w6057 = w6053 ^ w6056 ;
  assign w6058 = \pi27 & \pi56 ;
  assign w6059 = \pi36 & \pi43 ;
  assign w6060 = \pi27 & \pi52 ;
  assign w6061 = \pi23 & \pi56 ;
  assign w6062 = ( w6059 & w6060 ) | ( w6059 & w6061 ) | ( w6060 & w6061 ) ;
  assign w6063 = w6059 ^ w6061 ;
  assign w6064 = w6060 ^ w6063 ;
  assign w6065 = w492 & w4299 ;
  assign w6066 = w5845 | w6065 ;
  assign w6067 = ( w5891 & w5913 ) | ( w5891 & w6066 ) | ( w5913 & w6066 ) ;
  assign w6068 = w6057 ^ w6067 ;
  assign w6069 = w6064 ^ w6068 ;
  assign w6070 = w6051 ^ w6069 ;
  assign w6071 = w6050 ^ w6070 ;
  assign w6072 = ( w5973 & w5979 ) | ( w5973 & w5985 ) | ( w5979 & w5985 ) ;
  assign w6073 = w5963 ^ w5971 ;
  assign w6074 = w5977 ^ w6073 ;
  assign w6075 = w6072 ^ w6074 ;
  assign w6076 = w6019 ^ w6075 ;
  assign w6077 = w6025 ^ w6076 ;
  assign w6078 = \pi18 & \pi61 ;
  assign w6079 = w6077 ^ w6078 ;
  assign w6080 = w6048 ^ w6071 ;
  assign w6081 = w6079 ^ w6080 ;
  assign w6082 = ( w5945 & w5946 ) | ( w5945 & w5989 ) | ( w5946 & w5989 ) ;
  assign w6083 = w6081 ^ w6082 ;
  assign w6084 = w6047 ^ w6083 ;
  assign w6085 = ( w5993 & w6012 ) | ( w5993 & w6039 ) | ( w6012 & w6039 ) ;
  assign w6086 = ( w5999 & w6000 ) | ( w5999 & w6010 ) | ( w6000 & w6010 ) ;
  assign w6087 = ( w6005 & w6007 ) | ( w6005 & w6008 ) | ( w6007 & w6008 ) ;
  assign w6088 = \pi26 & \pi53 ;
  assign w6089 = \pi25 & \pi54 ;
  assign w6090 = \pi24 & \pi55 ;
  assign w6091 = ( w6088 & w6089 ) | ( w6088 & w6090 ) | ( w6089 & w6090 ) ;
  assign w6092 = w6088 ^ w6090 ;
  assign w6093 = w6089 ^ w6092 ;
  assign w6094 = \pi39 & \pi40 ;
  assign w6095 = \pi38 & \pi41 ;
  assign w6096 = \pi37 & \pi42 ;
  assign w6097 = ( w6094 & w6095 ) | ( w6094 & w6096 ) | ( w6095 & w6096 ) ;
  assign w6098 = w6094 ^ w6096 ;
  assign w6099 = w6095 ^ w6098 ;
  assign w6100 = \pi40 & \pi62 ;
  assign w6101 = \pi28 & \pi51 ;
  assign w6102 = \pi17 & \pi62 ;
  assign w6103 = ( \pi40 & w6101 ) | ( \pi40 & w6102 ) | ( w6101 & w6102 ) ;
  assign w6104 = \pi40 ^ w6102 ;
  assign w6105 = w6101 ^ w6104 ;
  assign w6106 = w6093 ^ w6099 ;
  assign w6107 = w6105 ^ w6106 ;
  assign w6108 = \pi21 & \pi58 ;
  assign w6109 = \pi20 & \pi59 ;
  assign w6110 = \pi19 & \pi60 ;
  assign w6111 = ( w6108 & w6109 ) | ( w6108 & w6110 ) | ( w6109 & w6110 ) ;
  assign w6112 = w6108 ^ w6110 ;
  assign w6113 = w6109 ^ w6112 ;
  assign w6114 = \pi30 & \pi49 ;
  assign w6115 = \pi29 & \pi50 ;
  assign w6116 = \pi22 & \pi57 ;
  assign w6117 = ( w6114 & w6115 ) | ( w6114 & w6116 ) | ( w6115 & w6116 ) ;
  assign w6118 = w6114 ^ w6116 ;
  assign w6119 = w6115 ^ w6118 ;
  assign w6120 = \pi33 & \pi46 ;
  assign w6121 = \pi32 & \pi47 ;
  assign w6122 = \pi31 & \pi48 ;
  assign w6123 = ( w6120 & w6121 ) | ( w6120 & w6122 ) | ( w6121 & w6122 ) ;
  assign w6124 = w6120 ^ w6122 ;
  assign w6125 = w6121 ^ w6124 ;
  assign w6126 = w6113 ^ w6119 ;
  assign w6127 = w6125 ^ w6126 ;
  assign w6128 = w6087 ^ w6107 ;
  assign w6129 = w6127 ^ w6128 ;
  assign w6130 = ( w5872 & w5897 ) | ( w5872 & w5925 ) | ( w5897 & w5925 ) ;
  assign w6131 = \pi38 & \pi39 ;
  assign w6132 = ( \pi39 & w6002 ) | ( \pi39 & w6131 ) | ( w6002 & w6131 ) ;
  assign w6133 = ( w5878 & w5919 ) | ( w5878 & w6132 ) | ( w5919 & w6132 ) ;
  assign w6134 = ( w5953 & w5959 ) | ( w5953 & w5965 ) | ( w5959 & w5965 ) ;
  assign w6135 = w6130 ^ w6133 ;
  assign w6136 = w6134 ^ w6135 ;
  assign w6137 = ( w5994 & w5996 ) | ( w5994 & w5997 ) | ( w5996 & w5997 ) ;
  assign w6138 = ( w6030 & w6034 ) | ( w6030 & w6035 ) | ( w6034 & w6035 ) ;
  assign w6139 = w6136 ^ w6138 ;
  assign w6140 = w6137 ^ w6139 ;
  assign w6141 = w6086 ^ w6140 ;
  assign w6142 = w6129 ^ w6141 ;
  assign w6143 = w6084 ^ w6085 ;
  assign w6144 = w6142 ^ w6143 ;
  assign w6145 = ( w5941 & w5943 ) | ( w5941 & w6042 ) | ( w5943 & w6042 ) ;
  assign w6146 = w6046 ^ w6145 ;
  assign w6147 = w6144 ^ w6146 ;
  assign w6148 = ( w6046 & w6144 ) | ( w6046 & w6145 ) | ( w6144 & w6145 ) ;
  assign w6149 = ( w6084 & w6085 ) | ( w6084 & w6142 ) | ( w6085 & w6142 ) ;
  assign w6150 = ( w6047 & w6081 ) | ( w6047 & w6082 ) | ( w6081 & w6082 ) ;
  assign w6151 = ( w6048 & w6071 ) | ( w6048 & w6079 ) | ( w6071 & w6079 ) ;
  assign w6152 = ( w6136 & w6137 ) | ( w6136 & w6138 ) | ( w6137 & w6138 ) ;
  assign w6153 = \pi29 & \pi63 ;
  assign w6154 = \pi33 & \pi47 ;
  assign w6155 = \pi29 & \pi51 ;
  assign w6156 = \pi17 & \pi63 ;
  assign w6157 = ( w6154 & w6155 ) | ( w6154 & w6156 ) | ( w6155 & w6156 ) ;
  assign w6158 = w6154 ^ w6156 ;
  assign w6159 = w6155 ^ w6158 ;
  assign w6160 = \pi36 & \pi44 ;
  assign w6161 = \pi35 & \pi45 ;
  assign w6162 = \pi34 & \pi46 ;
  assign w6163 = ( w6160 & w6161 ) | ( w6160 & w6162 ) | ( w6161 & w6162 ) ;
  assign w6164 = w6160 ^ w6162 ;
  assign w6165 = w6161 ^ w6164 ;
  assign w6166 = \pi19 & \pi61 ;
  assign w6167 = ( \pi18 & \pi62 ) | ( \pi18 & ~w6103 ) | ( \pi62 & ~w6103 ) ;
  assign w6168 = w6166 ^ w6167 ;
  assign w6169 = w6103 & w6168 ;
  assign w6170 = \pi18 & \pi62 ;
  assign w6171 = w6103 ^ w6170 ;
  assign w6172 = w6166 ^ w6171 ;
  assign w6173 = w6159 ^ w6172 ;
  assign w6174 = w6165 ^ w6173 ;
  assign w6175 = \pi20 & \pi60 ;
  assign w6176 = \pi22 & \pi58 ;
  assign w6177 = w6175 ^ w6176 ;
  assign w6178 = \pi21 & \pi59 ;
  assign w6179 = w6177 ^ w6178 ;
  assign w6180 = \pi32 & \pi48 ;
  assign w6181 = \pi31 & \pi49 ;
  assign w6182 = \pi30 & \pi50 ;
  assign w6183 = ( w6180 & w6181 ) | ( w6180 & w6182 ) | ( w6181 & w6182 ) ;
  assign w6184 = w6180 ^ w6182 ;
  assign w6185 = w6181 ^ w6184 ;
  assign w6186 = w6097 ^ w6179 ;
  assign w6187 = w6185 ^ w6186 ;
  assign w6188 = \pi26 & \pi54 ;
  assign w6189 = \pi24 & \pi56 ;
  assign w6190 = \pi23 & \pi57 ;
  assign w6191 = ( w6188 & w6189 ) | ( w6188 & w6190 ) | ( w6189 & w6190 ) ;
  assign w6192 = w6188 ^ w6190 ;
  assign w6193 = w6189 ^ w6192 ;
  assign w6194 = \pi38 & \pi42 ;
  assign w6195 = \pi37 & \pi43 ;
  assign w6196 = \pi25 & \pi55 ;
  assign w6197 = ( w6194 & w6195 ) | ( w6194 & w6196 ) | ( w6195 & w6196 ) ;
  assign w6198 = w6194 ^ w6196 ;
  assign w6199 = w6195 ^ w6198 ;
  assign w6200 = \pi28 & \pi52 ;
  assign w6201 = \pi27 & \pi53 ;
  assign w6202 = ( w1851 & w6200 ) | ( w1851 & w6201 ) | ( w6200 & w6201 ) ;
  assign w6203 = w1851 ^ w6201 ;
  assign w6204 = w6200 ^ w6203 ;
  assign w6205 = w6193 ^ w6204 ;
  assign w6206 = w6199 ^ w6205 ;
  assign w6207 = w6174 ^ w6206 ;
  assign w6208 = w6187 ^ w6207 ;
  assign w6209 = w6151 ^ w6152 ;
  assign w6210 = w6208 ^ w6209 ;
  assign w6211 = ( w6086 & w6129 ) | ( w6086 & w6140 ) | ( w6129 & w6140 ) ;
  assign w6212 = ( w5951 & w5957 ) | ( w5951 & w5983 ) | ( w5957 & w5983 ) ;
  assign w6213 = ( w5963 & w5971 ) | ( w5963 & w5977 ) | ( w5971 & w5977 ) ;
  assign w6214 = ( w6019 & w6025 ) | ( w6019 & w6078 ) | ( w6025 & w6078 ) ;
  assign w6215 = w6212 ^ w6214 ;
  assign w6216 = w6213 ^ w6215 ;
  assign w6217 = ( w6050 & w6051 ) | ( w6050 & w6069 ) | ( w6051 & w6069 ) ;
  assign w6218 = w6019 ^ w6025 ;
  assign w6219 = w6078 ^ w6218 ;
  assign w6220 = ( w6072 & w6074 ) | ( w6072 & w6219 ) | ( w6074 & w6219 ) ;
  assign w6221 = w6216 ^ w6217 ;
  assign w6222 = w6220 ^ w6221 ;
  assign w6223 = ( w6087 & w6107 ) | ( w6087 & w6127 ) | ( w6107 & w6127 ) ;
  assign w6224 = w6055 ^ w6062 ;
  assign w6225 = w6091 ^ w6224 ;
  assign w6226 = ( w6057 & w6064 ) | ( w6057 & w6067 ) | ( w6064 & w6067 ) ;
  assign w6227 = ( w6130 & w6133 ) | ( w6130 & w6134 ) | ( w6133 & w6134 ) ;
  assign w6228 = w6226 ^ w6227 ;
  assign w6229 = w6225 ^ w6228 ;
  assign w6230 = w6111 ^ w6117 ;
  assign w6231 = w6123 ^ w6230 ;
  assign w6232 = ( w6093 & w6099 ) | ( w6093 & w6105 ) | ( w6099 & w6105 ) ;
  assign w6233 = ( w6113 & w6119 ) | ( w6113 & w6125 ) | ( w6119 & w6125 ) ;
  assign w6234 = w6231 ^ w6232 ;
  assign w6235 = w6233 ^ w6234 ;
  assign w6236 = w6223 ^ w6229 ;
  assign w6237 = w6235 ^ w6236 ;
  assign w6238 = w6211 ^ w6222 ;
  assign w6239 = w6237 ^ w6238 ;
  assign w6240 = w6150 ^ w6210 ;
  assign w6241 = w6239 ^ w6240 ;
  assign w6242 = w6149 | w6241 ;
  assign w6243 = w6149 & w6241 ;
  assign w6244 = w6242 & ~w6243 ;
  assign w6245 = w6148 ^ w6244 ;
  assign w6246 = ( w6148 & w6242 ) | ( w6148 & w6243 ) | ( w6242 & w6243 ) ;
  assign w6247 = w6243 | w6246 ;
  assign w6248 = ( w6211 & w6222 ) | ( w6211 & w6237 ) | ( w6222 & w6237 ) ;
  assign w6249 = ( w6223 & w6229 ) | ( w6223 & w6235 ) | ( w6229 & w6235 ) ;
  assign w6250 = ( w6216 & w6217 ) | ( w6216 & w6220 ) | ( w6217 & w6220 ) ;
  assign w6251 = \pi25 & \pi56 ;
  assign w6252 = \pi23 & \pi58 ;
  assign w6253 = \pi22 & \pi59 ;
  assign w6254 = ( w6251 & w6252 ) | ( w6251 & w6253 ) | ( w6252 & w6253 ) ;
  assign w6255 = w6251 ^ w6253 ;
  assign w6256 = w6252 ^ w6255 ;
  assign w6257 = \pi34 & \pi47 ;
  assign w6258 = \pi33 & \pi48 ;
  assign w6259 = \pi24 & \pi57 ;
  assign w6260 = ( w6257 & w6258 ) | ( w6257 & w6259 ) | ( w6258 & w6259 ) ;
  assign w6261 = w6257 ^ w6259 ;
  assign w6262 = w6258 ^ w6261 ;
  assign w6263 = ~\pi40 & \pi41 ;
  assign w6264 = w6256 ^ w6263 ;
  assign w6265 = w6262 ^ w6264 ;
  assign w6266 = \pi19 & \pi62 ;
  assign w6267 = w6265 ^ w6266 ;
  assign w6268 = ( w6212 & w6213 ) | ( w6212 & w6214 ) | ( w6213 & w6214 ) ;
  assign w6269 = \pi21 & \pi60 ;
  assign w6270 = \pi20 & \pi61 ;
  assign w6271 = \pi18 & \pi63 ;
  assign w6272 = ( w6269 & w6270 ) | ( w6269 & w6271 ) | ( w6270 & w6271 ) ;
  assign w6273 = w6269 ^ w6271 ;
  assign w6274 = w6270 ^ w6273 ;
  assign w6275 = \pi37 & \pi44 ;
  assign w6276 = \pi36 & \pi45 ;
  assign w6277 = \pi35 & \pi46 ;
  assign w6278 = ( w6275 & w6276 ) | ( w6275 & w6277 ) | ( w6276 & w6277 ) ;
  assign w6279 = w6275 ^ w6277 ;
  assign w6280 = w6276 ^ w6279 ;
  assign w6281 = \pi29 & \pi52 ;
  assign w6282 = \pi28 & \pi53 ;
  assign w6283 = \pi26 & \pi55 ;
  assign w6284 = ( w6281 & w6282 ) | ( w6281 & w6283 ) | ( w6282 & w6283 ) ;
  assign w6285 = w6281 ^ w6283 ;
  assign w6286 = w6282 ^ w6285 ;
  assign w6287 = w6274 ^ w6280 ;
  assign w6288 = w6286 ^ w6287 ;
  assign w6289 = w6267 ^ w6268 ;
  assign w6290 = w6288 ^ w6289 ;
  assign w6291 = w6249 ^ w6250 ;
  assign w6292 = w6290 ^ w6291 ;
  assign w6293 = ( w6151 & w6152 ) | ( w6151 & w6208 ) | ( w6152 & w6208 ) ;
  assign w6294 = ( w6111 & w6117 ) | ( w6111 & w6123 ) | ( w6117 & w6123 ) ;
  assign w6295 = \pi27 & \pi54 ;
  assign w6296 = \pi39 & \pi42 ;
  assign w6297 = \pi38 & \pi43 ;
  assign w6298 = ( w6295 & w6296 ) | ( w6295 & w6297 ) | ( w6296 & w6297 ) ;
  assign w6299 = w6295 ^ w6297 ;
  assign w6300 = w6296 ^ w6299 ;
  assign w6301 = ( w6055 & w6062 ) | ( w6055 & w6091 ) | ( w6062 & w6091 ) ;
  assign w6302 = w6294 ^ w6300 ;
  assign w6303 = w6301 ^ w6302 ;
  assign w6304 = ( w6225 & w6226 ) | ( w6225 & w6227 ) | ( w6226 & w6227 ) ;
  assign w6305 = ( w6231 & w6232 ) | ( w6231 & w6233 ) | ( w6232 & w6233 ) ;
  assign w6306 = w6304 ^ w6305 ;
  assign w6307 = \pi32 & \pi49 ;
  assign w6308 = \pi31 & \pi50 ;
  assign w6309 = \pi30 & \pi51 ;
  assign w6310 = ( w6307 & w6308 ) | ( w6307 & w6309 ) | ( w6308 & w6309 ) ;
  assign w6311 = w6307 ^ w6309 ;
  assign w6312 = w6308 ^ w6311 ;
  assign w6313 = ~\pi18 & w4390 ;
  assign w6314 = ( w4390 & w6169 ) | ( w4390 & ~w6313 ) | ( w6169 & ~w6313 ) ;
  assign w6315 = ( \pi19 & w6169 ) | ( \pi19 & w6314 ) | ( w6169 & w6314 ) ;
  assign w6316 = w6163 ^ w6312 ;
  assign w6317 = w6315 ^ w6316 ;
  assign w6318 = ( w6175 & w6176 ) | ( w6175 & w6178 ) | ( w6176 & w6178 ) ;
  assign w6319 = w6157 ^ w6183 ;
  assign w6320 = w6318 ^ w6319 ;
  assign w6321 = ( w6159 & w6165 ) | ( w6159 & w6172 ) | ( w6165 & w6172 ) ;
  assign w6322 = w6317 ^ w6321 ;
  assign w6323 = w6320 ^ w6322 ;
  assign w6324 = ( w6174 & w6187 ) | ( w6174 & w6206 ) | ( w6187 & w6206 ) ;
  assign w6325 = w6191 ^ w6202 ;
  assign w6326 = w6197 ^ w6325 ;
  assign w6327 = ( w6193 & w6199 ) | ( w6193 & w6204 ) | ( w6199 & w6204 ) ;
  assign w6328 = ( w6097 & w6179 ) | ( w6097 & w6185 ) | ( w6179 & w6185 ) ;
  assign w6329 = w6326 ^ w6327 ;
  assign w6330 = w6328 ^ w6329 ;
  assign w6331 = w6323 ^ w6324 ;
  assign w6332 = w6330 ^ w6331 ;
  assign w6333 = w6303 ^ w6332 ;
  assign w6334 = w6293 ^ w6333 ;
  assign w6335 = w6306 ^ w6334 ;
  assign w6336 = w6248 ^ w6335 ;
  assign w6337 = w6292 ^ w6336 ;
  assign w6338 = ( w6150 & w6210 ) | ( w6150 & w6239 ) | ( w6210 & w6239 ) ;
  assign w6339 = w6247 ^ w6337 ;
  assign w6340 = w6338 ^ w6339 ;
  assign w6341 = ( w6247 & w6337 ) | ( w6247 & w6338 ) | ( w6337 & w6338 ) ;
  assign w6342 = ( w6248 & w6292 ) | ( w6248 & w6335 ) | ( w6292 & w6335 ) ;
  assign w6343 = w6303 ^ w6306 ;
  assign w6344 = ( w6293 & w6332 ) | ( w6293 & w6343 ) | ( w6332 & w6343 ) ;
  assign w6345 = ( w6323 & w6324 ) | ( w6323 & w6330 ) | ( w6324 & w6330 ) ;
  assign w6346 = ( w6303 & w6304 ) | ( w6303 & w6305 ) | ( w6304 & w6305 ) ;
  assign w6347 = \pi31 & \pi51 ;
  assign w6348 = \pi21 & \pi61 ;
  assign w6349 = \pi20 & \pi62 ;
  assign w6350 = ( w6347 & w6348 ) | ( w6347 & w6349 ) | ( w6348 & w6349 ) ;
  assign w6351 = w6347 ^ w6349 ;
  assign w6352 = w6348 ^ w6351 ;
  assign w6353 = \pi34 & \pi48 ;
  assign w6354 = \pi33 & \pi49 ;
  assign w6355 = \pi32 & \pi50 ;
  assign w6356 = ( w6353 & w6354 ) | ( w6353 & w6355 ) | ( w6354 & w6355 ) ;
  assign w6357 = w6353 ^ w6355 ;
  assign w6358 = w6354 ^ w6357 ;
  assign w6359 = \pi24 & \pi58 ;
  assign w6360 = \pi23 & \pi59 ;
  assign w6361 = \pi22 & \pi60 ;
  assign w6362 = ( w6359 & w6360 ) | ( w6359 & w6361 ) | ( w6360 & w6361 ) ;
  assign w6363 = w6359 ^ w6361 ;
  assign w6364 = w6360 ^ w6363 ;
  assign w6365 = w6352 ^ w6358 ;
  assign w6366 = w6364 ^ w6365 ;
  assign w6367 = ( w6294 & w6300 ) | ( w6294 & w6301 ) | ( w6300 & w6301 ) ;
  assign w6368 = \pi39 & \pi43 ;
  assign w6369 = \pi38 & \pi44 ;
  assign w6370 = \pi26 & \pi56 ;
  assign w6371 = ( w6368 & w6369 ) | ( w6368 & w6370 ) | ( w6369 & w6370 ) ;
  assign w6372 = w6368 ^ w6370 ;
  assign w6373 = w6369 ^ w6372 ;
  assign w6374 = \pi30 & \pi52 ;
  assign w6375 = \pi29 & \pi53 ;
  assign w6376 = ( w2959 & w6374 ) | ( w2959 & w6375 ) | ( w6374 & w6375 ) ;
  assign w6377 = w2959 ^ w6375 ;
  assign w6378 = w6374 ^ w6377 ;
  assign w6379 = \pi37 & \pi47 ;
  assign w6380 = \pi37 & \pi45 ;
  assign w6381 = \pi36 & \pi46 ;
  assign w6382 = \pi35 & \pi47 ;
  assign w6383 = ( w6380 & w6381 ) | ( w6380 & w6382 ) | ( w6381 & w6382 ) ;
  assign w6384 = w6380 ^ w6382 ;
  assign w6385 = w6381 ^ w6384 ;
  assign w6386 = w6373 ^ w6378 ;
  assign w6387 = w6385 ^ w6386 ;
  assign w6388 = w6367 ^ w6387 ;
  assign w6389 = w6366 ^ w6388 ;
  assign w6390 = w6345 ^ w6346 ;
  assign w6391 = w6389 ^ w6390 ;
  assign w6392 = ( w6249 & w6250 ) | ( w6249 & w6290 ) | ( w6250 & w6290 ) ;
  assign w6393 = ( w6157 & w6183 ) | ( w6157 & w6318 ) | ( w6183 & w6318 ) ;
  assign w6394 = \pi28 & \pi54 ;
  assign w6395 = \pi25 & \pi57 ;
  assign w6396 = ( w3648 & w6394 ) | ( w3648 & w6395 ) | ( w6394 & w6395 ) ;
  assign w6397 = w6394 ^ w6395 ;
  assign w6398 = w3648 ^ w6397 ;
  assign w6399 = ( w6191 & w6197 ) | ( w6191 & w6202 ) | ( w6197 & w6202 ) ;
  assign w6400 = w6393 ^ w6399 ;
  assign w6401 = w6398 ^ w6400 ;
  assign w6402 = ( w6317 & w6320 ) | ( w6317 & w6321 ) | ( w6320 & w6321 ) ;
  assign w6403 = ( w6326 & w6327 ) | ( w6326 & w6328 ) | ( w6327 & w6328 ) ;
  assign w6404 = w6402 ^ w6403 ;
  assign w6405 = ( w6267 & w6268 ) | ( w6267 & w6288 ) | ( w6268 & w6288 ) ;
  assign w6406 = w6260 ^ w6284 ;
  assign w6407 = w6310 ^ w6406 ;
  assign w6408 = w6254 ^ w6272 ;
  assign w6409 = w6278 ^ w6408 ;
  assign w6410 = ( w6274 & w6280 ) | ( w6274 & w6286 ) | ( w6280 & w6286 ) ;
  assign w6411 = w6407 ^ w6409 ;
  assign w6412 = w6410 ^ w6411 ;
  assign w6413 = \pi18 | w6169 ;
  assign w6414 = ( \pi19 & w6169 ) | ( \pi19 & w6413 ) | ( w6169 & w6413 ) ;
  assign w6415 = ( w4390 & w6169 ) | ( w4390 & w6414 ) | ( w6169 & w6414 ) ;
  assign w6416 = ( w6163 & w6312 ) | ( w6163 & w6415 ) | ( w6312 & w6415 ) ;
  assign w6417 = w6263 ^ w6266 ;
  assign w6418 = ( w6256 & w6262 ) | ( w6256 & w6417 ) | ( w6262 & w6417 ) ;
  assign w6419 = \pi19 & \pi63 ;
  assign w6420 = w6298 ^ w6419 ;
  assign w6421 = ~\pi40 & \pi62 ;
  assign w6422 = \pi19 & w6421 ;
  assign w6423 = ( \pi40 & \pi41 ) | ( \pi40 & w6422 ) | ( \pi41 & w6422 ) ;
  assign w6424 = w6420 ^ w6423 ;
  assign w6425 = w6416 ^ w6424 ;
  assign w6426 = w6418 ^ w6425 ;
  assign w6427 = w6405 ^ w6426 ;
  assign w6428 = w6412 ^ w6427 ;
  assign w6429 = w6401 ^ w6428 ;
  assign w6430 = w6392 ^ w6429 ;
  assign w6431 = w6404 ^ w6430 ;
  assign w6432 = w6344 ^ w6431 ;
  assign w6433 = w6391 ^ w6432 ;
  assign w6434 = w6341 ^ w6342 ;
  assign w6435 = w6433 ^ w6434 ;
  assign w6436 = ( w6344 & w6391 ) | ( w6344 & w6431 ) | ( w6391 & w6431 ) ;
  assign w6437 = ( w6366 & w6367 ) | ( w6366 & w6387 ) | ( w6367 & w6387 ) ;
  assign w6438 = ( w6407 & w6409 ) | ( w6407 & w6410 ) | ( w6409 & w6410 ) ;
  assign w6439 = w6362 ^ w6371 ;
  assign w6440 = w6383 ^ w6439 ;
  assign w6441 = w6350 ^ w6356 ;
  assign w6442 = w6396 ^ w6441 ;
  assign w6443 = ( w6373 & w6378 ) | ( w6373 & w6385 ) | ( w6378 & w6385 ) ;
  assign w6444 = w6440 ^ w6443 ;
  assign w6445 = w6442 ^ w6444 ;
  assign w6446 = w6437 ^ w6445 ;
  assign w6447 = w6438 ^ w6446 ;
  assign w6448 = ( w6345 & w6346 ) | ( w6345 & w6389 ) | ( w6346 & w6389 ) ;
  assign w6449 = ( w6260 & w6284 ) | ( w6260 & w6310 ) | ( w6284 & w6310 ) ;
  assign w6450 = ( w6254 & w6272 ) | ( w6254 & w6278 ) | ( w6272 & w6278 ) ;
  assign w6451 = ( w6352 & w6358 ) | ( w6352 & w6364 ) | ( w6358 & w6364 ) ;
  assign w6452 = w6449 ^ w6450 ;
  assign w6453 = w6451 ^ w6452 ;
  assign w6454 = \pi24 & \pi59 ;
  assign w6455 = ( \pi23 & \pi60 ) | ( \pi23 & ~w6376 ) | ( \pi60 & ~w6376 ) ;
  assign w6456 = w6454 ^ w6455 ;
  assign w6457 = w6376 & w6456 ;
  assign w6458 = \pi23 & \pi60 ;
  assign w6459 = w6376 ^ w6458 ;
  assign w6460 = w6454 ^ w6459 ;
  assign w6461 = \pi31 & \pi52 ;
  assign w6462 = \pi30 & \pi53 ;
  assign w6463 = \pi28 & \pi55 ;
  assign w6464 = ( w6461 & w6462 ) | ( w6461 & w6463 ) | ( w6462 & w6463 ) ;
  assign w6465 = w6461 ^ w6463 ;
  assign w6466 = w6462 ^ w6465 ;
  assign w6467 = \pi40 & \pi41 ;
  assign w6468 = w6298 & w6467 ;
  assign w6469 = ( \pi41 & \pi62 ) | ( \pi41 & w6467 ) | ( \pi62 & w6467 ) ;
  assign w6470 = ( \pi63 & w6298 ) | ( \pi63 & w6469 ) | ( w6298 & w6469 ) ;
  assign w6471 = ( \pi19 & w6468 ) | ( \pi19 & w6470 ) | ( w6468 & w6470 ) ;
  assign w6472 = w6460 ^ w6471 ;
  assign w6473 = w6466 ^ w6472 ;
  assign w6474 = ( w6416 & w6418 ) | ( w6416 & w6424 ) | ( w6418 & w6424 ) ;
  assign w6475 = w6473 ^ w6474 ;
  assign w6476 = w6453 ^ w6475 ;
  assign w6477 = w6447 ^ w6448 ;
  assign w6478 = w6476 ^ w6477 ;
  assign w6479 = w6401 ^ w6404 ;
  assign w6480 = ( w6392 & w6428 ) | ( w6392 & w6479 ) | ( w6428 & w6479 ) ;
  assign w6481 = ( w6405 & w6412 ) | ( w6405 & w6426 ) | ( w6412 & w6426 ) ;
  assign w6482 = ( w6401 & w6402 ) | ( w6401 & w6403 ) | ( w6402 & w6403 ) ;
  assign w6483 = \pi40 & \pi43 ;
  assign w6484 = \pi39 & \pi44 ;
  assign w6485 = \pi29 & \pi54 ;
  assign w6486 = ( w6483 & w6484 ) | ( w6483 & w6485 ) | ( w6484 & w6485 ) ;
  assign w6487 = w6483 ^ w6485 ;
  assign w6488 = w6484 ^ w6487 ;
  assign w6489 = \pi35 & \pi48 ;
  assign w6490 = \pi34 & \pi49 ;
  assign w6491 = \pi33 & \pi50 ;
  assign w6492 = ( w6489 & w6490 ) | ( w6489 & w6491 ) | ( w6490 & w6491 ) ;
  assign w6493 = w6489 ^ w6491 ;
  assign w6494 = w6490 ^ w6493 ;
  assign w6495 = ~\pi41 & \pi42 ;
  assign w6496 = w6488 ^ w6495 ;
  assign w6497 = w6494 ^ w6496 ;
  assign w6498 = \pi21 & \pi62 ;
  assign w6499 = w6497 ^ w6498 ;
  assign w6500 = ( w6393 & w6398 ) | ( w6393 & w6399 ) | ( w6398 & w6399 ) ;
  assign w6501 = \pi32 & \pi51 ;
  assign w6502 = \pi26 & \pi57 ;
  assign w6503 = \pi25 & \pi58 ;
  assign w6504 = ( w6501 & w6502 ) | ( w6501 & w6503 ) | ( w6502 & w6503 ) ;
  assign w6505 = w6501 ^ w6503 ;
  assign w6506 = w6502 ^ w6505 ;
  assign w6507 = \pi38 & \pi45 ;
  assign w6508 = \pi37 & \pi46 ;
  assign w6509 = \pi36 & \pi47 ;
  assign w6510 = ( w6507 & w6508 ) | ( w6507 & w6509 ) | ( w6508 & w6509 ) ;
  assign w6511 = w6507 ^ w6509 ;
  assign w6512 = w6508 ^ w6511 ;
  assign w6513 = \pi22 & \pi61 ;
  assign w6514 = \pi20 & \pi63 ;
  assign w6515 = ( w6058 & w6513 ) | ( w6058 & w6514 ) | ( w6513 & w6514 ) ;
  assign w6516 = w6058 ^ w6514 ;
  assign w6517 = w6513 ^ w6516 ;
  assign w6518 = w6506 ^ w6517 ;
  assign w6519 = w6512 ^ w6518 ;
  assign w6520 = w6500 ^ w6519 ;
  assign w6521 = w6499 ^ w6520 ;
  assign w6522 = w6481 ^ w6482 ;
  assign w6523 = w6521 ^ w6522 ;
  assign w6524 = w6478 ^ w6480 ;
  assign w6525 = w6523 ^ w6524 ;
  assign w6526 = ( w6341 & w6342 ) | ( w6341 & w6433 ) | ( w6342 & w6433 ) ;
  assign w6527 = w6436 ^ w6526 ;
  assign w6528 = w6525 ^ w6527 ;
  assign w6529 = ( w6436 & w6525 ) | ( w6436 & w6526 ) | ( w6525 & w6526 ) ;
  assign w6530 = ( w6478 & w6480 ) | ( w6478 & w6523 ) | ( w6480 & w6523 ) ;
  assign w6531 = ( w6447 & w6448 ) | ( w6447 & w6476 ) | ( w6448 & w6476 ) ;
  assign w6532 = \pi32 & \pi52 ;
  assign w6533 = \pi31 & \pi53 ;
  assign w6534 = \pi26 & \pi58 ;
  assign w6535 = ( w6532 & w6533 ) | ( w6532 & w6534 ) | ( w6533 & w6534 ) ;
  assign w6536 = w6532 ^ w6534 ;
  assign w6537 = w6533 ^ w6536 ;
  assign w6538 = ~\pi23 & w4299 ;
  assign w6539 = ( w4299 & w6457 ) | ( w4299 & ~w6538 ) | ( w6457 & ~w6538 ) ;
  assign w6540 = ( \pi24 & w6457 ) | ( \pi24 & w6539 ) | ( w6457 & w6539 ) ;
  assign w6541 = w6515 ^ w6537 ;
  assign w6542 = w6540 ^ w6541 ;
  assign w6543 = ( w6460 & w6466 ) | ( w6460 & w6471 ) | ( w6466 & w6471 ) ;
  assign w6544 = ( w6449 & w6450 ) | ( w6449 & w6451 ) | ( w6450 & w6451 ) ;
  assign w6545 = w6542 ^ w6543 ;
  assign w6546 = w6544 ^ w6545 ;
  assign w6547 = ( w6453 & w6473 ) | ( w6453 & w6474 ) | ( w6473 & w6474 ) ;
  assign w6548 = w6546 ^ w6547 ;
  assign w6549 = \pi23 & \pi61 ;
  assign w6550 = \pi22 & \pi62 ;
  assign w6551 = \pi21 & \pi63 ;
  assign w6552 = ( w6549 & w6550 ) | ( w6549 & w6551 ) | ( w6550 & w6551 ) ;
  assign w6553 = w6549 ^ w6551 ;
  assign w6554 = w6550 ^ w6553 ;
  assign w6555 = \pi33 & \pi51 ;
  assign w6556 = \pi25 & \pi59 ;
  assign w6557 = \pi24 & \pi60 ;
  assign w6558 = ( w6555 & w6556 ) | ( w6555 & w6557 ) | ( w6556 & w6557 ) ;
  assign w6559 = w6555 ^ w6557 ;
  assign w6560 = w6556 ^ w6559 ;
  assign w6561 = \pi36 & \pi48 ;
  assign w6562 = \pi35 & \pi49 ;
  assign w6563 = \pi34 & \pi50 ;
  assign w6564 = ( w6561 & w6562 ) | ( w6561 & w6563 ) | ( w6562 & w6563 ) ;
  assign w6565 = w6561 ^ w6563 ;
  assign w6566 = w6562 ^ w6565 ;
  assign w6567 = w6554 ^ w6560 ;
  assign w6568 = w6566 ^ w6567 ;
  assign w6569 = \pi38 & \pi56 ;
  assign w6570 = \pi38 & \pi46 ;
  assign w6571 = \pi29 & \pi55 ;
  assign w6572 = \pi28 & \pi56 ;
  assign w6573 = ( w6570 & w6571 ) | ( w6570 & w6572 ) | ( w6571 & w6572 ) ;
  assign w6574 = w6570 ^ w6572 ;
  assign w6575 = w6571 ^ w6574 ;
  assign w6576 = \pi41 & \pi43 ;
  assign w6577 = \pi40 & \pi44 ;
  assign w6578 = \pi39 & \pi45 ;
  assign w6579 = ( w6576 & w6577 ) | ( w6576 & w6578 ) | ( w6577 & w6578 ) ;
  assign w6580 = w6576 ^ w6578 ;
  assign w6581 = w6577 ^ w6580 ;
  assign w6582 = \pi30 & \pi54 ;
  assign w6583 = \pi27 & \pi57 ;
  assign w6584 = ( w6379 & w6582 ) | ( w6379 & w6583 ) | ( w6582 & w6583 ) ;
  assign w6585 = w6379 ^ w6583 ;
  assign w6586 = w6582 ^ w6585 ;
  assign w6587 = w6575 ^ w6586 ;
  assign w6588 = w6581 ^ w6587 ;
  assign w6589 = w6492 ^ w6504 ;
  assign w6590 = w6510 ^ w6589 ;
  assign w6591 = ( w6362 & w6371 ) | ( w6362 & w6383 ) | ( w6371 & w6383 ) ;
  assign w6592 = ( w6350 & w6356 ) | ( w6350 & w6396 ) | ( w6356 & w6396 ) ;
  assign w6593 = w6590 ^ w6591 ;
  assign w6594 = w6592 ^ w6593 ;
  assign w6595 = w6588 ^ w6594 ;
  assign w6596 = w6568 ^ w6595 ;
  assign w6597 = w6548 & w6596 ;
  assign w6598 = w6548 | w6596 ;
  assign w6599 = ( w6481 & w6482 ) | ( w6481 & w6521 ) | ( w6482 & w6521 ) ;
  assign w6600 = ( w6437 & w6438 ) | ( w6437 & w6445 ) | ( w6438 & w6445 ) ;
  assign w6601 = w6599 ^ w6600 ;
  assign w6602 = ( w6499 & w6500 ) | ( w6499 & w6519 ) | ( w6500 & w6519 ) ;
  assign w6603 = ( w6440 & w6442 ) | ( w6440 & w6443 ) | ( w6442 & w6443 ) ;
  assign w6604 = w6464 ^ w6486 ;
  assign w6605 = ( \pi21 & \pi41 ) | ( \pi21 & \pi62 ) | ( \pi41 & \pi62 ) ;
  assign w6606 = ~\pi41 & w6605 ;
  assign w6607 = ( \pi41 & \pi42 ) | ( \pi41 & w6606 ) | ( \pi42 & w6606 ) ;
  assign w6608 = w6604 ^ w6607 ;
  assign w6609 = ( w6506 & w6512 ) | ( w6506 & w6517 ) | ( w6512 & w6517 ) ;
  assign w6610 = w6495 ^ w6498 ;
  assign w6611 = ( w6488 & w6494 ) | ( w6488 & w6610 ) | ( w6494 & w6610 ) ;
  assign w6612 = w6608 ^ w6609 ;
  assign w6613 = w6611 ^ w6612 ;
  assign w6614 = w6602 ^ w6603 ;
  assign w6615 = w6613 ^ w6614 ;
  assign w6616 = ~w6597 & w6598 ;
  assign w6617 = w6531 ^ w6615 ;
  assign w6618 = w6601 ^ w6617 ;
  assign w6619 = w6616 ^ w6618 ;
  assign w6620 = w6529 ^ w6530 ;
  assign w6621 = w6619 ^ w6620 ;
  assign w6622 = ( w6529 & w6530 ) | ( w6529 & w6619 ) | ( w6530 & w6619 ) ;
  assign w6623 = w6601 ^ w6615 ;
  assign w6624 = ( w6531 & w6616 ) | ( w6531 & w6623 ) | ( w6616 & w6623 ) ;
  assign w6625 = ( w6599 & w6600 ) | ( w6599 & w6615 ) | ( w6600 & w6615 ) ;
  assign w6626 = \pi35 & \pi50 ;
  assign w6627 = \pi28 & \pi57 ;
  assign w6628 = \pi22 & \pi63 ;
  assign w6629 = ( w6626 & w6627 ) | ( w6626 & w6628 ) | ( w6627 & w6628 ) ;
  assign w6630 = w6626 ^ w6628 ;
  assign w6631 = w6627 ^ w6630 ;
  assign w6632 = \pi34 & \pi51 ;
  assign w6633 = \pi33 & \pi52 ;
  assign w6634 = \pi32 & \pi53 ;
  assign w6635 = ( w6632 & w6633 ) | ( w6632 & w6634 ) | ( w6633 & w6634 ) ;
  assign w6636 = w6632 ^ w6634 ;
  assign w6637 = w6633 ^ w6636 ;
  assign w6638 = \pi41 & \pi44 ;
  assign w6639 = \pi40 & \pi45 ;
  assign w6640 = \pi39 & \pi46 ;
  assign w6641 = ( w6638 & w6639 ) | ( w6638 & w6640 ) | ( w6639 & w6640 ) ;
  assign w6642 = w6638 ^ w6640 ;
  assign w6643 = w6639 ^ w6642 ;
  assign w6644 = w6631 ^ w6637 ;
  assign w6645 = w6643 ^ w6644 ;
  assign w6646 = \pi23 & \pi62 ;
  assign w6647 = \pi42 & ~w6646 ;
  assign w6648 = ( \pi43 & w6646 ) | ( \pi43 & w6647 ) | ( w6646 & w6647 ) ;
  assign w6649 = \pi38 & \pi47 ;
  assign w6650 = \pi37 & \pi48 ;
  assign w6651 = \pi36 & \pi49 ;
  assign w6652 = ( w6649 & w6650 ) | ( w6649 & w6651 ) | ( w6650 & w6651 ) ;
  assign w6653 = w6649 ^ w6651 ;
  assign w6654 = w6650 ^ w6653 ;
  assign w6655 = \pi31 & \pi54 ;
  assign w6656 = \pi30 & \pi55 ;
  assign w6657 = \pi29 & \pi56 ;
  assign w6658 = ( w6655 & w6656 ) | ( w6655 & w6657 ) | ( w6656 & w6657 ) ;
  assign w6659 = w6655 ^ w6657 ;
  assign w6660 = w6656 ^ w6659 ;
  assign w6661 = ~\pi42 & \pi43 ;
  assign w6662 = w6654 ^ w6661 ;
  assign w6663 = w6660 ^ w6662 ;
  assign w6664 = w6646 ^ w6663 ;
  assign w6665 = ( w6608 & w6609 ) | ( w6608 & w6611 ) | ( w6609 & w6611 ) ;
  assign w6666 = w6645 ^ w6665 ;
  assign w6667 = w6664 ^ w6666 ;
  assign w6668 = ( w6590 & w6591 ) | ( w6590 & w6592 ) | ( w6591 & w6592 ) ;
  assign w6669 = \pi27 & \pi58 ;
  assign w6670 = \pi26 & \pi59 ;
  assign w6671 = \pi25 & \pi60 ;
  assign w6672 = ( w6669 & w6670 ) | ( w6669 & w6671 ) | ( w6670 & w6671 ) ;
  assign w6673 = w6669 ^ w6671 ;
  assign w6674 = w6670 ^ w6673 ;
  assign w6675 = w6535 ^ w6584 ;
  assign w6676 = w6674 ^ w6675 ;
  assign w6677 = w6573 ^ w6579 ;
  assign w6678 = \pi24 & \pi61 ;
  assign w6679 = w6677 ^ w6678 ;
  assign w6680 = ( w6668 & w6676 ) | ( w6668 & w6679 ) | ( w6676 & w6679 ) ;
  assign w6681 = w6668 ^ w6676 ;
  assign w6682 = w6573 ^ w6681 ;
  assign w6683 = w6579 ^ w6682 ;
  assign w6684 = w6678 ^ w6683 ;
  assign w6685 = w6552 ^ w6558 ;
  assign w6686 = w6564 ^ w6685 ;
  assign w6687 = ( w6575 & w6581 ) | ( w6575 & w6586 ) | ( w6581 & w6586 ) ;
  assign w6688 = ( w6554 & w6560 ) | ( w6554 & w6566 ) | ( w6560 & w6566 ) ;
  assign w6689 = w6686 ^ w6687 ;
  assign w6690 = w6688 ^ w6689 ;
  assign w6691 = w6667 ^ w6684 ;
  assign w6692 = w6690 ^ w6691 ;
  assign w6693 = ( w6602 & w6603 ) | ( w6602 & w6613 ) | ( w6603 & w6613 ) ;
  assign w6694 = ( w6492 & w6504 ) | ( w6492 & w6510 ) | ( w6504 & w6510 ) ;
  assign w6695 = \pi41 & \pi42 ;
  assign w6696 = ( \pi42 & w6605 ) | ( \pi42 & w6695 ) | ( w6605 & w6695 ) ;
  assign w6697 = ( w6464 & w6486 ) | ( w6464 & w6696 ) | ( w6486 & w6696 ) ;
  assign w6698 = \pi23 | w6457 ;
  assign w6699 = ( \pi24 & w6457 ) | ( \pi24 & w6698 ) | ( w6457 & w6698 ) ;
  assign w6700 = ( w4299 & w6457 ) | ( w4299 & w6699 ) | ( w6457 & w6699 ) ;
  assign w6701 = ( w6515 & w6537 ) | ( w6515 & w6700 ) | ( w6537 & w6700 ) ;
  assign w6702 = w6694 ^ w6701 ;
  assign w6703 = w6697 ^ w6702 ;
  assign w6704 = ( w6542 & w6543 ) | ( w6542 & w6544 ) | ( w6543 & w6544 ) ;
  assign w6705 = ( w6568 & w6588 ) | ( w6568 & w6594 ) | ( w6588 & w6594 ) ;
  assign w6706 = w6703 ^ w6704 ;
  assign w6707 = w6705 ^ w6706 ;
  assign w6708 = ( w6546 & w6547 ) | ( w6546 & w6596 ) | ( w6547 & w6596 ) ;
  assign w6709 = w6693 ^ w6707 ;
  assign w6710 = w6708 ^ w6709 ;
  assign w6711 = w6625 ^ w6710 ;
  assign w6712 = w6692 ^ w6711 ;
  assign w6713 = w6622 ^ w6624 ;
  assign w6714 = w6712 ^ w6713 ;
  assign w6715 = ( w6622 & w6624 ) | ( w6622 & w6712 ) | ( w6624 & w6712 ) ;
  assign w6716 = ( w6625 & w6692 ) | ( w6625 & w6710 ) | ( w6692 & w6710 ) ;
  assign w6717 = ( w6693 & w6707 ) | ( w6693 & w6708 ) | ( w6707 & w6708 ) ;
  assign w6718 = ( w6535 & w6584 ) | ( w6535 & w6674 ) | ( w6584 & w6674 ) ;
  assign w6719 = ( w6631 & w6637 ) | ( w6631 & w6643 ) | ( w6637 & w6643 ) ;
  assign w6720 = w6646 ^ w6661 ;
  assign w6721 = ( w6654 & w6660 ) | ( w6654 & w6720 ) | ( w6660 & w6720 ) ;
  assign w6722 = w6718 ^ w6719 ;
  assign w6723 = w6721 ^ w6722 ;
  assign w6724 = ( w6694 & w6697 ) | ( w6694 & w6701 ) | ( w6697 & w6701 ) ;
  assign w6725 = w6641 ^ w6652 ;
  assign w6726 = w6658 ^ w6725 ;
  assign w6727 = w6629 ^ w6635 ;
  assign w6728 = w6672 ^ w6727 ;
  assign w6729 = w6724 ^ w6726 ;
  assign w6730 = w6728 ^ w6729 ;
  assign w6731 = ( w6686 & w6687 ) | ( w6686 & w6688 ) | ( w6687 & w6688 ) ;
  assign w6732 = \pi37 & \pi49 ;
  assign w6733 = \pi36 & \pi50 ;
  assign w6734 = \pi23 & \pi63 ;
  assign w6735 = ( w6732 & w6733 ) | ( w6732 & w6734 ) | ( w6733 & w6734 ) ;
  assign w6736 = w6732 ^ w6734 ;
  assign w6737 = w6733 ^ w6736 ;
  assign w6738 = \pi35 & \pi51 ;
  assign w6739 = \pi34 & \pi52 ;
  assign w6740 = \pi33 & \pi53 ;
  assign w6741 = ( w6738 & w6739 ) | ( w6738 & w6740 ) | ( w6739 & w6740 ) ;
  assign w6742 = w6738 ^ w6740 ;
  assign w6743 = w6739 ^ w6742 ;
  assign w6744 = \pi31 & \pi55 ;
  assign w6745 = \pi29 & \pi57 ;
  assign w6746 = ( w3176 & w6744 ) | ( w3176 & w6745 ) | ( w6744 & w6745 ) ;
  assign w6747 = w3176 ^ w6745 ;
  assign w6748 = w6744 ^ w6747 ;
  assign w6749 = w6737 ^ w6748 ;
  assign w6750 = w6743 ^ w6749 ;
  assign w6751 = \pi28 & \pi58 ;
  assign w6752 = \pi27 & \pi59 ;
  assign w6753 = \pi26 & \pi60 ;
  assign w6754 = ( w6751 & w6752 ) | ( w6751 & w6753 ) | ( w6752 & w6753 ) ;
  assign w6755 = w6751 ^ w6753 ;
  assign w6756 = w6752 ^ w6755 ;
  assign w6757 = \pi32 & \pi54 ;
  assign w6758 = \pi42 & \pi44 ;
  assign w6759 = \pi41 & \pi45 ;
  assign w6760 = ( w6757 & w6758 ) | ( w6757 & w6759 ) | ( w6758 & w6759 ) ;
  assign w6761 = w6757 ^ w6759 ;
  assign w6762 = w6758 ^ w6761 ;
  assign w6763 = \pi40 & \pi46 ;
  assign w6764 = \pi39 & \pi47 ;
  assign w6765 = \pi30 & \pi56 ;
  assign w6766 = ( w6763 & w6764 ) | ( w6763 & w6765 ) | ( w6764 & w6765 ) ;
  assign w6767 = w6763 ^ w6765 ;
  assign w6768 = w6764 ^ w6767 ;
  assign w6769 = w6756 ^ w6762 ;
  assign w6770 = w6768 ^ w6769 ;
  assign w6771 = w6731 ^ w6750 ;
  assign w6772 = w6770 ^ w6771 ;
  assign w6773 = w6730 ^ w6772 ;
  assign w6774 = w6723 ^ w6773 ;
  assign w6775 = ( w6667 & w6684 ) | ( w6667 & w6690 ) | ( w6684 & w6690 ) ;
  assign w6776 = ( w6703 & w6704 ) | ( w6703 & w6705 ) | ( w6704 & w6705 ) ;
  assign w6777 = \pi25 & \pi61 ;
  assign w6778 = \pi24 & \pi62 ;
  assign w6779 = w6648 ^ w6778 ;
  assign w6780 = w6777 ^ w6779 ;
  assign w6781 = ( w6552 & w6558 ) | ( w6552 & w6564 ) | ( w6558 & w6564 ) ;
  assign w6782 = ( w6573 & w6579 ) | ( w6573 & w6678 ) | ( w6579 & w6678 ) ;
  assign w6783 = w6780 ^ w6782 ;
  assign w6784 = w6781 ^ w6783 ;
  assign w6785 = ( w6645 & w6664 ) | ( w6645 & w6665 ) | ( w6664 & w6665 ) ;
  assign w6786 = w6680 ^ w6785 ;
  assign w6787 = w6784 ^ w6786 ;
  assign w6788 = w6775 ^ w6776 ;
  assign w6789 = w6787 ^ w6788 ;
  assign w6790 = w6717 ^ w6774 ;
  assign w6791 = w6789 ^ w6790 ;
  assign w6792 = w6716 | w6791 ;
  assign w6793 = w6716 & w6791 ;
  assign w6794 = w6792 & ~w6793 ;
  assign w6795 = w6715 ^ w6794 ;
  assign w6796 = ( w6715 & w6792 ) | ( w6715 & w6793 ) | ( w6792 & w6793 ) ;
  assign w6797 = w6793 | w6796 ;
  assign w6798 = ( w6717 & w6774 ) | ( w6717 & w6789 ) | ( w6774 & w6789 ) ;
  assign w6799 = ( w6731 & w6750 ) | ( w6731 & w6770 ) | ( w6750 & w6770 ) ;
  assign w6800 = ( w6641 & w6652 ) | ( w6641 & w6658 ) | ( w6652 & w6658 ) ;
  assign w6801 = ( w6737 & w6743 ) | ( w6737 & w6748 ) | ( w6743 & w6748 ) ;
  assign w6802 = ( w6756 & w6762 ) | ( w6756 & w6768 ) | ( w6762 & w6768 ) ;
  assign w6803 = w6801 ^ w6802 ;
  assign w6804 = w6800 ^ w6803 ;
  assign w6805 = ( w6680 & w6784 ) | ( w6680 & w6785 ) | ( w6784 & w6785 ) ;
  assign w6806 = w6799 ^ w6805 ;
  assign w6807 = w6804 ^ w6806 ;
  assign w6808 = ( w6775 & w6776 ) | ( w6775 & w6787 ) | ( w6776 & w6787 ) ;
  assign w6809 = ( w6724 & w6726 ) | ( w6724 & w6728 ) | ( w6726 & w6728 ) ;
  assign w6810 = ( w6718 & w6719 ) | ( w6718 & w6721 ) | ( w6719 & w6721 ) ;
  assign w6811 = w6809 ^ w6810 ;
  assign w6812 = ( w6780 & w6781 ) | ( w6780 & w6782 ) | ( w6781 & w6782 ) ;
  assign w6813 = w6746 ^ w6760 ;
  assign w6814 = w6766 ^ w6813 ;
  assign w6815 = w6735 ^ w6741 ;
  assign w6816 = w6754 ^ w6815 ;
  assign w6817 = w6812 ^ w6814 ;
  assign w6818 = w6816 ^ w6817 ;
  assign w6819 = ( w6723 & w6730 ) | ( w6723 & w6772 ) | ( w6730 & w6772 ) ;
  assign w6820 = \pi40 & \pi47 ;
  assign w6821 = \pi33 & \pi54 ;
  assign w6822 = \pi31 & \pi56 ;
  assign w6823 = ( w6820 & w6821 ) | ( w6820 & w6822 ) | ( w6821 & w6822 ) ;
  assign w6824 = w6820 ^ w6822 ;
  assign w6825 = w6821 ^ w6824 ;
  assign w6826 = ( w6629 & w6635 ) | ( w6629 & w6672 ) | ( w6635 & w6672 ) ;
  assign w6827 = ~\pi43 & \pi44 ;
  assign w6828 = w6826 ^ w6827 ;
  assign w6829 = w6825 ^ w6828 ;
  assign w6830 = \pi25 & \pi62 ;
  assign w6831 = w6829 ^ w6830 ;
  assign w6832 = \pi27 & \pi60 ;
  assign w6833 = \pi26 & \pi61 ;
  assign w6834 = \pi24 & \pi63 ;
  assign w6835 = ( w6832 & w6833 ) | ( w6832 & w6834 ) | ( w6833 & w6834 ) ;
  assign w6836 = w6832 ^ w6834 ;
  assign w6837 = w6833 ^ w6836 ;
  assign w6838 = \pi39 & \pi48 ;
  assign w6839 = \pi38 & \pi49 ;
  assign w6840 = \pi37 & \pi50 ;
  assign w6841 = ( w6838 & w6839 ) | ( w6838 & w6840 ) | ( w6839 & w6840 ) ;
  assign w6842 = w6838 ^ w6840 ;
  assign w6843 = w6839 ^ w6842 ;
  assign w6844 = \pi42 & \pi45 ;
  assign w6845 = \pi41 & \pi46 ;
  assign w6846 = \pi32 & \pi55 ;
  assign w6847 = ( w6844 & w6845 ) | ( w6844 & w6846 ) | ( w6845 & w6846 ) ;
  assign w6848 = w6844 ^ w6846 ;
  assign w6849 = w6845 ^ w6848 ;
  assign w6850 = w6837 ^ w6843 ;
  assign w6851 = w6849 ^ w6850 ;
  assign w6852 = \pi34 & \pi59 ;
  assign w6853 = \pi34 & \pi53 ;
  assign w6854 = \pi30 & \pi57 ;
  assign w6855 = \pi28 & \pi59 ;
  assign w6856 = ( w6853 & w6854 ) | ( w6853 & w6855 ) | ( w6854 & w6855 ) ;
  assign w6857 = w6853 ^ w6855 ;
  assign w6858 = w6854 ^ w6857 ;
  assign w6859 = ( w6648 & w6777 ) | ( w6648 & w6778 ) | ( w6777 & w6778 ) ;
  assign w6860 = \pi36 & \pi51 ;
  assign w6861 = \pi35 & \pi52 ;
  assign w6862 = \pi29 & \pi58 ;
  assign w6863 = ( w6860 & w6861 ) | ( w6860 & w6862 ) | ( w6861 & w6862 ) ;
  assign w6864 = w6860 ^ w6862 ;
  assign w6865 = w6861 ^ w6864 ;
  assign w6866 = w6858 ^ w6859 ;
  assign w6867 = w6865 ^ w6866 ;
  assign w6868 = w6831 ^ w6867 ;
  assign w6869 = w6851 ^ w6868 ;
  assign w6870 = w6818 ^ w6869 ;
  assign w6871 = w6811 ^ w6870 ;
  assign w6872 = w6819 ^ w6871 ;
  assign w6873 = w6807 ^ w6872 ;
  assign w6874 = w6808 ^ w6873 ;
  assign w6875 = w6797 ^ w6874 ;
  assign w6876 = w6798 ^ w6875 ;
  assign w6877 = ( w6807 & w6808 ) | ( w6807 & w6872 ) | ( w6808 & w6872 ) ;
  assign w6878 = ( w6799 & w6804 ) | ( w6799 & w6805 ) | ( w6804 & w6805 ) ;
  assign w6879 = \pi28 & \pi60 ;
  assign w6880 = \pi27 & \pi61 ;
  assign w6881 = \pi26 & \pi62 ;
  assign w6882 = ( w6879 & w6880 ) | ( w6879 & w6881 ) | ( w6880 & w6881 ) ;
  assign w6883 = w6879 ^ w6881 ;
  assign w6884 = w6880 ^ w6883 ;
  assign w6885 = \pi42 & \pi46 ;
  assign w6886 = \pi41 & \pi47 ;
  assign w6887 = \pi31 & \pi57 ;
  assign w6888 = ( w6885 & w6886 ) | ( w6885 & w6887 ) | ( w6886 & w6887 ) ;
  assign w6889 = w6885 ^ w6887 ;
  assign w6890 = w6886 ^ w6889 ;
  assign w6891 = \pi37 & \pi51 ;
  assign w6892 = \pi36 & \pi52 ;
  assign w6893 = \pi35 & \pi53 ;
  assign w6894 = ( w6891 & w6892 ) | ( w6891 & w6893 ) | ( w6892 & w6893 ) ;
  assign w6895 = w6891 ^ w6893 ;
  assign w6896 = w6892 ^ w6895 ;
  assign w6897 = w6884 ^ w6890 ;
  assign w6898 = w6896 ^ w6897 ;
  assign w6899 = \pi39 & \pi49 ;
  assign w6900 = \pi38 & \pi50 ;
  assign w6901 = ( w4082 & w6899 ) | ( w4082 & w6900 ) | ( w6899 & w6900 ) ;
  assign w6902 = w4082 ^ w6899 ;
  assign w6903 = w6900 ^ w6902 ;
  assign w6904 = \pi40 & \pi48 ;
  assign w6905 = \pi32 & \pi56 ;
  assign w6906 = \pi30 & \pi58 ;
  assign w6907 = ( w6904 & w6905 ) | ( w6904 & w6906 ) | ( w6905 & w6906 ) ;
  assign w6908 = w6904 ^ w6906 ;
  assign w6909 = w6905 ^ w6908 ;
  assign w6910 = ( w6746 & w6760 ) | ( w6746 & w6766 ) | ( w6760 & w6766 ) ;
  assign w6911 = w6903 ^ w6910 ;
  assign w6912 = w6909 ^ w6911 ;
  assign w6913 = \pi25 & \pi63 ;
  assign w6914 = w6847 ^ w6913 ;
  assign w6915 = ~\pi43 & \pi62 ;
  assign w6916 = \pi25 & w6915 ;
  assign w6917 = ( \pi43 & \pi44 ) | ( \pi43 & w6916 ) | ( \pi44 & w6916 ) ;
  assign w6918 = w6914 ^ w6917 ;
  assign w6919 = w6898 ^ w6912 ;
  assign w6920 = w6918 ^ w6919 ;
  assign w6921 = ( w6812 & w6814 ) | ( w6812 & w6816 ) | ( w6814 & w6816 ) ;
  assign w6922 = ( w6800 & w6801 ) | ( w6800 & w6802 ) | ( w6801 & w6802 ) ;
  assign w6923 = w6835 ^ w6841 ;
  assign w6924 = w6856 ^ w6923 ;
  assign w6925 = \pi43 & \pi45 ;
  assign w6926 = \pi34 & \pi54 ;
  assign w6927 = \pi33 & \pi55 ;
  assign w6928 = ( w6925 & w6926 ) | ( w6925 & w6927 ) | ( w6926 & w6927 ) ;
  assign w6929 = w6925 ^ w6927 ;
  assign w6930 = w6926 ^ w6929 ;
  assign w6931 = w6823 ^ w6863 ;
  assign w6932 = w6930 ^ w6931 ;
  assign w6933 = w6827 ^ w6830 ;
  assign w6934 = ( w6825 & w6826 ) | ( w6825 & w6933 ) | ( w6826 & w6933 ) ;
  assign w6935 = w6924 ^ w6934 ;
  assign w6936 = w6932 ^ w6935 ;
  assign w6937 = w6921 ^ w6922 ;
  assign w6938 = w6936 ^ w6937 ;
  assign w6939 = w6878 ^ w6920 ;
  assign w6940 = w6938 ^ w6939 ;
  assign w6941 = w6811 ^ w6818 ;
  assign w6942 = ( w6819 & w6869 ) | ( w6819 & w6941 ) | ( w6869 & w6941 ) ;
  assign w6943 = ( w6809 & w6810 ) | ( w6809 & w6818 ) | ( w6810 & w6818 ) ;
  assign w6944 = ( w6735 & w6741 ) | ( w6735 & w6754 ) | ( w6741 & w6754 ) ;
  assign w6945 = ( w6858 & w6859 ) | ( w6858 & w6865 ) | ( w6859 & w6865 ) ;
  assign w6946 = ( w6837 & w6843 ) | ( w6837 & w6849 ) | ( w6843 & w6849 ) ;
  assign w6947 = w6944 ^ w6945 ;
  assign w6948 = w6946 ^ w6947 ;
  assign w6949 = ( w6831 & w6851 ) | ( w6831 & w6867 ) | ( w6851 & w6867 ) ;
  assign w6950 = w6943 ^ w6948 ;
  assign w6951 = w6949 ^ w6950 ;
  assign w6952 = w6940 ^ w6942 ;
  assign w6953 = w6951 ^ w6952 ;
  assign w6954 = ( w6797 & w6798 ) | ( w6797 & w6874 ) | ( w6798 & w6874 ) ;
  assign w6955 = w6877 ^ w6954 ;
  assign w6956 = w6953 ^ w6955 ;
  assign w6957 = ( w6940 & w6942 ) | ( w6940 & w6951 ) | ( w6942 & w6951 ) ;
  assign w6958 = ( w6943 & w6948 ) | ( w6943 & w6949 ) | ( w6948 & w6949 ) ;
  assign w6959 = \pi41 & \pi48 ;
  assign w6960 = \pi35 & \pi54 ;
  assign w6961 = \pi33 & \pi56 ;
  assign w6962 = ( w6959 & w6960 ) | ( w6959 & w6961 ) | ( w6960 & w6961 ) ;
  assign w6963 = w6959 ^ w6961 ;
  assign w6964 = w6960 ^ w6963 ;
  assign w6965 = \pi38 & \pi51 ;
  assign w6966 = \pi37 & \pi52 ;
  assign w6967 = \pi36 & \pi53 ;
  assign w6968 = ( w6965 & w6966 ) | ( w6965 & w6967 ) | ( w6966 & w6967 ) ;
  assign w6969 = w6965 ^ w6967 ;
  assign w6970 = w6966 ^ w6969 ;
  assign w6971 = \pi32 & \pi57 ;
  assign w6972 = \pi31 & \pi58 ;
  assign w6973 = \pi30 & \pi59 ;
  assign w6974 = ( w6971 & w6972 ) | ( w6971 & w6973 ) | ( w6972 & w6973 ) ;
  assign w6975 = w6971 ^ w6973 ;
  assign w6976 = w6972 ^ w6975 ;
  assign w6977 = w6964 ^ w6970 ;
  assign w6978 = w6976 ^ w6977 ;
  assign w6979 = w6882 ^ w6894 ;
  assign w6980 = w6907 ^ w6979 ;
  assign w6981 = \pi43 & \pi46 ;
  assign w6982 = \pi42 & \pi47 ;
  assign w6983 = \pi34 & \pi55 ;
  assign w6984 = ( w6981 & w6982 ) | ( w6981 & w6983 ) | ( w6982 & w6983 ) ;
  assign w6985 = w6981 ^ w6983 ;
  assign w6986 = w6982 ^ w6985 ;
  assign w6987 = \pi29 & \pi60 ;
  assign w6988 = ( \pi28 & \pi61 ) | ( \pi28 & ~w6928 ) | ( \pi61 & ~w6928 ) ;
  assign w6989 = w6987 ^ w6988 ;
  assign w6990 = w6928 & w6989 ;
  assign w6991 = \pi28 & \pi61 ;
  assign w6992 = w6928 ^ w6991 ;
  assign w6993 = w6987 ^ w6992 ;
  assign w6994 = ~\pi44 & \pi45 ;
  assign w6995 = w6993 ^ w6994 ;
  assign w6996 = w6986 ^ w6995 ;
  assign w6997 = \pi27 & \pi62 ;
  assign w6998 = w6996 ^ w6997 ;
  assign w6999 = w6978 ^ w6998 ;
  assign w7000 = w6980 ^ w6999 ;
  assign w7001 = ( w6835 & w6841 ) | ( w6835 & w6856 ) | ( w6841 & w6856 ) ;
  assign w7002 = \pi43 & \pi44 ;
  assign w7003 = w6847 & w7002 ;
  assign w7004 = ( \pi44 & \pi62 ) | ( \pi44 & w7002 ) | ( \pi62 & w7002 ) ;
  assign w7005 = ( \pi63 & w6847 ) | ( \pi63 & w7004 ) | ( w6847 & w7004 ) ;
  assign w7006 = ( \pi25 & w7003 ) | ( \pi25 & w7005 ) | ( w7003 & w7005 ) ;
  assign w7007 = ( w6823 & w6863 ) | ( w6823 & w6930 ) | ( w6863 & w6930 ) ;
  assign w7008 = w7001 ^ w7006 ;
  assign w7009 = w7007 ^ w7008 ;
  assign w7010 = ( w6944 & w6945 ) | ( w6944 & w6946 ) | ( w6945 & w6946 ) ;
  assign w7011 = ( w6924 & w6932 ) | ( w6924 & w6934 ) | ( w6932 & w6934 ) ;
  assign w7012 = w7010 ^ w7011 ;
  assign w7013 = w7009 ^ w7012 ;
  assign w7014 = w6958 ^ w7013 ;
  assign w7015 = w7000 ^ w7014 ;
  assign w7016 = ( w6878 & w6920 ) | ( w6878 & w6938 ) | ( w6920 & w6938 ) ;
  assign w7017 = ( w6921 & w6922 ) | ( w6921 & w6936 ) | ( w6922 & w6936 ) ;
  assign w7018 = ( w6898 & w6912 ) | ( w6898 & w6918 ) | ( w6912 & w6918 ) ;
  assign w7019 = ( w6903 & w6909 ) | ( w6903 & w6910 ) | ( w6909 & w6910 ) ;
  assign w7020 = ( w6884 & w6890 ) | ( w6884 & w6896 ) | ( w6890 & w6896 ) ;
  assign w7021 = \pi40 & \pi49 ;
  assign w7022 = \pi39 & \pi50 ;
  assign w7023 = \pi26 & \pi63 ;
  assign w7024 = ( w7021 & w7022 ) | ( w7021 & w7023 ) | ( w7022 & w7023 ) ;
  assign w7025 = w7021 ^ w7023 ;
  assign w7026 = w7022 ^ w7025 ;
  assign w7027 = w6888 ^ w6901 ;
  assign w7028 = w7026 ^ w7027 ;
  assign w7029 = w7019 ^ w7020 ;
  assign w7030 = w7028 ^ w7029 ;
  assign w7031 = w7017 ^ w7018 ;
  assign w7032 = w7030 ^ w7031 ;
  assign w7033 = w7015 ^ w7016 ;
  assign w7034 = w7032 ^ w7033 ;
  assign w7035 = ( w6877 & w6953 ) | ( w6877 & w6954 ) | ( w6953 & w6954 ) ;
  assign w7036 = w7034 ^ w7035 ;
  assign w7037 = w6957 ^ w7036 ;
  assign w7038 = ( w6957 & w7034 ) | ( w6957 & w7035 ) | ( w7034 & w7035 ) ;
  assign w7039 = ( w7015 & w7016 ) | ( w7015 & w7032 ) | ( w7016 & w7032 ) ;
  assign w7040 = ( w7009 & w7010 ) | ( w7009 & w7011 ) | ( w7010 & w7011 ) ;
  assign w7041 = ( w6978 & w6980 ) | ( w6978 & w6998 ) | ( w6980 & w6998 ) ;
  assign w7042 = w6962 ^ w6984 ;
  assign w7043 = ( \pi27 & \pi44 ) | ( \pi27 & \pi62 ) | ( \pi44 & \pi62 ) ;
  assign w7044 = ~\pi44 & w7043 ;
  assign w7045 = ( \pi44 & \pi45 ) | ( \pi44 & w7044 ) | ( \pi45 & w7044 ) ;
  assign w7046 = w7042 ^ w7045 ;
  assign w7047 = w6994 ^ w6997 ;
  assign w7048 = ( w6986 & w6993 ) | ( w6986 & w7047 ) | ( w6993 & w7047 ) ;
  assign w7049 = ( w6964 & w6970 ) | ( w6964 & w6976 ) | ( w6970 & w6976 ) ;
  assign w7050 = w7046 ^ w7048 ;
  assign w7051 = w7049 ^ w7050 ;
  assign w7052 = w7040 ^ w7041 ;
  assign w7053 = w7051 ^ w7052 ;
  assign w7054 = ( w6958 & w7000 ) | ( w6958 & w7013 ) | ( w7000 & w7013 ) ;
  assign w7055 = ( w7017 & w7018 ) | ( w7017 & w7030 ) | ( w7018 & w7030 ) ;
  assign w7056 = w6968 ^ w6974 ;
  assign w7057 = w7024 ^ w7056 ;
  assign w7058 = ( w7001 & w7006 ) | ( w7001 & w7007 ) | ( w7006 & w7007 ) ;
  assign w7059 = w7057 ^ w7058 ;
  assign w7060 = \pi35 & \pi55 ;
  assign w7061 = \pi34 & \pi56 ;
  assign w7062 = \pi33 & \pi57 ;
  assign w7063 = ( w7060 & w7061 ) | ( w7060 & w7062 ) | ( w7061 & w7062 ) ;
  assign w7064 = w7060 ^ w7062 ;
  assign w7065 = w7061 ^ w7064 ;
  assign w7066 = \pi38 & \pi52 ;
  assign w7067 = \pi37 & \pi53 ;
  assign w7068 = \pi36 & \pi54 ;
  assign w7069 = ( w7066 & w7067 ) | ( w7066 & w7068 ) | ( w7067 & w7068 ) ;
  assign w7070 = w7066 ^ w7068 ;
  assign w7071 = w7067 ^ w7070 ;
  assign w7072 = \pi44 & \pi46 ;
  assign w7073 = \pi43 & \pi47 ;
  assign w7074 = \pi42 & \pi48 ;
  assign w7075 = ( w7072 & w7073 ) | ( w7072 & w7074 ) | ( w7073 & w7074 ) ;
  assign w7076 = w7072 ^ w7074 ;
  assign w7077 = w7073 ^ w7076 ;
  assign w7078 = w7065 ^ w7071 ;
  assign w7079 = w7077 ^ w7078 ;
  assign w7080 = ( w7019 & w7020 ) | ( w7019 & w7028 ) | ( w7020 & w7028 ) ;
  assign w7081 = ( w6882 & w6894 ) | ( w6882 & w6907 ) | ( w6894 & w6907 ) ;
  assign w7082 = \pi41 & \pi49 ;
  assign w7083 = \pi40 & \pi50 ;
  assign w7084 = \pi39 & \pi51 ;
  assign w7085 = ( w7082 & w7083 ) | ( w7082 & w7084 ) | ( w7083 & w7084 ) ;
  assign w7086 = w7082 ^ w7084 ;
  assign w7087 = w7083 ^ w7086 ;
  assign w7088 = ( w6888 & w6901 ) | ( w6888 & w7026 ) | ( w6901 & w7026 ) ;
  assign w7089 = w7081 ^ w7088 ;
  assign w7090 = w7087 ^ w7089 ;
  assign w7091 = \pi29 & \pi61 ;
  assign w7092 = \pi28 & \pi62 ;
  assign w7093 = \pi27 & \pi63 ;
  assign w7094 = ( w7091 & w7092 ) | ( w7091 & w7093 ) | ( w7092 & w7093 ) ;
  assign w7095 = w7091 ^ w7093 ;
  assign w7096 = w7092 ^ w7095 ;
  assign w7097 = \pi30 & \pi60 ;
  assign w7098 = \pi32 & \pi58 ;
  assign w7099 = w7097 ^ w7098 ;
  assign w7100 = \pi31 & \pi59 ;
  assign w7101 = w7099 ^ w7100 ;
  assign w7102 = ~\pi28 & w4300 ;
  assign w7103 = ( w4300 & w6990 ) | ( w4300 & ~w7102 ) | ( w6990 & ~w7102 ) ;
  assign w7104 = ( \pi29 & w6990 ) | ( \pi29 & w7103 ) | ( w6990 & w7103 ) ;
  assign w7105 = w7096 ^ w7101 ;
  assign w7106 = w7104 ^ w7105 ;
  assign w7107 = w7080 ^ w7090 ;
  assign w7108 = w7106 ^ w7107 ;
  assign w7109 = w7059 ^ w7079 ;
  assign w7110 = w7055 ^ w7109 ;
  assign w7111 = w7108 ^ w7110 ;
  assign w7112 = w7054 ^ w7111 ;
  assign w7113 = w7053 ^ w7112 ;
  assign w7114 = w7039 | w7113 ;
  assign w7115 = w7039 & w7113 ;
  assign w7116 = w7114 & ~w7115 ;
  assign w7117 = w7038 ^ w7116 ;
  assign w7118 = ( w7038 & w7114 ) | ( w7038 & w7115 ) | ( w7114 & w7115 ) ;
  assign w7119 = w7115 | w7118 ;
  assign w7120 = ( w7053 & w7054 ) | ( w7053 & w7111 ) | ( w7054 & w7111 ) ;
  assign w7121 = \pi44 & \pi45 ;
  assign w7122 = ( \pi45 & w7043 ) | ( \pi45 & w7121 ) | ( w7043 & w7121 ) ;
  assign w7123 = ( w6962 & w6984 ) | ( w6962 & w7122 ) | ( w6984 & w7122 ) ;
  assign w7124 = \pi36 & \pi55 ;
  assign w7125 = \pi34 & \pi57 ;
  assign w7126 = ( w3615 & w7124 ) | ( w3615 & w7125 ) | ( w7124 & w7125 ) ;
  assign w7127 = w3615 ^ w7125 ;
  assign w7128 = w7124 ^ w7127 ;
  assign w7129 = ( w6968 & w6974 ) | ( w6968 & w7024 ) | ( w6974 & w7024 ) ;
  assign w7130 = w7123 ^ w7128 ;
  assign w7131 = w7129 ^ w7130 ;
  assign w7132 = ( w7046 & w7048 ) | ( w7046 & w7049 ) | ( w7048 & w7049 ) ;
  assign w7133 = \pi33 & \pi58 ;
  assign w7134 = \pi32 & \pi59 ;
  assign w7135 = \pi31 & \pi60 ;
  assign w7136 = ( w7133 & w7134 ) | ( w7133 & w7135 ) | ( w7134 & w7135 ) ;
  assign w7137 = w7133 ^ w7135 ;
  assign w7138 = w7134 ^ w7137 ;
  assign w7139 = \pi39 & \pi52 ;
  assign w7140 = \pi38 & \pi53 ;
  assign w7141 = \pi37 & \pi54 ;
  assign w7142 = ( w7139 & w7140 ) | ( w7139 & w7141 ) | ( w7140 & w7141 ) ;
  assign w7143 = w7139 ^ w7141 ;
  assign w7144 = w7140 ^ w7143 ;
  assign w7145 = w7085 ^ w7138 ;
  assign w7146 = w7144 ^ w7145 ;
  assign w7147 = w7132 ^ w7146 ;
  assign w7148 = ( w7097 & w7098 ) | ( w7097 & w7100 ) | ( w7098 & w7100 ) ;
  assign w7149 = w7069 ^ w7094 ;
  assign w7150 = w7148 ^ w7149 ;
  assign w7151 = ( w7081 & w7087 ) | ( w7081 & w7088 ) | ( w7087 & w7088 ) ;
  assign w7152 = \pi41 & \pi50 ;
  assign w7153 = \pi40 & \pi51 ;
  assign w7154 = \pi28 & \pi63 ;
  assign w7155 = ( w7152 & w7153 ) | ( w7152 & w7154 ) | ( w7153 & w7154 ) ;
  assign w7156 = w7152 ^ w7154 ;
  assign w7157 = w7153 ^ w7156 ;
  assign w7158 = \pi44 & \pi47 ;
  assign w7159 = \pi43 & \pi48 ;
  assign w7160 = \pi35 & \pi56 ;
  assign w7161 = ( w7158 & w7159 ) | ( w7158 & w7160 ) | ( w7159 & w7160 ) ;
  assign w7162 = w7158 ^ w7160 ;
  assign w7163 = w7159 ^ w7162 ;
  assign w7164 = \pi29 & \pi62 ;
  assign w7165 = \pi45 & ~w7164 ;
  assign w7166 = ( \pi46 & w7164 ) | ( \pi46 & w7165 ) | ( w7164 & w7165 ) ;
  assign w7167 = ~\pi45 & \pi46 ;
  assign w7168 = w7157 ^ w7167 ;
  assign w7169 = w7163 ^ w7168 ;
  assign w7170 = w7164 ^ w7169 ;
  assign w7171 = w7150 ^ w7151 ;
  assign w7172 = w7170 ^ w7171 ;
  assign w7173 = ( w7040 & w7041 ) | ( w7040 & w7051 ) | ( w7041 & w7051 ) ;
  assign w7174 = w7131 ^ w7172 ;
  assign w7175 = w7173 ^ w7174 ;
  assign w7176 = w7147 ^ w7175 ;
  assign w7177 = ( w7055 & w7108 ) | ( w7055 & w7109 ) | ( w7108 & w7109 ) ;
  assign w7178 = ( w7080 & w7090 ) | ( w7080 & w7106 ) | ( w7090 & w7106 ) ;
  assign w7179 = ( w7057 & w7058 ) | ( w7057 & w7079 ) | ( w7058 & w7079 ) ;
  assign w7180 = \pi28 | w6990 ;
  assign w7181 = ( \pi29 & w6990 ) | ( \pi29 & w7180 ) | ( w6990 & w7180 ) ;
  assign w7182 = ( w4300 & w6990 ) | ( w4300 & w7181 ) | ( w6990 & w7181 ) ;
  assign w7183 = ( w7096 & w7101 ) | ( w7096 & w7182 ) | ( w7101 & w7182 ) ;
  assign w7184 = ( w7065 & w7071 ) | ( w7065 & w7077 ) | ( w7071 & w7077 ) ;
  assign w7185 = w7183 ^ w7184 ;
  assign w7186 = w7063 ^ w7185 ;
  assign w7187 = w7075 ^ w7186 ;
  assign w7188 = \pi30 & \pi61 ;
  assign w7189 = w7187 ^ w7188 ;
  assign w7190 = w7178 ^ w7179 ;
  assign w7191 = w7189 ^ w7190 ;
  assign w7192 = w7176 ^ w7177 ;
  assign w7193 = w7191 ^ w7192 ;
  assign w7194 = w7119 ^ w7120 ;
  assign w7195 = w7193 ^ w7194 ;
  assign w7196 = ( w7119 & w7120 ) | ( w7119 & w7193 ) | ( w7120 & w7193 ) ;
  assign w7197 = ( w7178 & w7179 ) | ( w7178 & w7189 ) | ( w7179 & w7189 ) ;
  assign w7198 = ( w7131 & w7132 ) | ( w7131 & w7146 ) | ( w7132 & w7146 ) ;
  assign w7199 = w7063 ^ w7075 ;
  assign w7200 = w7188 ^ w7199 ;
  assign w7201 = ( w7183 & w7184 ) | ( w7183 & w7200 ) | ( w7184 & w7200 ) ;
  assign w7202 = \pi31 & \pi61 ;
  assign w7203 = ( \pi30 & \pi62 ) | ( \pi30 & ~w7166 ) | ( \pi62 & ~w7166 ) ;
  assign w7204 = w7202 ^ w7203 ;
  assign w7205 = w7166 & w7204 ;
  assign w7206 = \pi30 & \pi62 ;
  assign w7207 = w7166 ^ w7206 ;
  assign w7208 = w7202 ^ w7207 ;
  assign w7209 = \pi41 & \pi51 ;
  assign w7210 = \pi40 & \pi52 ;
  assign w7211 = \pi39 & \pi53 ;
  assign w7212 = ( w7209 & w7210 ) | ( w7209 & w7211 ) | ( w7210 & w7211 ) ;
  assign w7213 = w7209 ^ w7211 ;
  assign w7214 = w7210 ^ w7213 ;
  assign w7215 = ( w7063 & w7075 ) | ( w7063 & w7188 ) | ( w7075 & w7188 ) ;
  assign w7216 = w7208 ^ w7215 ;
  assign w7217 = w7214 ^ w7216 ;
  assign w7218 = \pi42 & \pi50 ;
  assign w7219 = \pi35 & \pi57 ;
  assign w7220 = \pi34 & \pi58 ;
  assign w7221 = ( w7218 & w7219 ) | ( w7218 & w7220 ) | ( w7219 & w7220 ) ;
  assign w7222 = w7218 ^ w7220 ;
  assign w7223 = w7219 ^ w7222 ;
  assign w7224 = \pi45 & \pi47 ;
  assign w7225 = \pi44 & \pi48 ;
  assign w7226 = \pi43 & \pi49 ;
  assign w7227 = ( w7224 & w7225 ) | ( w7224 & w7226 ) | ( w7225 & w7226 ) ;
  assign w7228 = w7224 ^ w7226 ;
  assign w7229 = w7225 ^ w7228 ;
  assign w7230 = \pi36 & \pi56 ;
  assign w7231 = \pi33 & \pi59 ;
  assign w7232 = ( w6153 & w7230 ) | ( w6153 & w7231 ) | ( w7230 & w7231 ) ;
  assign w7233 = w6153 ^ w7231 ;
  assign w7234 = w7230 ^ w7233 ;
  assign w7235 = w7223 ^ w7234 ;
  assign w7236 = w7229 ^ w7235 ;
  assign w7237 = w7201 ^ w7217 ;
  assign w7238 = w7236 ^ w7237 ;
  assign w7239 = w7197 ^ w7198 ;
  assign w7240 = w7238 ^ w7239 ;
  assign w7241 = w7131 ^ w7147 ;
  assign w7242 = ( w7172 & w7173 ) | ( w7172 & w7241 ) | ( w7173 & w7241 ) ;
  assign w7243 = ( w7085 & w7138 ) | ( w7085 & w7144 ) | ( w7138 & w7144 ) ;
  assign w7244 = ( w7069 & w7094 ) | ( w7069 & w7148 ) | ( w7094 & w7148 ) ;
  assign w7245 = w7164 ^ w7167 ;
  assign w7246 = ( w7157 & w7163 ) | ( w7157 & w7245 ) | ( w7163 & w7245 ) ;
  assign w7247 = w7243 ^ w7244 ;
  assign w7248 = w7246 ^ w7247 ;
  assign w7249 = ( w7150 & w7151 ) | ( w7150 & w7170 ) | ( w7151 & w7170 ) ;
  assign w7250 = ( w7123 & w7128 ) | ( w7123 & w7129 ) | ( w7128 & w7129 ) ;
  assign w7251 = w7136 ^ w7142 ;
  assign w7252 = w7155 ^ w7251 ;
  assign w7253 = \pi38 & \pi54 ;
  assign w7254 = \pi37 & \pi55 ;
  assign w7255 = \pi32 & \pi60 ;
  assign w7256 = ( w7253 & w7254 ) | ( w7253 & w7255 ) | ( w7254 & w7255 ) ;
  assign w7257 = w7253 ^ w7255 ;
  assign w7258 = w7254 ^ w7257 ;
  assign w7259 = w7126 ^ w7161 ;
  assign w7260 = w7258 ^ w7259 ;
  assign w7261 = w7250 ^ w7260 ;
  assign w7262 = w7252 ^ w7261 ;
  assign w7263 = w7249 ^ w7262 ;
  assign w7264 = w7248 ^ w7263 ;
  assign w7265 = w7240 ^ w7242 ;
  assign w7266 = w7264 ^ w7265 ;
  assign w7267 = ( w7176 & w7177 ) | ( w7176 & w7191 ) | ( w7177 & w7191 ) ;
  assign w7268 = w7266 | w7267 ;
  assign w7269 = w7266 & w7267 ;
  assign w7270 = w7268 & ~w7269 ;
  assign w7271 = w7196 ^ w7270 ;
  assign w7272 = ( w7196 & w7268 ) | ( w7196 & w7269 ) | ( w7268 & w7269 ) ;
  assign w7273 = w7269 | w7272 ;
  assign w7274 = ( w7240 & w7242 ) | ( w7240 & w7264 ) | ( w7242 & w7264 ) ;
  assign w7275 = ( w7197 & w7198 ) | ( w7197 & w7238 ) | ( w7198 & w7238 ) ;
  assign w7276 = ( w7126 & w7161 ) | ( w7126 & w7258 ) | ( w7161 & w7258 ) ;
  assign w7277 = ( w7136 & w7142 ) | ( w7136 & w7155 ) | ( w7142 & w7155 ) ;
  assign w7278 = ( w7223 & w7229 ) | ( w7223 & w7234 ) | ( w7229 & w7234 ) ;
  assign w7279 = w7276 ^ w7278 ;
  assign w7280 = w7277 ^ w7279 ;
  assign w7281 = ( w7250 & w7252 ) | ( w7250 & w7260 ) | ( w7252 & w7260 ) ;
  assign w7282 = ( w7208 & w7214 ) | ( w7208 & w7215 ) | ( w7214 & w7215 ) ;
  assign w7283 = w7212 ^ w7221 ;
  assign w7284 = w7227 ^ w7283 ;
  assign w7285 = w7232 ^ w7256 ;
  assign w7286 = w1335 | w7205 ;
  assign w7287 = ( w4390 & w7205 ) | ( w4390 & w7286 ) | ( w7205 & w7286 ) ;
  assign w7288 = w7285 ^ w7287 ;
  assign w7289 = w7282 ^ w7284 ;
  assign w7290 = w7288 ^ w7289 ;
  assign w7291 = w7280 ^ w7281 ;
  assign w7292 = w7290 ^ w7291 ;
  assign w7293 = ( w7248 & w7249 ) | ( w7248 & w7262 ) | ( w7249 & w7262 ) ;
  assign w7294 = ( w7201 & w7217 ) | ( w7201 & w7236 ) | ( w7217 & w7236 ) ;
  assign w7295 = ( w7243 & w7244 ) | ( w7243 & w7246 ) | ( w7244 & w7246 ) ;
  assign w7296 = \pi33 & \pi60 ;
  assign w7297 = \pi32 & \pi61 ;
  assign w7298 = \pi30 & \pi63 ;
  assign w7299 = ( w7296 & w7297 ) | ( w7296 & w7298 ) | ( w7297 & w7298 ) ;
  assign w7300 = w7296 ^ w7298 ;
  assign w7301 = w7297 ^ w7300 ;
  assign w7302 = \pi39 & \pi54 ;
  assign w7303 = \pi36 & \pi57 ;
  assign w7304 = \pi35 & \pi58 ;
  assign w7305 = ( w7302 & w7303 ) | ( w7302 & w7304 ) | ( w7303 & w7304 ) ;
  assign w7306 = w7302 ^ w7304 ;
  assign w7307 = w7303 ^ w7306 ;
  assign w7308 = \pi41 & \pi52 ;
  assign w7309 = \pi40 & \pi53 ;
  assign w7310 = ( w6852 & w7308 ) | ( w6852 & w7309 ) | ( w7308 & w7309 ) ;
  assign w7311 = w6852 ^ w7309 ;
  assign w7312 = w7308 ^ w7311 ;
  assign w7313 = w7301 ^ w7312 ;
  assign w7314 = w7307 ^ w7313 ;
  assign w7315 = \pi45 & \pi48 ;
  assign w7316 = \pi38 & \pi55 ;
  assign w7317 = \pi37 & \pi56 ;
  assign w7318 = ( w7315 & w7316 ) | ( w7315 & w7317 ) | ( w7316 & w7317 ) ;
  assign w7319 = w7315 ^ w7317 ;
  assign w7320 = w7316 ^ w7319 ;
  assign w7321 = \pi44 & \pi49 ;
  assign w7322 = \pi43 & \pi50 ;
  assign w7323 = \pi42 & \pi51 ;
  assign w7324 = ( w7321 & w7322 ) | ( w7321 & w7323 ) | ( w7322 & w7323 ) ;
  assign w7325 = w7321 ^ w7323 ;
  assign w7326 = w7322 ^ w7325 ;
  assign w7327 = ~\pi46 & \pi47 ;
  assign w7328 = w7320 ^ w7327 ;
  assign w7329 = w7326 ^ w7328 ;
  assign w7330 = \pi31 & \pi62 ;
  assign w7331 = w7329 ^ w7330 ;
  assign w7332 = w7295 ^ w7314 ;
  assign w7333 = w7331 ^ w7332 ;
  assign w7334 = w7293 ^ w7294 ;
  assign w7335 = w7333 ^ w7334 ;
  assign w7336 = w7275 ^ w7335 ;
  assign w7337 = w7292 ^ w7336 ;
  assign w7338 = w7273 ^ w7274 ;
  assign w7339 = w7337 ^ w7338 ;
  assign w7340 = ( w7293 & w7294 ) | ( w7293 & w7333 ) | ( w7294 & w7333 ) ;
  assign w7341 = ( w7295 & w7314 ) | ( w7295 & w7331 ) | ( w7314 & w7331 ) ;
  assign w7342 = w1335 & w4390 ;
  assign w7343 = w7205 | w7342 ;
  assign w7344 = ( w7232 & w7256 ) | ( w7232 & w7343 ) | ( w7256 & w7343 ) ;
  assign w7345 = ( w7212 & w7221 ) | ( w7212 & w7227 ) | ( w7221 & w7227 ) ;
  assign w7346 = ( w7301 & w7307 ) | ( w7301 & w7312 ) | ( w7307 & w7312 ) ;
  assign w7347 = w7344 ^ w7345 ;
  assign w7348 = w7346 ^ w7347 ;
  assign w7349 = ( w7282 & w7284 ) | ( w7282 & w7288 ) | ( w7284 & w7288 ) ;
  assign w7350 = w7341 ^ w7348 ;
  assign w7351 = w7349 ^ w7350 ;
  assign w7352 = \pi44 & \pi50 ;
  assign w7353 = \pi43 & \pi51 ;
  assign w7354 = \pi36 & \pi58 ;
  assign w7355 = ( w7352 & w7353 ) | ( w7352 & w7354 ) | ( w7353 & w7354 ) ;
  assign w7356 = w7352 ^ w7354 ;
  assign w7357 = w7353 ^ w7356 ;
  assign w7358 = \pi42 & \pi52 ;
  assign w7359 = \pi41 & \pi53 ;
  assign w7360 = \pi40 & \pi54 ;
  assign w7361 = ( w7358 & w7359 ) | ( w7358 & w7360 ) | ( w7359 & w7360 ) ;
  assign w7362 = w7358 ^ w7360 ;
  assign w7363 = w7359 ^ w7362 ;
  assign w7364 = \pi46 & \pi48 ;
  assign w7365 = \pi45 & \pi49 ;
  assign w7366 = ( w6569 & w7364 ) | ( w6569 & w7365 ) | ( w7364 & w7365 ) ;
  assign w7367 = w6569 ^ w7365 ;
  assign w7368 = w7364 ^ w7367 ;
  assign w7369 = w7357 ^ w7368 ;
  assign w7370 = w7363 ^ w7369 ;
  assign w7371 = ( w7276 & w7277 ) | ( w7276 & w7278 ) | ( w7277 & w7278 ) ;
  assign w7372 = w7370 ^ w7371 ;
  assign w7373 = \pi59 & \pi62 ;
  assign w7374 = \pi35 & \pi59 ;
  assign w7375 = \pi33 & \pi61 ;
  assign w7376 = \pi32 & \pi62 ;
  assign w7377 = ( w7374 & w7375 ) | ( w7374 & w7376 ) | ( w7375 & w7376 ) ;
  assign w7378 = w7374 ^ w7376 ;
  assign w7379 = w7375 ^ w7378 ;
  assign w7380 = \pi39 & \pi55 ;
  assign w7381 = \pi37 & \pi57 ;
  assign w7382 = \pi34 & \pi60 ;
  assign w7383 = ( w7380 & w7381 ) | ( w7380 & w7382 ) | ( w7381 & w7382 ) ;
  assign w7384 = w7380 ^ w7382 ;
  assign w7385 = w7381 ^ w7384 ;
  assign w7386 = w7324 ^ w7379 ;
  assign w7387 = w7385 ^ w7386 ;
  assign w7388 = ( w7280 & w7281 ) | ( w7280 & w7290 ) | ( w7281 & w7290 ) ;
  assign w7389 = \pi31 & \pi63 ;
  assign w7390 = w7318 ^ w7389 ;
  assign w7391 = ~\pi46 & \pi62 ;
  assign w7392 = \pi31 & w7391 ;
  assign w7393 = ( \pi46 & \pi47 ) | ( \pi46 & w7392 ) | ( \pi47 & w7392 ) ;
  assign w7394 = w7390 ^ w7393 ;
  assign w7395 = w7327 ^ w7330 ;
  assign w7396 = ( w7320 & w7326 ) | ( w7320 & w7395 ) | ( w7326 & w7395 ) ;
  assign w7397 = w7299 ^ w7310 ;
  assign w7398 = w7305 ^ w7397 ;
  assign w7399 = w7394 ^ w7398 ;
  assign w7400 = w7396 ^ w7399 ;
  assign w7401 = w7387 ^ w7400 ;
  assign w7402 = w7372 ^ w7401 ;
  assign w7403 = w7388 ^ w7402 ;
  assign w7404 = w7340 ^ w7403 ;
  assign w7405 = w7351 ^ w7404 ;
  assign w7406 = ( w7275 & w7292 ) | ( w7275 & w7335 ) | ( w7292 & w7335 ) ;
  assign w7407 = ( w7273 & w7274 ) | ( w7273 & w7337 ) | ( w7274 & w7337 ) ;
  assign w7408 = w7406 ^ w7407 ;
  assign w7409 = w7405 ^ w7408 ;
  assign w7410 = w7372 ^ w7387 ;
  assign w7411 = ( w7388 & w7400 ) | ( w7388 & w7410 ) | ( w7400 & w7410 ) ;
  assign w7412 = ( w7370 & w7371 ) | ( w7370 & w7387 ) | ( w7371 & w7387 ) ;
  assign w7413 = \pi36 & \pi59 ;
  assign w7414 = ( \pi35 & \pi60 ) | ( \pi35 & ~w7366 ) | ( \pi60 & ~w7366 ) ;
  assign w7415 = w7413 ^ w7414 ;
  assign w7416 = w7366 & w7415 ;
  assign w7417 = \pi35 & \pi60 ;
  assign w7418 = w7366 ^ w7417 ;
  assign w7419 = w7413 ^ w7418 ;
  assign w7420 = \pi46 & \pi47 ;
  assign w7421 = w7318 & w7420 ;
  assign w7422 = ( \pi47 & \pi62 ) | ( \pi47 & w7420 ) | ( \pi62 & w7420 ) ;
  assign w7423 = ( \pi63 & w7318 ) | ( \pi63 & w7422 ) | ( w7318 & w7422 ) ;
  assign w7424 = ( \pi31 & w7421 ) | ( \pi31 & w7423 ) | ( w7421 & w7423 ) ;
  assign w7425 = ( w7299 & w7305 ) | ( w7299 & w7310 ) | ( w7305 & w7310 ) ;
  assign w7426 = w7419 ^ w7425 ;
  assign w7427 = w7424 ^ w7426 ;
  assign w7428 = ( w7394 & w7396 ) | ( w7394 & w7398 ) | ( w7396 & w7398 ) ;
  assign w7429 = w7412 ^ w7427 ;
  assign w7430 = w7428 ^ w7429 ;
  assign w7431 = \pi46 & \pi49 ;
  assign w7432 = \pi45 & \pi50 ;
  assign w7433 = \pi39 & \pi56 ;
  assign w7434 = ( w7431 & w7432 ) | ( w7431 & w7433 ) | ( w7432 & w7433 ) ;
  assign w7435 = w7431 ^ w7433 ;
  assign w7436 = w7432 ^ w7435 ;
  assign w7437 = \pi44 & \pi51 ;
  assign w7438 = \pi43 & \pi52 ;
  assign w7439 = \pi42 & \pi53 ;
  assign w7440 = ( w7437 & w7438 ) | ( w7437 & w7439 ) | ( w7438 & w7439 ) ;
  assign w7441 = w7437 ^ w7439 ;
  assign w7442 = w7438 ^ w7441 ;
  assign w7443 = ~\pi47 & \pi48 ;
  assign w7444 = w7436 ^ w7443 ;
  assign w7445 = w7442 ^ w7444 ;
  assign w7446 = \pi33 & \pi62 ;
  assign w7447 = w7445 ^ w7446 ;
  assign w7448 = ( w7344 & w7345 ) | ( w7344 & w7346 ) | ( w7345 & w7346 ) ;
  assign w7449 = \pi41 & \pi54 ;
  assign w7450 = \pi34 & \pi61 ;
  assign w7451 = \pi32 & \pi63 ;
  assign w7452 = ( w7449 & w7450 ) | ( w7449 & w7451 ) | ( w7450 & w7451 ) ;
  assign w7453 = w7449 ^ w7451 ;
  assign w7454 = w7450 ^ w7453 ;
  assign w7455 = \pi40 & \pi55 ;
  assign w7456 = \pi38 & \pi57 ;
  assign w7457 = \pi37 & \pi58 ;
  assign w7458 = ( w7455 & w7456 ) | ( w7455 & w7457 ) | ( w7456 & w7457 ) ;
  assign w7459 = w7455 ^ w7457 ;
  assign w7460 = w7456 ^ w7459 ;
  assign w7461 = w7355 ^ w7454 ;
  assign w7462 = w7460 ^ w7461 ;
  assign w7463 = w7447 ^ w7448 ;
  assign w7464 = w7462 ^ w7463 ;
  assign w7465 = ( w7341 & w7348 ) | ( w7341 & w7349 ) | ( w7348 & w7349 ) ;
  assign w7466 = w7361 ^ w7377 ;
  assign w7467 = w7383 ^ w7466 ;
  assign w7468 = ( w7357 & w7363 ) | ( w7357 & w7368 ) | ( w7363 & w7368 ) ;
  assign w7469 = ( w7324 & w7379 ) | ( w7324 & w7385 ) | ( w7379 & w7385 ) ;
  assign w7470 = w7467 ^ w7468 ;
  assign w7471 = w7469 ^ w7470 ;
  assign w7472 = w7464 ^ w7465 ;
  assign w7473 = w7471 ^ w7472 ;
  assign w7474 = w7411 ^ w7430 ;
  assign w7475 = w7473 ^ w7474 ;
  assign w7476 = ( w7340 & w7351 ) | ( w7340 & w7403 ) | ( w7351 & w7403 ) ;
  assign w7477 = ( w7405 & w7406 ) | ( w7405 & w7407 ) | ( w7406 & w7407 ) ;
  assign w7478 = w7475 ^ w7477 ;
  assign w7479 = w7476 ^ w7478 ;
  assign w7480 = ( w7475 & w7476 ) | ( w7475 & w7477 ) | ( w7476 & w7477 ) ;
  assign w7481 = ( w7411 & w7430 ) | ( w7411 & w7473 ) | ( w7430 & w7473 ) ;
  assign w7482 = ( w7447 & w7448 ) | ( w7447 & w7462 ) | ( w7448 & w7462 ) ;
  assign w7483 = \pi40 & \pi56 ;
  assign w7484 = \pi37 & \pi59 ;
  assign w7485 = \pi36 & \pi60 ;
  assign w7486 = ( w7483 & w7484 ) | ( w7483 & w7485 ) | ( w7484 & w7485 ) ;
  assign w7487 = w7483 ^ w7485 ;
  assign w7488 = w7484 ^ w7487 ;
  assign w7489 = \pi39 & \pi57 ;
  assign w7490 = \pi38 & \pi58 ;
  assign w7491 = ( w3945 & w7489 ) | ( w3945 & w7490 ) | ( w7489 & w7490 ) ;
  assign w7492 = w3945 ^ w7490 ;
  assign w7493 = w7489 ^ w7492 ;
  assign w7494 = \pi47 & \pi49 ;
  assign w7495 = \pi46 & \pi50 ;
  assign w7496 = \pi45 & \pi51 ;
  assign w7497 = ( w7494 & w7495 ) | ( w7494 & w7496 ) | ( w7495 & w7496 ) ;
  assign w7498 = w7494 ^ w7496 ;
  assign w7499 = w7495 ^ w7498 ;
  assign w7500 = w7488 ^ w7493 ;
  assign w7501 = w7499 ^ w7500 ;
  assign w7502 = ( w7467 & w7468 ) | ( w7467 & w7469 ) | ( w7468 & w7469 ) ;
  assign w7503 = w7482 ^ w7502 ;
  assign w7504 = w7501 ^ w7503 ;
  assign w7505 = ( w7464 & w7465 ) | ( w7464 & w7471 ) | ( w7465 & w7471 ) ;
  assign w7506 = ( w7412 & w7427 ) | ( w7412 & w7428 ) | ( w7427 & w7428 ) ;
  assign w7507 = w7434 ^ w7440 ;
  assign w7508 = ( \pi33 & \pi47 ) | ( \pi33 & \pi62 ) | ( \pi47 & \pi62 ) ;
  assign w7509 = ~\pi47 & w7508 ;
  assign w7510 = ( \pi47 & \pi48 ) | ( \pi47 & w7509 ) | ( \pi48 & w7509 ) ;
  assign w7511 = w7507 ^ w7510 ;
  assign w7512 = ( w7355 & w7454 ) | ( w7355 & w7460 ) | ( w7454 & w7460 ) ;
  assign w7513 = w7443 ^ w7446 ;
  assign w7514 = ( w7436 & w7442 ) | ( w7436 & w7513 ) | ( w7442 & w7513 ) ;
  assign w7515 = w7511 ^ w7512 ;
  assign w7516 = w7514 ^ w7515 ;
  assign w7517 = \pi35 & \pi61 ;
  assign w7518 = \pi34 & \pi62 ;
  assign w7519 = \pi33 & \pi63 ;
  assign w7520 = ( w7517 & w7518 ) | ( w7517 & w7519 ) | ( w7518 & w7519 ) ;
  assign w7521 = w7517 ^ w7519 ;
  assign w7522 = w7518 ^ w7521 ;
  assign w7523 = \pi43 & \pi53 ;
  assign w7524 = \pi42 & \pi54 ;
  assign w7525 = \pi41 & \pi55 ;
  assign w7526 = ( w7523 & w7524 ) | ( w7523 & w7525 ) | ( w7524 & w7525 ) ;
  assign w7527 = w7523 ^ w7525 ;
  assign w7528 = w7524 ^ w7527 ;
  assign w7529 = ( w7361 & w7377 ) | ( w7361 & w7383 ) | ( w7377 & w7383 ) ;
  assign w7530 = w7522 ^ w7529 ;
  assign w7531 = w7528 ^ w7530 ;
  assign w7532 = w7452 ^ w7458 ;
  assign w7533 = w4299 | w7416 ;
  assign w7534 = ( w1779 & w7416 ) | ( w1779 & w7533 ) | ( w7416 & w7533 ) ;
  assign w7535 = w7532 ^ w7534 ;
  assign w7536 = ( w7419 & w7424 ) | ( w7419 & w7425 ) | ( w7424 & w7425 ) ;
  assign w7537 = w7535 ^ w7536 ;
  assign w7538 = w7531 ^ w7537 ;
  assign w7539 = w7506 ^ w7538 ;
  assign w7540 = w7516 ^ w7539 ;
  assign w7541 = w7504 ^ w7540 ;
  assign w7542 = w7505 ^ w7541 ;
  assign w7543 = w7481 | w7542 ;
  assign w7544 = w7481 & w7542 ;
  assign w7545 = w7543 & ~w7544 ;
  assign w7546 = w7480 ^ w7545 ;
  assign w7547 = ( w7480 & w7543 ) | ( w7480 & w7544 ) | ( w7543 & w7544 ) ;
  assign w7548 = w7544 | w7547 ;
  assign w7549 = ( w7504 & w7505 ) | ( w7504 & w7540 ) | ( w7505 & w7540 ) ;
  assign w7550 = ( w7482 & w7501 ) | ( w7482 & w7502 ) | ( w7501 & w7502 ) ;
  assign w7551 = ( w7488 & w7493 ) | ( w7488 & w7499 ) | ( w7493 & w7499 ) ;
  assign w7552 = w1779 & w4299 ;
  assign w7553 = w7416 | w7552 ;
  assign w7554 = ( w7452 & w7458 ) | ( w7452 & w7553 ) | ( w7458 & w7553 ) ;
  assign w7555 = w7551 ^ w7554 ;
  assign w7556 = w7491 ^ w7555 ;
  assign w7557 = w7497 ^ w7556 ;
  assign w7558 = \pi36 & \pi61 ;
  assign w7559 = w7557 ^ w7558 ;
  assign w7560 = \pi35 & \pi62 ;
  assign w7561 = \pi48 & ~w7560 ;
  assign w7562 = ( \pi49 & w7560 ) | ( \pi49 & w7561 ) | ( w7560 & w7561 ) ;
  assign w7563 = \pi47 & \pi50 ;
  assign w7564 = \pi46 & \pi51 ;
  assign w7565 = \pi40 & \pi57 ;
  assign w7566 = ( w7563 & w7564 ) | ( w7563 & w7565 ) | ( w7564 & w7565 ) ;
  assign w7567 = w7563 ^ w7565 ;
  assign w7568 = w7564 ^ w7567 ;
  assign w7569 = \pi47 & \pi48 ;
  assign w7570 = ( \pi48 & w7508 ) | ( \pi48 & w7569 ) | ( w7508 & w7569 ) ;
  assign w7571 = ( w7434 & w7440 ) | ( w7434 & w7570 ) | ( w7440 & w7570 ) ;
  assign w7572 = ~\pi48 & \pi49 ;
  assign w7573 = w7571 ^ w7572 ;
  assign w7574 = w7568 ^ w7573 ;
  assign w7575 = w7560 ^ w7574 ;
  assign w7576 = w7486 ^ w7520 ;
  assign w7577 = w7526 ^ w7576 ;
  assign w7578 = ( w7522 & w7528 ) | ( w7522 & w7529 ) | ( w7528 & w7529 ) ;
  assign w7579 = w7575 ^ w7578 ;
  assign w7580 = w7577 ^ w7579 ;
  assign w7581 = w7550 ^ w7559 ;
  assign w7582 = w7580 ^ w7581 ;
  assign w7583 = ( w7531 & w7535 ) | ( w7531 & w7536 ) | ( w7535 & w7536 ) ;
  assign w7584 = \pi34 & \pi63 ;
  assign w7585 = \pi42 & \pi55 ;
  assign w7586 = \pi41 & \pi56 ;
  assign w7587 = ( w7584 & w7585 ) | ( w7584 & w7586 ) | ( w7585 & w7586 ) ;
  assign w7588 = w7584 ^ w7586 ;
  assign w7589 = w7585 ^ w7588 ;
  assign w7590 = \pi39 & \pi58 ;
  assign w7591 = \pi38 & \pi59 ;
  assign w7592 = \pi37 & \pi60 ;
  assign w7593 = ( w7590 & w7591 ) | ( w7590 & w7592 ) | ( w7591 & w7592 ) ;
  assign w7594 = w7590 ^ w7592 ;
  assign w7595 = w7591 ^ w7594 ;
  assign w7596 = \pi45 & \pi52 ;
  assign w7597 = \pi44 & \pi53 ;
  assign w7598 = \pi43 & \pi54 ;
  assign w7599 = ( w7596 & w7597 ) | ( w7596 & w7598 ) | ( w7597 & w7598 ) ;
  assign w7600 = w7596 ^ w7598 ;
  assign w7601 = w7597 ^ w7600 ;
  assign w7602 = w7589 ^ w7595 ;
  assign w7603 = w7601 ^ w7602 ;
  assign w7604 = ( w7511 & w7512 ) | ( w7511 & w7514 ) | ( w7512 & w7514 ) ;
  assign w7605 = w7583 ^ w7603 ;
  assign w7606 = w7604 ^ w7605 ;
  assign w7607 = ( w7506 & w7516 ) | ( w7506 & w7538 ) | ( w7516 & w7538 ) ;
  assign w7608 = w7582 ^ w7607 ;
  assign w7609 = w7606 ^ w7608 ;
  assign w7610 = w7548 ^ w7549 ;
  assign w7611 = w7609 ^ w7610 ;
  assign w7612 = ( w7582 & w7606 ) | ( w7582 & w7607 ) | ( w7606 & w7607 ) ;
  assign w7613 = ( w7583 & w7603 ) | ( w7583 & w7604 ) | ( w7603 & w7604 ) ;
  assign w7614 = ( w7486 & w7520 ) | ( w7486 & w7526 ) | ( w7520 & w7526 ) ;
  assign w7615 = ( w7589 & w7595 ) | ( w7589 & w7601 ) | ( w7595 & w7601 ) ;
  assign w7616 = ( w7491 & w7497 ) | ( w7491 & w7558 ) | ( w7497 & w7558 ) ;
  assign w7617 = w7615 ^ w7616 ;
  assign w7618 = w7614 ^ w7617 ;
  assign w7619 = w7587 ^ w7593 ;
  assign w7620 = w7599 ^ w7619 ;
  assign w7621 = w7560 ^ w7572 ;
  assign w7622 = ( w7568 & w7571 ) | ( w7568 & w7621 ) | ( w7571 & w7621 ) ;
  assign w7623 = \pi45 & \pi53 ;
  assign w7624 = \pi40 & \pi58 ;
  assign w7625 = \pi39 & \pi59 ;
  assign w7626 = ( w7623 & w7624 ) | ( w7623 & w7625 ) | ( w7624 & w7625 ) ;
  assign w7627 = w7623 ^ w7625 ;
  assign w7628 = w7624 ^ w7627 ;
  assign w7629 = \pi48 & \pi50 ;
  assign w7630 = \pi47 & \pi51 ;
  assign w7631 = \pi46 & \pi52 ;
  assign w7632 = ( w7629 & w7630 ) | ( w7629 & w7631 ) | ( w7630 & w7631 ) ;
  assign w7633 = w7629 ^ w7631 ;
  assign w7634 = w7630 ^ w7633 ;
  assign w7635 = \pi37 & \pi61 ;
  assign w7636 = \pi36 & \pi62 ;
  assign w7637 = w7562 ^ w7636 ;
  assign w7638 = w7635 ^ w7637 ;
  assign w7639 = w7628 ^ w7638 ;
  assign w7640 = w7634 ^ w7639 ;
  assign w7641 = w7620 ^ w7622 ;
  assign w7642 = w7640 ^ w7641 ;
  assign w7643 = ( w7613 & w7618 ) | ( w7613 & w7642 ) | ( w7618 & w7642 ) ;
  assign w7644 = w7613 ^ w7618 ;
  assign w7645 = w7642 ^ w7644 ;
  assign w7646 = ( w7550 & w7559 ) | ( w7550 & w7580 ) | ( w7559 & w7580 ) ;
  assign w7647 = ( w7575 & w7577 ) | ( w7575 & w7578 ) | ( w7577 & w7578 ) ;
  assign w7648 = \pi35 & \pi63 ;
  assign w7649 = \pi44 & \pi54 ;
  assign w7650 = w7648 ^ w7649 ;
  assign w7651 = \pi43 & \pi55 ;
  assign w7652 = w7650 ^ w7651 ;
  assign w7653 = \pi42 & \pi56 ;
  assign w7654 = \pi41 & \pi57 ;
  assign w7655 = \pi38 & \pi60 ;
  assign w7656 = ( w7653 & w7654 ) | ( w7653 & w7655 ) | ( w7654 & w7655 ) ;
  assign w7657 = w7653 ^ w7655 ;
  assign w7658 = w7654 ^ w7657 ;
  assign w7659 = w7566 ^ w7652 ;
  assign w7660 = w7658 ^ w7659 ;
  assign w7661 = w7491 ^ w7497 ;
  assign w7662 = w7558 ^ w7661 ;
  assign w7663 = ( w7551 & w7554 ) | ( w7551 & w7662 ) | ( w7554 & w7662 ) ;
  assign w7664 = w7647 ^ w7663 ;
  assign w7665 = w7660 ^ w7664 ;
  assign w7666 = w7645 ^ w7646 ;
  assign w7667 = w7665 ^ w7666 ;
  assign w7668 = ( w7548 & w7549 ) | ( w7548 & w7609 ) | ( w7549 & w7609 ) ;
  assign w7669 = w7612 ^ w7668 ;
  assign w7670 = w7667 ^ w7669 ;
  assign w7671 = ( w7645 & w7646 ) | ( w7645 & w7665 ) | ( w7646 & w7665 ) ;
  assign w7672 = ( w7647 & w7660 ) | ( w7647 & w7663 ) | ( w7660 & w7663 ) ;
  assign w7673 = ( w7587 & w7593 ) | ( w7587 & w7599 ) | ( w7593 & w7599 ) ;
  assign w7674 = ( w7566 & w7652 ) | ( w7566 & w7658 ) | ( w7652 & w7658 ) ;
  assign w7675 = ~\pi49 & \pi50 ;
  assign w7676 = w7673 ^ w7675 ;
  assign w7677 = w7674 ^ w7676 ;
  assign w7678 = \pi37 & \pi62 ;
  assign w7679 = w7677 ^ w7678 ;
  assign w7680 = ( w7562 & w7635 ) | ( w7562 & w7636 ) | ( w7635 & w7636 ) ;
  assign w7681 = \pi39 & \pi60 ;
  assign w7682 = \pi38 & \pi61 ;
  assign w7683 = \pi36 & \pi63 ;
  assign w7684 = ( w7681 & w7682 ) | ( w7681 & w7683 ) | ( w7682 & w7683 ) ;
  assign w7685 = w7681 ^ w7683 ;
  assign w7686 = w7682 ^ w7685 ;
  assign w7687 = w7656 ^ w7680 ;
  assign w7688 = w7686 ^ w7687 ;
  assign w7689 = ( w7648 & w7649 ) | ( w7648 & w7651 ) | ( w7649 & w7651 ) ;
  assign w7690 = w7626 ^ w7632 ;
  assign w7691 = w7689 ^ w7690 ;
  assign w7692 = ( w7628 & w7634 ) | ( w7628 & w7638 ) | ( w7634 & w7638 ) ;
  assign w7693 = w7688 ^ w7692 ;
  assign w7694 = w7691 ^ w7693 ;
  assign w7695 = w7672 ^ w7679 ;
  assign w7696 = w7694 ^ w7695 ;
  assign w7697 = \pi44 & \pi55 ;
  assign w7698 = \pi41 & \pi58 ;
  assign w7699 = \pi40 & \pi59 ;
  assign w7700 = ( w7697 & w7698 ) | ( w7697 & w7699 ) | ( w7698 & w7699 ) ;
  assign w7701 = w7697 ^ w7699 ;
  assign w7702 = w7698 ^ w7701 ;
  assign w7703 = \pi47 & \pi52 ;
  assign w7704 = \pi46 & \pi53 ;
  assign w7705 = \pi45 & \pi54 ;
  assign w7706 = ( w7703 & w7704 ) | ( w7703 & w7705 ) | ( w7704 & w7705 ) ;
  assign w7707 = w7703 ^ w7705 ;
  assign w7708 = w7704 ^ w7707 ;
  assign w7709 = \pi48 & \pi51 ;
  assign w7710 = \pi43 & \pi56 ;
  assign w7711 = \pi42 & \pi57 ;
  assign w7712 = ( w7709 & w7710 ) | ( w7709 & w7711 ) | ( w7710 & w7711 ) ;
  assign w7713 = w7709 ^ w7711 ;
  assign w7714 = w7710 ^ w7713 ;
  assign w7715 = w7702 ^ w7714 ;
  assign w7716 = w7708 ^ w7715 ;
  assign w7717 = ( w7614 & w7615 ) | ( w7614 & w7616 ) | ( w7615 & w7616 ) ;
  assign w7718 = ( w7620 & w7622 ) | ( w7620 & w7640 ) | ( w7622 & w7640 ) ;
  assign w7719 = w7717 ^ w7718 ;
  assign w7720 = w7716 ^ w7719 ;
  assign w7721 = w7643 ^ w7696 ;
  assign w7722 = w7720 ^ w7721 ;
  assign w7723 = ( w7612 & w7667 ) | ( w7612 & w7668 ) | ( w7667 & w7668 ) ;
  assign w7724 = w7671 ^ w7723 ;
  assign w7725 = w7722 ^ w7724 ;
  assign w7726 = ( w7671 & w7722 ) | ( w7671 & w7723 ) | ( w7722 & w7723 ) ;
  assign w7727 = ( w7643 & w7696 ) | ( w7643 & w7720 ) | ( w7696 & w7720 ) ;
  assign w7728 = ( w7626 & w7632 ) | ( w7626 & w7689 ) | ( w7632 & w7689 ) ;
  assign w7729 = \pi49 & \pi51 ;
  assign w7730 = \pi48 & \pi52 ;
  assign w7731 = \pi47 & \pi53 ;
  assign w7732 = ( w7729 & w7730 ) | ( w7729 & w7731 ) | ( w7730 & w7731 ) ;
  assign w7733 = w7729 ^ w7731 ;
  assign w7734 = w7730 ^ w7733 ;
  assign w7735 = ( w7656 & w7680 ) | ( w7656 & w7686 ) | ( w7680 & w7686 ) ;
  assign w7736 = w7728 ^ w7735 ;
  assign w7737 = w7734 ^ w7736 ;
  assign w7738 = ( w7716 & w7717 ) | ( w7716 & w7718 ) | ( w7717 & w7718 ) ;
  assign w7739 = w7684 ^ w7700 ;
  assign w7740 = w7706 ^ w7739 ;
  assign w7741 = ( w7702 & w7708 ) | ( w7702 & w7714 ) | ( w7708 & w7714 ) ;
  assign w7742 = \pi37 & \pi63 ;
  assign w7743 = w7712 ^ w7742 ;
  assign w7744 = ~\pi49 & \pi62 ;
  assign w7745 = \pi37 & w7744 ;
  assign w7746 = ( \pi49 & \pi50 ) | ( \pi49 & w7745 ) | ( \pi50 & w7745 ) ;
  assign w7747 = w7743 ^ w7746 ;
  assign w7748 = w7741 ^ w7747 ;
  assign w7749 = w7740 ^ w7748 ;
  assign w7750 = w7737 ^ w7738 ;
  assign w7751 = w7749 ^ w7750 ;
  assign w7752 = ( w7672 & w7679 ) | ( w7672 & w7694 ) | ( w7679 & w7694 ) ;
  assign w7753 = \pi40 & \pi60 ;
  assign w7754 = \pi39 & \pi61 ;
  assign w7755 = \pi38 & \pi62 ;
  assign w7756 = ( w7753 & w7754 ) | ( w7753 & w7755 ) | ( w7754 & w7755 ) ;
  assign w7757 = w7753 ^ w7755 ;
  assign w7758 = w7754 ^ w7757 ;
  assign w7759 = \pi45 & \pi55 ;
  assign w7760 = \pi44 & \pi56 ;
  assign w7761 = \pi43 & \pi57 ;
  assign w7762 = ( w7759 & w7760 ) | ( w7759 & w7761 ) | ( w7760 & w7761 ) ;
  assign w7763 = w7759 ^ w7761 ;
  assign w7764 = w7760 ^ w7763 ;
  assign w7765 = \pi42 & \pi58 ;
  assign w7766 = \pi41 & \pi59 ;
  assign w7767 = ( w4259 & w7765 ) | ( w4259 & w7766 ) | ( w7765 & w7766 ) ;
  assign w7768 = w4259 ^ w7766 ;
  assign w7769 = w7765 ^ w7768 ;
  assign w7770 = w7758 ^ w7769 ;
  assign w7771 = w7764 ^ w7770 ;
  assign w7772 = w7675 ^ w7678 ;
  assign w7773 = ( w7673 & w7674 ) | ( w7673 & w7772 ) | ( w7674 & w7772 ) ;
  assign w7774 = ( w7688 & w7691 ) | ( w7688 & w7692 ) | ( w7691 & w7692 ) ;
  assign w7775 = w7773 ^ w7774 ;
  assign w7776 = w7771 ^ w7775 ;
  assign w7777 = w7751 ^ w7752 ;
  assign w7778 = w7776 ^ w7777 ;
  assign w7779 = w7727 & w7778 ;
  assign w7780 = w7727 | w7778 ;
  assign w7781 = ~w7779 & w7780 ;
  assign w7782 = w7726 ^ w7781 ;
  assign w7783 = ( w7726 & w7779 ) | ( w7726 & w7780 ) | ( w7779 & w7780 ) ;
  assign w7784 = w7779 | w7783 ;
  assign w7785 = ( w7751 & w7752 ) | ( w7751 & w7776 ) | ( w7752 & w7776 ) ;
  assign w7786 = ( w7737 & w7738 ) | ( w7737 & w7749 ) | ( w7738 & w7749 ) ;
  assign w7787 = \pi47 & \pi54 ;
  assign w7788 = \pi46 & \pi55 ;
  assign w7789 = \pi38 & \pi63 ;
  assign w7790 = ( w7787 & w7788 ) | ( w7787 & w7789 ) | ( w7788 & w7789 ) ;
  assign w7791 = w7787 ^ w7789 ;
  assign w7792 = w7788 ^ w7791 ;
  assign w7793 = \pi45 & \pi56 ;
  assign w7794 = \pi43 & \pi58 ;
  assign w7795 = \pi42 & \pi59 ;
  assign w7796 = ( w7793 & w7794 ) | ( w7793 & w7795 ) | ( w7794 & w7795 ) ;
  assign w7797 = w7793 ^ w7795 ;
  assign w7798 = w7794 ^ w7797 ;
  assign w7799 = \pi49 & \pi52 ;
  assign w7800 = \pi48 & \pi53 ;
  assign w7801 = \pi44 & \pi57 ;
  assign w7802 = ( w7799 & w7800 ) | ( w7799 & w7801 ) | ( w7800 & w7801 ) ;
  assign w7803 = w7799 ^ w7801 ;
  assign w7804 = w7800 ^ w7803 ;
  assign w7805 = w7792 ^ w7798 ;
  assign w7806 = w7804 ^ w7805 ;
  assign w7807 = ( w7728 & w7734 ) | ( w7728 & w7735 ) | ( w7734 & w7735 ) ;
  assign w7808 = w7806 ^ w7807 ;
  assign w7809 = \pi49 & \pi50 ;
  assign w7810 = w7712 & w7809 ;
  assign w7811 = ( \pi50 & \pi62 ) | ( \pi50 & w7809 ) | ( \pi62 & w7809 ) ;
  assign w7812 = ( \pi63 & w7712 ) | ( \pi63 & w7811 ) | ( w7712 & w7811 ) ;
  assign w7813 = ( \pi37 & w7810 ) | ( \pi37 & w7812 ) | ( w7810 & w7812 ) ;
  assign w7814 = \pi41 & \pi60 ;
  assign w7815 = ( \pi40 & \pi61 ) | ( \pi40 & ~w7732 ) | ( \pi61 & ~w7732 ) ;
  assign w7816 = w7814 ^ w7815 ;
  assign w7817 = w7732 & w7816 ;
  assign w7818 = \pi40 & \pi61 ;
  assign w7819 = w7732 ^ w7818 ;
  assign w7820 = w7814 ^ w7819 ;
  assign w7821 = ~\pi50 & \pi51 ;
  assign w7822 = w7813 ^ w7821 ;
  assign w7823 = w7820 ^ w7822 ;
  assign w7824 = \pi39 & \pi62 ;
  assign w7825 = w7823 ^ w7824 ;
  assign w7826 = ( w7771 & w7773 ) | ( w7771 & w7774 ) | ( w7773 & w7774 ) ;
  assign w7827 = ( w7740 & w7741 ) | ( w7740 & w7747 ) | ( w7741 & w7747 ) ;
  assign w7828 = w7756 ^ w7767 ;
  assign w7829 = w7762 ^ w7828 ;
  assign w7830 = ( w7758 & w7764 ) | ( w7758 & w7769 ) | ( w7764 & w7769 ) ;
  assign w7831 = ( w7684 & w7700 ) | ( w7684 & w7706 ) | ( w7700 & w7706 ) ;
  assign w7832 = w7829 ^ w7830 ;
  assign w7833 = w7831 ^ w7832 ;
  assign w7834 = w7826 ^ w7827 ;
  assign w7835 = w7833 ^ w7834 ;
  assign w7836 = w7808 ^ w7825 ;
  assign w7837 = w7786 ^ w7836 ;
  assign w7838 = w7835 ^ w7837 ;
  assign w7839 = w7784 ^ w7785 ;
  assign w7840 = w7838 ^ w7839 ;
  assign w7841 = ( w7784 & w7785 ) | ( w7784 & w7838 ) | ( w7785 & w7838 ) ;
  assign w7842 = ( w7786 & w7835 ) | ( w7786 & w7836 ) | ( w7835 & w7836 ) ;
  assign w7843 = ( w7826 & w7827 ) | ( w7826 & w7833 ) | ( w7827 & w7833 ) ;
  assign w7844 = \pi42 & \pi60 ;
  assign w7845 = \pi41 & \pi61 ;
  assign w7846 = \pi39 & \pi63 ;
  assign w7847 = ( w7844 & w7845 ) | ( w7844 & w7846 ) | ( w7845 & w7846 ) ;
  assign w7848 = w7844 ^ w7846 ;
  assign w7849 = w7845 ^ w7848 ;
  assign w7850 = ~\pi40 & w4300 ;
  assign w7851 = ( w4300 & w7817 ) | ( w4300 & ~w7850 ) | ( w7817 & ~w7850 ) ;
  assign w7852 = ( \pi41 & w7817 ) | ( \pi41 & w7851 ) | ( w7817 & w7851 ) ;
  assign w7853 = w7796 ^ w7849 ;
  assign w7854 = w7852 ^ w7853 ;
  assign w7855 = w7821 ^ w7824 ;
  assign w7856 = ( w7813 & w7820 ) | ( w7813 & w7855 ) | ( w7820 & w7855 ) ;
  assign w7857 = w7854 ^ w7856 ;
  assign w7858 = \pi44 & \pi58 ;
  assign w7859 = \pi43 & \pi59 ;
  assign w7860 = ( w6100 & w7858 ) | ( w6100 & w7859 ) | ( w7858 & w7859 ) ;
  assign w7861 = w6100 ^ w7859 ;
  assign w7862 = w7858 ^ w7861 ;
  assign w7863 = \pi47 & \pi55 ;
  assign w7864 = \pi46 & \pi56 ;
  assign w7865 = \pi45 & \pi57 ;
  assign w7866 = ( w7863 & w7864 ) | ( w7863 & w7865 ) | ( w7864 & w7865 ) ;
  assign w7867 = w7863 ^ w7865 ;
  assign w7868 = w7864 ^ w7867 ;
  assign w7869 = \pi50 & \pi52 ;
  assign w7870 = \pi49 & \pi53 ;
  assign w7871 = \pi48 & \pi54 ;
  assign w7872 = ( w7869 & w7870 ) | ( w7869 & w7871 ) | ( w7870 & w7871 ) ;
  assign w7873 = w7869 ^ w7871 ;
  assign w7874 = w7870 ^ w7873 ;
  assign w7875 = w7862 ^ w7868 ;
  assign w7876 = w7874 ^ w7875 ;
  assign w7877 = w7790 ^ w7802 ;
  assign w7878 = ( \pi39 & \pi50 ) | ( \pi39 & \pi62 ) | ( \pi50 & \pi62 ) ;
  assign w7879 = ~\pi50 & w7878 ;
  assign w7880 = ( \pi50 & \pi51 ) | ( \pi50 & w7879 ) | ( \pi51 & w7879 ) ;
  assign w7881 = w7877 ^ w7880 ;
  assign w7882 = ( w7756 & w7762 ) | ( w7756 & w7767 ) | ( w7762 & w7767 ) ;
  assign w7883 = ( w7792 & w7798 ) | ( w7792 & w7804 ) | ( w7798 & w7804 ) ;
  assign w7884 = w7881 ^ w7882 ;
  assign w7885 = w7883 ^ w7884 ;
  assign w7886 = ( w7806 & w7807 ) | ( w7806 & w7825 ) | ( w7807 & w7825 ) ;
  assign w7887 = ( w7829 & w7830 ) | ( w7829 & w7831 ) | ( w7830 & w7831 ) ;
  assign w7888 = w7886 ^ w7887 ;
  assign w7889 = w7857 ^ w7888 ;
  assign w7890 = w7843 ^ w7885 ;
  assign w7891 = w7876 ^ w7890 ;
  assign w7892 = w7889 ^ w7891 ;
  assign w7893 = w7842 | w7892 ;
  assign w7894 = w7842 & w7892 ;
  assign w7895 = w7893 & ~w7894 ;
  assign w7896 = w7841 ^ w7895 ;
  assign w7897 = ( w7841 & w7893 ) | ( w7841 & w7894 ) | ( w7893 & w7894 ) ;
  assign w7898 = w7894 | w7897 ;
  assign w7899 = ( w7885 & w7886 ) | ( w7885 & w7887 ) | ( w7886 & w7887 ) ;
  assign w7900 = \pi47 & \pi56 ;
  assign w7901 = \pi46 & \pi57 ;
  assign w7902 = \pi43 & \pi60 ;
  assign w7903 = ( w7900 & w7901 ) | ( w7900 & w7902 ) | ( w7901 & w7902 ) ;
  assign w7904 = w7900 ^ w7902 ;
  assign w7905 = w7901 ^ w7904 ;
  assign w7906 = \pi50 & \pi53 ;
  assign w7907 = \pi49 & \pi54 ;
  assign w7908 = \pi48 & \pi55 ;
  assign w7909 = ( w7906 & w7907 ) | ( w7906 & w7908 ) | ( w7907 & w7908 ) ;
  assign w7910 = w7906 ^ w7908 ;
  assign w7911 = w7907 ^ w7910 ;
  assign w7912 = ~\pi51 & \pi52 ;
  assign w7913 = w7905 ^ w7912 ;
  assign w7914 = w7911 ^ w7913 ;
  assign w7915 = \pi41 & \pi62 ;
  assign w7916 = w7914 ^ w7915 ;
  assign w7917 = \pi45 & \pi58 ;
  assign w7918 = \pi44 & \pi59 ;
  assign w7919 = \pi42 & \pi61 ;
  assign w7920 = ( w7917 & w7918 ) | ( w7917 & w7919 ) | ( w7918 & w7919 ) ;
  assign w7921 = w7917 ^ w7919 ;
  assign w7922 = w7918 ^ w7921 ;
  assign w7923 = w7847 ^ w7860 ;
  assign w7924 = w7922 ^ w7923 ;
  assign w7925 = w7916 ^ w7924 ;
  assign w7926 = w7866 ^ w7925 ;
  assign w7927 = w7872 ^ w7926 ;
  assign w7928 = \pi40 & \pi63 ;
  assign w7929 = w7927 ^ w7928 ;
  assign w7930 = \pi40 | w7817 ;
  assign w7931 = ( \pi41 & w7817 ) | ( \pi41 & w7930 ) | ( w7817 & w7930 ) ;
  assign w7932 = ( w4300 & w7817 ) | ( w4300 & w7931 ) | ( w7817 & w7931 ) ;
  assign w7933 = ( w7796 & w7849 ) | ( w7796 & w7932 ) | ( w7849 & w7932 ) ;
  assign w7934 = \pi50 & \pi51 ;
  assign w7935 = ( \pi51 & w7878 ) | ( \pi51 & w7934 ) | ( w7878 & w7934 ) ;
  assign w7936 = ( w7790 & w7802 ) | ( w7790 & w7935 ) | ( w7802 & w7935 ) ;
  assign w7937 = ( w7862 & w7868 ) | ( w7862 & w7874 ) | ( w7868 & w7874 ) ;
  assign w7938 = w7933 ^ w7937 ;
  assign w7939 = w7936 ^ w7938 ;
  assign w7940 = ( w7854 & w7856 ) | ( w7854 & w7876 ) | ( w7856 & w7876 ) ;
  assign w7941 = ( w7881 & w7882 ) | ( w7881 & w7883 ) | ( w7882 & w7883 ) ;
  assign w7942 = w7939 ^ w7940 ;
  assign w7943 = w7941 ^ w7942 ;
  assign w7944 = w7899 ^ w7943 ;
  assign w7945 = w7929 ^ w7944 ;
  assign w7946 = w7857 ^ w7876 ;
  assign w7947 = w7885 ^ w7888 ;
  assign w7948 = ( w7843 & w7946 ) | ( w7843 & w7947 ) | ( w7946 & w7947 ) ;
  assign w7949 = w7898 ^ w7945 ;
  assign w7950 = w7948 ^ w7949 ;
  assign w7951 = ( w7898 & w7945 ) | ( w7898 & w7948 ) | ( w7945 & w7948 ) ;
  assign w7952 = ( w7899 & w7929 ) | ( w7899 & w7943 ) | ( w7929 & w7943 ) ;
  assign w7953 = ( w7939 & w7940 ) | ( w7939 & w7941 ) | ( w7940 & w7941 ) ;
  assign w7954 = w7903 ^ w7909 ;
  assign w7955 = w7920 ^ w7954 ;
  assign w7956 = w7912 ^ w7915 ;
  assign w7957 = ( w7905 & w7911 ) | ( w7905 & w7956 ) | ( w7911 & w7956 ) ;
  assign w7958 = w7955 ^ w7957 ;
  assign w7959 = \pi45 & \pi59 ;
  assign w7960 = \pi44 & \pi60 ;
  assign w7961 = \pi43 & \pi61 ;
  assign w7962 = ( w7959 & w7960 ) | ( w7959 & w7961 ) | ( w7960 & w7961 ) ;
  assign w7963 = w7959 ^ w7961 ;
  assign w7964 = w7960 ^ w7963 ;
  assign w7965 = \pi48 & \pi56 ;
  assign w7966 = \pi47 & \pi57 ;
  assign w7967 = \pi46 & \pi58 ;
  assign w7968 = ( w7965 & w7966 ) | ( w7965 & w7967 ) | ( w7966 & w7967 ) ;
  assign w7969 = w7965 ^ w7967 ;
  assign w7970 = w7966 ^ w7969 ;
  assign w7971 = \pi51 & \pi53 ;
  assign w7972 = \pi50 & \pi54 ;
  assign w7973 = \pi49 & \pi55 ;
  assign w7974 = ( w7971 & w7972 ) | ( w7971 & w7973 ) | ( w7972 & w7973 ) ;
  assign w7975 = w7971 ^ w7973 ;
  assign w7976 = w7972 ^ w7975 ;
  assign w7977 = w7964 ^ w7970 ;
  assign w7978 = w7976 ^ w7977 ;
  assign w7979 = w7866 ^ w7872 ;
  assign w7980 = w7928 ^ w7979 ;
  assign w7981 = ( w7916 & w7924 ) | ( w7916 & w7980 ) | ( w7924 & w7980 ) ;
  assign w7982 = ( w7933 & w7936 ) | ( w7933 & w7937 ) | ( w7936 & w7937 ) ;
  assign w7983 = \pi42 & \pi62 ;
  assign w7984 = \pi52 & \pi62 ;
  assign w7985 = ( ~\pi51 & \pi63 ) | ( ~\pi51 & w7984 ) | ( \pi63 & w7984 ) ;
  assign w7986 = ( \pi41 & \pi51 ) | ( \pi41 & w7985 ) | ( \pi51 & w7985 ) ;
  assign w7987 = ( ~\pi41 & w7984 ) | ( ~\pi41 & w7985 ) | ( w7984 & w7985 ) ;
  assign w7988 = ( ~\pi41 & \pi51 ) | ( ~\pi41 & w7985 ) | ( \pi51 & w7985 ) ;
  assign w7989 = ( \pi52 & w7987 ) | ( \pi52 & w7988 ) | ( w7987 & w7988 ) ;
  assign w7990 = w7985 ^ w7989 ;
  assign w7991 = \pi52 ^ \pi63 ;
  assign w7992 = \pi41 & ~w7991 ;
  assign w7993 = ( w7986 & w7990 ) | ( w7986 & ~w7992 ) | ( w7990 & ~w7992 ) ;
  assign w7994 = w7983 ^ w7993 ;
  assign w7995 = ( w7847 & w7860 ) | ( w7847 & w7922 ) | ( w7860 & w7922 ) ;
  assign w7996 = ( w7866 & w7872 ) | ( w7866 & w7928 ) | ( w7872 & w7928 ) ;
  assign w7997 = w7995 ^ w7996 ;
  assign w7998 = w7994 ^ w7997 ;
  assign w7999 = w7981 ^ w7982 ;
  assign w8000 = w7998 ^ w7999 ;
  assign w8001 = w7958 ^ w7978 ;
  assign w8002 = w7953 ^ w8001 ;
  assign w8003 = w8000 ^ w8002 ;
  assign w8004 = w7951 ^ w7952 ;
  assign w8005 = w8003 ^ w8004 ;
  assign w8006 = w7962 ^ w7968 ;
  assign w8007 = w7974 ^ w8006 ;
  assign w8008 = ( w7964 & w7970 ) | ( w7964 & w7976 ) | ( w7970 & w7976 ) ;
  assign w8009 = ( w7994 & w7995 ) | ( w7994 & w7996 ) | ( w7995 & w7996 ) ;
  assign w8010 = w8007 ^ w8009 ;
  assign w8011 = w8008 ^ w8010 ;
  assign w8012 = ( w7981 & w7982 ) | ( w7981 & w7998 ) | ( w7982 & w7998 ) ;
  assign w8013 = ( w7955 & w7957 ) | ( w7955 & w7978 ) | ( w7957 & w7978 ) ;
  assign w8014 = \pi51 & \pi54 ;
  assign w8015 = \pi50 & \pi55 ;
  assign w8016 = \pi49 & \pi56 ;
  assign w8017 = ( w8014 & w8015 ) | ( w8014 & w8016 ) | ( w8015 & w8016 ) ;
  assign w8018 = w8014 ^ w8016 ;
  assign w8019 = w8015 ^ w8018 ;
  assign w8020 = ( w7903 & w7909 ) | ( w7903 & w7920 ) | ( w7909 & w7920 ) ;
  assign w8021 = ~\pi52 & \pi53 ;
  assign w8022 = w8020 ^ w8021 ;
  assign w8023 = w8019 ^ w8022 ;
  assign w8024 = \pi43 & \pi62 ;
  assign w8025 = w8023 ^ w8024 ;
  assign w8026 = \pi45 & \pi60 ;
  assign w8027 = \pi44 & \pi61 ;
  assign w8028 = \pi42 & \pi63 ;
  assign w8029 = ( w8026 & w8027 ) | ( w8026 & w8028 ) | ( w8027 & w8028 ) ;
  assign w8030 = w8026 ^ w8028 ;
  assign w8031 = w8027 ^ w8030 ;
  assign w8032 = \pi41 & \pi63 ;
  assign w8033 = ( \pi41 & \pi51 ) | ( \pi41 & \pi62 ) | ( \pi51 & \pi62 ) ;
  assign w8034 = \pi52 & w8033 ;
  assign w8035 = ( w7983 & w8032 ) | ( w7983 & w8034 ) | ( w8032 & w8034 ) ;
  assign w8036 = \pi48 & \pi57 ;
  assign w8037 = \pi47 & \pi58 ;
  assign w8038 = \pi46 & \pi59 ;
  assign w8039 = ( w8036 & w8037 ) | ( w8036 & w8038 ) | ( w8037 & w8038 ) ;
  assign w8040 = w8036 ^ w8038 ;
  assign w8041 = w8037 ^ w8040 ;
  assign w8042 = w8031 ^ w8035 ;
  assign w8043 = w8041 ^ w8042 ;
  assign w8044 = w8013 ^ w8025 ;
  assign w8045 = w8043 ^ w8044 ;
  assign w8046 = w8011 ^ w8012 ;
  assign w8047 = w8045 ^ w8046 ;
  assign w8048 = ( w7953 & w8000 ) | ( w7953 & w8001 ) | ( w8000 & w8001 ) ;
  assign w8049 = ( w7951 & w7952 ) | ( w7951 & w8003 ) | ( w7952 & w8003 ) ;
  assign w8050 = w8048 ^ w8049 ;
  assign w8051 = w8047 ^ w8050 ;
  assign w8052 = ( w8047 & w8048 ) | ( w8047 & w8049 ) | ( w8048 & w8049 ) ;
  assign w8053 = ( w8011 & w8012 ) | ( w8011 & w8045 ) | ( w8012 & w8045 ) ;
  assign w8054 = ( w8007 & w8008 ) | ( w8007 & w8009 ) | ( w8008 & w8009 ) ;
  assign w8055 = \pi49 & \pi57 ;
  assign w8056 = \pi48 & \pi58 ;
  assign w8057 = \pi47 & \pi59 ;
  assign w8058 = ( w8055 & w8056 ) | ( w8055 & w8057 ) | ( w8056 & w8057 ) ;
  assign w8059 = w8055 ^ w8057 ;
  assign w8060 = w8056 ^ w8059 ;
  assign w8061 = \pi52 & \pi54 ;
  assign w8062 = \pi51 & \pi55 ;
  assign w8063 = \pi50 & \pi56 ;
  assign w8064 = ( w8061 & w8062 ) | ( w8061 & w8063 ) | ( w8062 & w8063 ) ;
  assign w8065 = w8061 ^ w8063 ;
  assign w8066 = w8062 ^ w8065 ;
  assign w8067 = ( w7962 & w7968 ) | ( w7962 & w7974 ) | ( w7968 & w7974 ) ;
  assign w8068 = w8060 ^ w8067 ;
  assign w8069 = w8066 ^ w8068 ;
  assign w8070 = \pi46 & \pi60 ;
  assign w8071 = \pi45 & \pi61 ;
  assign w8072 = \pi44 & \pi62 ;
  assign w8073 = ( w8070 & w8071 ) | ( w8070 & w8072 ) | ( w8071 & w8072 ) ;
  assign w8074 = w8070 ^ w8072 ;
  assign w8075 = w8071 ^ w8074 ;
  assign w8076 = w8029 ^ w8039 ;
  assign w8077 = w8075 ^ w8076 ;
  assign w8078 = ( w8054 & w8069 ) | ( w8054 & w8077 ) | ( w8069 & w8077 ) ;
  assign w8079 = w8054 ^ w8069 ;
  assign w8080 = w8077 ^ w8079 ;
  assign w8081 = \pi43 & \pi63 ;
  assign w8082 = w8017 ^ w8081 ;
  assign w8083 = ~\pi52 & \pi62 ;
  assign w8084 = \pi43 & w8083 ;
  assign w8085 = ( \pi52 & \pi53 ) | ( \pi52 & w8084 ) | ( \pi53 & w8084 ) ;
  assign w8086 = w8082 ^ w8085 ;
  assign w8087 = ( w8031 & w8035 ) | ( w8031 & w8041 ) | ( w8035 & w8041 ) ;
  assign w8088 = w8021 ^ w8024 ;
  assign w8089 = ( w8019 & w8020 ) | ( w8019 & w8088 ) | ( w8020 & w8088 ) ;
  assign w8090 = w8086 ^ w8089 ;
  assign w8091 = w8087 ^ w8090 ;
  assign w8092 = ( w8013 & w8025 ) | ( w8013 & w8043 ) | ( w8025 & w8043 ) ;
  assign w8093 = w8080 ^ w8091 ;
  assign w8094 = w8092 ^ w8093 ;
  assign w8095 = w8053 & w8094 ;
  assign w8096 = w8053 | w8094 ;
  assign w8097 = ~w8095 & w8096 ;
  assign w8098 = w8052 ^ w8097 ;
  assign w8099 = ( w8052 & w8095 ) | ( w8052 & w8096 ) | ( w8095 & w8096 ) ;
  assign w8100 = w8095 | w8099 ;
  assign w8101 = ( w8080 & w8091 ) | ( w8080 & w8092 ) | ( w8091 & w8092 ) ;
  assign w8102 = ( w8086 & w8087 ) | ( w8086 & w8089 ) | ( w8087 & w8089 ) ;
  assign w8103 = \pi49 & \pi58 ;
  assign w8104 = \pi48 & \pi59 ;
  assign w8105 = \pi44 & \pi63 ;
  assign w8106 = ( w8103 & w8104 ) | ( w8103 & w8105 ) | ( w8104 & w8105 ) ;
  assign w8107 = w8103 ^ w8105 ;
  assign w8108 = w8104 ^ w8107 ;
  assign w8109 = w8058 ^ w8073 ;
  assign w8110 = w8108 ^ w8109 ;
  assign w8111 = \pi52 & \pi55 ;
  assign w8112 = \pi51 & \pi56 ;
  assign w8113 = \pi50 & \pi57 ;
  assign w8114 = ( w8111 & w8112 ) | ( w8111 & w8113 ) | ( w8112 & w8113 ) ;
  assign w8115 = w8111 ^ w8113 ;
  assign w8116 = w8112 ^ w8115 ;
  assign w8117 = \pi47 & \pi60 ;
  assign w8118 = \pi46 & \pi61 ;
  assign w8119 = w8064 ^ w8118 ;
  assign w8120 = w8117 ^ w8119 ;
  assign w8121 = ~\pi53 & \pi54 ;
  assign w8122 = w8120 ^ w8121 ;
  assign w8123 = w8116 ^ w8122 ;
  assign w8124 = \pi45 & \pi62 ;
  assign w8125 = w8123 ^ w8124 ;
  assign w8126 = w8102 ^ w8125 ;
  assign w8127 = w8110 ^ w8126 ;
  assign w8128 = ( w8029 & w8039 ) | ( w8029 & w8075 ) | ( w8039 & w8075 ) ;
  assign w8129 = \pi52 & \pi53 ;
  assign w8130 = w8017 & w8129 ;
  assign w8131 = ( \pi53 & \pi62 ) | ( \pi53 & w8129 ) | ( \pi62 & w8129 ) ;
  assign w8132 = ( \pi63 & w8017 ) | ( \pi63 & w8131 ) | ( w8017 & w8131 ) ;
  assign w8133 = ( \pi43 & w8130 ) | ( \pi43 & w8132 ) | ( w8130 & w8132 ) ;
  assign w8134 = ( w8060 & w8066 ) | ( w8060 & w8067 ) | ( w8066 & w8067 ) ;
  assign w8135 = w8128 ^ w8134 ;
  assign w8136 = w8133 ^ w8135 ;
  assign w8137 = w8078 ^ w8127 ;
  assign w8138 = w8136 ^ w8137 ;
  assign w8139 = w8100 ^ w8101 ;
  assign w8140 = w8138 ^ w8139 ;
  assign w8141 = ( w8100 & w8101 ) | ( w8100 & w8138 ) | ( w8101 & w8138 ) ;
  assign w8142 = ( w8078 & w8127 ) | ( w8078 & w8136 ) | ( w8127 & w8136 ) ;
  assign w8143 = ( w8058 & w8073 ) | ( w8058 & w8108 ) | ( w8073 & w8108 ) ;
  assign w8144 = \pi53 & \pi55 ;
  assign w8145 = \pi52 & \pi56 ;
  assign w8146 = \pi51 & \pi57 ;
  assign w8147 = ( w8144 & w8145 ) | ( w8144 & w8146 ) | ( w8145 & w8146 ) ;
  assign w8148 = w8144 ^ w8146 ;
  assign w8149 = w8145 ^ w8148 ;
  assign w8150 = w8121 ^ w8124 ;
  assign w8151 = ( w8116 & w8120 ) | ( w8116 & w8150 ) | ( w8120 & w8150 ) ;
  assign w8152 = w8143 ^ w8151 ;
  assign w8153 = w8149 ^ w8152 ;
  assign w8154 = ( w8102 & w8110 ) | ( w8102 & w8125 ) | ( w8110 & w8125 ) ;
  assign w8155 = w8106 ^ w8114 ;
  assign w8156 = ( \pi45 & \pi53 ) | ( \pi45 & \pi62 ) | ( \pi53 & \pi62 ) ;
  assign w8157 = ~\pi53 & w8156 ;
  assign w8158 = ( \pi53 & \pi54 ) | ( \pi53 & w8157 ) | ( \pi54 & w8157 ) ;
  assign w8159 = w8155 ^ w8158 ;
  assign w8160 = ( w8128 & w8133 ) | ( w8128 & w8134 ) | ( w8133 & w8134 ) ;
  assign w8161 = w8159 ^ w8160 ;
  assign w8162 = \pi47 & \pi61 ;
  assign w8163 = \pi46 & \pi62 ;
  assign w8164 = \pi45 & \pi63 ;
  assign w8165 = ( w8162 & w8163 ) | ( w8162 & w8164 ) | ( w8163 & w8164 ) ;
  assign w8166 = w8162 ^ w8164 ;
  assign w8167 = w8163 ^ w8166 ;
  assign w8168 = ( w8064 & w8117 ) | ( w8064 & w8118 ) | ( w8117 & w8118 ) ;
  assign w8169 = \pi50 & \pi58 ;
  assign w8170 = \pi49 & \pi59 ;
  assign w8171 = \pi48 & \pi60 ;
  assign w8172 = ( w8169 & w8170 ) | ( w8169 & w8171 ) | ( w8170 & w8171 ) ;
  assign w8173 = w8169 ^ w8171 ;
  assign w8174 = w8170 ^ w8173 ;
  assign w8175 = w8167 ^ w8168 ;
  assign w8176 = w8174 ^ w8175 ;
  assign w8177 = w8153 ^ w8176 ;
  assign w8178 = w8154 ^ w8177 ;
  assign w8179 = w8161 ^ w8178 ;
  assign w8180 = w8142 | w8179 ;
  assign w8181 = w8142 & w8179 ;
  assign w8182 = w8180 & ~w8181 ;
  assign w8183 = w8141 ^ w8182 ;
  assign w8184 = ( w8141 & w8180 ) | ( w8141 & w8181 ) | ( w8180 & w8181 ) ;
  assign w8185 = w8181 | w8184 ;
  assign w8186 = ( \pi54 & w3491 ) | ( \pi54 & w8156 ) | ( w3491 & w8156 ) ;
  assign w8187 = ( w8106 & w8114 ) | ( w8106 & w8186 ) | ( w8114 & w8186 ) ;
  assign w8188 = ( w8167 & w8168 ) | ( w8167 & w8174 ) | ( w8168 & w8174 ) ;
  assign w8189 = ~\pi54 & \pi55 ;
  assign w8190 = w8188 ^ w8189 ;
  assign w8191 = w8187 ^ w8190 ;
  assign w8192 = \pi47 & \pi62 ;
  assign w8193 = w8191 ^ w8192 ;
  assign w8194 = ( w8159 & w8160 ) | ( w8159 & w8176 ) | ( w8160 & w8176 ) ;
  assign w8195 = ( w8143 & w8149 ) | ( w8143 & w8151 ) | ( w8149 & w8151 ) ;
  assign w8196 = \pi46 & \pi63 ;
  assign w8197 = w8147 ^ w8172 ;
  assign w8198 = w8195 ^ w8197 ;
  assign w8199 = w8196 ^ w8198 ;
  assign w8200 = \pi50 & \pi59 ;
  assign w8201 = \pi49 & \pi60 ;
  assign w8202 = \pi48 & \pi61 ;
  assign w8203 = ( w8200 & w8201 ) | ( w8200 & w8202 ) | ( w8201 & w8202 ) ;
  assign w8204 = w8200 ^ w8202 ;
  assign w8205 = w8201 ^ w8204 ;
  assign w8206 = \pi53 & \pi56 ;
  assign w8207 = \pi52 & \pi57 ;
  assign w8208 = \pi51 & \pi58 ;
  assign w8209 = ( w8206 & w8207 ) | ( w8206 & w8208 ) | ( w8207 & w8208 ) ;
  assign w8210 = w8206 ^ w8208 ;
  assign w8211 = w8207 ^ w8210 ;
  assign w8212 = w8165 ^ w8205 ;
  assign w8213 = w8211 ^ w8212 ;
  assign w8214 = w8193 ^ w8213 ;
  assign w8215 = w8194 ^ w8214 ;
  assign w8216 = w8199 ^ w8215 ;
  assign w8217 = w8161 ^ w8176 ;
  assign w8218 = ( w8153 & w8154 ) | ( w8153 & w8217 ) | ( w8154 & w8217 ) ;
  assign w8219 = w8185 ^ w8216 ;
  assign w8220 = w8218 ^ w8219 ;
  assign w8221 = ( w8185 & w8216 ) | ( w8185 & w8218 ) | ( w8216 & w8218 ) ;
  assign w8222 = w8199 ^ w8213 ;
  assign w8223 = ( w8193 & w8194 ) | ( w8193 & w8222 ) | ( w8194 & w8222 ) ;
  assign w8224 = \pi51 & \pi59 ;
  assign w8225 = \pi50 & \pi60 ;
  assign w8226 = \pi49 & \pi61 ;
  assign w8227 = ( w8224 & w8225 ) | ( w8224 & w8226 ) | ( w8225 & w8226 ) ;
  assign w8228 = w8224 ^ w8226 ;
  assign w8229 = w8225 ^ w8228 ;
  assign w8230 = w8203 ^ w8209 ;
  assign w8231 = w8229 ^ w8230 ;
  assign w8232 = ( w8165 & w8205 ) | ( w8165 & w8211 ) | ( w8205 & w8211 ) ;
  assign w8233 = w8189 ^ w8192 ;
  assign w8234 = ( w8187 & w8188 ) | ( w8187 & w8233 ) | ( w8188 & w8233 ) ;
  assign w8235 = w8231 ^ w8234 ;
  assign w8236 = w8232 ^ w8235 ;
  assign w8237 = \pi54 & \pi56 ;
  assign w8238 = \pi53 & \pi57 ;
  assign w8239 = \pi52 & \pi58 ;
  assign w8240 = ( w8237 & w8238 ) | ( w8237 & w8239 ) | ( w8238 & w8239 ) ;
  assign w8241 = w8237 ^ w8239 ;
  assign w8242 = w8238 ^ w8241 ;
  assign w8243 = \pi48 & \pi62 ;
  assign w8244 = \pi55 & \pi62 ;
  assign w8245 = ( ~\pi54 & \pi63 ) | ( ~\pi54 & w8244 ) | ( \pi63 & w8244 ) ;
  assign w8246 = ( \pi47 & \pi54 ) | ( \pi47 & w8245 ) | ( \pi54 & w8245 ) ;
  assign w8247 = ( ~\pi47 & w8244 ) | ( ~\pi47 & w8245 ) | ( w8244 & w8245 ) ;
  assign w8248 = ( ~\pi47 & \pi54 ) | ( ~\pi47 & w8245 ) | ( \pi54 & w8245 ) ;
  assign w8249 = ( \pi55 & w8247 ) | ( \pi55 & w8248 ) | ( w8247 & w8248 ) ;
  assign w8250 = w8245 ^ w8249 ;
  assign w8251 = \pi55 ^ \pi63 ;
  assign w8252 = \pi47 & ~w8251 ;
  assign w8253 = ( w8246 & w8250 ) | ( w8246 & ~w8252 ) | ( w8250 & ~w8252 ) ;
  assign w8254 = w8243 ^ w8253 ;
  assign w8255 = ( w8147 & w8172 ) | ( w8147 & w8196 ) | ( w8172 & w8196 ) ;
  assign w8256 = w8242 ^ w8255 ;
  assign w8257 = w8254 ^ w8256 ;
  assign w8258 = w8196 ^ w8197 ;
  assign w8259 = ( w8195 & w8213 ) | ( w8195 & w8258 ) | ( w8213 & w8258 ) ;
  assign w8260 = w8236 ^ w8259 ;
  assign w8261 = w8257 ^ w8260 ;
  assign w8262 = w8221 ^ w8223 ;
  assign w8263 = w8261 ^ w8262 ;
  assign w8264 = ( w8221 & w8223 ) | ( w8221 & w8261 ) | ( w8223 & w8261 ) ;
  assign w8265 = ( w8236 & w8257 ) | ( w8236 & w8259 ) | ( w8257 & w8259 ) ;
  assign w8266 = \pi47 & \pi63 ;
  assign w8267 = ( \pi47 & \pi54 ) | ( \pi47 & \pi62 ) | ( \pi54 & \pi62 ) ;
  assign w8268 = \pi55 & w8267 ;
  assign w8269 = ( w8243 & w8266 ) | ( w8243 & w8268 ) | ( w8266 & w8268 ) ;
  assign w8270 = w8227 ^ w8240 ;
  assign w8271 = w8269 ^ w8270 ;
  assign w8272 = ( w8203 & w8209 ) | ( w8203 & w8229 ) | ( w8209 & w8229 ) ;
  assign w8273 = ( w8242 & w8254 ) | ( w8242 & w8255 ) | ( w8254 & w8255 ) ;
  assign w8274 = w8271 ^ w8272 ;
  assign w8275 = w8273 ^ w8274 ;
  assign w8276 = \pi51 & \pi60 ;
  assign w8277 = \pi50 & \pi61 ;
  assign w8278 = \pi48 & \pi63 ;
  assign w8279 = ( w8276 & w8277 ) | ( w8276 & w8278 ) | ( w8277 & w8278 ) ;
  assign w8280 = w8276 ^ w8278 ;
  assign w8281 = w8277 ^ w8280 ;
  assign w8282 = \pi54 & \pi57 ;
  assign w8283 = \pi53 & \pi58 ;
  assign w8284 = \pi52 & \pi59 ;
  assign w8285 = ( w8282 & w8283 ) | ( w8282 & w8284 ) | ( w8283 & w8284 ) ;
  assign w8286 = w8282 ^ w8284 ;
  assign w8287 = w8283 ^ w8286 ;
  assign w8288 = ~\pi55 & \pi56 ;
  assign w8289 = w8281 ^ w8288 ;
  assign w8290 = w8287 ^ w8289 ;
  assign w8291 = \pi49 & \pi62 ;
  assign w8292 = w8290 ^ w8291 ;
  assign w8293 = ( w8231 & w8232 ) | ( w8231 & w8234 ) | ( w8232 & w8234 ) ;
  assign w8294 = w8275 ^ w8293 ;
  assign w8295 = w8292 ^ w8294 ;
  assign w8296 = w8264 ^ w8265 ;
  assign w8297 = w8295 ^ w8296 ;
  assign w8298 = ( w8264 & w8265 ) | ( w8264 & w8295 ) | ( w8265 & w8295 ) ;
  assign w8299 = ( w8275 & w8292 ) | ( w8275 & w8293 ) | ( w8292 & w8293 ) ;
  assign w8300 = ( w8271 & w8272 ) | ( w8271 & w8273 ) | ( w8272 & w8273 ) ;
  assign w8301 = \pi52 & \pi60 ;
  assign w8302 = \pi51 & \pi61 ;
  assign w8303 = \pi49 & \pi63 ;
  assign w8304 = ( w8301 & w8302 ) | ( w8301 & w8303 ) | ( w8302 & w8303 ) ;
  assign w8305 = w8301 ^ w8303 ;
  assign w8306 = w8302 ^ w8305 ;
  assign w8307 = \pi55 & \pi57 ;
  assign w8308 = \pi54 & \pi58 ;
  assign w8309 = \pi53 & \pi59 ;
  assign w8310 = ( w8307 & w8308 ) | ( w8307 & w8309 ) | ( w8308 & w8309 ) ;
  assign w8311 = w8307 ^ w8309 ;
  assign w8312 = w8308 ^ w8311 ;
  assign w8313 = w8279 ^ w8306 ;
  assign w8314 = w8312 ^ w8313 ;
  assign w8315 = \pi50 & \pi62 ;
  assign w8316 = w8285 ^ w8315 ;
  assign w8317 = \pi49 & ~\pi55 ;
  assign w8318 = \pi62 & w8317 ;
  assign w8319 = ( \pi55 & \pi56 ) | ( \pi55 & w8318 ) | ( \pi56 & w8318 ) ;
  assign w8320 = w8316 ^ w8319 ;
  assign w8321 = ( w8227 & w8240 ) | ( w8227 & w8269 ) | ( w8240 & w8269 ) ;
  assign w8322 = w8288 ^ w8291 ;
  assign w8323 = ( w8281 & w8287 ) | ( w8281 & w8322 ) | ( w8287 & w8322 ) ;
  assign w8324 = w8320 ^ w8321 ;
  assign w8325 = w8323 ^ w8324 ;
  assign w8326 = w8300 ^ w8325 ;
  assign w8327 = w8314 ^ w8326 ;
  assign w8328 = w8298 ^ w8299 ;
  assign w8329 = w8327 ^ w8328 ;
  assign w8330 = ( w8298 & w8299 ) | ( w8298 & w8327 ) | ( w8299 & w8327 ) ;
  assign w8331 = ( w8300 & w8314 ) | ( w8300 & w8325 ) | ( w8314 & w8325 ) ;
  assign w8332 = \pi53 & \pi60 ;
  assign w8333 = \pi52 & \pi61 ;
  assign w8334 = w8310 ^ w8333 ;
  assign w8335 = w8332 ^ w8334 ;
  assign w8336 = \pi55 & \pi56 ;
  assign w8337 = w8285 & w8336 ;
  assign w8338 = ( \pi49 & \pi56 ) | ( \pi49 & w8336 ) | ( \pi56 & w8336 ) ;
  assign w8339 = ( \pi50 & w8285 ) | ( \pi50 & w8338 ) | ( w8285 & w8338 ) ;
  assign w8340 = ( \pi62 & w8337 ) | ( \pi62 & w8339 ) | ( w8337 & w8339 ) ;
  assign w8341 = ( w8279 & w8306 ) | ( w8279 & w8312 ) | ( w8306 & w8312 ) ;
  assign w8342 = w8335 ^ w8340 ;
  assign w8343 = w8341 ^ w8342 ;
  assign w8344 = ( w8320 & w8321 ) | ( w8320 & w8323 ) | ( w8321 & w8323 ) ;
  assign w8345 = \pi55 & \pi58 ;
  assign w8346 = \pi54 & \pi59 ;
  assign w8347 = \pi50 & \pi63 ;
  assign w8348 = ( w8345 & w8346 ) | ( w8345 & w8347 ) | ( w8346 & w8347 ) ;
  assign w8349 = w8345 ^ w8347 ;
  assign w8350 = w8346 ^ w8349 ;
  assign w8351 = ~\pi56 & \pi57 ;
  assign w8352 = w8304 ^ w8351 ;
  assign w8353 = w8350 ^ w8352 ;
  assign w8354 = \pi51 & \pi62 ;
  assign w8355 = w8353 ^ w8354 ;
  assign w8356 = w8343 ^ w8344 ;
  assign w8357 = w8355 ^ w8356 ;
  assign w8358 = w8330 ^ w8331 ;
  assign w8359 = w8357 ^ w8358 ;
  assign w8360 = ( w8330 & w8331 ) | ( w8330 & w8357 ) | ( w8331 & w8357 ) ;
  assign w8361 = ( w8343 & w8344 ) | ( w8343 & w8355 ) | ( w8344 & w8355 ) ;
  assign w8362 = ( w8310 & w8332 ) | ( w8310 & w8333 ) | ( w8332 & w8333 ) ;
  assign w8363 = w8348 ^ w8362 ;
  assign w8364 = ( \pi51 & \pi56 ) | ( \pi51 & \pi62 ) | ( \pi56 & \pi62 ) ;
  assign w8365 = ~\pi56 & w8364 ;
  assign w8366 = ( \pi56 & \pi57 ) | ( \pi56 & w8365 ) | ( \pi57 & w8365 ) ;
  assign w8367 = w8363 ^ w8366 ;
  assign w8368 = ( w8335 & w8340 ) | ( w8335 & w8341 ) | ( w8340 & w8341 ) ;
  assign w8369 = \pi53 & \pi61 ;
  assign w8370 = \pi51 & \pi63 ;
  assign w8371 = ( w7984 & w8369 ) | ( w7984 & w8370 ) | ( w8369 & w8370 ) ;
  assign w8372 = w8369 ^ w8370 ;
  assign w8373 = w7984 ^ w8372 ;
  assign w8374 = \pi56 & \pi58 ;
  assign w8375 = \pi55 & \pi59 ;
  assign w8376 = \pi54 & \pi60 ;
  assign w8377 = ( w8374 & w8375 ) | ( w8374 & w8376 ) | ( w8375 & w8376 ) ;
  assign w8378 = w8374 ^ w8376 ;
  assign w8379 = w8375 ^ w8378 ;
  assign w8380 = w8351 ^ w8354 ;
  assign w8381 = ( w8304 & w8350 ) | ( w8304 & w8380 ) | ( w8350 & w8380 ) ;
  assign w8382 = w8373 ^ w8381 ;
  assign w8383 = w8379 ^ w8382 ;
  assign w8384 = w8367 ^ w8368 ;
  assign w8385 = w8383 ^ w8384 ;
  assign w8386 = w8360 ^ w8361 ;
  assign w8387 = w8385 ^ w8386 ;
  assign w8388 = ( w8360 & w8361 ) | ( w8360 & w8385 ) | ( w8361 & w8385 ) ;
  assign w8389 = ( w8367 & w8368 ) | ( w8367 & w8383 ) | ( w8368 & w8383 ) ;
  assign w8390 = \pi56 & \pi59 ;
  assign w8391 = \pi55 & \pi60 ;
  assign w8392 = \pi54 & \pi61 ;
  assign w8393 = ( w8390 & w8391 ) | ( w8390 & w8392 ) | ( w8391 & w8392 ) ;
  assign w8394 = w8390 ^ w8392 ;
  assign w8395 = w8391 ^ w8394 ;
  assign w8396 = \pi56 & \pi57 ;
  assign w8397 = ( \pi57 & w8364 ) | ( \pi57 & w8396 ) | ( w8364 & w8396 ) ;
  assign w8398 = ( w8348 & w8362 ) | ( w8348 & w8397 ) | ( w8362 & w8397 ) ;
  assign w8399 = ~\pi57 & \pi58 ;
  assign w8400 = w8398 ^ w8399 ;
  assign w8401 = w8395 ^ w8400 ;
  assign w8402 = \pi53 & \pi62 ;
  assign w8403 = w8401 ^ w8402 ;
  assign w8404 = ( w8373 & w8379 ) | ( w8373 & w8381 ) | ( w8379 & w8381 ) ;
  assign w8405 = w8403 ^ w8404 ;
  assign w8406 = w8371 ^ w8405 ;
  assign w8407 = w8377 ^ w8406 ;
  assign w8408 = \pi52 & \pi63 ;
  assign w8409 = w8407 ^ w8408 ;
  assign w8410 = w8388 ^ w8409 ;
  assign w8411 = w8389 ^ w8410 ;
  assign w8412 = ( w8388 & w8389 ) | ( w8388 & w8409 ) | ( w8389 & w8409 ) ;
  assign w8413 = w8399 ^ w8402 ;
  assign w8414 = ( w8395 & w8398 ) | ( w8395 & w8413 ) | ( w8398 & w8413 ) ;
  assign w8415 = ( \pi57 & \pi58 ) | ( \pi57 & w8402 ) | ( \pi58 & w8402 ) ;
  assign w8416 = ( \pi54 & ~\pi58 ) | ( \pi54 & \pi62 ) | ( ~\pi58 & \pi62 ) ;
  assign w8417 = ( \pi53 & ~\pi58 ) | ( \pi53 & \pi63 ) | ( ~\pi58 & \pi63 ) ;
  assign w8418 = w8416 ^ w8417 ;
  assign w8419 = w8415 & w8418 ;
  assign w8420 = \pi54 & \pi62 ;
  assign w8421 = \pi58 & \pi62 ;
  assign w8422 = ( ~\pi57 & \pi63 ) | ( ~\pi57 & w8421 ) | ( \pi63 & w8421 ) ;
  assign w8423 = ( \pi53 & \pi57 ) | ( \pi53 & w8422 ) | ( \pi57 & w8422 ) ;
  assign w8424 = ( ~\pi53 & w8421 ) | ( ~\pi53 & w8422 ) | ( w8421 & w8422 ) ;
  assign w8425 = ( ~\pi53 & \pi57 ) | ( ~\pi53 & w8422 ) | ( \pi57 & w8422 ) ;
  assign w8426 = ( \pi58 & w8424 ) | ( \pi58 & w8425 ) | ( w8424 & w8425 ) ;
  assign w8427 = w8422 ^ w8426 ;
  assign w8428 = \pi58 ^ \pi63 ;
  assign w8429 = \pi53 & ~w8428 ;
  assign w8430 = ( w8423 & w8427 ) | ( w8423 & ~w8429 ) | ( w8427 & ~w8429 ) ;
  assign w8431 = w8420 ^ w8430 ;
  assign w8432 = \pi57 & \pi59 ;
  assign w8433 = \pi56 & \pi60 ;
  assign w8434 = \pi55 & \pi61 ;
  assign w8435 = ( w8432 & w8433 ) | ( w8432 & w8434 ) | ( w8433 & w8434 ) ;
  assign w8436 = w8432 ^ w8434 ;
  assign w8437 = w8433 ^ w8436 ;
  assign w8438 = w8393 ^ w8431 ;
  assign w8439 = w8437 ^ w8438 ;
  assign w8440 = ( w8371 & w8377 ) | ( w8371 & w8408 ) | ( w8377 & w8408 ) ;
  assign w8441 = w8414 ^ w8440 ;
  assign w8442 = w8439 ^ w8441 ;
  assign w8443 = w8371 ^ w8377 ;
  assign w8444 = w8408 ^ w8443 ;
  assign w8445 = ( w8403 & w8404 ) | ( w8403 & w8444 ) | ( w8404 & w8444 ) ;
  assign w8446 = w8412 ^ w8442 ;
  assign w8447 = w8445 ^ w8446 ;
  assign w8448 = ( w8412 & w8442 ) | ( w8412 & w8445 ) | ( w8442 & w8445 ) ;
  assign w8449 = ( w8414 & w8439 ) | ( w8414 & w8440 ) | ( w8439 & w8440 ) ;
  assign w8450 = \pi57 & \pi60 ;
  assign w8451 = \pi56 & \pi61 ;
  assign w8452 = \pi54 & \pi63 ;
  assign w8453 = ( w8450 & w8451 ) | ( w8450 & w8452 ) | ( w8451 & w8452 ) ;
  assign w8454 = w8450 ^ w8452 ;
  assign w8455 = w8451 ^ w8454 ;
  assign w8456 = ~\pi62 & w3491 ;
  assign w8457 = ( w3491 & w8419 ) | ( w3491 & ~w8456 ) | ( w8419 & ~w8456 ) ;
  assign w8458 = ( \pi63 & w8419 ) | ( \pi63 & w8457 ) | ( w8419 & w8457 ) ;
  assign w8459 = w8435 ^ w8455 ;
  assign w8460 = w8458 ^ w8459 ;
  assign w8461 = ( w8393 & w8431 ) | ( w8393 & w8437 ) | ( w8431 & w8437 ) ;
  assign w8462 = ~\pi58 & \pi59 ;
  assign w8463 = w8460 ^ w8462 ;
  assign w8464 = w8461 ^ w8463 ;
  assign w8465 = w8244 ^ w8464 ;
  assign w8466 = w8448 ^ w8449 ;
  assign w8467 = w8465 ^ w8466 ;
  assign w8468 = ( \pi55 & w4068 ) | ( \pi55 & ~w7373 ) | ( w4068 & ~w7373 ) ;
  assign w8469 = \pi63 ^ w8468 ;
  assign w8470 = \pi55 & ~w8469 ;
  assign w8471 = w4068 ^ w8453 ;
  assign w8472 = w8470 ^ w8471 ;
  assign w8473 = \pi62 | w8419 ;
  assign w8474 = ( \pi63 & w8419 ) | ( \pi63 & w8473 ) | ( w8419 & w8473 ) ;
  assign w8475 = ( w3491 & w8419 ) | ( w3491 & w8474 ) | ( w8419 & w8474 ) ;
  assign w8476 = ( w8435 & w8455 ) | ( w8435 & w8475 ) | ( w8455 & w8475 ) ;
  assign w8477 = \pi58 & \pi60 ;
  assign w8478 = \pi57 & \pi61 ;
  assign w8479 = \pi56 & \pi62 ;
  assign w8480 = ( w8477 & w8478 ) | ( w8477 & w8479 ) | ( w8478 & w8479 ) ;
  assign w8481 = w8477 ^ w8479 ;
  assign w8482 = w8478 ^ w8481 ;
  assign w8483 = w8472 ^ w8476 ;
  assign w8484 = w8482 ^ w8483 ;
  assign w8485 = w8244 ^ w8462 ;
  assign w8486 = ( w8460 & w8461 ) | ( w8460 & w8485 ) | ( w8461 & w8485 ) ;
  assign w8487 = ( w8448 & w8449 ) | ( w8448 & w8465 ) | ( w8449 & w8465 ) ;
  assign w8488 = w8484 ^ w8487 ;
  assign w8489 = w8486 ^ w8488 ;
  assign w8490 = \pi58 & \pi61 ;
  assign w8491 = \pi56 & \pi63 ;
  assign w8492 = w8480 ^ w8491 ;
  assign w8493 = w8490 ^ w8492 ;
  assign w8494 = \pi55 & \pi63 ;
  assign w8495 = ~\pi55 & w7373 ;
  assign w8496 = ( w4068 & w7373 ) | ( w4068 & ~w8495 ) | ( w7373 & ~w8495 ) ;
  assign w8497 = ( w8453 & w8494 ) | ( w8453 & w8496 ) | ( w8494 & w8496 ) ;
  assign w8498 = ~\pi59 & \pi60 ;
  assign w8499 = w8493 ^ w8498 ;
  assign w8500 = w8497 ^ w8499 ;
  assign w8501 = \pi57 & \pi62 ;
  assign w8502 = w8500 ^ w8501 ;
  assign w8503 = ( w8472 & w8476 ) | ( w8472 & w8482 ) | ( w8476 & w8482 ) ;
  assign w8504 = ( w8484 & w8486 ) | ( w8484 & w8487 ) | ( w8486 & w8487 ) ;
  assign w8505 = w8502 ^ w8504 ;
  assign w8506 = w8503 ^ w8505 ;
  assign w8507 = ( w8502 & w8503 ) | ( w8502 & w8504 ) | ( w8503 & w8504 ) ;
  assign w8508 = w8498 ^ w8501 ;
  assign w8509 = ( w8493 & w8497 ) | ( w8493 & w8508 ) | ( w8497 & w8508 ) ;
  assign w8510 = ( w8480 & w8490 ) | ( w8480 & w8491 ) | ( w8490 & w8491 ) ;
  assign w8511 = \pi59 & \pi61 ;
  assign w8512 = \pi57 & \pi63 ;
  assign w8513 = ( w8421 & w8511 ) | ( w8421 & w8512 ) | ( w8511 & w8512 ) ;
  assign w8514 = w8511 ^ w8512 ;
  assign w8515 = w8421 ^ w8514 ;
  assign w8516 = w8510 ^ w8515 ;
  assign w8517 = ( \pi57 & \pi59 ) | ( \pi57 & \pi62 ) | ( \pi59 & \pi62 ) ;
  assign w8518 = ~\pi59 & w8517 ;
  assign w8519 = ( \pi59 & \pi60 ) | ( \pi59 & w8518 ) | ( \pi60 & w8518 ) ;
  assign w8520 = w8516 ^ w8519 ;
  assign w8521 = w8507 ^ w8509 ;
  assign w8522 = w8520 ^ w8521 ;
  assign w8523 = \pi58 & \pi63 ;
  assign w8524 = w8513 ^ w8523 ;
  assign w8525 = ( \pi60 & w4299 ) | ( \pi60 & w8517 ) | ( w4299 & w8517 ) ;
  assign w8526 = ( w8510 & w8515 ) | ( w8510 & w8525 ) | ( w8515 & w8525 ) ;
  assign w8527 = ( w8507 & w8509 ) | ( w8507 & w8520 ) | ( w8509 & w8520 ) ;
  assign w8528 = w8526 ^ w8527 ;
  assign w8529 = w8524 ^ w8528 ;
  assign w8530 = w7373 ^ w8529 ;
  assign w8531 = ~\pi60 & \pi61 ;
  assign w8532 = w8530 ^ w8531 ;
  assign w8533 = w7373 ^ w8524 ;
  assign w8534 = w8531 ^ w8533 ;
  assign w8535 = ( w8526 & w8527 ) | ( w8526 & w8534 ) | ( w8527 & w8534 ) ;
  assign w8536 = \pi59 & ~\pi63 ;
  assign w8537 = ( \pi59 & \pi60 ) | ( \pi59 & ~\pi61 ) | ( \pi60 & ~\pi61 ) ;
  assign w8538 = ( \pi59 & ~\pi62 ) | ( \pi59 & w8537 ) | ( ~\pi62 & w8537 ) ;
  assign w8539 = \pi60 ^ w8538 ;
  assign w8540 = \pi61 ^ \pi62 ;
  assign w8541 = \pi59 ^ w8540 ;
  assign w8542 = ( w8538 & w8539 ) | ( w8538 & w8541 ) | ( w8539 & w8541 ) ;
  assign w8543 = w8536 ^ w8542 ;
  assign w8544 = w7373 ^ w8531 ;
  assign w8545 = ( w8513 & w8523 ) | ( w8513 & w8544 ) | ( w8523 & w8544 ) ;
  assign w8546 = w8535 ^ w8545 ;
  assign w8547 = w8543 ^ w8546 ;
  assign w8548 = ( w8535 & w8543 ) | ( w8535 & w8545 ) | ( w8543 & w8545 ) ;
  assign w8549 = ( \pi62 & \pi63 ) | ( \pi62 & ~w8548 ) | ( \pi63 & ~w8548 ) ;
  assign w8550 = \pi59 & \pi63 ;
  assign w8551 = ( ~\pi62 & \pi63 ) | ( ~\pi62 & w8548 ) | ( \pi63 & w8548 ) ;
  assign w8552 = ( \pi60 & w8550 ) | ( \pi60 & ~w8551 ) | ( w8550 & ~w8551 ) ;
  assign w8553 = ( \pi63 & ~w8549 ) | ( \pi63 & w8552 ) | ( ~w8549 & w8552 ) ;
  assign w8554 = \pi60 ^ w8553 ;
  assign w8555 = \pi62 | w8550 ;
  assign w8556 = ( \pi61 & ~w8548 ) | ( \pi61 & w8555 ) | ( ~w8548 & w8555 ) ;
  assign w8557 = \pi60 ^ w8550 ;
  assign w8558 = ( \pi61 & ~w8548 ) | ( \pi61 & w8557 ) | ( ~w8548 & w8557 ) ;
  assign w8559 = w8556 & ~w8558 ;
  assign w8560 = \pi60 | \pi63 ;
  assign w8561 = ~\pi62 & w8548 ;
  assign w8562 = ~w8560 & w8561 ;
  assign w8563 = w8559 | w8562 ;
  assign w8564 = w8554 | w8563 ;
  assign w8565 = ( \pi59 & ~\pi62 ) | ( \pi59 & w8548 ) | ( ~\pi62 & w8548 ) ;
  assign w8566 = ( \pi60 & \pi62 ) | ( \pi60 & w8548 ) | ( \pi62 & w8548 ) ;
  assign w8567 = w8565 & w8566 ;
  assign w8568 = ( \pi59 & \pi61 ) | ( \pi59 & \pi62 ) | ( \pi61 & \pi62 ) ;
  assign w8569 = w4300 & w8568 ;
  assign w8570 = ( \pi63 & w8567 ) | ( \pi63 & w8569 ) | ( w8567 & w8569 ) ;
  assign w8571 = \pi63 & w8570 ;
  assign w8572 = ( \pi60 & ~\pi62 ) | ( \pi60 & \pi63 ) | ( ~\pi62 & \pi63 ) ;
  assign w8573 = ( \pi60 & ~\pi61 ) | ( \pi60 & \pi62 ) | ( ~\pi61 & \pi62 ) ;
  assign w8574 = ~w8572 & w8573 ;
  assign w8575 = ( w8548 & w8571 ) | ( w8548 & w8574 ) | ( w8571 & w8574 ) ;
  assign w8576 = w8571 | w8575 ;
  assign w8577 = \pi62 ^ \pi63 ;
  assign w8578 = ~\pi61 & w8577 ;
  assign w8579 = \pi60 & \pi62 ;
  assign w8580 = ( ~\pi61 & w8578 ) | ( ~\pi61 & w8579 ) | ( w8578 & w8579 ) ;
  assign w8581 = w8576 ^ w8580 ;
  assign w8582 = w8577 ^ w8581 ;
  assign w8583 = ( \pi62 & \pi63 ) | ( \pi62 & ~w8576 ) | ( \pi63 & ~w8576 ) ;
  assign w8584 = ( \pi62 & \pi63 ) | ( \pi62 & ~w8583 ) | ( \pi63 & ~w8583 ) ;
  assign w8585 = \pi60 & w8576 ;
  assign w8586 = w8583 & w8585 ;
  assign w8587 = ( \pi61 & w8584 ) | ( \pi61 & w8586 ) | ( w8584 & w8586 ) ;
  assign w8588 = ~\pi62 & \pi63 ;
  assign w8589 = w8587 ^ w8588 ;
  assign w8590 = ( \pi62 & \pi63 ) | ( \pi62 & w8587 ) | ( \pi63 & w8587 ) ;
  assign w8591 = \pi63 & w8590 ;
  assign \po000 = \pi00 ;
  assign \po001 = zero ;
  assign \po002 = w65 ;
  assign \po003 = w67 ;
  assign \po004 = w71 ;
  assign \po005 = w76 ;
  assign \po006 = w86 ;
  assign \po007 = w100 ;
  assign \po008 = w120 ;
  assign \po009 = w139 ;
  assign \po010 = w160 ;
  assign \po011 = w186 ;
  assign \po012 = w213 ;
  assign \po013 = w241 ;
  assign \po014 = w266 ;
  assign \po015 = w298 ;
  assign \po016 = w330 ;
  assign \po017 = w363 ;
  assign \po018 = w403 ;
  assign \po019 = w441 ;
  assign \po020 = w482 ;
  assign \po021 = w528 ;
  assign \po022 = w575 ;
  assign \po023 = w625 ;
  assign \po024 = w679 ;
  assign \po025 = w733 ;
  assign \po026 = w785 ;
  assign \po027 = w838 ;
  assign \po028 = w892 ;
  assign \po029 = w948 ;
  assign \po030 = w1012 ;
  assign \po031 = w1072 ;
  assign \po032 = w1141 ;
  assign \po033 = w1210 ;
  assign \po034 = w1280 ;
  assign \po035 = w1350 ;
  assign \po036 = w1428 ;
  assign \po037 = w1500 ;
  assign \po038 = w1578 ;
  assign \po039 = w1660 ;
  assign \po040 = w1742 ;
  assign \po041 = w1830 ;
  assign \po042 = w1916 ;
  assign \po043 = w2007 ;
  assign \po044 = w2098 ;
  assign \po045 = w2192 ;
  assign \po046 = w2285 ;
  assign \po047 = w2378 ;
  assign \po048 = w2476 ;
  assign \po049 = w2576 ;
  assign \po050 = w2678 ;
  assign \po051 = w2785 ;
  assign \po052 = w2891 ;
  assign \po053 = w3004 ;
  assign \po054 = w3115 ;
  assign \po055 = w3223 ;
  assign \po056 = w3331 ;
  assign \po057 = w3443 ;
  assign \po058 = w3565 ;
  assign \po059 = w3690 ;
  assign \po060 = w3814 ;
  assign \po061 = w3934 ;
  assign \po062 = w4064 ;
  assign \po063 = w4194 ;
  assign \po064 = w4324 ;
  assign \po065 = w4451 ;
  assign \po066 = w4581 ;
  assign \po067 = w4703 ;
  assign \po068 = w4827 ;
  assign \po069 = w4944 ;
  assign \po070 = w5061 ;
  assign \po071 = w5182 ;
  assign \po072 = w5295 ;
  assign \po073 = w5406 ;
  assign \po074 = w5516 ;
  assign \po075 = w5624 ;
  assign \po076 = w5728 ;
  assign \po077 = w5838 ;
  assign \po078 = w5940 ;
  assign \po079 = w6044 ;
  assign \po080 = w6147 ;
  assign \po081 = w6245 ;
  assign \po082 = w6340 ;
  assign \po083 = w6435 ;
  assign \po084 = w6528 ;
  assign \po085 = w6621 ;
  assign \po086 = w6714 ;
  assign \po087 = w6795 ;
  assign \po088 = w6876 ;
  assign \po089 = w6956 ;
  assign \po090 = w7037 ;
  assign \po091 = w7117 ;
  assign \po092 = w7195 ;
  assign \po093 = w7271 ;
  assign \po094 = w7339 ;
  assign \po095 = w7409 ;
  assign \po096 = w7479 ;
  assign \po097 = w7546 ;
  assign \po098 = w7611 ;
  assign \po099 = w7670 ;
  assign \po100 = w7725 ;
  assign \po101 = w7782 ;
  assign \po102 = w7840 ;
  assign \po103 = w7896 ;
  assign \po104 = w7950 ;
  assign \po105 = w8005 ;
  assign \po106 = w8051 ;
  assign \po107 = w8098 ;
  assign \po108 = w8140 ;
  assign \po109 = w8183 ;
  assign \po110 = w8220 ;
  assign \po111 = w8263 ;
  assign \po112 = w8297 ;
  assign \po113 = w8329 ;
  assign \po114 = w8359 ;
  assign \po115 = w8387 ;
  assign \po116 = w8411 ;
  assign \po117 = w8447 ;
  assign \po118 = w8467 ;
  assign \po119 = w8489 ;
  assign \po120 = w8506 ;
  assign \po121 = w8522 ;
  assign \po122 = w8532 ;
  assign \po123 = w8547 ;
  assign \po124 = w8564 ;
  assign \po125 = w8582 ;
  assign \po126 = w8589 ;
  assign \po127 = w8591 ;
endmodule
