module ctrl( \pi0 , \pi1 , \pi2 , \pi3 , \pi4 , \pi5 , \pi6 , \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po24 , \po25 );
  input \pi0 , \pi1 , \pi2 , \pi3 , \pi4 , \pi5 , \pi6 ;
  output \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po23 , \po24 , \po25 ;
  wire zero , w8 , w9 , w10 , w11 , w12 , w13 , w14 , w15 , w16 , w17 , w18 , w19 , w20 , w21 , w22 , w23 , w24 , w25 , w26 , w27 , w28 , w29 , w30 , w31 , w32 , w33 , w34 , w35 , w36 , w37 , w38 , w39 , w40 , w41 , w42 , w43 , w44 , w45 , w46 , w47 , w48 , w49 , w50 , w51 , w52 , w53 , w54 , w55 , w56 , w57 , w58 , w59 , w60 , w61 , w62 , w63 , w64 , w65 , w66 , w67 , w68 , w69 , w70 , w71 , w72 , w73 , w74 , w75 , w76 , w77 , w78 , w79 , w80 , w81 , w82 , w83 , w84 , w85 , w86 , w87 , w88 , w89 , w90 , w91 , w92 , w93 , w94 , w95 , w96 , w97 , w98 , w99 , w100 , w101 , w102 , w103 , w104 , w105 , w106 , w107 , w108 , w109 , w110 , w111 , w112 , w113 , w114 , w115 , w116 , w117 , w118 , w119 , w120 , w121 , w122 ;
  assign zero = 0;
  assign w8 = \pi0 & \pi3 ;
  assign w9 = \pi4 & w8 ;
  assign w10 = ( \pi1 & \pi2 ) | ( \pi1 & \pi3 ) | ( \pi2 & \pi3 ) ;
  assign w11 = \pi3 ^ \pi4 ;
  assign w12 = ( w9 & w10 ) | ( w9 & ~w11 ) | ( w10 & ~w11 ) ;
  assign w13 = \pi2 | \pi4 ;
  assign w14 = ~\pi0 & \pi4 ;
  assign w15 = ( ~\pi3 & w13 ) | ( ~\pi3 & w14 ) | ( w13 & w14 ) ;
  assign w16 = \pi1 ^ \pi3 ;
  assign w17 = ( \pi2 & \pi4 ) | ( \pi2 & ~w16 ) | ( \pi4 & ~w16 ) ;
  assign w18 = w15 & ~w17 ;
  assign w19 = ( \pi1 & \pi3 ) | ( \pi1 & \pi4 ) | ( \pi3 & \pi4 ) ;
  assign w20 = ( \pi0 & \pi1 ) | ( \pi0 & \pi3 ) | ( \pi1 & \pi3 ) ;
  assign w21 = ( \pi2 & \pi4 ) | ( \pi2 & w20 ) | ( \pi4 & w20 ) ;
  assign w22 = w19 & ~w21 ;
  assign w23 = ( \pi0 & \pi1 ) | ( \pi0 & \pi4 ) | ( \pi1 & \pi4 ) ;
  assign w24 = \pi3 ^ w23 ;
  assign w25 = ( \pi1 & ~\pi2 ) | ( \pi1 & w24 ) | ( ~\pi2 & w24 ) ;
  assign w26 = ~\pi3 & \pi4 ;
  assign w27 = ( ~\pi1 & w25 ) | ( ~\pi1 & w26 ) | ( w25 & w26 ) ;
  assign w28 = \pi5 & \pi6 ;
  assign w29 = \pi4 | w28 ;
  assign w30 = ( \pi3 & w28 ) | ( \pi3 & ~w29 ) | ( w28 & ~w29 ) ;
  assign w31 = \pi0 & ~\pi4 ;
  assign w32 = \pi1 & \pi3 ;
  assign w33 = ( ~\pi0 & \pi4 ) | ( ~\pi0 & \pi6 ) | ( \pi4 & \pi6 ) ;
  assign w34 = \pi5 & w33 ;
  assign w35 = ( ~\pi4 & w32 ) | ( ~\pi4 & w34 ) | ( w32 & w34 ) ;
  assign w36 = ( \pi4 & w31 ) | ( \pi4 & w35 ) | ( w31 & w35 ) ;
  assign w37 = \pi0 & w26 ;
  assign w38 = \pi2 ^ w37 ;
  assign w39 = ( w36 & w37 ) | ( w36 & ~w38 ) | ( w37 & ~w38 ) ;
  assign w40 = ( \pi3 & ~\pi4 ) | ( \pi3 & \pi6 ) | ( ~\pi4 & \pi6 ) ;
  assign w41 = ( \pi1 & \pi2 ) | ( \pi1 & w40 ) | ( \pi2 & w40 ) ;
  assign w42 = ~\pi2 & \pi3 ;
  assign w43 = ( w26 & w41 ) | ( w26 & w42 ) | ( w41 & w42 ) ;
  assign w44 = \pi0 & \pi1 ;
  assign w45 = ( \pi2 & \pi3 ) | ( \pi2 & w44 ) | ( \pi3 & w44 ) ;
  assign w46 = \pi3 & w45 ;
  assign w47 = \pi4 ^ w45 ;
  assign w48 = \pi3 ^ w47 ;
  assign w49 = ( ~\pi2 & w46 ) | ( ~\pi2 & w48 ) | ( w46 & w48 ) ;
  assign w50 = ( ~\pi0 & \pi4 ) | ( ~\pi0 & w26 ) | ( \pi4 & w26 ) ;
  assign w51 = ( \pi1 & ~\pi3 ) | ( \pi1 & w50 ) | ( ~\pi3 & w50 ) ;
  assign w52 = ( \pi2 & \pi4 ) | ( \pi2 & w51 ) | ( \pi4 & w51 ) ;
  assign w53 = w50 ^ w52 ;
  assign w54 = ( \pi2 & ~\pi3 ) | ( \pi2 & \pi4 ) | ( ~\pi3 & \pi4 ) ;
  assign w55 = ( \pi1 & \pi3 ) | ( \pi1 & ~\pi4 ) | ( \pi3 & ~\pi4 ) ;
  assign w56 = ( \pi0 & \pi2 ) | ( \pi0 & ~w55 ) | ( \pi2 & ~w55 ) ;
  assign w57 = ( \pi1 & w55 ) | ( \pi1 & ~w56 ) | ( w55 & ~w56 ) ;
  assign w58 = w54 & w57 ;
  assign w59 = \pi0 | \pi4 ;
  assign w60 = ( ~\pi1 & \pi2 ) | ( ~\pi1 & \pi4 ) | ( \pi2 & \pi4 ) ;
  assign w61 = ( ~\pi0 & w59 ) | ( ~\pi0 & w60 ) | ( w59 & w60 ) ;
  assign w62 = ( \pi2 & ~\pi3 ) | ( \pi2 & w61 ) | ( ~\pi3 & w61 ) ;
  assign w63 = w60 ^ w62 ;
  assign w64 = ( \pi0 & \pi2 ) | ( \pi0 & ~\pi3 ) | ( \pi2 & ~\pi3 ) ;
  assign w65 = \pi4 & w64 ;
  assign w66 = ( ~\pi1 & \pi4 ) | ( ~\pi1 & w65 ) | ( \pi4 & w65 ) ;
  assign w67 = \pi3 ^ w66 ;
  assign w68 = ( ~\pi2 & w65 ) | ( ~\pi2 & w67 ) | ( w65 & w67 ) ;
  assign w69 = ( \pi0 & ~\pi1 ) | ( \pi0 & \pi2 ) | ( ~\pi1 & \pi2 ) ;
  assign w70 = \pi1 | w69 ;
  assign w71 = ( ~\pi3 & \pi4 ) | ( ~\pi3 & w70 ) | ( \pi4 & w70 ) ;
  assign w72 = \pi3 | w71 ;
  assign w73 = \pi2 ^ \pi3 ;
  assign w74 = \pi1 | \pi3 ;
  assign w75 = ( \pi4 & w73 ) | ( \pi4 & w74 ) | ( w73 & w74 ) ;
  assign w76 = \pi4 | w75 ;
  assign w77 = ( \pi0 & w75 ) | ( \pi0 & w76 ) | ( w75 & w76 ) ;
  assign w78 = ( ~\pi0 & \pi2 ) | ( ~\pi0 & \pi3 ) | ( \pi2 & \pi3 ) ;
  assign w79 = \pi2 & ~\pi4 ;
  assign w80 = ~w78 & w79 ;
  assign w81 = ( \pi0 & \pi2 ) | ( \pi0 & \pi3 ) | ( \pi2 & \pi3 ) ;
  assign w82 = w79 & ~w81 ;
  assign w83 = ( ~\pi0 & \pi1 ) | ( ~\pi0 & \pi2 ) | ( \pi1 & \pi2 ) ;
  assign w84 = ~\pi1 & w83 ;
  assign w85 = ( \pi3 & \pi4 ) | ( \pi3 & ~w84 ) | ( \pi4 & ~w84 ) ;
  assign w86 = \pi3 & ~w85 ;
  assign w87 = ( \pi0 & \pi1 ) | ( \pi0 & \pi2 ) | ( \pi1 & \pi2 ) ;
  assign w88 = ~\pi1 & w87 ;
  assign w89 = ( \pi3 & \pi4 ) | ( \pi3 & ~w88 ) | ( \pi4 & ~w88 ) ;
  assign w90 = \pi3 & ~w89 ;
  assign w91 = \pi1 & w69 ;
  assign w92 = ( \pi3 & \pi4 ) | ( \pi3 & ~w91 ) | ( \pi4 & ~w91 ) ;
  assign w93 = \pi3 & ~w92 ;
  assign w94 = ( \pi0 & \pi1 ) | ( \pi0 & ~\pi2 ) | ( \pi1 & ~\pi2 ) ;
  assign w95 = \pi1 & ~w94 ;
  assign w96 = ( \pi3 & \pi4 ) | ( \pi3 & ~w95 ) | ( \pi4 & ~w95 ) ;
  assign w97 = \pi3 & ~w96 ;
  assign w98 = ( \pi2 & \pi3 ) | ( \pi2 & ~\pi4 ) | ( \pi3 & ~\pi4 ) ;
  assign w99 = ~\pi3 & w98 ;
  assign w100 = ( \pi0 & \pi1 ) | ( \pi0 & ~\pi3 ) | ( \pi1 & ~\pi3 ) ;
  assign w101 = ~\pi5 & w100 ;
  assign w102 = ( \pi0 & \pi2 ) | ( \pi0 & ~w101 ) | ( \pi2 & ~w101 ) ;
  assign w103 = ( ~\pi4 & w100 ) | ( ~\pi4 & w102 ) | ( w100 & w102 ) ;
  assign w104 = \pi2 ^ w103 ;
  assign w105 = \pi3 & w104 ;
  assign w106 = ( \pi0 & \pi1 ) | ( \pi0 & ~\pi4 ) | ( \pi1 & ~\pi4 ) ;
  assign w107 = ( \pi4 & \pi5 ) | ( \pi4 & \pi6 ) | ( \pi5 & \pi6 ) ;
  assign w108 = ~\pi6 & w107 ;
  assign w109 = ( ~\pi1 & \pi3 ) | ( ~\pi1 & w108 ) | ( \pi3 & w108 ) ;
  assign w110 = w106 & w109 ;
  assign w111 = ~\pi2 & w110 ;
  assign w112 = w30 & w44 ;
  assign w113 = \pi2 ^ w112 ;
  assign w114 = ( \pi2 & ~\pi4 ) | ( \pi2 & w44 ) | ( ~\pi4 & w44 ) ;
  assign w115 = \pi3 & ~w114 ;
  assign w116 = ( w112 & w113 ) | ( w112 & w115 ) | ( w113 & w115 ) ;
  assign w117 = ( ~\pi0 & \pi1 ) | ( ~\pi0 & \pi4 ) | ( \pi1 & \pi4 ) ;
  assign w118 = \pi3 | w83 ;
  assign w119 = w117 & ~w118 ;
  assign w120 = ~\pi1 & w94 ;
  assign w121 = ( \pi3 & \pi4 ) | ( \pi3 & w120 ) | ( \pi4 & w120 ) ;
  assign w122 = ~\pi3 & w121 ;
  assign \po00 = w12 ;
  assign \po01 = w18 ;
  assign \po02 = w22 ;
  assign \po03 = w27 ;
  assign \po04 = w39 ;
  assign \po05 = w43 ;
  assign \po06 = w49 ;
  assign \po07 = w53 ;
  assign \po08 = w58 ;
  assign \po09 = w63 ;
  assign \po10 = w68 ;
  assign \po11 = ~w72 ;
  assign \po12 = w77 ;
  assign \po13 = w80 ;
  assign \po14 = w82 ;
  assign \po15 = w86 ;
  assign \po16 = w90 ;
  assign \po17 = w93 ;
  assign \po18 = w97 ;
  assign \po19 = w99 ;
  assign \po20 = w105 ;
  assign \po21 = w111 ;
  assign \po22 = w116 ;
  assign \po24 = w119 ;
  assign \po25 = w122 ;
endmodule
