module sin( \pi00 , \pi01 , \pi02 , \pi03 , \pi04 , \pi05 , \pi06 , \pi07 , \pi08 , \pi09 , \pi10 , \pi11 , \pi12 , \pi13 , \pi14 , \pi15 , \pi16 , \pi17 , \pi18 , \pi19 , \pi20 , \pi21 , \pi22 , \pi23 , \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po23 , \po24 );
  input \pi00 , \pi01 , \pi02 , \pi03 , \pi04 , \pi05 , \pi06 , \pi07 , \pi08 , \pi09 , \pi10 , \pi11 , \pi12 , \pi13 , \pi14 , \pi15 , \pi16 , \pi17 , \pi18 , \pi19 , \pi20 , \pi21 , \pi22 , \pi23 ;
  output \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po23 , \po24 ;
  wire zero , w25 , w26 , w27 , w28 , w29 , w30 , w31 , w32 , w33 , w34 , w35 , w36 , w37 , w38 , w39 , w40 , w41 , w42 , w43 , w44 , w45 , w46 , w47 , w48 , w49 , w50 , w51 , w52 , w53 , w54 , w55 , w56 , w57 , w58 , w59 , w60 , w61 , w62 , w63 , w64 , w65 , w66 , w67 , w68 , w69 , w70 , w71 , w72 , w73 , w74 , w75 , w76 , w77 , w78 , w79 , w80 , w81 , w82 , w83 , w84 , w85 , w86 , w87 , w88 , w89 , w90 , w91 , w92 , w93 , w94 , w95 , w96 , w97 , w98 , w99 , w100 , w101 , w102 , w103 , w104 , w105 , w106 , w107 , w108 , w109 , w110 , w111 , w112 , w113 , w114 , w115 , w116 , w117 , w118 , w119 , w120 , w121 , w122 , w123 , w124 , w125 , w126 , w127 , w128 , w129 , w130 , w131 , w132 , w133 , w134 , w135 , w136 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w146 , w147 , w148 , w149 , w150 , w151 , w152 , w153 , w154 , w155 , w156 , w157 , w158 , w159 , w160 , w161 , w162 , w163 , w164 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w174 , w175 , w176 , w177 , w178 , w179 , w180 , w181 , w182 , w183 , w184 , w185 , w186 , w187 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w203 , w204 , w205 , w206 , w207 , w208 , w209 , w210 , w211 , w212 , w213 , w214 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w224 , w225 , w226 , w227 , w228 , w229 , w230 , w231 , w232 , w233 , w234 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w250 , w251 , w252 , w253 , w254 , w255 , w256 , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 , w2495 , w2496 , w2497 , w2498 , w2499 , w2500 , w2501 , w2502 , w2503 , w2504 , w2505 , w2506 , w2507 , w2508 , w2509 , w2510 , w2511 , w2512 , w2513 , w2514 , w2515 , w2516 , w2517 , w2518 , w2519 , w2520 , w2521 , w2522 , w2523 , w2524 , w2525 , w2526 , w2527 , w2528 , w2529 , w2530 , w2531 , w2532 , w2533 , w2534 , w2535 , w2536 , w2537 , w2538 , w2539 , w2540 , w2541 , w2542 , w2543 , w2544 , w2545 , w2546 , w2547 , w2548 , w2549 , w2550 , w2551 , w2552 , w2553 , w2554 , w2555 , w2556 , w2557 , w2558 , w2559 , w2560 , w2561 , w2562 , w2563 , w2564 , w2565 , w2566 , w2567 , w2568 , w2569 , w2570 , w2571 , w2572 , w2573 , w2574 , w2575 , w2576 , w2577 , w2578 , w2579 , w2580 , w2581 , w2582 , w2583 , w2584 , w2585 , w2586 , w2587 , w2588 , w2589 , w2590 , w2591 , w2592 , w2593 , w2594 , w2595 , w2596 , w2597 , w2598 , w2599 , w2600 , w2601 , w2602 , w2603 , w2604 , w2605 , w2606 , w2607 , w2608 , w2609 , w2610 , w2611 , w2612 , w2613 , w2614 , w2615 , w2616 , w2617 , w2618 , w2619 , w2620 , w2621 , w2622 , w2623 , w2624 , w2625 , w2626 , w2627 , w2628 , w2629 , w2630 , w2631 , w2632 , w2633 , w2634 , w2635 , w2636 , w2637 , w2638 , w2639 , w2640 , w2641 , w2642 , w2643 , w2644 , w2645 , w2646 , w2647 , w2648 , w2649 , w2650 , w2651 , w2652 , w2653 , w2654 , w2655 , w2656 , w2657 , w2658 , w2659 , w2660 , w2661 , w2662 , w2663 , w2664 , w2665 , w2666 , w2667 , w2668 , w2669 , w2670 , w2671 , w2672 , w2673 , w2674 , w2675 , w2676 , w2677 , w2678 , w2679 , w2680 , w2681 , w2682 , w2683 , w2684 , w2685 , w2686 , w2687 , w2688 , w2689 , w2690 , w2691 , w2692 , w2693 , w2694 , w2695 , w2696 , w2697 , w2698 , w2699 , w2700 , w2701 , w2702 , w2703 , w2704 , w2705 , w2706 , w2707 , w2708 , w2709 , w2710 , w2711 , w2712 , w2713 , w2714 , w2715 , w2716 , w2717 , w2718 , w2719 , w2720 , w2721 , w2722 , w2723 , w2724 , w2725 , w2726 , w2727 , w2728 , w2729 , w2730 , w2731 , w2732 , w2733 , w2734 , w2735 , w2736 , w2737 , w2738 , w2739 , w2740 , w2741 , w2742 , w2743 , w2744 , w2745 , w2746 , w2747 , w2748 , w2749 , w2750 , w2751 , w2752 , w2753 , w2754 , w2755 , w2756 , w2757 , w2758 , w2759 , w2760 , w2761 , w2762 , w2763 , w2764 , w2765 , w2766 , w2767 , w2768 , w2769 , w2770 , w2771 , w2772 , w2773 , w2774 , w2775 , w2776 , w2777 , w2778 , w2779 , w2780 , w2781 , w2782 , w2783 , w2784 , w2785 , w2786 , w2787 , w2788 , w2789 , w2790 , w2791 , w2792 , w2793 , w2794 , w2795 , w2796 , w2797 , w2798 , w2799 , w2800 , w2801 , w2802 , w2803 , w2804 , w2805 , w2806 , w2807 , w2808 , w2809 , w2810 , w2811 , w2812 , w2813 , w2814 , w2815 , w2816 , w2817 , w2818 , w2819 , w2820 , w2821 , w2822 , w2823 , w2824 , w2825 , w2826 , w2827 , w2828 , w2829 , w2830 , w2831 , w2832 , w2833 , w2834 , w2835 , w2836 , w2837 , w2838 , w2839 , w2840 , w2841 , w2842 , w2843 , w2844 , w2845 , w2846 , w2847 , w2848 , w2849 , w2850 , w2851 , w2852 , w2853 , w2854 , w2855 , w2856 , w2857 , w2858 , w2859 , w2860 , w2861 , w2862 , w2863 , w2864 , w2865 , w2866 , w2867 , w2868 , w2869 , w2870 , w2871 , w2872 , w2873 , w2874 , w2875 , w2876 , w2877 , w2878 , w2879 , w2880 , w2881 , w2882 , w2883 , w2884 , w2885 , w2886 , w2887 , w2888 , w2889 , w2890 , w2891 , w2892 , w2893 , w2894 , w2895 , w2896 , w2897 , w2898 , w2899 , w2900 , w2901 , w2902 , w2903 , w2904 , w2905 , w2906 , w2907 , w2908 , w2909 , w2910 , w2911 , w2912 , w2913 , w2914 , w2915 , w2916 , w2917 , w2918 , w2919 , w2920 , w2921 , w2922 , w2923 , w2924 , w2925 , w2926 , w2927 , w2928 , w2929 , w2930 , w2931 , w2932 , w2933 , w2934 , w2935 , w2936 , w2937 , w2938 , w2939 , w2940 , w2941 , w2942 , w2943 , w2944 , w2945 , w2946 , w2947 , w2948 , w2949 , w2950 , w2951 , w2952 , w2953 , w2954 , w2955 , w2956 , w2957 , w2958 , w2959 , w2960 , w2961 , w2962 , w2963 , w2964 , w2965 , w2966 , w2967 , w2968 , w2969 , w2970 , w2971 , w2972 , w2973 , w2974 , w2975 , w2976 , w2977 , w2978 , w2979 , w2980 , w2981 , w2982 , w2983 , w2984 , w2985 , w2986 , w2987 , w2988 , w2989 , w2990 , w2991 , w2992 , w2993 , w2994 , w2995 , w2996 , w2997 , w2998 , w2999 , w3000 , w3001 , w3002 , w3003 , w3004 , w3005 , w3006 , w3007 , w3008 , w3009 , w3010 , w3011 , w3012 , w3013 , w3014 , w3015 , w3016 , w3017 , w3018 , w3019 , w3020 , w3021 , w3022 , w3023 , w3024 , w3025 , w3026 , w3027 , w3028 , w3029 , w3030 , w3031 , w3032 , w3033 , w3034 , w3035 , w3036 , w3037 , w3038 , w3039 , w3040 , w3041 , w3042 , w3043 , w3044 , w3045 , w3046 , w3047 , w3048 , w3049 , w3050 , w3051 , w3052 , w3053 , w3054 , w3055 , w3056 , w3057 , w3058 , w3059 , w3060 , w3061 , w3062 , w3063 , w3064 , w3065 , w3066 , w3067 , w3068 , w3069 , w3070 , w3071 , w3072 , w3073 , w3074 , w3075 , w3076 , w3077 , w3078 , w3079 , w3080 , w3081 , w3082 , w3083 , w3084 , w3085 , w3086 , w3087 , w3088 , w3089 , w3090 , w3091 , w3092 , w3093 , w3094 , w3095 , w3096 , w3097 , w3098 , w3099 , w3100 , w3101 , w3102 , w3103 , w3104 , w3105 , w3106 , w3107 , w3108 , w3109 , w3110 , w3111 , w3112 , w3113 , w3114 , w3115 , w3116 , w3117 , w3118 , w3119 , w3120 , w3121 , w3122 , w3123 , w3124 , w3125 , w3126 , w3127 , w3128 , w3129 , w3130 , w3131 , w3132 , w3133 , w3134 , w3135 , w3136 , w3137 , w3138 , w3139 , w3140 , w3141 , w3142 , w3143 , w3144 , w3145 , w3146 , w3147 , w3148 , w3149 , w3150 , w3151 , w3152 , w3153 , w3154 , w3155 , w3156 , w3157 , w3158 , w3159 , w3160 , w3161 , w3162 , w3163 , w3164 , w3165 , w3166 , w3167 , w3168 , w3169 , w3170 , w3171 , w3172 , w3173 , w3174 , w3175 , w3176 , w3177 , w3178 , w3179 , w3180 , w3181 , w3182 , w3183 , w3184 , w3185 , w3186 , w3187 , w3188 , w3189 , w3190 , w3191 , w3192 , w3193 , w3194 , w3195 , w3196 , w3197 , w3198 , w3199 , w3200 , w3201 , w3202 , w3203 , w3204 , w3205 , w3206 , w3207 , w3208 , w3209 , w3210 , w3211 , w3212 , w3213 , w3214 , w3215 , w3216 , w3217 , w3218 , w3219 , w3220 , w3221 , w3222 , w3223 , w3224 , w3225 , w3226 , w3227 , w3228 , w3229 , w3230 , w3231 , w3232 , w3233 , w3234 , w3235 , w3236 , w3237 , w3238 , w3239 , w3240 , w3241 , w3242 , w3243 , w3244 , w3245 , w3246 , w3247 , w3248 , w3249 , w3250 , w3251 , w3252 , w3253 , w3254 , w3255 , w3256 , w3257 , w3258 , w3259 , w3260 , w3261 , w3262 , w3263 , w3264 , w3265 , w3266 , w3267 , w3268 , w3269 , w3270 , w3271 , w3272 , w3273 , w3274 , w3275 , w3276 , w3277 , w3278 , w3279 , w3280 , w3281 , w3282 , w3283 , w3284 , w3285 , w3286 , w3287 , w3288 , w3289 , w3290 , w3291 , w3292 , w3293 , w3294 , w3295 , w3296 , w3297 , w3298 , w3299 , w3300 , w3301 , w3302 , w3303 , w3304 , w3305 , w3306 , w3307 , w3308 , w3309 , w3310 , w3311 , w3312 , w3313 , w3314 , w3315 , w3316 , w3317 , w3318 , w3319 , w3320 , w3321 , w3322 , w3323 , w3324 , w3325 , w3326 , w3327 , w3328 , w3329 , w3330 , w3331 , w3332 , w3333 , w3334 , w3335 , w3336 , w3337 , w3338 , w3339 , w3340 , w3341 , w3342 , w3343 , w3344 , w3345 , w3346 , w3347 , w3348 , w3349 , w3350 , w3351 , w3352 , w3353 , w3354 , w3355 , w3356 , w3357 , w3358 , w3359 , w3360 , w3361 , w3362 , w3363 , w3364 , w3365 , w3366 , w3367 , w3368 , w3369 , w3370 , w3371 , w3372 , w3373 , w3374 , w3375 , w3376 , w3377 , w3378 , w3379 , w3380 , w3381 , w3382 , w3383 , w3384 , w3385 , w3386 , w3387 , w3388 , w3389 , w3390 , w3391 , w3392 , w3393 , w3394 , w3395 , w3396 , w3397 , w3398 , w3399 , w3400 , w3401 , w3402 , w3403 , w3404 , w3405 , w3406 , w3407 , w3408 , w3409 , w3410 , w3411 , w3412 , w3413 , w3414 , w3415 , w3416 , w3417 , w3418 , w3419 , w3420 , w3421 , w3422 , w3423 , w3424 , w3425 , w3426 , w3427 , w3428 , w3429 , w3430 , w3431 , w3432 , w3433 , w3434 , w3435 , w3436 , w3437 , w3438 , w3439 , w3440 , w3441 , w3442 , w3443 , w3444 , w3445 , w3446 , w3447 , w3448 , w3449 , w3450 , w3451 , w3452 , w3453 , w3454 , w3455 , w3456 , w3457 , w3458 , w3459 , w3460 , w3461 , w3462 , w3463 , w3464 , w3465 , w3466 , w3467 , w3468 , w3469 , w3470 , w3471 , w3472 , w3473 , w3474 , w3475 , w3476 , w3477 , w3478 , w3479 , w3480 , w3481 , w3482 , w3483 , w3484 , w3485 , w3486 , w3487 , w3488 , w3489 , w3490 , w3491 , w3492 , w3493 , w3494 , w3495 , w3496 , w3497 , w3498 , w3499 , w3500 , w3501 , w3502 , w3503 , w3504 , w3505 , w3506 , w3507 , w3508 , w3509 , w3510 , w3511 , w3512 , w3513 , w3514 , w3515 , w3516 , w3517 , w3518 , w3519 , w3520 , w3521 , w3522 , w3523 , w3524 , w3525 , w3526 , w3527 , w3528 , w3529 , w3530 , w3531 , w3532 , w3533 , w3534 , w3535 , w3536 , w3537 , w3538 , w3539 , w3540 , w3541 , w3542 , w3543 , w3544 , w3545 , w3546 , w3547 , w3548 , w3549 , w3550 , w3551 , w3552 , w3553 , w3554 , w3555 , w3556 , w3557 , w3558 , w3559 , w3560 , w3561 , w3562 , w3563 , w3564 , w3565 , w3566 , w3567 , w3568 , w3569 , w3570 , w3571 , w3572 , w3573 , w3574 , w3575 , w3576 , w3577 , w3578 , w3579 , w3580 , w3581 , w3582 , w3583 , w3584 , w3585 , w3586 , w3587 , w3588 , w3589 , w3590 , w3591 , w3592 , w3593 , w3594 , w3595 , w3596 , w3597 , w3598 , w3599 , w3600 , w3601 , w3602 , w3603 , w3604 , w3605 , w3606 , w3607 , w3608 , w3609 , w3610 , w3611 , w3612 , w3613 , w3614 , w3615 , w3616 , w3617 , w3618 , w3619 , w3620 , w3621 , w3622 , w3623 , w3624 , w3625 , w3626 , w3627 , w3628 , w3629 , w3630 , w3631 , w3632 , w3633 , w3634 , w3635 , w3636 , w3637 , w3638 , w3639 , w3640 , w3641 , w3642 , w3643 , w3644 , w3645 , w3646 , w3647 , w3648 , w3649 , w3650 , w3651 , w3652 , w3653 , w3654 , w3655 , w3656 , w3657 , w3658 , w3659 , w3660 , w3661 , w3662 , w3663 , w3664 , w3665 , w3666 , w3667 , w3668 , w3669 , w3670 , w3671 , w3672 , w3673 , w3674 , w3675 , w3676 , w3677 , w3678 , w3679 , w3680 , w3681 , w3682 , w3683 , w3684 , w3685 , w3686 , w3687 , w3688 , w3689 , w3690 , w3691 , w3692 , w3693 , w3694 , w3695 , w3696 , w3697 , w3698 , w3699 , w3700 , w3701 , w3702 , w3703 , w3704 , w3705 , w3706 , w3707 , w3708 , w3709 , w3710 , w3711 , w3712 , w3713 , w3714 , w3715 , w3716 , w3717 , w3718 , w3719 , w3720 , w3721 , w3722 , w3723 , w3724 , w3725 , w3726 , w3727 , w3728 , w3729 , w3730 , w3731 , w3732 , w3733 , w3734 , w3735 , w3736 , w3737 , w3738 , w3739 , w3740 , w3741 , w3742 , w3743 , w3744 , w3745 , w3746 , w3747 , w3748 , w3749 , w3750 , w3751 , w3752 , w3753 , w3754 , w3755 , w3756 , w3757 , w3758 , w3759 , w3760 , w3761 , w3762 , w3763 , w3764 , w3765 , w3766 , w3767 , w3768 , w3769 , w3770 , w3771 , w3772 , w3773 , w3774 , w3775 , w3776 , w3777 , w3778 , w3779 , w3780 , w3781 , w3782 , w3783 , w3784 , w3785 , w3786 , w3787 , w3788 , w3789 , w3790 , w3791 , w3792 , w3793 , w3794 , w3795 , w3796 , w3797 , w3798 , w3799 , w3800 , w3801 , w3802 , w3803 , w3804 , w3805 , w3806 , w3807 , w3808 , w3809 , w3810 , w3811 , w3812 , w3813 , w3814 , w3815 , w3816 , w3817 , w3818 , w3819 , w3820 , w3821 , w3822 , w3823 , w3824 , w3825 , w3826 , w3827 , w3828 , w3829 , w3830 , w3831 , w3832 , w3833 , w3834 , w3835 , w3836 , w3837 , w3838 , w3839 , w3840 , w3841 , w3842 , w3843 , w3844 , w3845 , w3846 , w3847 , w3848 , w3849 ;
  assign zero = 0;
  assign w25 = ( \pi02 & \pi03 ) | ( \pi02 & ~\pi04 ) | ( \pi03 & ~\pi04 ) ;
  assign w26 = \pi00 | \pi01 ;
  assign w27 = ( ~\pi01 & \pi04 ) | ( ~\pi01 & \pi05 ) | ( \pi04 & \pi05 ) ;
  assign w28 = w26 | w27 ;
  assign w29 = w25 | w28 ;
  assign w30 = \pi08 | \pi09 ;
  assign w31 = \pi06 | w30 ;
  assign w32 = ( ~\pi06 & \pi07 ) | ( ~\pi06 & w29 ) | ( \pi07 & w29 ) ;
  assign w33 = w31 | w32 ;
  assign w34 = \pi10 | w33 ;
  assign w35 = \pi13 | \pi14 ;
  assign w36 = \pi11 | w35 ;
  assign w37 = ( ~\pi11 & \pi12 ) | ( ~\pi11 & w34 ) | ( \pi12 & w34 ) ;
  assign w38 = w36 | w37 ;
  assign w39 = \pi15 | w38 ;
  assign w40 = \pi18 | \pi19 ;
  assign w41 = \pi16 | w40 ;
  assign w42 = ( ~\pi16 & \pi17 ) | ( ~\pi16 & w39 ) | ( \pi17 & w39 ) ;
  assign w43 = w41 | w42 ;
  assign w44 = ( ~\pi20 & \pi21 ) | ( ~\pi20 & w43 ) | ( \pi21 & w43 ) ;
  assign w45 = \pi20 | w44 ;
  assign w46 = ~\pi22 & w38 ;
  assign w47 = \pi15 ^ w46 ;
  assign w48 = ~\pi22 & w43 ;
  assign w49 = ( \pi20 & \pi21 ) | ( \pi20 & ~w48 ) | ( \pi21 & ~w48 ) ;
  assign w50 = w48 ^ w49 ;
  assign w51 = w47 | w50 ;
  assign w52 = ( \pi16 & \pi17 ) | ( \pi16 & \pi18 ) | ( \pi17 & \pi18 ) ;
  assign w53 = ~\pi18 & w39 ;
  assign w54 = ( ~\pi16 & \pi19 ) | ( ~\pi16 & w53 ) | ( \pi19 & w53 ) ;
  assign w55 = ( \pi17 & ~\pi22 ) | ( \pi17 & w53 ) | ( ~\pi22 & w53 ) ;
  assign w56 = ( w52 & ~w54 ) | ( w52 & w55 ) | ( ~w54 & w55 ) ;
  assign w57 = w52 ^ w56 ;
  assign w58 = ~w51 & w57 ;
  assign w59 = \pi16 ^ \pi18 ;
  assign w60 = ( \pi19 & ~\pi22 ) | ( \pi19 & w59 ) | ( ~\pi22 & w59 ) ;
  assign w61 = ( \pi22 & ~w39 ) | ( \pi22 & w59 ) | ( ~w39 & w59 ) ;
  assign w62 = ( \pi17 & \pi18 ) | ( \pi17 & ~w61 ) | ( \pi18 & ~w61 ) ;
  assign w63 = \pi18 ^ w62 ;
  assign w64 = ( ~\pi19 & \pi22 ) | ( ~\pi19 & w63 ) | ( \pi22 & w63 ) ;
  assign w65 = w60 & w64 ;
  assign w66 = \pi21 & w43 ;
  assign w67 = ( \pi20 & w47 ) | ( \pi20 & w66 ) | ( w47 & w66 ) ;
  assign w68 = \pi21 ^ \pi22 ;
  assign w69 = ( \pi20 & w66 ) | ( \pi20 & w68 ) | ( w66 & w68 ) ;
  assign w70 = ~w67 & w69 ;
  assign w71 = w65 & w70 ;
  assign w72 = ~\pi22 & w39 ;
  assign w73 = ( ~\pi16 & \pi17 ) | ( ~\pi16 & \pi19 ) | ( \pi17 & \pi19 ) ;
  assign w74 = ( ~\pi17 & w72 ) | ( ~\pi17 & w73 ) | ( w72 & w73 ) ;
  assign w75 = ( ~\pi18 & w72 ) | ( ~\pi18 & w74 ) | ( w72 & w74 ) ;
  assign w76 = w72 ^ w75 ;
  assign w77 = w70 & w76 ;
  assign w78 = ( \pi20 & ~w47 ) | ( \pi20 & w66 ) | ( ~w47 & w66 ) ;
  assign w79 = w69 & ~w78 ;
  assign w80 = ( \pi19 & \pi22 ) | ( \pi19 & ~w59 ) | ( \pi22 & ~w59 ) ;
  assign w81 = ( \pi19 & \pi22 ) | ( \pi19 & w63 ) | ( \pi22 & w63 ) ;
  assign w82 = ~w80 & w81 ;
  assign w83 = w79 & w82 ;
  assign w84 = ( ~\pi20 & \pi21 ) | ( ~\pi20 & w48 ) | ( \pi21 & w48 ) ;
  assign w85 = w48 ^ w84 ;
  assign w86 = w47 & w85 ;
  assign w87 = \pi17 & w39 ;
  assign w88 = \pi16 ^ w87 ;
  assign w89 = ( \pi16 & ~\pi17 ) | ( \pi16 & w39 ) | ( ~\pi17 & w39 ) ;
  assign w90 = ( \pi18 & \pi19 ) | ( \pi18 & w89 ) | ( \pi19 & w89 ) ;
  assign w91 = ( \pi18 & ~\pi22 ) | ( \pi18 & w90 ) | ( ~\pi22 & w90 ) ;
  assign w92 = w90 ^ w91 ;
  assign w93 = w88 & w92 ;
  assign w94 = w86 & w93 ;
  assign w95 = ~\pi21 & w43 ;
  assign w96 = ( \pi20 & ~w47 ) | ( \pi20 & w95 ) | ( ~w47 & w95 ) ;
  assign w97 = ( \pi20 & ~w68 ) | ( \pi20 & w95 ) | ( ~w68 & w95 ) ;
  assign w98 = ~w96 & w97 ;
  assign w99 = ( \pi16 & \pi17 ) | ( \pi16 & ~\pi18 ) | ( \pi17 & ~\pi18 ) ;
  assign w100 = \pi18 & w39 ;
  assign w101 = ( ~\pi16 & \pi19 ) | ( ~\pi16 & w100 ) | ( \pi19 & w100 ) ;
  assign w102 = ( \pi17 & ~\pi22 ) | ( \pi17 & w100 ) | ( ~\pi22 & w100 ) ;
  assign w103 = ( w99 & ~w101 ) | ( w99 & w102 ) | ( ~w101 & w102 ) ;
  assign w104 = w99 ^ w103 ;
  assign w105 = w98 & w104 ;
  assign w106 = ( \pi20 & w47 ) | ( \pi20 & w95 ) | ( w47 & w95 ) ;
  assign w107 = w97 & ~w106 ;
  assign w108 = w57 & w107 ;
  assign w109 = w47 & ~w50 ;
  assign w110 = ( \pi16 & \pi19 ) | ( \pi16 & ~w53 ) | ( \pi19 & ~w53 ) ;
  assign w111 = ( w52 & w55 ) | ( w52 & w110 ) | ( w55 & w110 ) ;
  assign w112 = w52 ^ w111 ;
  assign w113 = w109 & w112 ;
  assign w114 = w57 & w86 ;
  assign w115 = w93 & w98 ;
  assign w116 = ~\pi17 & w39 ;
  assign w117 = \pi16 ^ w116 ;
  assign w118 = ( \pi16 & \pi17 ) | ( \pi16 & w39 ) | ( \pi17 & w39 ) ;
  assign w119 = ( \pi18 & \pi19 ) | ( \pi18 & ~w118 ) | ( \pi19 & ~w118 ) ;
  assign w120 = ( \pi18 & \pi22 ) | ( \pi18 & w119 ) | ( \pi22 & w119 ) ;
  assign w121 = w119 ^ w120 ;
  assign w122 = w117 & w121 ;
  assign w123 = w98 & w122 ;
  assign w124 = w107 & w122 ;
  assign w125 = w93 & w107 ;
  assign w126 = w107 & w112 ;
  assign w127 = w125 | w126 ;
  assign w128 = w57 & w70 ;
  assign w129 = ( ~\pi18 & \pi19 ) | ( ~\pi18 & w89 ) | ( \pi19 & w89 ) ;
  assign w130 = ( \pi18 & \pi22 ) | ( \pi18 & ~w129 ) | ( \pi22 & ~w129 ) ;
  assign w131 = w129 ^ w130 ;
  assign w132 = w88 & ~w131 ;
  assign w133 = w107 & w132 ;
  assign w134 = w57 & w79 ;
  assign w135 = ( \pi18 & \pi19 ) | ( \pi18 & ~w89 ) | ( \pi19 & ~w89 ) ;
  assign w136 = ( \pi18 & \pi22 ) | ( \pi18 & w135 ) | ( \pi22 & w135 ) ;
  assign w137 = w135 ^ w136 ;
  assign w138 = w88 & w137 ;
  assign w139 = w70 & w138 ;
  assign w140 = w134 | w139 ;
  assign w141 = w104 & w107 ;
  assign w142 = ( \pi18 & \pi19 ) | ( \pi18 & w118 ) | ( \pi19 & w118 ) ;
  assign w143 = ( \pi18 & ~\pi22 ) | ( \pi18 & w142 ) | ( ~\pi22 & w142 ) ;
  assign w144 = w142 ^ w143 ;
  assign w145 = w117 & w144 ;
  assign w146 = w107 & w145 ;
  assign w147 = w141 | w146 ;
  assign w148 = w109 & w122 ;
  assign w149 = w57 & w98 ;
  assign w150 = w148 | w149 ;
  assign w151 = ( ~w128 & w147 ) | ( ~w128 & w150 ) | ( w147 & w150 ) ;
  assign w152 = w127 | w140 ;
  assign w153 = ( w128 & w133 ) | ( w128 & ~w140 ) | ( w133 & ~w140 ) ;
  assign w154 = w152 | w153 ;
  assign w155 = w151 | w154 ;
  assign w156 = ( w114 & w115 ) | ( w114 & ~w123 ) | ( w115 & ~w123 ) ;
  assign w157 = w113 | w155 ;
  assign w158 = ( ~w113 & w123 ) | ( ~w113 & w124 ) | ( w123 & w124 ) ;
  assign w159 = w157 | w158 ;
  assign w160 = w156 | w159 ;
  assign w161 = w70 & w132 ;
  assign w162 = w86 & w145 ;
  assign w163 = ~w51 & w145 ;
  assign w164 = w79 & w93 ;
  assign w165 = ( \pi16 & ~\pi17 ) | ( \pi16 & \pi19 ) | ( ~\pi17 & \pi19 ) ;
  assign w166 = ( \pi17 & ~w72 ) | ( \pi17 & w165 ) | ( ~w72 & w165 ) ;
  assign w167 = ( \pi18 & ~w72 ) | ( \pi18 & w166 ) | ( ~w72 & w166 ) ;
  assign w168 = w72 ^ w167 ;
  assign w169 = w79 & ~w168 ;
  assign w170 = ~w47 & w85 ;
  assign w171 = w145 & w170 ;
  assign w172 = w65 & w98 ;
  assign w173 = w98 & w132 ;
  assign w174 = w82 & w170 ;
  assign w175 = w65 & w107 ;
  assign w176 = ( w172 & w173 ) | ( w172 & ~w174 ) | ( w173 & ~w174 ) ;
  assign w177 = w169 | w171 ;
  assign w178 = ( ~w171 & w174 ) | ( ~w171 & w175 ) | ( w174 & w175 ) ;
  assign w179 = w177 | w178 ;
  assign w180 = w176 | w179 ;
  assign w181 = ( ~w163 & w164 ) | ( ~w163 & w180 ) | ( w164 & w180 ) ;
  assign w182 = w163 | w181 ;
  assign w183 = w65 & w86 ;
  assign w184 = ( \pi18 & ~\pi19 ) | ( \pi18 & w118 ) | ( ~\pi19 & w118 ) ;
  assign w185 = ( \pi18 & ~\pi22 ) | ( \pi18 & w184 ) | ( ~\pi22 & w184 ) ;
  assign w186 = w184 ^ w185 ;
  assign w187 = w117 & w186 ;
  assign w188 = w107 & w187 ;
  assign w189 = w183 | w188 ;
  assign w190 = w70 & w145 ;
  assign w191 = w82 & w86 ;
  assign w192 = w86 & w104 ;
  assign w193 = ( \pi18 & ~\pi19 ) | ( \pi18 & w89 ) | ( ~\pi19 & w89 ) ;
  assign w194 = ( \pi18 & ~\pi22 ) | ( \pi18 & w193 ) | ( ~\pi22 & w193 ) ;
  assign w195 = w193 ^ w194 ;
  assign w196 = w88 & w195 ;
  assign w197 = w98 & w196 ;
  assign w198 = ( ~\pi18 & \pi19 ) | ( ~\pi18 & w118 ) | ( \pi19 & w118 ) ;
  assign w199 = ( \pi18 & \pi22 ) | ( \pi18 & ~w198 ) | ( \pi22 & ~w198 ) ;
  assign w200 = w198 ^ w199 ;
  assign w201 = w117 & ~w200 ;
  assign w202 = w107 & w201 ;
  assign w203 = w197 | w202 ;
  assign w204 = w191 | w203 ;
  assign w205 = ( w190 & ~w191 ) | ( w190 & w192 ) | ( ~w191 & w192 ) ;
  assign w206 = w204 | w205 ;
  assign w207 = w161 | w162 ;
  assign w208 = w189 | w207 ;
  assign w209 = ( w182 & ~w189 ) | ( w182 & w206 ) | ( ~w189 & w206 ) ;
  assign w210 = w208 | w209 ;
  assign w211 = ( \pi16 & \pi19 ) | ( \pi16 & ~w100 ) | ( \pi19 & ~w100 ) ;
  assign w212 = ( w99 & w102 ) | ( w99 & w211 ) | ( w102 & w211 ) ;
  assign w213 = w99 ^ w212 ;
  assign w214 = w79 & w213 ;
  assign w215 = w86 & w112 ;
  assign w216 = w107 & w138 ;
  assign w217 = ( w214 & ~w215 ) | ( w214 & w216 ) | ( ~w215 & w216 ) ;
  assign w218 = w215 | w217 ;
  assign w219 = w109 & w138 ;
  assign w220 = w79 & w201 ;
  assign w221 = ~w168 & w170 ;
  assign w222 = w98 & ~w168 ;
  assign w223 = w82 & w109 ;
  assign w224 = w70 & w104 ;
  assign w225 = w86 & w138 ;
  assign w226 = w65 & w170 ;
  assign w227 = w98 & w187 ;
  assign w228 = w98 & w112 ;
  assign w229 = w98 & w138 ;
  assign w230 = w107 & w196 ;
  assign w231 = w93 & w109 ;
  assign w232 = w79 & w104 ;
  assign w233 = w86 & w132 ;
  assign w234 = w57 & w170 ;
  assign w235 = w98 & w145 ;
  assign w236 = w76 & w98 ;
  assign w237 = ( w233 & w234 ) | ( w233 & ~w235 ) | ( w234 & ~w235 ) ;
  assign w238 = w231 | w232 ;
  assign w239 = ( ~w232 & w235 ) | ( ~w232 & w236 ) | ( w235 & w236 ) ;
  assign w240 = w238 | w239 ;
  assign w241 = w237 | w240 ;
  assign w242 = w79 & w187 ;
  assign w243 = w57 & w109 ;
  assign w244 = w109 & w187 ;
  assign w245 = w109 & w213 ;
  assign w246 = ( w242 & w243 ) | ( w242 & ~w244 ) | ( w243 & ~w244 ) ;
  assign w247 = w230 | w241 ;
  assign w248 = ( ~w230 & w244 ) | ( ~w230 & w245 ) | ( w244 & w245 ) ;
  assign w249 = w247 | w248 ;
  assign w250 = w246 | w249 ;
  assign w251 = ( w226 & w227 ) | ( w226 & ~w228 ) | ( w227 & ~w228 ) ;
  assign w252 = w225 | w250 ;
  assign w253 = ( ~w225 & w228 ) | ( ~w225 & w229 ) | ( w228 & w229 ) ;
  assign w254 = w252 | w253 ;
  assign w255 = w251 | w254 ;
  assign w256 = ( ~w223 & w224 ) | ( ~w223 & w255 ) | ( w224 & w255 ) ;
  assign w257 = w223 | w256 ;
  assign w258 = w221 | w222 ;
  assign w259 = w219 | w258 ;
  assign w260 = ( ~w219 & w220 ) | ( ~w219 & w257 ) | ( w220 & w257 ) ;
  assign w261 = w259 | w260 ;
  assign w262 = w170 & w196 ;
  assign w263 = w86 & w201 ;
  assign w264 = w262 | w263 ;
  assign w265 = w76 & w170 ;
  assign w266 = ~w51 & w196 ;
  assign w267 = w265 | w266 ;
  assign w268 = w218 | w267 ;
  assign w269 = ( ~w218 & w261 ) | ( ~w218 & w264 ) | ( w261 & w264 ) ;
  assign w270 = w268 | w269 ;
  assign w271 = ( w94 & ~w105 ) | ( w94 & w210 ) | ( ~w105 & w210 ) ;
  assign w272 = w160 | w270 ;
  assign w273 = ( w105 & w108 ) | ( w105 & ~w160 ) | ( w108 & ~w160 ) ;
  assign w274 = w272 | w273 ;
  assign w275 = w271 | w274 ;
  assign w276 = w77 | w83 ;
  assign w277 = w58 | w276 ;
  assign w278 = ( ~w58 & w71 ) | ( ~w58 & w275 ) | ( w71 & w275 ) ;
  assign w279 = w277 | w278 ;
  assign w280 = ( \pi01 & \pi02 ) | ( \pi01 & ~\pi03 ) | ( \pi02 & ~\pi03 ) ;
  assign w281 = \pi04 & ~\pi22 ;
  assign w282 = ( ~\pi22 & w280 ) | ( ~\pi22 & w281 ) | ( w280 & w281 ) ;
  assign w283 = ( \pi00 & ~\pi03 ) | ( \pi00 & w282 ) | ( ~\pi03 & w282 ) ;
  assign w284 = ( \pi03 & ~\pi22 ) | ( \pi03 & w283 ) | ( ~\pi22 & w283 ) ;
  assign w285 = \pi05 ^ w284 ;
  assign w286 = \pi00 & ~\pi22 ;
  assign w287 = \pi01 | \pi02 ;
  assign w288 = ( ~\pi00 & \pi03 ) | ( ~\pi00 & w287 ) | ( \pi03 & w287 ) ;
  assign w289 = ( ~\pi22 & w286 ) | ( ~\pi22 & w288 ) | ( w286 & w288 ) ;
  assign w290 = \pi04 ^ w289 ;
  assign w291 = \pi00 & ~\pi01 ;
  assign w292 = ( \pi01 & ~\pi02 ) | ( \pi01 & w291 ) | ( ~\pi02 & w291 ) ;
  assign w293 = ( \pi02 & ~\pi22 ) | ( \pi02 & w292 ) | ( ~\pi22 & w292 ) ;
  assign w294 = \pi03 ^ w293 ;
  assign w295 = ~\pi00 & \pi01 ;
  assign w296 = ( \pi00 & ~\pi22 ) | ( \pi00 & w295 ) | ( ~\pi22 & w295 ) ;
  assign w297 = \pi02 ^ w296 ;
  assign w298 = w294 ^ w297 ;
  assign w299 = w285 ^ w290 ;
  assign w300 = w298 & ~w299 ;
  assign w301 = w109 & w145 ;
  assign w302 = w65 & w79 ;
  assign w303 = w76 & w79 ;
  assign w304 = w93 & w170 ;
  assign w305 = w86 & w213 ;
  assign w306 = w219 | w305 ;
  assign w307 = w79 & w112 ;
  assign w308 = ( w123 & w174 ) | ( w123 & ~w175 ) | ( w174 & ~w175 ) ;
  assign w309 = w71 | w306 ;
  assign w310 = ( ~w71 & w175 ) | ( ~w71 & w307 ) | ( w175 & w307 ) ;
  assign w311 = w309 | w310 ;
  assign w312 = w308 | w311 ;
  assign w313 = ( w301 & w302 ) | ( w301 & ~w303 ) | ( w302 & ~w303 ) ;
  assign w314 = w191 | w312 ;
  assign w315 = ( ~w191 & w303 ) | ( ~w191 & w304 ) | ( w303 & w304 ) ;
  assign w316 = w314 | w315 ;
  assign w317 = w313 | w316 ;
  assign w318 = w170 & w201 ;
  assign w319 = w86 & w122 ;
  assign w320 = w229 | w319 ;
  assign w321 = w70 & w187 ;
  assign w322 = w98 & w213 ;
  assign w323 = ( w108 & ~w215 ) | ( w108 & w322 ) | ( ~w215 & w322 ) ;
  assign w324 = w215 | w323 ;
  assign w325 = ( w77 & w220 ) | ( w77 & ~w318 ) | ( w220 & ~w318 ) ;
  assign w326 = w320 | w324 ;
  assign w327 = ( w318 & w321 ) | ( w318 & ~w324 ) | ( w321 & ~w324 ) ;
  assign w328 = w326 | w327 ;
  assign w329 = w325 | w328 ;
  assign w330 = w51 | w168 ;
  assign w331 = ~w94 & w330 ;
  assign w332 = ~w51 & w138 ;
  assign w333 = w122 & w170 ;
  assign w334 = w107 & w213 ;
  assign w335 = w138 & w170 ;
  assign w336 = ( w332 & w333 ) | ( w332 & ~w334 ) | ( w333 & ~w334 ) ;
  assign w337 = w163 | w263 ;
  assign w338 = ( ~w263 & w334 ) | ( ~w263 & w335 ) | ( w334 & w335 ) ;
  assign w339 = w337 | w338 ;
  assign w340 = w336 | w339 ;
  assign w341 = w70 & w196 ;
  assign w342 = w76 & w86 ;
  assign w343 = w76 & w107 ;
  assign w344 = w342 | w343 ;
  assign w345 = w188 | w344 ;
  assign w346 = ( w172 & ~w188 ) | ( w172 & w341 ) | ( ~w188 & w341 ) ;
  assign w347 = w345 | w346 ;
  assign w348 = w65 & w109 ;
  assign w349 = w170 & w187 ;
  assign w350 = w348 | w349 ;
  assign w351 = w109 & ~w168 ;
  assign w352 = w70 & w201 ;
  assign w353 = w112 & w170 ;
  assign w354 = w104 & w170 ;
  assign w355 = ~w51 & w76 ;
  assign w356 = w234 | w355 ;
  assign w357 = w224 | w356 ;
  assign w358 = ( w192 & ~w224 ) | ( w192 & w225 ) | ( ~w224 & w225 ) ;
  assign w359 = w357 | w358 ;
  assign w360 = w70 & ~w168 ;
  assign w361 = w70 & w122 ;
  assign w362 = w70 & w213 ;
  assign w363 = w70 & w82 ;
  assign w364 = w86 & w187 ;
  assign w365 = w79 & w138 ;
  assign w366 = ( w362 & w363 ) | ( w362 & ~w364 ) | ( w363 & ~w364 ) ;
  assign w367 = w360 | w361 ;
  assign w368 = ( ~w361 & w364 ) | ( ~w361 & w365 ) | ( w364 & w365 ) ;
  assign w369 = w367 | w368 ;
  assign w370 = w366 | w369 ;
  assign w371 = ~w51 & w201 ;
  assign w372 = ~w51 & w104 ;
  assign w373 = w105 | w372 ;
  assign w374 = w170 & w213 ;
  assign w375 = w58 | w223 ;
  assign w376 = ( ~w371 & w373 ) | ( ~w371 & w375 ) | ( w373 & w375 ) ;
  assign w377 = w359 | w370 ;
  assign w378 = ( ~w370 & w371 ) | ( ~w370 & w374 ) | ( w371 & w374 ) ;
  assign w379 = w377 | w378 ;
  assign w380 = w376 | w379 ;
  assign w381 = w171 | w231 ;
  assign w382 = w114 | w381 ;
  assign w383 = ( ~w114 & w134 ) | ( ~w114 & w380 ) | ( w134 & w380 ) ;
  assign w384 = w382 | w383 ;
  assign w385 = ( ~w150 & w354 ) | ( ~w150 & w384 ) | ( w354 & w384 ) ;
  assign w386 = w150 | w385 ;
  assign w387 = ( w141 & w351 ) | ( w141 & ~w352 ) | ( w351 & ~w352 ) ;
  assign w388 = w267 | w386 ;
  assign w389 = ( ~w267 & w352 ) | ( ~w267 & w353 ) | ( w352 & w353 ) ;
  assign w390 = w388 | w389 ;
  assign w391 = w387 | w390 ;
  assign w392 = ( w331 & ~w340 ) | ( w331 & w347 ) | ( ~w340 & w347 ) ;
  assign w393 = w329 | w391 ;
  assign w394 = ( ~w329 & w347 ) | ( ~w329 & w350 ) | ( w347 & w350 ) ;
  assign w395 = w393 | w394 ;
  assign w396 = w392 & ~w395 ;
  assign w397 = w216 | w317 ;
  assign w398 = ( ~w115 & w317 ) | ( ~w115 & w396 ) | ( w317 & w396 ) ;
  assign w399 = ~w397 & w398 ;
  assign w400 = w98 & w201 ;
  assign w401 = w215 | w333 ;
  assign w402 = ( w171 & ~w216 ) | ( w171 & w401 ) | ( ~w216 & w401 ) ;
  assign w403 = w127 | w320 ;
  assign w404 = ( w216 & ~w320 ) | ( w216 & w343 ) | ( ~w320 & w343 ) ;
  assign w405 = w403 | w404 ;
  assign w406 = w402 | w405 ;
  assign w407 = w236 | w354 ;
  assign w408 = w162 | w407 ;
  assign w409 = ( ~w162 & w192 ) | ( ~w162 & w406 ) | ( w192 & w406 ) ;
  assign w410 = w408 | w409 ;
  assign w411 = w82 & w98 ;
  assign w412 = w82 & w107 ;
  assign w413 = w228 | w412 ;
  assign w414 = ( w124 & ~w228 ) | ( w124 & w304 ) | ( ~w228 & w304 ) ;
  assign w415 = w413 | w414 ;
  assign w416 = ( w123 & w265 ) | ( w123 & ~w342 ) | ( w265 & ~w342 ) ;
  assign w417 = w94 | w415 ;
  assign w418 = ( ~w94 & w342 ) | ( ~w94 & w411 ) | ( w342 & w411 ) ;
  assign w419 = w417 | w418 ;
  assign w420 = w416 | w419 ;
  assign w421 = w107 & ~w168 ;
  assign w422 = w132 & w170 ;
  assign w423 = w227 | w233 ;
  assign w424 = w189 | w423 ;
  assign w425 = ( w105 & w147 ) | ( w105 & ~w189 ) | ( w147 & ~w189 ) ;
  assign w426 = w424 | w425 ;
  assign w427 = ( ~w226 & w422 ) | ( ~w226 & w426 ) | ( w422 & w426 ) ;
  assign w428 = w226 | w427 ;
  assign w429 = ( w133 & w230 ) | ( w133 & ~w263 ) | ( w230 & ~w263 ) ;
  assign w430 = w420 | w428 ;
  assign w431 = ( w263 & ~w420 ) | ( w263 & w421 ) | ( ~w420 & w421 ) ;
  assign w432 = w430 | w431 ;
  assign w433 = w429 | w432 ;
  assign w434 = w173 | w222 ;
  assign w435 = w108 | w434 ;
  assign w436 = ( ~w108 & w115 ) | ( ~w108 & w433 ) | ( w115 & w433 ) ;
  assign w437 = w435 | w436 ;
  assign w438 = w149 | w197 ;
  assign w439 = ( w175 & w234 ) | ( w175 & ~w235 ) | ( w234 & ~w235 ) ;
  assign w440 = w114 | w172 ;
  assign w441 = ( ~w172 & w235 ) | ( ~w172 & w318 ) | ( w235 & w318 ) ;
  assign w442 = w440 | w441 ;
  assign w443 = w439 | w442 ;
  assign w444 = ( ~w202 & w438 ) | ( ~w202 & w443 ) | ( w438 & w443 ) ;
  assign w445 = w410 | w437 ;
  assign w446 = ( w202 & w334 ) | ( w202 & ~w410 ) | ( w334 & ~w410 ) ;
  assign w447 = w445 | w446 ;
  assign w448 = w444 | w447 ;
  assign w449 = ( ~w322 & w400 ) | ( ~w322 & w448 ) | ( w400 & w448 ) ;
  assign w450 = w322 | w449 ;
  assign w451 = ~w51 & w93 ;
  assign w452 = w86 & ~w168 ;
  assign w453 = w79 & w145 ;
  assign w454 = w190 | w453 ;
  assign w455 = w79 & w132 ;
  assign w456 = ( w161 & ~w302 ) | ( w161 & w455 ) | ( ~w302 & w455 ) ;
  assign w457 = w302 | w456 ;
  assign w458 = ( w134 & w454 ) | ( w134 & ~w457 ) | ( w454 & ~w457 ) ;
  assign w459 = w457 | w458 ;
  assign w460 = w262 | w349 ;
  assign w461 = w220 | w460 ;
  assign w462 = ( w128 & ~w220 ) | ( w128 & w232 ) | ( ~w220 & w232 ) ;
  assign w463 = w461 | w462 ;
  assign w464 = w86 & w196 ;
  assign w465 = ( w353 & w364 ) | ( w353 & ~w374 ) | ( w364 & ~w374 ) ;
  assign w466 = w305 | w352 ;
  assign w467 = ( ~w352 & w374 ) | ( ~w352 & w464 ) | ( w374 & w464 ) ;
  assign w468 = w466 | w467 ;
  assign w469 = w465 | w468 ;
  assign w470 = ( w71 & ~w221 ) | ( w71 & w469 ) | ( ~w221 & w469 ) ;
  assign w471 = w459 | w463 ;
  assign w472 = ( w221 & w452 ) | ( w221 & ~w463 ) | ( w452 & ~w463 ) ;
  assign w473 = w471 | w472 ;
  assign w474 = w470 | w473 ;
  assign w475 = w76 & w109 ;
  assign w476 = w104 & w109 ;
  assign w477 = ~w51 & w65 ;
  assign w478 = w109 & w201 ;
  assign w479 = ~w51 & w132 ;
  assign w480 = w174 | w335 ;
  assign w481 = w243 | w360 ;
  assign w482 = w191 | w225 ;
  assign w483 = w169 | w482 ;
  assign w484 = w109 & w132 ;
  assign w485 = ( w58 & ~w348 ) | ( w58 & w481 ) | ( ~w348 & w481 ) ;
  assign w486 = w480 | w483 ;
  assign w487 = ( w348 & ~w480 ) | ( w348 & w484 ) | ( ~w480 & w484 ) ;
  assign w488 = w486 | w487 ;
  assign w489 = w485 | w488 ;
  assign w490 = w371 | w479 ;
  assign w491 = ( ~w371 & w478 ) | ( ~w371 & w489 ) | ( w478 & w489 ) ;
  assign w492 = w490 | w491 ;
  assign w493 = w476 | w477 ;
  assign w494 = w163 | w493 ;
  assign w495 = ( ~w163 & w301 ) | ( ~w163 & w492 ) | ( w301 & w492 ) ;
  assign w496 = w494 | w495 ;
  assign w497 = ( w231 & w372 ) | ( w231 & ~w451 ) | ( w372 & ~w451 ) ;
  assign w498 = w474 | w496 ;
  assign w499 = ( w451 & ~w474 ) | ( w451 & w475 ) | ( ~w474 & w475 ) ;
  assign w500 = w498 | w499 ;
  assign w501 = w497 | w500 ;
  assign w502 = w79 & w196 ;
  assign w503 = w362 | w502 ;
  assign w504 = w321 | w503 ;
  assign w505 = ( w83 & ~w321 ) | ( w83 & w341 ) | ( ~w321 & w341 ) ;
  assign w506 = w504 | w505 ;
  assign w507 = w214 | w363 ;
  assign w508 = ( ~w214 & w242 ) | ( ~w214 & w506 ) | ( w242 & w506 ) ;
  assign w509 = w507 | w508 ;
  assign w510 = w70 & w93 ;
  assign w511 = w79 & w122 ;
  assign w512 = w224 | w511 ;
  assign w513 = w70 & w112 ;
  assign w514 = w365 | w513 ;
  assign w515 = w307 | w514 ;
  assign w516 = ( ~w307 & w361 ) | ( ~w307 & w512 ) | ( w361 & w512 ) ;
  assign w517 = w515 | w516 ;
  assign w518 = w303 | w510 ;
  assign w519 = w77 | w518 ;
  assign w520 = ( ~w77 & w164 ) | ( ~w77 & w517 ) | ( w164 & w517 ) ;
  assign w521 = w519 | w520 ;
  assign w522 = w482 | w521 ;
  assign w523 = ( w474 & w480 ) | ( w474 & ~w521 ) | ( w480 & ~w521 ) ;
  assign w524 = w522 | w523 ;
  assign w525 = ( w139 & ~w509 ) | ( w139 & w524 ) | ( ~w509 & w524 ) ;
  assign w526 = w509 | w525 ;
  assign w527 = w501 & w526 ;
  assign w528 = ~\pi22 & w34 ;
  assign w529 = \pi11 | \pi12 ;
  assign w530 = ( \pi13 & ~w34 ) | ( \pi13 & w529 ) | ( ~w34 & w529 ) ;
  assign w531 = ( ~\pi22 & w528 ) | ( ~\pi22 & w530 ) | ( w528 & w530 ) ;
  assign w532 = \pi14 ^ w531 ;
  assign w533 = ~\pi11 & w34 ;
  assign w534 = ( \pi11 & ~\pi12 ) | ( \pi11 & w533 ) | ( ~\pi12 & w533 ) ;
  assign w535 = ( \pi12 & ~\pi22 ) | ( \pi12 & w534 ) | ( ~\pi22 & w534 ) ;
  assign w536 = \pi13 ^ w535 ;
  assign w537 = w501 ^ w526 ;
  assign w538 = ( ~w450 & w501 ) | ( ~w450 & w526 ) | ( w501 & w526 ) ;
  assign w539 = ~w450 & w538 ;
  assign w540 = w450 & ~w527 ;
  assign w541 = ( w450 & w526 ) | ( w450 & ~w532 ) | ( w526 & ~w532 ) ;
  assign w542 = ( w450 & w501 ) | ( w450 & w541 ) | ( w501 & w541 ) ;
  assign w543 = w527 ^ w542 ;
  assign w544 = ~w51 & w122 ;
  assign w545 = ~w51 & w213 ;
  assign w546 = ~w51 & w112 ;
  assign w547 = w371 | w546 ;
  assign w548 = w229 | w547 ;
  assign w549 = ( w216 & ~w229 ) | ( w216 & w245 ) | ( ~w229 & w245 ) ;
  assign w550 = w548 | w549 ;
  assign w551 = ( w233 & ~w301 ) | ( w233 & w422 ) | ( ~w301 & w422 ) ;
  assign w552 = w301 | w551 ;
  assign w553 = ( w242 & ~w244 ) | ( w242 & w478 ) | ( ~w244 & w478 ) ;
  assign w554 = w244 | w553 ;
  assign w555 = w235 | w400 ;
  assign w556 = w554 | w555 ;
  assign w557 = ( w105 & w552 ) | ( w105 & ~w554 ) | ( w552 & ~w554 ) ;
  assign w558 = w556 | w557 ;
  assign w559 = ( w108 & ~w353 ) | ( w108 & w550 ) | ( ~w353 & w550 ) ;
  assign w560 = w182 | w558 ;
  assign w561 = ( w353 & w545 ) | ( w353 & ~w558 ) | ( w545 & ~w558 ) ;
  assign w562 = w560 | w561 ;
  assign w563 = w559 | w562 ;
  assign w564 = ( w220 & w228 ) | ( w220 & ~w343 ) | ( w228 & ~w343 ) ;
  assign w565 = w162 | w191 ;
  assign w566 = ( ~w191 & w343 ) | ( ~w191 & w364 ) | ( w343 & w364 ) ;
  assign w567 = w565 | w566 ;
  assign w568 = w564 | w567 ;
  assign w569 = w477 | w568 ;
  assign w570 = w476 | w510 ;
  assign w571 = w83 | w570 ;
  assign w572 = ( w77 & ~w83 ) | ( w77 & w202 ) | ( ~w83 & w202 ) ;
  assign w573 = w571 | w572 ;
  assign w574 = w335 | w455 ;
  assign w575 = ( w226 & ~w335 ) | ( w226 & w349 ) | ( ~w335 & w349 ) ;
  assign w576 = w574 | w575 ;
  assign w577 = ( w303 & ~w352 ) | ( w303 & w360 ) | ( ~w352 & w360 ) ;
  assign w578 = w352 | w577 ;
  assign w579 = ( w160 & ~w236 ) | ( w160 & w363 ) | ( ~w236 & w363 ) ;
  assign w580 = w236 | w579 ;
  assign w581 = ~w51 & w187 ;
  assign w582 = ( ~w183 & w576 ) | ( ~w183 & w578 ) | ( w576 & w578 ) ;
  assign w583 = w573 | w580 ;
  assign w584 = ( w183 & ~w573 ) | ( w183 & w581 ) | ( ~w573 & w581 ) ;
  assign w585 = w583 | w584 ;
  assign w586 = w582 | w585 ;
  assign w587 = w359 | w544 ;
  assign w588 = w563 | w587 ;
  assign w589 = ( ~w563 & w569 ) | ( ~w563 & w586 ) | ( w569 & w586 ) ;
  assign w590 = w588 | w589 ;
  assign w591 = ~w51 & w82 ;
  assign w592 = ( w115 & w169 ) | ( w115 & ~w228 ) | ( w169 & ~w228 ) ;
  assign w593 = w127 | w375 ;
  assign w594 = ( w228 & w303 ) | ( w228 & ~w375 ) | ( w303 & ~w375 ) ;
  assign w595 = w593 | w594 ;
  assign w596 = w592 | w595 ;
  assign w597 = ( ~w513 & w546 ) | ( ~w513 & w596 ) | ( w546 & w596 ) ;
  assign w598 = w513 | w597 ;
  assign w599 = ( w77 & ~w230 ) | ( w77 & w343 ) | ( ~w230 & w343 ) ;
  assign w600 = w230 | w599 ;
  assign w601 = w322 | w411 ;
  assign w602 = ( w148 & w235 ) | ( w148 & ~w335 ) | ( w235 & ~w335 ) ;
  assign w603 = w481 | w601 ;
  assign w604 = ( w335 & w353 ) | ( w335 & ~w601 ) | ( w353 & ~w601 ) ;
  assign w605 = w603 | w604 ;
  assign w606 = w602 | w605 ;
  assign w607 = ( ~w188 & w438 ) | ( ~w188 & w512 ) | ( w438 & w512 ) ;
  assign w608 = w147 | w606 ;
  assign w609 = ( ~w147 & w188 ) | ( ~w147 & w412 ) | ( w188 & w412 ) ;
  assign w610 = w608 | w609 ;
  assign w611 = w607 | w610 ;
  assign w612 = w332 | w361 ;
  assign w613 = w108 | w612 ;
  assign w614 = ( ~w108 & w225 ) | ( ~w108 & w611 ) | ( w225 & w611 ) ;
  assign w615 = w613 | w614 ;
  assign w616 = ( ~w355 & w400 ) | ( ~w355 & w615 ) | ( w400 & w615 ) ;
  assign w617 = w355 | w616 ;
  assign w618 = w216 | w222 ;
  assign w619 = w123 | w618 ;
  assign w620 = ( ~w123 & w164 ) | ( ~w123 & w617 ) | ( w164 & w617 ) ;
  assign w621 = w619 | w620 ;
  assign w622 = w598 | w600 ;
  assign w623 = ( w350 & ~w598 ) | ( w350 & w621 ) | ( ~w598 & w621 ) ;
  assign w624 = w622 | w623 ;
  assign w625 = w452 | w591 ;
  assign w626 = w191 | w625 ;
  assign w627 = ( ~w191 & w219 ) | ( ~w191 & w624 ) | ( w219 & w624 ) ;
  assign w628 = w626 | w627 ;
  assign w629 = w318 | w421 ;
  assign w630 = ( w173 & w202 ) | ( w173 & ~w305 ) | ( w202 & ~w305 ) ;
  assign w631 = w172 | w629 ;
  assign w632 = ( ~w172 & w305 ) | ( ~w172 & w510 ) | ( w305 & w510 ) ;
  assign w633 = w631 | w632 ;
  assign w634 = w630 | w633 ;
  assign w635 = w307 | w634 ;
  assign w636 = w221 | w479 ;
  assign w637 = w334 | w374 ;
  assign w638 = w105 | w637 ;
  assign w639 = ( ~w105 & w133 ) | ( ~w105 & w264 ) | ( w133 & w264 ) ;
  assign w640 = w638 | w639 ;
  assign w641 = w113 | w478 ;
  assign w642 = ( ~w113 & w229 ) | ( ~w113 & w640 ) | ( w229 & w640 ) ;
  assign w643 = w641 | w642 ;
  assign w644 = ( ~w227 & w464 ) | ( ~w227 & w643 ) | ( w464 & w643 ) ;
  assign w645 = w227 | w644 ;
  assign w646 = ( w174 & w175 ) | ( w174 & ~w236 ) | ( w175 & ~w236 ) ;
  assign w647 = w124 | w645 ;
  assign w648 = ( ~w124 & w236 ) | ( ~w124 & w484 ) | ( w236 & w484 ) ;
  assign w649 = w647 | w648 ;
  assign w650 = w646 | w649 ;
  assign w651 = ( ~w635 & w636 ) | ( ~w635 & w650 ) | ( w636 & w650 ) ;
  assign w652 = w635 | w651 ;
  assign w653 = ( w364 & w365 ) | ( w364 & ~w371 ) | ( w365 & ~w371 ) ;
  assign w654 = w628 | w652 ;
  assign w655 = ( w371 & w544 ) | ( w371 & ~w652 ) | ( w544 & ~w652 ) ;
  assign w656 = w654 | w655 ;
  assign w657 = w653 | w656 ;
  assign w658 = ( ~w501 & w590 ) | ( ~w501 & w657 ) | ( w590 & w657 ) ;
  assign w659 = w501 & ~w658 ;
  assign w660 = \pi11 ^ w528 ;
  assign w661 = w450 & w660 ;
  assign w662 = \pi11 & ~w34 ;
  assign w663 = ( ~\pi22 & w34 ) | ( ~\pi22 & w662 ) | ( w34 & w662 ) ;
  assign w664 = \pi12 ^ w663 ;
  assign w665 = ( ~w659 & w660 ) | ( ~w659 & w664 ) | ( w660 & w664 ) ;
  assign w666 = w450 & w665 ;
  assign w667 = ( w501 & w526 ) | ( w501 & w536 ) | ( w526 & w536 ) ;
  assign w668 = ( w450 & ~w536 ) | ( w450 & w667 ) | ( ~w536 & w667 ) ;
  assign w669 = ( w501 & w526 ) | ( w501 & w532 ) | ( w526 & w532 ) ;
  assign w670 = w668 ^ w669 ;
  assign w671 = w590 & w657 ;
  assign w672 = ( w501 & ~w532 ) | ( w501 & w657 ) | ( ~w532 & w657 ) ;
  assign w673 = ( w501 & w590 ) | ( w501 & w672 ) | ( w590 & w672 ) ;
  assign w674 = w671 ^ w673 ;
  assign w675 = ( w501 & w526 ) | ( w501 & w664 ) | ( w526 & w664 ) ;
  assign w676 = ( w450 & ~w664 ) | ( w450 & w675 ) | ( ~w664 & w675 ) ;
  assign w677 = w667 ^ w676 ;
  assign w678 = ( ~w661 & w674 ) | ( ~w661 & w677 ) | ( w674 & w677 ) ;
  assign w679 = w660 ^ w664 ;
  assign w680 = w450 & w679 ;
  assign w681 = w659 ^ w680 ;
  assign w682 = ( w670 & w678 ) | ( w670 & ~w681 ) | ( w678 & ~w681 ) ;
  assign w683 = ( w230 & w363 ) | ( w230 & ~w421 ) | ( w363 & ~w421 ) ;
  assign w684 = w161 | w227 ;
  assign w685 = ( ~w227 & w421 ) | ( ~w227 & w477 ) | ( w421 & w477 ) ;
  assign w686 = w684 | w685 ;
  assign w687 = w683 | w686 ;
  assign w688 = ( ~w351 & w372 ) | ( ~w351 & w687 ) | ( w372 & w687 ) ;
  assign w689 = w351 | w688 ;
  assign w690 = w109 & w196 ;
  assign w691 = w162 | w690 ;
  assign w692 = ( w94 & ~w162 ) | ( w94 & w224 ) | ( ~w162 & w224 ) ;
  assign w693 = w691 | w692 ;
  assign w694 = ( w355 & w502 ) | ( w355 & ~w510 ) | ( w502 & ~w510 ) ;
  assign w695 = w243 | w343 ;
  assign w696 = ( ~w343 & w510 ) | ( ~w343 & w513 ) | ( w510 & w513 ) ;
  assign w697 = w695 | w696 ;
  assign w698 = w694 | w697 ;
  assign w699 = ( w125 & ~w302 ) | ( w125 & w698 ) | ( ~w302 & w698 ) ;
  assign w700 = w483 | w693 ;
  assign w701 = ( w302 & w511 ) | ( w302 & ~w693 ) | ( w511 & ~w693 ) ;
  assign w702 = w700 | w701 ;
  assign w703 = w699 | w702 ;
  assign w704 = w58 | w245 ;
  assign w705 = ( ~w58 & w214 ) | ( ~w58 & w703 ) | ( w214 & w703 ) ;
  assign w706 = w704 | w705 ;
  assign w707 = w113 | w303 ;
  assign w708 = ( w226 & w236 ) | ( w226 & ~w353 ) | ( w236 & ~w353 ) ;
  assign w709 = w124 | w139 ;
  assign w710 = ( ~w139 & w353 ) | ( ~w139 & w354 ) | ( w353 & w354 ) ;
  assign w711 = w709 | w710 ;
  assign w712 = w708 | w711 ;
  assign w713 = w220 | w479 ;
  assign w714 = ( w174 & ~w219 ) | ( w174 & w713 ) | ( ~w219 & w713 ) ;
  assign w715 = w707 | w712 ;
  assign w716 = ( w219 & w223 ) | ( w219 & ~w712 ) | ( w223 & ~w712 ) ;
  assign w717 = w715 | w716 ;
  assign w718 = w714 | w717 ;
  assign w719 = ( w188 & w265 ) | ( w188 & ~w451 ) | ( w265 & ~w451 ) ;
  assign w720 = w128 | w718 ;
  assign w721 = ( ~w128 & w451 ) | ( ~w128 & w544 ) | ( w451 & w544 ) ;
  assign w722 = w720 | w721 ;
  assign w723 = w719 | w722 ;
  assign w724 = ( w319 & w321 ) | ( w319 & ~w453 ) | ( w321 & ~w453 ) ;
  assign w725 = w123 | w163 ;
  assign w726 = ( ~w163 & w453 ) | ( ~w163 & w478 ) | ( w453 & w478 ) ;
  assign w727 = w725 | w726 ;
  assign w728 = w724 | w727 ;
  assign w729 = ( w262 & w305 ) | ( w262 & ~w307 ) | ( w305 & ~w307 ) ;
  assign w730 = w222 | w233 ;
  assign w731 = ( ~w233 & w307 ) | ( ~w233 & w411 ) | ( w307 & w411 ) ;
  assign w732 = w730 | w731 ;
  assign w733 = w729 | w732 ;
  assign w734 = ( w689 & w728 ) | ( w689 & ~w733 ) | ( w728 & ~w733 ) ;
  assign w735 = w706 | w723 ;
  assign w736 = ( w412 & ~w723 ) | ( w412 & w733 ) | ( ~w723 & w733 ) ;
  assign w737 = w735 | w736 ;
  assign w738 = w734 | w737 ;
  assign w739 = w114 | w244 ;
  assign w740 = ( ~w114 & w234 ) | ( ~w114 & w738 ) | ( w234 & w738 ) ;
  assign w741 = w739 | w740 ;
  assign w742 = w234 | w484 ;
  assign w743 = ( w161 & ~w234 ) | ( w161 & w244 ) | ( ~w234 & w244 ) ;
  assign w744 = w742 | w743 ;
  assign w745 = w183 | w352 ;
  assign w746 = ( w164 & ~w183 ) | ( w164 & w231 ) | ( ~w183 & w231 ) ;
  assign w747 = w745 | w746 ;
  assign w748 = ( w173 & w175 ) | ( w173 & ~w220 ) | ( w175 & ~w220 ) ;
  assign w749 = w71 | w115 ;
  assign w750 = ( ~w115 & w220 ) | ( ~w115 & w477 ) | ( w220 & w477 ) ;
  assign w751 = w749 | w750 ;
  assign w752 = w748 | w751 ;
  assign w753 = ( w105 & w227 ) | ( w105 & ~w334 ) | ( w227 & ~w334 ) ;
  assign w754 = w747 | w752 ;
  assign w755 = ( w334 & w374 ) | ( w334 & ~w752 ) | ( w374 & ~w752 ) ;
  assign w756 = w754 | w755 ;
  assign w757 = w753 | w756 ;
  assign w758 = ( w114 & w321 ) | ( w114 & ~w354 ) | ( w321 & ~w354 ) ;
  assign w759 = w58 | w757 ;
  assign w760 = ( ~w58 & w354 ) | ( ~w58 & w422 ) | ( w354 & w422 ) ;
  assign w761 = w759 | w760 ;
  assign w762 = w758 | w761 ;
  assign w763 = w464 | w581 ;
  assign w764 = w266 | w372 ;
  assign w765 = w306 | w764 ;
  assign w766 = ( w140 & ~w306 ) | ( w140 & w763 ) | ( ~w306 & w763 ) ;
  assign w767 = w765 | w766 ;
  assign w768 = ( ~w214 & w302 ) | ( ~w214 & w767 ) | ( w302 & w767 ) ;
  assign w769 = w214 | w768 ;
  assign w770 = w342 | w769 ;
  assign w771 = ( w133 & w617 ) | ( w133 & ~w769 ) | ( w617 & ~w769 ) ;
  assign w772 = w770 | w771 ;
  assign w773 = ( w94 & w172 ) | ( w94 & ~w233 ) | ( w172 & ~w233 ) ;
  assign w774 = w762 | w772 ;
  assign w775 = ( w233 & w304 ) | ( w233 & ~w762 ) | ( w304 & ~w762 ) ;
  assign w776 = w774 | w775 ;
  assign w777 = w773 | w776 ;
  assign w778 = w169 | w202 ;
  assign w779 = w744 | w778 ;
  assign w780 = ( w83 & ~w744 ) | ( w83 & w777 ) | ( ~w744 & w777 ) ;
  assign w781 = w779 | w780 ;
  assign w782 = w301 | w690 ;
  assign w783 = ( ~w301 & w362 ) | ( ~w301 & w781 ) | ( w362 & w781 ) ;
  assign w784 = w782 | w783 ;
  assign w785 = ( ~w590 & w741 ) | ( ~w590 & w784 ) | ( w741 & w784 ) ;
  assign w786 = w590 & ~w785 ;
  assign w787 = ~\pi22 & w29 ;
  assign w788 = \pi06 | \pi07 ;
  assign w789 = ( \pi08 & ~w29 ) | ( \pi08 & w788 ) | ( ~w29 & w788 ) ;
  assign w790 = ( ~\pi22 & w787 ) | ( ~\pi22 & w789 ) | ( w787 & w789 ) ;
  assign w791 = \pi09 ^ w790 ;
  assign w792 = w450 & w791 ;
  assign w793 = ~\pi22 & w33 ;
  assign w794 = \pi10 ^ w793 ;
  assign w795 = ( ~w786 & w791 ) | ( ~w786 & w794 ) | ( w791 & w794 ) ;
  assign w796 = w450 & w795 ;
  assign w797 = ( w536 & w590 ) | ( w536 & w657 ) | ( w590 & w657 ) ;
  assign w798 = ( w501 & ~w536 ) | ( w501 & w797 ) | ( ~w536 & w797 ) ;
  assign w799 = ( w532 & w590 ) | ( w532 & w657 ) | ( w590 & w657 ) ;
  assign w800 = w798 ^ w799 ;
  assign w801 = ( w501 & w526 ) | ( w501 & w660 ) | ( w526 & w660 ) ;
  assign w802 = ( w450 & ~w660 ) | ( w450 & w801 ) | ( ~w660 & w801 ) ;
  assign w803 = w675 ^ w802 ;
  assign w804 = w741 ^ w784 ;
  assign w805 = ~w590 & w785 ;
  assign w806 = w741 & w784 ;
  assign w807 = ( ~w532 & w590 ) | ( ~w532 & w784 ) | ( w590 & w784 ) ;
  assign w808 = ( w590 & w741 ) | ( w590 & w807 ) | ( w741 & w807 ) ;
  assign w809 = w806 ^ w808 ;
  assign w810 = ( w590 & w657 ) | ( w590 & w664 ) | ( w657 & w664 ) ;
  assign w811 = ( w501 & ~w664 ) | ( w501 & w810 ) | ( ~w664 & w810 ) ;
  assign w812 = w797 ^ w811 ;
  assign w813 = ( ~w792 & w809 ) | ( ~w792 & w812 ) | ( w809 & w812 ) ;
  assign w814 = ( w800 & w803 ) | ( w800 & w813 ) | ( w803 & w813 ) ;
  assign w815 = w661 ^ w674 ;
  assign w816 = w677 ^ w815 ;
  assign w817 = ( w796 & w814 ) | ( w796 & ~w816 ) | ( w814 & ~w816 ) ;
  assign w818 = w678 ^ w681 ;
  assign w819 = w670 ^ w818 ;
  assign w820 = ( w501 & w526 ) | ( w501 & w794 ) | ( w526 & w794 ) ;
  assign w821 = ( w450 & ~w794 ) | ( w450 & w820 ) | ( ~w794 & w820 ) ;
  assign w822 = w801 ^ w821 ;
  assign w823 = w161 | w452 ;
  assign w824 = ( w133 & w245 ) | ( w133 & ~w301 ) | ( w245 & ~w301 ) ;
  assign w825 = w128 | w823 ;
  assign w826 = ( ~w128 & w301 ) | ( ~w128 & w544 ) | ( w301 & w544 ) ;
  assign w827 = w825 | w826 ;
  assign w828 = w824 | w827 ;
  assign w829 = w354 | w477 ;
  assign w830 = w230 | w829 ;
  assign w831 = ( w171 & ~w230 ) | ( w171 & w351 ) | ( ~w230 & w351 ) ;
  assign w832 = w830 | w831 ;
  assign w833 = ( w71 & ~w146 ) | ( w71 & w832 ) | ( ~w146 & w832 ) ;
  assign w834 = w329 | w828 ;
  assign w835 = ( w146 & w307 ) | ( w146 & ~w828 ) | ( w307 & ~w828 ) ;
  assign w836 = w834 | w835 ;
  assign w837 = w833 | w836 ;
  assign w838 = ( w183 & w202 ) | ( w183 & ~w502 ) | ( w202 & ~w502 ) ;
  assign w839 = w148 | w837 ;
  assign w840 = ( ~w148 & w502 ) | ( ~w148 & w511 ) | ( w502 & w511 ) ;
  assign w841 = w839 | w840 ;
  assign w842 = w838 | w841 ;
  assign w843 = w374 | w475 ;
  assign w844 = ( w352 & ~w374 ) | ( w352 & w451 ) | ( ~w374 & w451 ) ;
  assign w845 = w843 | w844 ;
  assign w846 = ( w224 & w265 ) | ( w224 & ~w342 ) | ( w265 & ~w342 ) ;
  assign w847 = w105 | w123 ;
  assign w848 = ( ~w123 & w342 ) | ( ~w123 & w581 ) | ( w342 & w581 ) ;
  assign w849 = w847 | w848 ;
  assign w850 = w846 | w849 ;
  assign w851 = w371 | w850 ;
  assign w852 = w333 | w510 ;
  assign w853 = w125 | w852 ;
  assign w854 = ( ~w125 & w173 ) | ( ~w125 & w554 ) | ( w173 & w554 ) ;
  assign w855 = w853 | w854 ;
  assign w856 = ( w139 & ~w227 ) | ( w139 & w845 ) | ( ~w227 & w845 ) ;
  assign w857 = w851 | w855 ;
  assign w858 = ( w227 & w304 ) | ( w227 & ~w855 ) | ( w304 & ~w855 ) ;
  assign w859 = w857 | w858 ;
  assign w860 = w856 | w859 ;
  assign w861 = ( w192 & w222 ) | ( w192 & ~w226 ) | ( w222 & ~w226 ) ;
  assign w862 = w114 | w174 ;
  assign w863 = ( ~w174 & w226 ) | ( ~w174 & w690 ) | ( w226 & w690 ) ;
  assign w864 = w862 | w863 ;
  assign w865 = w861 | w864 ;
  assign w866 = w348 | w865 ;
  assign w867 = ( w190 & ~w243 ) | ( w190 & w400 ) | ( ~w243 & w400 ) ;
  assign w868 = w243 | w867 ;
  assign w869 = ( w149 & ~w355 ) | ( w149 & w411 ) | ( ~w355 & w411 ) ;
  assign w870 = w355 | w869 ;
  assign w871 = ( w162 & w191 ) | ( w162 & ~w228 ) | ( w191 & ~w228 ) ;
  assign w872 = w83 | w870 ;
  assign w873 = ( ~w83 & w228 ) | ( ~w83 & w341 ) | ( w228 & w341 ) ;
  assign w874 = w872 | w873 ;
  assign w875 = w871 | w874 ;
  assign w876 = ( w331 & w866 ) | ( w331 & w875 ) | ( w866 & w875 ) ;
  assign w877 = w842 | w860 ;
  assign w878 = ( w331 & w860 ) | ( w331 & ~w868 ) | ( w860 & ~w868 ) ;
  assign w879 = ~w877 & w878 ;
  assign w880 = ~w876 & w879 ;
  assign w881 = w305 | w545 ;
  assign w882 = w263 | w881 ;
  assign w883 = ( w263 & ~w266 ) | ( w263 & w880 ) | ( ~w266 & w880 ) ;
  assign w884 = ~w882 & w883 ;
  assign w885 = ( w226 & w354 ) | ( w226 & ~w364 ) | ( w354 & ~w364 ) ;
  assign w886 = w149 | w164 ;
  assign w887 = ( ~w164 & w364 ) | ( ~w164 & w453 ) | ( w364 & w453 ) ;
  assign w888 = w886 | w887 ;
  assign w889 = w885 | w888 ;
  assign w890 = w242 | w363 ;
  assign w891 = ( ~w242 & w361 ) | ( ~w242 & w889 ) | ( w361 & w889 ) ;
  assign w892 = w890 | w891 ;
  assign w893 = ( w114 & ~w265 ) | ( w114 & w372 ) | ( ~w265 & w372 ) ;
  assign w894 = w265 | w893 ;
  assign w895 = w476 | w478 ;
  assign w896 = ( w133 & w321 ) | ( w133 & ~w333 ) | ( w321 & ~w333 ) ;
  assign w897 = w894 | w895 ;
  assign w898 = ( w333 & w452 ) | ( w333 & ~w895 ) | ( w452 & ~w895 ) ;
  assign w899 = w897 | w898 ;
  assign w900 = w896 | w899 ;
  assign w901 = w190 | w307 ;
  assign w902 = w163 | w191 ;
  assign w903 = ( ~w163 & w171 ) | ( ~w163 & w901 ) | ( w171 & w901 ) ;
  assign w904 = w902 | w903 ;
  assign w905 = w230 | w412 ;
  assign w906 = w236 | w422 ;
  assign w907 = ( ~w236 & w400 ) | ( ~w236 & w905 ) | ( w400 & w905 ) ;
  assign w908 = w906 | w907 ;
  assign w909 = w175 | w455 ;
  assign w910 = ( w108 & ~w175 ) | ( w108 & w202 ) | ( ~w175 & w202 ) ;
  assign w911 = w909 | w910 ;
  assign w912 = ( ~w173 & w845 ) | ( ~w173 & w911 ) | ( w845 & w911 ) ;
  assign w913 = w264 | w908 ;
  assign w914 = ( w173 & ~w264 ) | ( w173 & w334 ) | ( ~w264 & w334 ) ;
  assign w915 = w913 | w914 ;
  assign w916 = w912 | w915 ;
  assign w917 = ( w169 & w228 ) | ( w169 & ~w231 ) | ( w228 & ~w231 ) ;
  assign w918 = w161 | w916 ;
  assign w919 = ( ~w161 & w231 ) | ( ~w161 & w234 ) | ( w231 & w234 ) ;
  assign w920 = w918 | w919 ;
  assign w921 = w917 | w920 ;
  assign w922 = w355 | w544 ;
  assign w923 = w172 | w922 ;
  assign w924 = ( ~w172 & w343 ) | ( ~w172 & w921 ) | ( w343 & w921 ) ;
  assign w925 = w923 | w924 ;
  assign w926 = ( w892 & w900 ) | ( w892 & ~w904 ) | ( w900 & ~w904 ) ;
  assign w927 = w606 | w925 ;
  assign w928 = ( w127 & ~w606 ) | ( w127 & w904 ) | ( ~w606 & w904 ) ;
  assign w929 = w927 | w928 ;
  assign w930 = w926 | w929 ;
  assign w931 = w304 | w510 ;
  assign w932 = ( ~w304 & w371 ) | ( ~w304 & w930 ) | ( w371 & w930 ) ;
  assign w933 = w931 | w932 ;
  assign w934 = ( w741 & w884 ) | ( w741 & ~w933 ) | ( w884 & ~w933 ) ;
  assign w935 = w741 & w934 ;
  assign w936 = \pi06 & ~w29 ;
  assign w937 = ( ~\pi22 & w29 ) | ( ~\pi22 & w936 ) | ( w29 & w936 ) ;
  assign w938 = \pi07 ^ w937 ;
  assign w939 = w450 & w938 ;
  assign w940 = ~\pi06 & w29 ;
  assign w941 = ( \pi06 & ~\pi07 ) | ( \pi06 & w940 ) | ( ~\pi07 & w940 ) ;
  assign w942 = ( \pi07 & ~\pi22 ) | ( \pi07 & w941 ) | ( ~\pi22 & w941 ) ;
  assign w943 = \pi08 ^ w942 ;
  assign w944 = ( ~w935 & w938 ) | ( ~w935 & w943 ) | ( w938 & w943 ) ;
  assign w945 = w450 & w944 ;
  assign w946 = ( w501 & w526 ) | ( w501 & w791 ) | ( w526 & w791 ) ;
  assign w947 = ( w450 & ~w791 ) | ( w450 & w946 ) | ( ~w791 & w946 ) ;
  assign w948 = w820 ^ w947 ;
  assign w949 = ( w536 & w741 ) | ( w536 & w784 ) | ( w741 & w784 ) ;
  assign w950 = ( ~w536 & w590 ) | ( ~w536 & w949 ) | ( w590 & w949 ) ;
  assign w951 = ( w532 & w741 ) | ( w532 & w784 ) | ( w741 & w784 ) ;
  assign w952 = w950 ^ w951 ;
  assign w953 = ( w590 & w657 ) | ( w590 & w660 ) | ( w657 & w660 ) ;
  assign w954 = ( w501 & ~w660 ) | ( w501 & w953 ) | ( ~w660 & w953 ) ;
  assign w955 = w810 ^ w954 ;
  assign w956 = ( w948 & w952 ) | ( w948 & w955 ) | ( w952 & w955 ) ;
  assign w957 = ( w822 & w945 ) | ( w822 & w956 ) | ( w945 & w956 ) ;
  assign w958 = w791 ^ w794 ;
  assign w959 = w450 & w958 ;
  assign w960 = w786 ^ w959 ;
  assign w961 = w800 ^ w813 ;
  assign w962 = w803 ^ w961 ;
  assign w963 = ( w957 & ~w960 ) | ( w957 & w962 ) | ( ~w960 & w962 ) ;
  assign w964 = w796 ^ w814 ;
  assign w965 = w816 ^ w964 ;
  assign w966 = ( w590 & w657 ) | ( w590 & w794 ) | ( w657 & w794 ) ;
  assign w967 = ( w501 & ~w794 ) | ( w501 & w966 ) | ( ~w794 & w966 ) ;
  assign w968 = w953 ^ w967 ;
  assign w969 = ( w501 & w526 ) | ( w501 & w943 ) | ( w526 & w943 ) ;
  assign w970 = ( w450 & ~w943 ) | ( w450 & w969 ) | ( ~w943 & w969 ) ;
  assign w971 = w946 ^ w970 ;
  assign w972 = ( w341 & ~w353 ) | ( w341 & w502 ) | ( ~w353 & w502 ) ;
  assign w973 = w353 | w972 ;
  assign w974 = w349 | w510 ;
  assign w975 = ( w172 & ~w349 ) | ( w172 & w479 ) | ( ~w349 & w479 ) ;
  assign w976 = w974 | w975 ;
  assign w977 = ( w234 & ~w452 ) | ( w234 & w976 ) | ( ~w452 & w976 ) ;
  assign w978 = w908 | w973 ;
  assign w979 = ( w452 & w545 ) | ( w452 & ~w973 ) | ( w545 & ~w973 ) ;
  assign w980 = w978 | w979 ;
  assign w981 = w977 | w980 ;
  assign w982 = ( w202 & w220 ) | ( w202 & ~w333 ) | ( w220 & ~w333 ) ;
  assign w983 = w140 | w981 ;
  assign w984 = ( ~w140 & w333 ) | ( ~w140 & w476 ) | ( w333 & w476 ) ;
  assign w985 = w983 | w984 ;
  assign w986 = w982 | w985 ;
  assign w987 = w192 | w354 ;
  assign w988 = ( w83 & ~w192 ) | ( w83 & w243 ) | ( ~w192 & w243 ) ;
  assign w989 = w987 | w988 ;
  assign w990 = ( w232 & w454 ) | ( w232 & ~w989 ) | ( w454 & ~w989 ) ;
  assign w991 = w989 | w990 ;
  assign w992 = ( w226 & w364 ) | ( w226 & ~w374 ) | ( w364 & ~w374 ) ;
  assign w993 = ( ~w222 & w374 ) | ( ~w222 & w475 ) | ( w374 & w475 ) ;
  assign w994 = w434 | w993 ;
  assign w995 = w992 | w994 ;
  assign w996 = w351 | w511 ;
  assign w997 = ( ~w351 & w362 ) | ( ~w351 & w995 ) | ( w362 & w995 ) ;
  assign w998 = w996 | w997 ;
  assign w999 = ( w126 & w231 ) | ( w126 & ~w342 ) | ( w231 & ~w342 ) ;
  assign w1000 = w550 | w601 ;
  assign w1001 = ( w342 & w591 ) | ( w342 & ~w601 ) | ( w591 & ~w601 ) ;
  assign w1002 = w1000 | w1001 ;
  assign w1003 = w999 | w1002 ;
  assign w1004 = ( w991 & w998 ) | ( w991 & ~w1003 ) | ( w998 & ~w1003 ) ;
  assign w1005 = w317 | w986 ;
  assign w1006 = ( w317 & w331 ) | ( w317 & ~w1003 ) | ( w331 & ~w1003 ) ;
  assign w1007 = ~w1005 & w1006 ;
  assign w1008 = ~w1004 & w1007 ;
  assign w1009 = ( w161 & w188 ) | ( w161 & ~w214 ) | ( w188 & ~w214 ) ;
  assign w1010 = ~w114 & w1008 ;
  assign w1011 = ( ~w114 & w214 ) | ( ~w114 & w544 ) | ( w214 & w544 ) ;
  assign w1012 = w1010 & ~w1011 ;
  assign w1013 = ~w1009 & w1012 ;
  assign w1014 = ( w231 & w305 ) | ( w231 & ~w464 ) | ( w305 & ~w464 ) ;
  assign w1015 = w94 | w172 ;
  assign w1016 = ( ~w172 & w464 ) | ( ~w172 & w591 ) | ( w464 & w591 ) ;
  assign w1017 = w1015 | w1016 ;
  assign w1018 = w1014 | w1017 ;
  assign w1019 = ( ~w228 & w400 ) | ( ~w228 & w1018 ) | ( w400 & w1018 ) ;
  assign w1020 = w228 | w1019 ;
  assign w1021 = ( w124 & ~w236 ) | ( w124 & w870 ) | ( ~w236 & w870 ) ;
  assign w1022 = w320 | w991 ;
  assign w1023 = ( w236 & ~w320 ) | ( w236 & w484 ) | ( ~w320 & w484 ) ;
  assign w1024 = w1022 | w1023 ;
  assign w1025 = w1021 | w1024 ;
  assign w1026 = ( w108 & w141 ) | ( w108 & ~w202 ) | ( w141 & ~w202 ) ;
  assign w1027 = w1020 | w1025 ;
  assign w1028 = ( w202 & w221 ) | ( w202 & ~w1020 ) | ( w221 & ~w1020 ) ;
  assign w1029 = w1027 | w1028 ;
  assign w1030 = w1026 | w1029 ;
  assign w1031 = w164 | w332 ;
  assign w1032 = ( ~w164 & w321 ) | ( ~w164 & w1030 ) | ( w321 & w1030 ) ;
  assign w1033 = w1031 | w1032 ;
  assign w1034 = ( w197 & w222 ) | ( w197 & ~w353 ) | ( w222 & ~w353 ) ;
  assign w1035 = w171 | w629 ;
  assign w1036 = ( ~w171 & w353 ) | ( ~w171 & w477 ) | ( w353 & w477 ) ;
  assign w1037 = w1035 | w1036 ;
  assign w1038 = w1034 | w1037 ;
  assign w1039 = w304 | w690 ;
  assign w1040 = ( ~w304 & w544 ) | ( ~w304 & w1038 ) | ( w544 & w1038 ) ;
  assign w1041 = w1039 | w1040 ;
  assign w1042 = ( ~w162 & w552 ) | ( ~w162 & w894 ) | ( w552 & w894 ) ;
  assign w1043 = w482 | w1041 ;
  assign w1044 = ( ~w162 & w330 ) | ( ~w162 & w482 ) | ( w330 & w482 ) ;
  assign w1045 = ~w1043 & w1044 ;
  assign w1046 = ~w1042 & w1045 ;
  assign w1047 = ( w223 & w266 ) | ( w223 & ~w342 ) | ( w266 & ~w342 ) ;
  assign w1048 = ~w148 & w1046 ;
  assign w1049 = ( ~w148 & w342 ) | ( ~w148 & w351 ) | ( w342 & w351 ) ;
  assign w1050 = w1048 & ~w1049 ;
  assign w1051 = ~w1047 & w1050 ;
  assign w1052 = w128 | w412 ;
  assign w1053 = ( w71 & ~w128 ) | ( w71 & w216 ) | ( ~w128 & w216 ) ;
  assign w1054 = w1052 | w1053 ;
  assign w1055 = ( w457 & w512 ) | ( w457 & ~w713 ) | ( w512 & ~w713 ) ;
  assign w1056 = w127 | w370 ;
  assign w1057 = ( ~w370 & w713 ) | ( ~w370 & w1054 ) | ( w713 & w1054 ) ;
  assign w1058 = w1056 | w1057 ;
  assign w1059 = w1055 | w1058 ;
  assign w1060 = ( w146 & ~w227 ) | ( w146 & w1059 ) | ( ~w227 & w1059 ) ;
  assign w1061 = ~w1033 & w1051 ;
  assign w1062 = ( w227 & w341 ) | ( w227 & w1051 ) | ( w341 & w1051 ) ;
  assign w1063 = w1061 & ~w1062 ;
  assign w1064 = ~w1060 & w1063 ;
  assign w1065 = ( ~w884 & w1013 ) | ( ~w884 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1066 = ~w884 & w1065 ;
  assign w1067 = \pi06 ^ w787 ;
  assign w1068 = w450 & w1067 ;
  assign w1069 = ( w1013 & ~w1066 ) | ( w1013 & w1068 ) | ( ~w1066 & w1068 ) ;
  assign w1070 = ( w968 & w971 ) | ( w968 & w1069 ) | ( w971 & w1069 ) ;
  assign w1071 = w884 ^ w933 ;
  assign w1072 = ~w884 & w933 ;
  assign w1073 = ( ~w532 & w741 ) | ( ~w532 & w933 ) | ( w741 & w933 ) ;
  assign w1074 = ( w741 & ~w884 ) | ( w741 & w1073 ) | ( ~w884 & w1073 ) ;
  assign w1075 = w1072 ^ w1074 ;
  assign w1076 = ( w664 & w741 ) | ( w664 & w784 ) | ( w741 & w784 ) ;
  assign w1077 = ( w590 & ~w664 ) | ( w590 & w1076 ) | ( ~w664 & w1076 ) ;
  assign w1078 = w949 ^ w1077 ;
  assign w1079 = ( ~w939 & w1075 ) | ( ~w939 & w1078 ) | ( w1075 & w1078 ) ;
  assign w1080 = w938 ^ w943 ;
  assign w1081 = w450 & w1080 ;
  assign w1082 = w935 ^ w1081 ;
  assign w1083 = ( w1070 & w1079 ) | ( w1070 & ~w1082 ) | ( w1079 & ~w1082 ) ;
  assign w1084 = w809 ^ w812 ;
  assign w1085 = w792 ^ w1084 ;
  assign w1086 = w945 ^ w956 ;
  assign w1087 = w822 ^ w1086 ;
  assign w1088 = ( w1083 & ~w1085 ) | ( w1083 & w1087 ) | ( ~w1085 & w1087 ) ;
  assign w1089 = w957 ^ w962 ;
  assign w1090 = w960 ^ w1089 ;
  assign w1091 = w1083 ^ w1087 ;
  assign w1092 = w1085 ^ w1091 ;
  assign w1093 = ( w536 & ~w884 ) | ( w536 & w933 ) | ( ~w884 & w933 ) ;
  assign w1094 = ( ~w536 & w741 ) | ( ~w536 & w1093 ) | ( w741 & w1093 ) ;
  assign w1095 = ( w532 & ~w884 ) | ( w532 & w933 ) | ( ~w884 & w933 ) ;
  assign w1096 = w1094 ^ w1095 ;
  assign w1097 = ( w590 & w657 ) | ( w590 & w791 ) | ( w657 & w791 ) ;
  assign w1098 = ( w501 & ~w791 ) | ( w501 & w1097 ) | ( ~w791 & w1097 ) ;
  assign w1099 = w966 ^ w1098 ;
  assign w1100 = ( w501 & w526 ) | ( w501 & w938 ) | ( w526 & w938 ) ;
  assign w1101 = ( w450 & ~w938 ) | ( w450 & w1100 ) | ( ~w938 & w1100 ) ;
  assign w1102 = w969 ^ w1101 ;
  assign w1103 = ( w1096 & w1099 ) | ( w1096 & w1102 ) | ( w1099 & w1102 ) ;
  assign w1104 = w939 ^ w1078 ;
  assign w1105 = w1075 ^ w1104 ;
  assign w1106 = w968 ^ w971 ;
  assign w1107 = w1069 ^ w1106 ;
  assign w1108 = ( w1103 & ~w1105 ) | ( w1103 & w1107 ) | ( ~w1105 & w1107 ) ;
  assign w1109 = w952 ^ w955 ;
  assign w1110 = w948 ^ w1109 ;
  assign w1111 = w1070 ^ w1079 ;
  assign w1112 = w1082 ^ w1111 ;
  assign w1113 = ( w1108 & w1110 ) | ( w1108 & ~w1112 ) | ( w1110 & ~w1112 ) ;
  assign w1114 = ( w660 & w741 ) | ( w660 & w784 ) | ( w741 & w784 ) ;
  assign w1115 = ( w590 & ~w660 ) | ( w590 & w1114 ) | ( ~w660 & w1114 ) ;
  assign w1116 = w1076 ^ w1115 ;
  assign w1117 = w1066 ^ w1068 ;
  assign w1118 = w1013 ^ w1117 ;
  assign w1119 = w1013 ^ w1064 ;
  assign w1120 = w884 & ~w1065 ;
  assign w1121 = w1013 | w1064 ;
  assign w1122 = ( w532 & w884 ) | ( w532 & w1064 ) | ( w884 & w1064 ) ;
  assign w1123 = ( w884 & w1013 ) | ( w884 & w1122 ) | ( w1013 & w1122 ) ;
  assign w1124 = w1121 ^ w1123 ;
  assign w1125 = w285 & w450 ;
  assign w1126 = ( ~w1013 & w1124 ) | ( ~w1013 & w1125 ) | ( w1124 & w1125 ) ;
  assign w1127 = ( w1116 & ~w1118 ) | ( w1116 & w1126 ) | ( ~w1118 & w1126 ) ;
  assign w1128 = ( w664 & ~w884 ) | ( w664 & w933 ) | ( ~w884 & w933 ) ;
  assign w1129 = ( ~w664 & w741 ) | ( ~w664 & w1128 ) | ( w741 & w1128 ) ;
  assign w1130 = w1093 ^ w1129 ;
  assign w1131 = ( w741 & w784 ) | ( w741 & w794 ) | ( w784 & w794 ) ;
  assign w1132 = ( w590 & ~w794 ) | ( w590 & w1131 ) | ( ~w794 & w1131 ) ;
  assign w1133 = w1114 ^ w1132 ;
  assign w1134 = ( w590 & w657 ) | ( w590 & w943 ) | ( w657 & w943 ) ;
  assign w1135 = ( w501 & ~w943 ) | ( w501 & w1134 ) | ( ~w943 & w1134 ) ;
  assign w1136 = w1097 ^ w1135 ;
  assign w1137 = ( w1130 & w1133 ) | ( w1130 & w1136 ) | ( w1133 & w1136 ) ;
  assign w1138 = w1096 ^ w1099 ;
  assign w1139 = w1102 ^ w1138 ;
  assign w1140 = ( w501 & w526 ) | ( w501 & w1067 ) | ( w526 & w1067 ) ;
  assign w1141 = ( w450 & ~w1067 ) | ( w450 & w1140 ) | ( ~w1067 & w1140 ) ;
  assign w1142 = w1100 ^ w1141 ;
  assign w1143 = ( ~w536 & w1013 ) | ( ~w536 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1144 = ( w536 & w884 ) | ( w536 & w1143 ) | ( w884 & w1143 ) ;
  assign w1145 = ( ~w532 & w1013 ) | ( ~w532 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1146 = w1144 ^ w1145 ;
  assign w1147 = w290 & w450 ;
  assign w1148 = ( ~w1013 & w1146 ) | ( ~w1013 & w1147 ) | ( w1146 & w1147 ) ;
  assign w1149 = ( w741 & w784 ) | ( w741 & w791 ) | ( w784 & w791 ) ;
  assign w1150 = ( w590 & ~w791 ) | ( w590 & w1149 ) | ( ~w791 & w1149 ) ;
  assign w1151 = w1131 ^ w1150 ;
  assign w1152 = ( w660 & ~w884 ) | ( w660 & w933 ) | ( ~w884 & w933 ) ;
  assign w1153 = ( ~w660 & w741 ) | ( ~w660 & w1152 ) | ( w741 & w1152 ) ;
  assign w1154 = w1128 ^ w1153 ;
  assign w1155 = ( w590 & w657 ) | ( w590 & w938 ) | ( w657 & w938 ) ;
  assign w1156 = ( w501 & ~w938 ) | ( w501 & w1155 ) | ( ~w938 & w1155 ) ;
  assign w1157 = w1134 ^ w1156 ;
  assign w1158 = ( w1151 & w1154 ) | ( w1151 & w1157 ) | ( w1154 & w1157 ) ;
  assign w1159 = ( w1142 & w1148 ) | ( w1142 & w1158 ) | ( w1148 & w1158 ) ;
  assign w1160 = ( w1137 & w1139 ) | ( w1137 & w1159 ) | ( w1139 & w1159 ) ;
  assign w1161 = w1103 ^ w1105 ;
  assign w1162 = w1107 ^ w1161 ;
  assign w1163 = ( w1127 & w1160 ) | ( w1127 & ~w1162 ) | ( w1160 & ~w1162 ) ;
  assign w1164 = w1108 ^ w1112 ;
  assign w1165 = w1110 ^ w1164 ;
  assign w1166 = w1160 ^ w1162 ;
  assign w1167 = w1127 ^ w1166 ;
  assign w1168 = w1124 ^ w1125 ;
  assign w1169 = w1013 ^ w1168 ;
  assign w1170 = w1133 ^ w1136 ;
  assign w1171 = w1130 ^ w1170 ;
  assign w1172 = ( w285 & w501 ) | ( w285 & w526 ) | ( w501 & w526 ) ;
  assign w1173 = ( ~w285 & w450 ) | ( ~w285 & w1172 ) | ( w450 & w1172 ) ;
  assign w1174 = w1140 ^ w1173 ;
  assign w1175 = ( w171 & w220 ) | ( w171 & ~w229 ) | ( w220 & ~w229 ) ;
  assign w1176 = w94 | w763 ;
  assign w1177 = ( ~w94 & w229 ) | ( ~w94 & w305 ) | ( w229 & w305 ) ;
  assign w1178 = w1176 | w1177 ;
  assign w1179 = w1175 | w1178 ;
  assign w1180 = w352 | w545 ;
  assign w1181 = ( ~w352 & w544 ) | ( ~w352 & w1179 ) | ( w544 & w1179 ) ;
  assign w1182 = w1180 | w1181 ;
  assign w1183 = ( w228 & ~w321 ) | ( w228 & w354 ) | ( ~w321 & w354 ) ;
  assign w1184 = w321 | w1183 ;
  assign w1185 = ( ~w114 & w636 ) | ( ~w114 & w1184 ) | ( w636 & w1184 ) ;
  assign w1186 = w438 | w576 ;
  assign w1187 = ( w114 & w265 ) | ( w114 & ~w576 ) | ( w265 & ~w576 ) ;
  assign w1188 = w1186 | w1187 ;
  assign w1189 = w1185 | w1188 ;
  assign w1190 = ( w242 & w343 ) | ( w242 & ~w371 ) | ( w343 & ~w371 ) ;
  assign w1191 = w222 | w1189 ;
  assign w1192 = ( ~w222 & w371 ) | ( ~w222 & w422 ) | ( w371 & w422 ) ;
  assign w1193 = w1191 | w1192 ;
  assign w1194 = w1190 | w1193 ;
  assign w1195 = w452 | w510 ;
  assign w1196 = w330 & ~w1195 ;
  assign w1197 = ( w169 & w330 ) | ( w169 & w364 ) | ( w330 & w364 ) ;
  assign w1198 = w1196 & ~w1197 ;
  assign w1199 = w348 | w360 ;
  assign w1200 = w148 | w1199 ;
  assign w1201 = ( w148 & ~w224 ) | ( w148 & w1198 ) | ( ~w224 & w1198 ) ;
  assign w1202 = ~w1200 & w1201 ;
  assign w1203 = ( w375 & ~w426 ) | ( w375 & w1202 ) | ( ~w426 & w1202 ) ;
  assign w1204 = w1182 | w1194 ;
  assign w1205 = ( w175 & w375 ) | ( w175 & ~w1194 ) | ( w375 & ~w1194 ) ;
  assign w1206 = w1204 | w1205 ;
  assign w1207 = w1203 & ~w1206 ;
  assign w1208 = ( w216 & w266 ) | ( w216 & ~w365 ) | ( w266 & ~w365 ) ;
  assign w1209 = ~w83 & w1207 ;
  assign w1210 = ( ~w83 & w365 ) | ( ~w83 & w591 ) | ( w365 & w591 ) ;
  assign w1211 = w1209 & ~w1210 ;
  assign w1212 = ~w1208 & w1211 ;
  assign w1213 = ~w219 & w1212 ;
  assign w1214 = ( w532 & w1013 ) | ( w532 & w1213 ) | ( w1013 & w1213 ) ;
  assign w1215 = w1013 | w1214 ;
  assign w1216 = ( ~w664 & w1013 ) | ( ~w664 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1217 = ( w664 & w884 ) | ( w664 & w1216 ) | ( w884 & w1216 ) ;
  assign w1218 = w1143 ^ w1217 ;
  assign w1219 = w294 & w450 ;
  assign w1220 = ( ~w1215 & w1218 ) | ( ~w1215 & w1219 ) | ( w1218 & w1219 ) ;
  assign w1221 = ( w741 & w784 ) | ( w741 & w943 ) | ( w784 & w943 ) ;
  assign w1222 = ( w590 & ~w943 ) | ( w590 & w1221 ) | ( ~w943 & w1221 ) ;
  assign w1223 = w1149 ^ w1222 ;
  assign w1224 = ( w794 & ~w884 ) | ( w794 & w933 ) | ( ~w884 & w933 ) ;
  assign w1225 = ( w741 & ~w794 ) | ( w741 & w1224 ) | ( ~w794 & w1224 ) ;
  assign w1226 = w1152 ^ w1225 ;
  assign w1227 = ( w590 & w657 ) | ( w590 & w1067 ) | ( w657 & w1067 ) ;
  assign w1228 = ( w501 & ~w1067 ) | ( w501 & w1227 ) | ( ~w1067 & w1227 ) ;
  assign w1229 = w1155 ^ w1228 ;
  assign w1230 = ( w1223 & w1226 ) | ( w1223 & w1229 ) | ( w1226 & w1229 ) ;
  assign w1231 = ( w1174 & w1220 ) | ( w1174 & w1230 ) | ( w1220 & w1230 ) ;
  assign w1232 = ( ~w1169 & w1171 ) | ( ~w1169 & w1231 ) | ( w1171 & w1231 ) ;
  assign w1233 = w1116 ^ w1118 ;
  assign w1234 = w1126 ^ w1233 ;
  assign w1235 = w1137 ^ w1159 ;
  assign w1236 = w1139 ^ w1235 ;
  assign w1237 = ( w1232 & ~w1234 ) | ( w1232 & w1236 ) | ( ~w1234 & w1236 ) ;
  assign w1238 = ~w536 & w1213 ;
  assign w1239 = w532 & ~w1213 ;
  assign w1240 = w1013 ^ w1239 ;
  assign w1241 = ( w1213 & ~w1238 ) | ( w1213 & w1240 ) | ( ~w1238 & w1240 ) ;
  assign w1242 = ( w294 & w501 ) | ( w294 & w526 ) | ( w501 & w526 ) ;
  assign w1243 = w450 & ~w1242 ;
  assign w1244 = ~w1241 & w1243 ;
  assign w1245 = ( w290 & w501 ) | ( w290 & w526 ) | ( w501 & w526 ) ;
  assign w1246 = ( ~w290 & w450 ) | ( ~w290 & w1245 ) | ( w450 & w1245 ) ;
  assign w1247 = w1172 ^ w1246 ;
  assign w1248 = ( w791 & ~w884 ) | ( w791 & w933 ) | ( ~w884 & w933 ) ;
  assign w1249 = ( w741 & ~w791 ) | ( w741 & w1248 ) | ( ~w791 & w1248 ) ;
  assign w1250 = w1224 ^ w1249 ;
  assign w1251 = ( w741 & w784 ) | ( w741 & w938 ) | ( w784 & w938 ) ;
  assign w1252 = ( w590 & ~w938 ) | ( w590 & w1251 ) | ( ~w938 & w1251 ) ;
  assign w1253 = w1221 ^ w1252 ;
  assign w1254 = ( w285 & w590 ) | ( w285 & w657 ) | ( w590 & w657 ) ;
  assign w1255 = ( ~w285 & w501 ) | ( ~w285 & w1254 ) | ( w501 & w1254 ) ;
  assign w1256 = w1227 ^ w1255 ;
  assign w1257 = ( w1250 & w1253 ) | ( w1250 & w1256 ) | ( w1253 & w1256 ) ;
  assign w1258 = ( w1244 & w1247 ) | ( w1244 & w1257 ) | ( w1247 & w1257 ) ;
  assign w1259 = w1146 ^ w1147 ;
  assign w1260 = w1013 ^ w1259 ;
  assign w1261 = w1151 ^ w1157 ;
  assign w1262 = w1154 ^ w1261 ;
  assign w1263 = ( w1258 & ~w1260 ) | ( w1258 & w1262 ) | ( ~w1260 & w1262 ) ;
  assign w1264 = w1142 ^ w1158 ;
  assign w1265 = w1148 ^ w1264 ;
  assign w1266 = w1171 ^ w1231 ;
  assign w1267 = w1169 ^ w1266 ;
  assign w1268 = ( w1263 & w1265 ) | ( w1263 & ~w1267 ) | ( w1265 & ~w1267 ) ;
  assign w1269 = w1232 ^ w1236 ;
  assign w1270 = w1234 ^ w1269 ;
  assign w1271 = ( ~w660 & w1013 ) | ( ~w660 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1272 = ( w660 & w884 ) | ( w660 & w1271 ) | ( w884 & w1271 ) ;
  assign w1273 = w1216 ^ w1272 ;
  assign w1274 = ( ~w294 & w450 ) | ( ~w294 & w1242 ) | ( w450 & w1242 ) ;
  assign w1275 = w1245 ^ w1274 ;
  assign w1276 = w1241 ^ w1243 ;
  assign w1277 = ( w1273 & w1275 ) | ( w1273 & ~w1276 ) | ( w1275 & ~w1276 ) ;
  assign w1278 = w1215 ^ w1219 ;
  assign w1279 = w1218 ^ w1278 ;
  assign w1280 = w1223 ^ w1229 ;
  assign w1281 = w1226 ^ w1280 ;
  assign w1282 = ( w1277 & ~w1279 ) | ( w1277 & w1281 ) | ( ~w1279 & w1281 ) ;
  assign w1283 = w1174 ^ w1230 ;
  assign w1284 = w1220 ^ w1283 ;
  assign w1285 = w1258 ^ w1262 ;
  assign w1286 = w1260 ^ w1285 ;
  assign w1287 = ( w1282 & w1284 ) | ( w1282 & ~w1286 ) | ( w1284 & ~w1286 ) ;
  assign w1288 = w1263 ^ w1267 ;
  assign w1289 = w1265 ^ w1288 ;
  assign w1290 = ~w660 & w1213 ;
  assign w1291 = w664 & ~w1213 ;
  assign w1292 = w1013 ^ w1291 ;
  assign w1293 = ( w1213 & ~w1290 ) | ( w1213 & w1292 ) | ( ~w1290 & w1292 ) ;
  assign w1294 = ( w294 & w590 ) | ( w294 & w657 ) | ( w590 & w657 ) ;
  assign w1295 = w501 & ~w1294 ;
  assign w1296 = ~w1293 & w1295 ;
  assign w1297 = ( ~w884 & w933 ) | ( ~w884 & w943 ) | ( w933 & w943 ) ;
  assign w1298 = ( w741 & ~w943 ) | ( w741 & w1297 ) | ( ~w943 & w1297 ) ;
  assign w1299 = w1248 ^ w1298 ;
  assign w1300 = ( w741 & w784 ) | ( w741 & w1067 ) | ( w784 & w1067 ) ;
  assign w1301 = ( w590 & ~w1067 ) | ( w590 & w1300 ) | ( ~w1067 & w1300 ) ;
  assign w1302 = w1251 ^ w1301 ;
  assign w1303 = ( w1296 & w1299 ) | ( w1296 & w1302 ) | ( w1299 & w1302 ) ;
  assign w1304 = ( w290 & w590 ) | ( w290 & w657 ) | ( w590 & w657 ) ;
  assign w1305 = ( ~w290 & w501 ) | ( ~w290 & w1304 ) | ( w501 & w1304 ) ;
  assign w1306 = w1254 ^ w1305 ;
  assign w1307 = ~w664 & w1213 ;
  assign w1308 = w536 & ~w1213 ;
  assign w1309 = w1013 ^ w1308 ;
  assign w1310 = ( w1213 & ~w1307 ) | ( w1213 & w1309 ) | ( ~w1307 & w1309 ) ;
  assign w1311 = ( ~w794 & w1013 ) | ( ~w794 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1312 = ( w794 & w884 ) | ( w794 & w1311 ) | ( w884 & w1311 ) ;
  assign w1313 = w1271 ^ w1312 ;
  assign w1314 = ( w1306 & ~w1310 ) | ( w1306 & w1313 ) | ( ~w1310 & w1313 ) ;
  assign w1315 = w1253 ^ w1256 ;
  assign w1316 = w1250 ^ w1315 ;
  assign w1317 = ( w1303 & w1314 ) | ( w1303 & w1316 ) | ( w1314 & w1316 ) ;
  assign w1318 = w1244 ^ w1257 ;
  assign w1319 = w1247 ^ w1318 ;
  assign w1320 = w1277 ^ w1281 ;
  assign w1321 = w1279 ^ w1320 ;
  assign w1322 = ( w1317 & w1319 ) | ( w1317 & ~w1321 ) | ( w1319 & ~w1321 ) ;
  assign w1323 = w1282 ^ w1286 ;
  assign w1324 = w1284 ^ w1323 ;
  assign w1325 = ( ~w884 & w933 ) | ( ~w884 & w938 ) | ( w933 & w938 ) ;
  assign w1326 = ( w741 & ~w938 ) | ( w741 & w1325 ) | ( ~w938 & w1325 ) ;
  assign w1327 = w1297 ^ w1326 ;
  assign w1328 = ( ~w791 & w1013 ) | ( ~w791 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1329 = ( w791 & w884 ) | ( w791 & w1328 ) | ( w884 & w1328 ) ;
  assign w1330 = w1311 ^ w1329 ;
  assign w1331 = ( w285 & w741 ) | ( w285 & w784 ) | ( w741 & w784 ) ;
  assign w1332 = ( ~w285 & w590 ) | ( ~w285 & w1331 ) | ( w590 & w1331 ) ;
  assign w1333 = w1300 ^ w1332 ;
  assign w1334 = ( w1327 & w1330 ) | ( w1327 & w1333 ) | ( w1330 & w1333 ) ;
  assign w1335 = w1296 ^ w1302 ;
  assign w1336 = w1299 ^ w1335 ;
  assign w1337 = w539 ^ w540 ;
  assign w1338 = ( ~w294 & w537 ) | ( ~w294 & w1337 ) | ( w537 & w1337 ) ;
  assign w1339 = w294 & w1338 ;
  assign w1340 = ( w1334 & w1336 ) | ( w1334 & w1339 ) | ( w1336 & w1339 ) ;
  assign w1341 = w1275 ^ w1276 ;
  assign w1342 = w1273 ^ w1341 ;
  assign w1343 = w1303 ^ w1314 ;
  assign w1344 = w1316 ^ w1343 ;
  assign w1345 = ( w1340 & ~w1342 ) | ( w1340 & w1344 ) | ( ~w1342 & w1344 ) ;
  assign w1346 = w1317 ^ w1319 ;
  assign w1347 = w1321 ^ w1346 ;
  assign w1348 = ~w794 & w1213 ;
  assign w1349 = w660 & ~w1213 ;
  assign w1350 = w1013 ^ w1349 ;
  assign w1351 = ( w1213 & ~w1348 ) | ( w1213 & w1350 ) | ( ~w1348 & w1350 ) ;
  assign w1352 = ( ~w943 & w1013 ) | ( ~w943 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1353 = ( w884 & w943 ) | ( w884 & w1352 ) | ( w943 & w1352 ) ;
  assign w1354 = w1328 ^ w1353 ;
  assign w1355 = ( ~w884 & w933 ) | ( ~w884 & w1067 ) | ( w933 & w1067 ) ;
  assign w1356 = ( w741 & ~w1067 ) | ( w741 & w1355 ) | ( ~w1067 & w1355 ) ;
  assign w1357 = w1325 ^ w1356 ;
  assign w1358 = ( ~w1351 & w1354 ) | ( ~w1351 & w1357 ) | ( w1354 & w1357 ) ;
  assign w1359 = ( ~w294 & w501 ) | ( ~w294 & w1294 ) | ( w501 & w1294 ) ;
  assign w1360 = w1304 ^ w1359 ;
  assign w1361 = w1293 ^ w1295 ;
  assign w1362 = ( w1358 & w1360 ) | ( w1358 & ~w1361 ) | ( w1360 & ~w1361 ) ;
  assign w1363 = w1306 ^ w1310 ;
  assign w1364 = w1313 ^ w1363 ;
  assign w1365 = ( ~w537 & w539 ) | ( ~w537 & w540 ) | ( w539 & w540 ) ;
  assign w1366 = ( w294 & w539 ) | ( w294 & w540 ) | ( w539 & w540 ) ;
  assign w1367 = ~w1365 & w1366 ;
  assign w1368 = w1336 ^ w1367 ;
  assign w1369 = w1334 ^ w1368 ;
  assign w1370 = ( w1362 & ~w1364 ) | ( w1362 & w1369 ) | ( ~w1364 & w1369 ) ;
  assign w1371 = ( w290 & w741 ) | ( w290 & w784 ) | ( w741 & w784 ) ;
  assign w1372 = ( ~w290 & w590 ) | ( ~w290 & w1371 ) | ( w590 & w1371 ) ;
  assign w1373 = w1331 ^ w1372 ;
  assign w1374 = ~w791 & w1213 ;
  assign w1375 = w794 & ~w1213 ;
  assign w1376 = w1013 ^ w1375 ;
  assign w1377 = ( w1213 & ~w1374 ) | ( w1213 & w1376 ) | ( ~w1374 & w1376 ) ;
  assign w1378 = ( w294 & w741 ) | ( w294 & w784 ) | ( w741 & w784 ) ;
  assign w1379 = w590 & ~w1378 ;
  assign w1380 = ~w1377 & w1379 ;
  assign w1381 = w590 ^ w657 ;
  assign w1382 = w294 & w1381 ;
  assign w1383 = ( w1373 & w1380 ) | ( w1373 & w1382 ) | ( w1380 & w1382 ) ;
  assign w1384 = w1327 ^ w1333 ;
  assign w1385 = w1330 ^ w1384 ;
  assign w1386 = w1360 ^ w1361 ;
  assign w1387 = w1358 ^ w1386 ;
  assign w1388 = ( ~w294 & w590 ) | ( ~w294 & w1378 ) | ( w590 & w1378 ) ;
  assign w1389 = w1371 ^ w1388 ;
  assign w1390 = ( ~w938 & w1013 ) | ( ~w938 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1391 = ( w884 & w938 ) | ( w884 & w1390 ) | ( w938 & w1390 ) ;
  assign w1392 = w1352 ^ w1391 ;
  assign w1393 = ( w285 & ~w884 ) | ( w285 & w933 ) | ( ~w884 & w933 ) ;
  assign w1394 = ( ~w285 & w741 ) | ( ~w285 & w1393 ) | ( w741 & w1393 ) ;
  assign w1395 = w1355 ^ w1394 ;
  assign w1396 = ( w1389 & w1392 ) | ( w1389 & w1395 ) | ( w1392 & w1395 ) ;
  assign w1397 = w1351 ^ w1357 ;
  assign w1398 = w1354 ^ w1397 ;
  assign w1399 = w1373 ^ w1380 ;
  assign w1400 = w1382 ^ w1399 ;
  assign w1401 = ( w1396 & ~w1398 ) | ( w1396 & w1400 ) | ( ~w1398 & w1400 ) ;
  assign w1402 = ~w938 & w1213 ;
  assign w1403 = w943 & ~w1213 ;
  assign w1404 = w1013 ^ w1403 ;
  assign w1405 = ( w1213 & ~w1402 ) | ( w1213 & w1404 ) | ( ~w1402 & w1404 ) ;
  assign w1406 = ( w294 & ~w884 ) | ( w294 & w933 ) | ( ~w884 & w933 ) ;
  assign w1407 = w741 & ~w1406 ;
  assign w1408 = ~w1405 & w1407 ;
  assign w1409 = ( ~w285 & w1013 ) | ( ~w285 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1410 = ( w285 & w884 ) | ( w285 & w1409 ) | ( w884 & w1409 ) ;
  assign w1411 = ( w1013 & w1064 ) | ( w1013 & ~w1067 ) | ( w1064 & ~w1067 ) ;
  assign w1412 = w1410 ^ w1411 ;
  assign w1413 = ( ~w294 & w741 ) | ( ~w294 & w1406 ) | ( w741 & w1406 ) ;
  assign w1414 = ( w290 & ~w884 ) | ( w290 & w933 ) | ( ~w884 & w933 ) ;
  assign w1415 = w1413 ^ w1414 ;
  assign w1416 = w1405 ^ w1407 ;
  assign w1417 = ( w1412 & w1415 ) | ( w1412 & ~w1416 ) | ( w1415 & ~w1416 ) ;
  assign w1418 = w786 ^ w805 ;
  assign w1419 = ( ~w294 & w804 ) | ( ~w294 & w1418 ) | ( w804 & w1418 ) ;
  assign w1420 = w294 & w1419 ;
  assign w1421 = ( w1408 & w1417 ) | ( w1408 & w1420 ) | ( w1417 & w1420 ) ;
  assign w1422 = ( ~w290 & w741 ) | ( ~w290 & w1414 ) | ( w741 & w1414 ) ;
  assign w1423 = w1393 ^ w1422 ;
  assign w1424 = ( w884 & w1067 ) | ( w884 & w1411 ) | ( w1067 & w1411 ) ;
  assign w1425 = w1390 ^ w1424 ;
  assign w1426 = ~w943 & w1213 ;
  assign w1427 = w791 & ~w1213 ;
  assign w1428 = w1013 ^ w1427 ;
  assign w1429 = ( w1213 & ~w1426 ) | ( w1213 & w1428 ) | ( ~w1426 & w1428 ) ;
  assign w1430 = ~w1067 & w1213 ;
  assign w1431 = w938 & ~w1213 ;
  assign w1432 = w1013 ^ w1431 ;
  assign w1433 = ( w1213 & ~w1430 ) | ( w1213 & w1432 ) | ( ~w1430 & w1432 ) ;
  assign w1434 = ( ~w290 & w1013 ) | ( ~w290 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1435 = ( w290 & w884 ) | ( w290 & w1434 ) | ( w884 & w1434 ) ;
  assign w1436 = w1409 ^ w1435 ;
  assign w1437 = ~w285 & w1213 ;
  assign w1438 = w1067 & ~w1213 ;
  assign w1439 = w1013 ^ w1438 ;
  assign w1440 = ( w1213 & ~w1437 ) | ( w1213 & w1439 ) | ( ~w1437 & w1439 ) ;
  assign w1441 = ( ~w294 & w1013 ) | ( ~w294 & w1064 ) | ( w1013 & w1064 ) ;
  assign w1442 = ~w884 & w1441 ;
  assign w1443 = ~w1440 & w1442 ;
  assign w1444 = ~w290 & w1213 ;
  assign w1445 = w285 & ~w1213 ;
  assign w1446 = w1013 ^ w1445 ;
  assign w1447 = ( w1213 & ~w1444 ) | ( w1213 & w1446 ) | ( ~w1444 & w1446 ) ;
  assign w1448 = w294 | w1013 ;
  assign w1449 = ( w290 & w1013 ) | ( w290 & ~w1213 ) | ( w1013 & ~w1213 ) ;
  assign w1450 = w1448 | w1449 ;
  assign w1451 = w1066 ^ w1120 ;
  assign w1452 = ( ~w294 & w1119 ) | ( ~w294 & w1451 ) | ( w1119 & w1451 ) ;
  assign w1453 = w294 & w1452 ;
  assign w1454 = ( w1447 & w1450 ) | ( w1447 & ~w1453 ) | ( w1450 & ~w1453 ) ;
  assign w1455 = w1440 ^ w1442 ;
  assign w1456 = w294 | w1119 ;
  assign w1457 = w1066 & ~w1456 ;
  assign w1458 = w1454 & w1455 ;
  assign w1459 = ( w1119 & w1120 ) | ( w1119 & w1456 ) | ( w1120 & w1456 ) ;
  assign w1460 = ( w1457 & ~w1458 ) | ( w1457 & w1459 ) | ( ~w1458 & w1459 ) ;
  assign w1461 = w290 & w1120 ;
  assign w1462 = ~w290 & w1066 ;
  assign w1463 = ( ~w1119 & w1460 ) | ( ~w1119 & w1462 ) | ( w1460 & w1462 ) ;
  assign w1464 = ( w1460 & w1461 ) | ( w1460 & w1463 ) | ( w1461 & w1463 ) ;
  assign w1465 = ( w1454 & w1455 ) | ( w1454 & ~w1464 ) | ( w1455 & ~w1464 ) ;
  assign w1466 = ~w1464 & w1465 ;
  assign w1467 = w294 & ~w1071 ;
  assign w1468 = w1433 ^ w1443 ;
  assign w1469 = w1436 ^ w1468 ;
  assign w1470 = ( w1466 & ~w1467 ) | ( w1466 & w1469 ) | ( ~w1467 & w1469 ) ;
  assign w1471 = ( ~w1433 & w1436 ) | ( ~w1433 & w1443 ) | ( w1436 & w1443 ) ;
  assign w1472 = w1415 ^ w1416 ;
  assign w1473 = w1412 ^ w1472 ;
  assign w1474 = ( w1470 & ~w1471 ) | ( w1470 & w1473 ) | ( ~w1471 & w1473 ) ;
  assign w1475 = ( w786 & ~w804 ) | ( w786 & w805 ) | ( ~w804 & w805 ) ;
  assign w1476 = ( w294 & w786 ) | ( w294 & w805 ) | ( w786 & w805 ) ;
  assign w1477 = ~w1475 & w1476 ;
  assign w1478 = w1417 ^ w1477 ;
  assign w1479 = w1408 ^ w1478 ;
  assign w1480 = w1423 ^ w1425 ;
  assign w1481 = w1429 ^ w1480 ;
  assign w1482 = ( w1474 & ~w1479 ) | ( w1474 & w1481 ) | ( ~w1479 & w1481 ) ;
  assign w1483 = w1389 ^ w1395 ;
  assign w1484 = w1392 ^ w1483 ;
  assign w1485 = w1377 ^ w1379 ;
  assign w1486 = ( w1423 & w1425 ) | ( w1423 & ~w1429 ) | ( w1425 & ~w1429 ) ;
  assign w1487 = w1396 ^ w1400 ;
  assign w1488 = w1398 ^ w1487 ;
  assign w1489 = ( w1421 & w1484 ) | ( w1421 & ~w1485 ) | ( w1484 & ~w1485 ) ;
  assign w1490 = ( w1421 & ~w1484 ) | ( w1421 & w1485 ) | ( ~w1484 & w1485 ) ;
  assign w1491 = ( ~w1421 & w1488 ) | ( ~w1421 & w1490 ) | ( w1488 & w1490 ) ;
  assign w1492 = ( w1482 & ~w1486 ) | ( w1482 & w1491 ) | ( ~w1486 & w1491 ) ;
  assign w1493 = ( w1488 & ~w1489 ) | ( w1488 & w1492 ) | ( ~w1489 & w1492 ) ;
  assign w1494 = w1362 ^ w1369 ;
  assign w1495 = w1364 ^ w1494 ;
  assign w1496 = ( w1383 & ~w1387 ) | ( w1383 & w1401 ) | ( ~w1387 & w1401 ) ;
  assign w1497 = ( ~w1383 & w1387 ) | ( ~w1383 & w1401 ) | ( w1387 & w1401 ) ;
  assign w1498 = ( ~w1401 & w1495 ) | ( ~w1401 & w1497 ) | ( w1495 & w1497 ) ;
  assign w1499 = ( ~w1385 & w1493 ) | ( ~w1385 & w1498 ) | ( w1493 & w1498 ) ;
  assign w1500 = ( w1495 & ~w1496 ) | ( w1495 & w1499 ) | ( ~w1496 & w1499 ) ;
  assign w1501 = w1340 ^ w1344 ;
  assign w1502 = w1342 ^ w1501 ;
  assign w1503 = ( ~w1370 & w1500 ) | ( ~w1370 & w1502 ) | ( w1500 & w1502 ) ;
  assign w1504 = ( ~w1345 & w1347 ) | ( ~w1345 & w1503 ) | ( w1347 & w1503 ) ;
  assign w1505 = ( ~w1322 & w1324 ) | ( ~w1322 & w1504 ) | ( w1324 & w1504 ) ;
  assign w1506 = ( ~w1287 & w1289 ) | ( ~w1287 & w1505 ) | ( w1289 & w1505 ) ;
  assign w1507 = ( ~w1268 & w1270 ) | ( ~w1268 & w1506 ) | ( w1270 & w1506 ) ;
  assign w1508 = ( w1167 & ~w1237 ) | ( w1167 & w1507 ) | ( ~w1237 & w1507 ) ;
  assign w1509 = ( ~w1163 & w1165 ) | ( ~w1163 & w1508 ) | ( w1165 & w1508 ) ;
  assign w1510 = ( w1092 & ~w1113 ) | ( w1092 & w1509 ) | ( ~w1113 & w1509 ) ;
  assign w1511 = ( ~w1088 & w1090 ) | ( ~w1088 & w1510 ) | ( w1090 & w1510 ) ;
  assign w1512 = ( ~w963 & w965 ) | ( ~w963 & w1511 ) | ( w965 & w1511 ) ;
  assign w1513 = ( ~w817 & w819 ) | ( ~w817 & w1512 ) | ( w819 & w1512 ) ;
  assign w1514 = w450 & w536 ;
  assign w1515 = w666 ^ w1513 ;
  assign w1516 = w682 ^ w1515 ;
  assign w1517 = ( ~w543 & w1514 ) | ( ~w543 & w1516 ) | ( w1514 & w1516 ) ;
  assign w1518 = ( w682 & ~w1513 ) | ( w682 & w1516 ) | ( ~w1513 & w1516 ) ;
  assign w1519 = w1517 ^ w1518 ;
  assign w1520 = w527 ^ w532 ;
  assign w1521 = w536 ^ w1520 ;
  assign w1522 = w450 & ~w1521 ;
  assign w1523 = w1519 ^ w1522 ;
  assign w1524 = ( w115 & ~w227 ) | ( w115 & w475 ) | ( ~w227 & w475 ) ;
  assign w1525 = w227 | w1524 ;
  assign w1526 = w348 | w362 ;
  assign w1527 = w332 | w1526 ;
  assign w1528 = ( w262 & ~w332 ) | ( w262 & w335 ) | ( ~w332 & w335 ) ;
  assign w1529 = w1527 | w1528 ;
  assign w1530 = w226 | w234 ;
  assign w1531 = w1529 | w1530 ;
  assign w1532 = ( w162 & w713 ) | ( w162 & ~w1529 ) | ( w713 & ~w1529 ) ;
  assign w1533 = w1531 | w1532 ;
  assign w1534 = w581 | w690 ;
  assign w1535 = w190 | w1534 ;
  assign w1536 = ( ~w190 & w214 ) | ( ~w190 & w1533 ) | ( w214 & w1533 ) ;
  assign w1537 = w1535 | w1536 ;
  assign w1538 = w360 | w421 ;
  assign w1539 = w222 | w1538 ;
  assign w1540 = ( w216 & ~w222 ) | ( w216 & w302 ) | ( ~w222 & w302 ) ;
  assign w1541 = w1539 | w1540 ;
  assign w1542 = w128 | w365 ;
  assign w1543 = ( w114 & ~w128 ) | ( w114 & w265 ) | ( ~w128 & w265 ) ;
  assign w1544 = w1542 | w1543 ;
  assign w1545 = ( ~w245 & w1541 ) | ( ~w245 & w1544 ) | ( w1541 & w1544 ) ;
  assign w1546 = w483 | w973 ;
  assign w1547 = ( w245 & w546 ) | ( w245 & ~w973 ) | ( w546 & ~w973 ) ;
  assign w1548 = w1546 | w1547 ;
  assign w1549 = w1545 | w1548 ;
  assign w1550 = w148 | w707 ;
  assign w1551 = ( ~w707 & w911 ) | ( ~w707 & w1549 ) | ( w911 & w1549 ) ;
  assign w1552 = w1550 | w1551 ;
  assign w1553 = ( ~w126 & w304 ) | ( ~w126 & w747 ) | ( w304 & w747 ) ;
  assign w1554 = w126 | w1553 ;
  assign w1555 = w464 | w545 ;
  assign w1556 = w139 | w1555 ;
  assign w1557 = ( ~w139 & w361 ) | ( ~w139 & w1554 ) | ( w361 & w1554 ) ;
  assign w1558 = w1556 | w1557 ;
  assign w1559 = ( ~w133 & w401 ) | ( ~w133 & w728 ) | ( w401 & w728 ) ;
  assign w1560 = w147 | w1558 ;
  assign w1561 = ( w133 & ~w147 ) | ( w133 & w342 ) | ( ~w147 & w342 ) ;
  assign w1562 = w1560 | w1561 ;
  assign w1563 = w1559 | w1562 ;
  assign w1564 = ( ~w236 & w1525 ) | ( ~w236 & w1537 ) | ( w1525 & w1537 ) ;
  assign w1565 = w1552 | w1563 ;
  assign w1566 = ( w236 & w334 ) | ( w236 & ~w1563 ) | ( w334 & ~w1563 ) ;
  assign w1567 = w1565 | w1566 ;
  assign w1568 = w1564 | w1567 ;
  assign w1569 = w371 | w511 ;
  assign w1570 = w174 | w1569 ;
  assign w1571 = ( ~w174 & w223 ) | ( ~w174 & w1568 ) | ( w223 & w1568 ) ;
  assign w1572 = w1570 | w1571 ;
  assign w1573 = w682 ^ w1513 ;
  assign w1574 = w666 ^ w1573 ;
  assign w1575 = w543 ^ w1574 ;
  assign w1576 = w1514 ^ w1575 ;
  assign w1577 = w173 | w477 ;
  assign w1578 = w128 | w1577 ;
  assign w1579 = ( w71 & ~w128 ) | ( w71 & w133 ) | ( ~w128 & w133 ) ;
  assign w1580 = w1578 | w1579 ;
  assign w1581 = ( w324 & ~w481 ) | ( w324 & w1580 ) | ( ~w481 & w1580 ) ;
  assign w1582 = w481 | w1581 ;
  assign w1583 = ( ~w629 & w892 ) | ( ~w629 & w1582 ) | ( w892 & w1582 ) ;
  assign w1584 = w598 | w986 ;
  assign w1585 = ( ~w598 & w629 ) | ( ~w598 & w693 ) | ( w629 & w693 ) ;
  assign w1586 = w1584 | w1585 ;
  assign w1587 = w1583 | w1586 ;
  assign w1588 = ( w244 & w302 ) | ( w244 & ~w362 ) | ( w302 & ~w362 ) ;
  assign w1589 = w163 | w1587 ;
  assign w1590 = ( ~w163 & w362 ) | ( ~w163 & w464 ) | ( w362 & w464 ) ;
  assign w1591 = w1589 | w1590 ;
  assign w1592 = w1588 | w1591 ;
  assign w1593 = w817 ^ w1512 ;
  assign w1594 = w819 ^ w1593 ;
  assign w1595 = ( w243 & w263 ) | ( w243 & ~w334 ) | ( w263 & ~w334 ) ;
  assign w1596 = w242 | w1544 ;
  assign w1597 = ( ~w242 & w334 ) | ( ~w242 & w335 ) | ( w334 & w335 ) ;
  assign w1598 = w1596 | w1597 ;
  assign w1599 = w1595 | w1598 ;
  assign w1600 = w629 | w1525 ;
  assign w1601 = w306 | w1600 ;
  assign w1602 = ( ~w306 & w359 ) | ( ~w306 & w1599 ) | ( w359 & w1599 ) ;
  assign w1603 = w1601 | w1602 ;
  assign w1604 = w233 | w400 ;
  assign w1605 = w214 | w1604 ;
  assign w1606 = ( ~w214 & w229 ) | ( ~w214 & w1603 ) | ( w229 & w1603 ) ;
  assign w1607 = w1605 | w1606 ;
  assign w1608 = ( w139 & w245 ) | ( w139 & ~w262 ) | ( w245 & ~w262 ) ;
  assign w1609 = w71 | w823 ;
  assign w1610 = ( ~w71 & w262 ) | ( ~w71 & w453 ) | ( w262 & w453 ) ;
  assign w1611 = w1609 | w1610 ;
  assign w1612 = w1608 | w1611 ;
  assign w1613 = ( w123 & w164 ) | ( w123 & ~w216 ) | ( w164 & ~w216 ) ;
  assign w1614 = w573 | w1612 ;
  assign w1615 = ( w216 & w222 ) | ( w216 & ~w573 ) | ( w222 & ~w573 ) ;
  assign w1616 = w1614 | w1615 ;
  assign w1617 = w1613 | w1616 ;
  assign w1618 = w422 | w690 ;
  assign w1619 = w94 | w1618 ;
  assign w1620 = ( ~w94 & w235 ) | ( ~w94 & w1617 ) | ( w235 & w1617 ) ;
  assign w1621 = w1619 | w1620 ;
  assign w1622 = ( w175 & ~w478 ) | ( w175 & w513 ) | ( ~w478 & w513 ) ;
  assign w1623 = w478 | w1622 ;
  assign w1624 = ( w307 & ~w319 ) | ( w307 & w451 ) | ( ~w319 & w451 ) ;
  assign w1625 = w319 | w1624 ;
  assign w1626 = w484 | w1625 ;
  assign w1627 = ( w348 & w1623 ) | ( w348 & ~w1625 ) | ( w1623 & ~w1625 ) ;
  assign w1628 = w1626 | w1627 ;
  assign w1629 = ( ~w150 & w569 ) | ( ~w150 & w1628 ) | ( w569 & w1628 ) ;
  assign w1630 = w1607 | w1621 ;
  assign w1631 = ( w150 & w636 ) | ( w150 & ~w1621 ) | ( w636 & ~w1621 ) ;
  assign w1632 = w1630 | w1631 ;
  assign w1633 = w1629 | w1632 ;
  assign w1634 = w322 | w546 ;
  assign w1635 = ( ~w322 & w342 ) | ( ~w322 & w1633 ) | ( w342 & w1633 ) ;
  assign w1636 = w1634 | w1635 ;
  assign w1637 = w963 ^ w1511 ;
  assign w1638 = w965 ^ w1637 ;
  assign w1639 = ( w125 & w171 ) | ( w125 & ~w188 ) | ( w171 & ~w188 ) ;
  assign w1640 = w457 | w1623 ;
  assign w1641 = ( w188 & w343 ) | ( w188 & ~w1623 ) | ( w343 & ~w1623 ) ;
  assign w1642 = w1640 | w1641 ;
  assign w1643 = w1639 | w1642 ;
  assign w1644 = ( w341 & w363 ) | ( w341 & ~w371 ) | ( w363 & ~w371 ) ;
  assign w1645 = w108 | w1643 ;
  assign w1646 = ( ~w108 & w371 ) | ( ~w108 & w591 ) | ( w371 & w591 ) ;
  assign w1647 = w1645 | w1646 ;
  assign w1648 = w1644 | w1647 ;
  assign w1649 = w146 | w301 ;
  assign w1650 = ( ~w146 & w223 ) | ( ~w146 & w1607 ) | ( w223 & w1607 ) ;
  assign w1651 = w1649 | w1650 ;
  assign w1652 = ( w244 & ~w453 ) | ( w244 & w1184 ) | ( ~w453 & w1184 ) ;
  assign w1653 = w331 & ~w1651 ;
  assign w1654 = ( w331 & w453 ) | ( w331 & w544 ) | ( w453 & w544 ) ;
  assign w1655 = w1653 & ~w1654 ;
  assign w1656 = ~w1652 & w1655 ;
  assign w1657 = ( ~w173 & w905 ) | ( ~w173 & w1648 ) | ( w905 & w1648 ) ;
  assign w1658 = ~w1558 & w1656 ;
  assign w1659 = ( w173 & w349 ) | ( w173 & ~w1558 ) | ( w349 & ~w1558 ) ;
  assign w1660 = w1658 & ~w1659 ;
  assign w1661 = ~w1657 & w1660 ;
  assign w1662 = w162 | w364 ;
  assign w1663 = ( w162 & ~w319 ) | ( w162 & w1661 ) | ( ~w319 & w1661 ) ;
  assign w1664 = ~w1662 & w1663 ;
  assign w1665 = w1088 ^ w1510 ;
  assign w1666 = w1090 ^ w1665 ;
  assign w1667 = ( w169 & w235 ) | ( w169 & ~w242 ) | ( w235 & ~w242 ) ;
  assign w1668 = w94 | w124 ;
  assign w1669 = ( ~w124 & w242 ) | ( ~w124 & w361 ) | ( w242 & w361 ) ;
  assign w1670 = w1668 | w1669 ;
  assign w1671 = w1667 | w1670 ;
  assign w1672 = ( ~w163 & w224 ) | ( ~w163 & w1671 ) | ( w224 & w1671 ) ;
  assign w1673 = w163 | w1672 ;
  assign w1674 = ( ~w231 & w373 ) | ( ~w231 & w636 ) | ( w373 & w636 ) ;
  assign w1675 = w127 | w866 ;
  assign w1676 = ( ~w127 & w231 ) | ( ~w127 & w591 ) | ( w231 & w591 ) ;
  assign w1677 = w1675 | w1676 ;
  assign w1678 = w1674 | w1677 ;
  assign w1679 = w453 | w464 ;
  assign w1680 = w343 | w1679 ;
  assign w1681 = ( ~w343 & w352 ) | ( ~w343 & w1678 ) | ( w352 & w1678 ) ;
  assign w1682 = w1680 | w1681 ;
  assign w1683 = ( ~w58 & w332 ) | ( ~w58 & w842 ) | ( w332 & w842 ) ;
  assign w1684 = w58 | w1683 ;
  assign w1685 = w236 | w476 ;
  assign w1686 = w219 | w1685 ;
  assign w1687 = ( w134 & ~w219 ) | ( w134 & w225 ) | ( ~w219 & w225 ) ;
  assign w1688 = w1686 | w1687 ;
  assign w1689 = ( ~w334 & w1673 ) | ( ~w334 & w1688 ) | ( w1673 & w1688 ) ;
  assign w1690 = w1682 | w1684 ;
  assign w1691 = ( w334 & w412 ) | ( w334 & ~w1682 ) | ( w412 & ~w1682 ) ;
  assign w1692 = w1690 | w1691 ;
  assign w1693 = w1689 | w1692 ;
  assign w1694 = ( w227 & w302 ) | ( w227 & ~w303 ) | ( w302 & ~w303 ) ;
  assign w1695 = w197 | w1693 ;
  assign w1696 = ( ~w197 & w303 ) | ( ~w197 & w455 ) | ( w303 & w455 ) ;
  assign w1697 = w1695 | w1696 ;
  assign w1698 = w1694 | w1697 ;
  assign w1699 = w451 | w1698 ;
  assign w1700 = w1092 ^ w1509 ;
  assign w1701 = w1113 ^ w1700 ;
  assign w1702 = ( w361 & w365 ) | ( w361 & ~w513 ) | ( w365 & ~w513 ) ;
  assign w1703 = w221 | w351 ;
  assign w1704 = ( ~w351 & w513 ) | ( ~w351 & w690 ) | ( w513 & w690 ) ;
  assign w1705 = w1703 | w1704 ;
  assign w1706 = w1702 | w1705 ;
  assign w1707 = w223 | w307 ;
  assign w1708 = w174 | w1707 ;
  assign w1709 = ( w71 & ~w174 ) | ( w71 & w219 ) | ( ~w174 & w219 ) ;
  assign w1710 = w1708 | w1709 ;
  assign w1711 = ( ~w125 & w333 ) | ( ~w125 & w1710 ) | ( w333 & w1710 ) ;
  assign w1712 = w125 | w1711 ;
  assign w1713 = w332 | w476 ;
  assign w1714 = w77 | w1713 ;
  assign w1715 = ( ~w77 & w164 ) | ( ~w77 & w1712 ) | ( w164 & w1712 ) ;
  assign w1716 = w1714 | w1715 ;
  assign w1717 = w124 | w134 ;
  assign w1718 = ( w58 & ~w245 ) | ( w58 & w353 ) | ( ~w245 & w353 ) ;
  assign w1719 = w245 | w1718 ;
  assign w1720 = w989 | w1719 ;
  assign w1721 = ( w438 & ~w989 ) | ( w438 & w1717 ) | ( ~w989 & w1717 ) ;
  assign w1722 = w1720 | w1721 ;
  assign w1723 = ( ~w320 & w851 ) | ( ~w320 & w1722 ) | ( w851 & w1722 ) ;
  assign w1724 = w921 | w1716 ;
  assign w1725 = ( w320 & w350 ) | ( w320 & ~w1716 ) | ( w350 & ~w1716 ) ;
  assign w1726 = w1724 | w1725 ;
  assign w1727 = w1723 | w1726 ;
  assign w1728 = w225 | w502 ;
  assign w1729 = w1706 | w1728 ;
  assign w1730 = ( w146 & ~w1706 ) | ( w146 & w1727 ) | ( ~w1706 & w1727 ) ;
  assign w1731 = w1729 | w1730 ;
  assign w1732 = w1163 ^ w1508 ;
  assign w1733 = w1165 ^ w1732 ;
  assign w1734 = ( w318 & w319 ) | ( w318 & ~w422 ) | ( w319 & ~w422 ) ;
  assign w1735 = w127 | w232 ;
  assign w1736 = ( ~w232 & w422 ) | ( ~w232 & w545 ) | ( w422 & w545 ) ;
  assign w1737 = w1735 | w1736 ;
  assign w1738 = w1734 | w1737 ;
  assign w1739 = w243 | w1738 ;
  assign w1740 = ( w263 & ~w455 ) | ( w263 & w546 ) | ( ~w455 & w546 ) ;
  assign w1741 = w455 | w1740 ;
  assign w1742 = ( w188 & w197 ) | ( w188 & ~w244 ) | ( w197 & ~w244 ) ;
  assign w1743 = w828 | w1741 ;
  assign w1744 = ( w244 & w333 ) | ( w244 & ~w1741 ) | ( w333 & ~w1741 ) ;
  assign w1745 = w1743 | w1744 ;
  assign w1746 = w1742 | w1745 ;
  assign w1747 = w353 | w510 ;
  assign w1748 = w191 | w1747 ;
  assign w1749 = ( ~w191 & w335 ) | ( ~w191 & w1746 ) | ( w335 & w1746 ) ;
  assign w1750 = w1748 | w1749 ;
  assign w1751 = ( w454 & ~w707 ) | ( w454 & w1739 ) | ( ~w707 & w1739 ) ;
  assign w1752 = w386 | w1750 ;
  assign w1753 = ( w202 & w707 ) | ( w202 & ~w1750 ) | ( w707 & ~w1750 ) ;
  assign w1754 = w1752 | w1753 ;
  assign w1755 = w1751 | w1754 ;
  assign w1756 = ( w229 & w352 ) | ( w229 & ~w400 ) | ( w352 & ~w400 ) ;
  assign w1757 = w162 | w1755 ;
  assign w1758 = ( ~w162 & w400 ) | ( ~w162 & w479 ) | ( w400 & w479 ) ;
  assign w1759 = w1757 | w1758 ;
  assign w1760 = w1756 | w1759 ;
  assign w1761 = w1167 ^ w1507 ;
  assign w1762 = w1237 ^ w1761 ;
  assign w1763 = w555 | w1625 ;
  assign w1764 = ( w105 & w823 ) | ( w105 & ~w1625 ) | ( w823 & ~w1625 ) ;
  assign w1765 = w1763 | w1764 ;
  assign w1766 = ( w77 & w231 ) | ( w77 & ~w332 ) | ( w231 & ~w332 ) ;
  assign w1767 = w415 | w1765 ;
  assign w1768 = ( w332 & w364 ) | ( w332 & ~w415 ) | ( w364 & ~w415 ) ;
  assign w1769 = w1767 | w1768 ;
  assign w1770 = w1766 | w1769 ;
  assign w1771 = ( w232 & w263 ) | ( w232 & ~w303 ) | ( w263 & ~w303 ) ;
  assign w1772 = w83 | w480 ;
  assign w1773 = ( ~w83 & w303 ) | ( ~w83 & w421 ) | ( w303 & w421 ) ;
  assign w1774 = w1772 | w1773 ;
  assign w1775 = w1771 | w1774 ;
  assign w1776 = w371 | w1775 ;
  assign w1777 = ( ~w183 & w911 ) | ( ~w183 & w1776 ) | ( w911 & w1776 ) ;
  assign w1778 = w706 | w1770 ;
  assign w1779 = ( w183 & w581 ) | ( w183 & ~w1770 ) | ( w581 & ~w1770 ) ;
  assign w1780 = w1778 | w1779 ;
  assign w1781 = w1777 | w1780 ;
  assign w1782 = ( w227 & w234 ) | ( w227 & ~w236 ) | ( w234 & ~w236 ) ;
  assign w1783 = w140 | w1781 ;
  assign w1784 = ( ~w140 & w236 ) | ( ~w140 & w342 ) | ( w236 & w342 ) ;
  assign w1785 = w1783 | w1784 ;
  assign w1786 = w1782 | w1785 ;
  assign w1787 = ( w266 & w301 ) | ( w266 & ~w348 ) | ( w301 & ~w348 ) ;
  assign w1788 = w242 | w1786 ;
  assign w1789 = ( ~w242 & w348 ) | ( ~w242 & w546 ) | ( w348 & w546 ) ;
  assign w1790 = w1788 | w1789 ;
  assign w1791 = w1787 | w1790 ;
  assign w1792 = w1268 ^ w1506 ;
  assign w1793 = w1270 ^ w1792 ;
  assign w1794 = w545 | w591 ;
  assign w1795 = w71 | w484 ;
  assign w1796 = ( ~w71 & w341 ) | ( ~w71 & w1794 ) | ( w341 & w1794 ) ;
  assign w1797 = w1795 | w1796 ;
  assign w1798 = w455 | w895 ;
  assign w1799 = ( w301 & ~w895 ) | ( w301 & w1797 ) | ( ~w895 & w1797 ) ;
  assign w1800 = w1798 | w1799 ;
  assign w1801 = ( w244 & ~w453 ) | ( w244 & w1706 ) | ( ~w453 & w1706 ) ;
  assign w1802 = w375 | w1800 ;
  assign w1803 = ( ~w375 & w453 ) | ( ~w375 & w544 ) | ( w453 & w544 ) ;
  assign w1804 = w1802 | w1803 ;
  assign w1805 = w1801 | w1804 ;
  assign w1806 = ( w231 & w362 ) | ( w231 & ~w363 ) | ( w362 & ~w363 ) ;
  assign w1807 = w845 | w1805 ;
  assign w1808 = ( w363 & w479 ) | ( w363 & ~w845 ) | ( w479 & ~w845 ) ;
  assign w1809 = w1807 | w1808 ;
  assign w1810 = w1806 | w1809 ;
  assign w1811 = w355 | w511 ;
  assign w1812 = ( w171 & w233 ) | ( w171 & ~w304 ) | ( w233 & ~w304 ) ;
  assign w1813 = w1776 | w1811 ;
  assign w1814 = ( w304 & w343 ) | ( w304 & ~w1811 ) | ( w343 & ~w1811 ) ;
  assign w1815 = w1813 | w1814 ;
  assign w1816 = w1812 | w1815 ;
  assign w1817 = ( w160 & w329 ) | ( w160 & ~w908 ) | ( w329 & ~w908 ) ;
  assign w1818 = w1810 | w1816 ;
  assign w1819 = ( w331 & ~w908 ) | ( w331 & w1816 ) | ( ~w908 & w1816 ) ;
  assign w1820 = ~w1818 & w1819 ;
  assign w1821 = ~w1817 & w1820 ;
  assign w1822 = ( w245 & w265 ) | ( w245 & ~w334 ) | ( w265 & ~w334 ) ;
  assign w1823 = ~w222 & w1821 ;
  assign w1824 = ( ~w222 & w334 ) | ( ~w222 & w364 ) | ( w334 & w364 ) ;
  assign w1825 = w1823 & ~w1824 ;
  assign w1826 = ~w1822 & w1825 ;
  assign w1827 = w1287 ^ w1505 ;
  assign w1828 = w1289 ^ w1827 ;
  assign w1829 = ( w235 & w342 ) | ( w235 & ~w352 ) | ( w342 & ~w352 ) ;
  assign w1830 = w126 | w146 ;
  assign w1831 = ( ~w146 & w352 ) | ( ~w146 & w546 ) | ( w352 & w546 ) ;
  assign w1832 = w1830 | w1831 ;
  assign w1833 = w1829 | w1832 ;
  assign w1834 = w365 | w374 ;
  assign w1835 = w173 | w1834 ;
  assign w1836 = ( w113 & ~w173 ) | ( w113 & w318 ) | ( ~w173 & w318 ) ;
  assign w1837 = w1835 | w1836 ;
  assign w1838 = w1833 | w1837 ;
  assign w1839 = ( w349 & w363 ) | ( w349 & ~w464 ) | ( w363 & ~w464 ) ;
  assign w1840 = w148 | w1838 ;
  assign w1841 = ( ~w148 & w464 ) | ( ~w148 & w544 ) | ( w464 & w544 ) ;
  assign w1842 = w1840 | w1841 ;
  assign w1843 = w1839 | w1842 ;
  assign w1844 = w301 | w455 ;
  assign w1845 = w264 | w1844 ;
  assign w1846 = ( ~w264 & w481 ) | ( ~w264 & w1716 ) | ( w481 & w1716 ) ;
  assign w1847 = w1845 | w1846 ;
  assign w1848 = ( w115 & ~w216 ) | ( w115 & w744 ) | ( ~w216 & w744 ) ;
  assign w1849 = w1843 | w1847 ;
  assign w1850 = ( w216 & w343 ) | ( w216 & ~w1843 ) | ( w343 & ~w1843 ) ;
  assign w1851 = w1849 | w1850 ;
  assign w1852 = w1848 | w1851 ;
  assign w1853 = ( w192 & w232 ) | ( w192 & ~w361 ) | ( w232 & ~w361 ) ;
  assign w1854 = w94 | w1852 ;
  assign w1855 = ( ~w94 & w361 ) | ( ~w94 & w451 ) | ( w361 & w451 ) ;
  assign w1856 = w1854 | w1855 ;
  assign w1857 = w1853 | w1856 ;
  assign w1858 = w1322 ^ w1504 ;
  assign w1859 = w1324 ^ w1858 ;
  assign w1860 = w1345 ^ w1503 ;
  assign w1861 = w1347 ^ w1860 ;
  assign w1862 = ( w233 & ~w262 ) | ( w233 & w976 ) | ( ~w262 & w976 ) ;
  assign w1863 = w375 | w832 ;
  assign w1864 = ( w262 & w305 ) | ( w262 & ~w832 ) | ( w305 & ~w832 ) ;
  assign w1865 = w1863 | w1864 ;
  assign w1866 = w1862 | w1865 ;
  assign w1867 = ( ~w192 & w693 ) | ( ~w192 & w1866 ) | ( w693 & w1866 ) ;
  assign w1868 = w1552 | w1770 ;
  assign w1869 = ( w192 & w422 ) | ( w192 & ~w1770 ) | ( w422 & ~w1770 ) ;
  assign w1870 = w1868 | w1869 ;
  assign w1871 = w1867 | w1870 ;
  assign w1872 = w190 | w591 ;
  assign w1873 = ( ~w190 & w362 ) | ( ~w190 & w1871 ) | ( w362 & w1871 ) ;
  assign w1874 = w1872 | w1873 ;
  assign w1875 = w1861 & ~w1874 ;
  assign w1876 = ( ~w1857 & w1859 ) | ( ~w1857 & w1875 ) | ( w1859 & w1875 ) ;
  assign w1877 = ( w1826 & w1828 ) | ( w1826 & w1876 ) | ( w1828 & w1876 ) ;
  assign w1878 = ( ~w1791 & w1793 ) | ( ~w1791 & w1877 ) | ( w1793 & w1877 ) ;
  assign w1879 = ( ~w1760 & w1762 ) | ( ~w1760 & w1878 ) | ( w1762 & w1878 ) ;
  assign w1880 = ( ~w1731 & w1733 ) | ( ~w1731 & w1879 ) | ( w1733 & w1879 ) ;
  assign w1881 = ( ~w1699 & w1701 ) | ( ~w1699 & w1880 ) | ( w1701 & w1880 ) ;
  assign w1882 = ( w1664 & w1666 ) | ( w1664 & w1881 ) | ( w1666 & w1881 ) ;
  assign w1883 = ( ~w1636 & w1638 ) | ( ~w1636 & w1882 ) | ( w1638 & w1882 ) ;
  assign w1884 = ( ~w1592 & w1594 ) | ( ~w1592 & w1883 ) | ( w1594 & w1883 ) ;
  assign w1885 = ( ~w1572 & w1576 ) | ( ~w1572 & w1884 ) | ( w1576 & w1884 ) ;
  assign w1886 = ( w399 & w1523 ) | ( w399 & w1885 ) | ( w1523 & w1885 ) ;
  assign w1887 = ( w188 & w220 ) | ( w188 & ~w235 ) | ( w220 & ~w235 ) ;
  assign w1888 = w115 | w175 ;
  assign w1889 = ( ~w175 & w235 ) | ( ~w175 & w412 ) | ( w235 & w412 ) ;
  assign w1890 = w1888 | w1889 ;
  assign w1891 = w1887 | w1890 ;
  assign w1892 = ( ~w171 & w372 ) | ( ~w171 & w1891 ) | ( w372 & w1891 ) ;
  assign w1893 = w171 | w1892 ;
  assign w1894 = w484 | w973 ;
  assign w1895 = ( w348 & ~w973 ) | ( w348 & w1716 ) | ( ~w973 & w1716 ) ;
  assign w1896 = w1894 | w1895 ;
  assign w1897 = ( ~w140 & w1194 ) | ( ~w140 & w1893 ) | ( w1194 & w1893 ) ;
  assign w1898 = w643 | w1896 ;
  assign w1899 = ( w140 & w304 ) | ( w140 & ~w643 ) | ( w304 & ~w643 ) ;
  assign w1900 = w1898 | w1899 ;
  assign w1901 = w1897 | w1900 ;
  assign w1902 = ( w231 & w400 ) | ( w231 & ~w544 ) | ( w400 & ~w544 ) ;
  assign w1903 = w190 | w1901 ;
  assign w1904 = ( ~w190 & w544 ) | ( ~w190 & w546 ) | ( w544 & w546 ) ;
  assign w1905 = w1903 | w1904 ;
  assign w1906 = w1902 | w1905 ;
  assign w1907 = w1886 & ~w1906 ;
  assign w1908 = w1886 ^ w1906 ;
  assign w1909 = ( w285 & ~w290 ) | ( w285 & w294 ) | ( ~w290 & w294 ) ;
  assign w1910 = ( w294 & w297 ) | ( w294 & w1909 ) | ( w297 & w1909 ) ;
  assign w1911 = w1909 ^ w1910 ;
  assign w1912 = w1576 ^ w1884 ;
  assign w1913 = w1572 ^ w1912 ;
  assign w1914 = w1523 ^ w1885 ;
  assign w1915 = w399 ^ w1914 ;
  assign w1916 = ( w290 & w294 ) | ( w290 & w297 ) | ( w294 & w297 ) ;
  assign w1917 = w290 ^ w1916 ;
  assign w1918 = w300 & w1908 ;
  assign w1919 = ( ~w1915 & w1917 ) | ( ~w1915 & w1918 ) | ( w1917 & w1918 ) ;
  assign w1920 = w1911 | w1919 ;
  assign w1921 = ( w1913 & w1919 ) | ( w1913 & w1920 ) | ( w1919 & w1920 ) ;
  assign w1922 = w1918 | w1921 ;
  assign w1923 = w298 & w299 ;
  assign w1924 = w1594 ^ w1883 ;
  assign w1925 = w1592 ^ w1924 ;
  assign w1926 = w1638 ^ w1882 ;
  assign w1927 = w1636 ^ w1926 ;
  assign w1928 = w1666 ^ w1881 ;
  assign w1929 = w1664 ^ w1928 ;
  assign w1930 = w1701 ^ w1880 ;
  assign w1931 = w1699 ^ w1930 ;
  assign w1932 = w1733 ^ w1879 ;
  assign w1933 = w1731 ^ w1932 ;
  assign w1934 = w1762 ^ w1878 ;
  assign w1935 = w1760 ^ w1934 ;
  assign w1936 = w1793 ^ w1877 ;
  assign w1937 = w1791 ^ w1936 ;
  assign w1938 = w1828 ^ w1876 ;
  assign w1939 = w1826 ^ w1938 ;
  assign w1940 = w1859 ^ w1875 ;
  assign w1941 = w1857 ^ w1940 ;
  assign w1942 = w1861 ^ w1874 ;
  assign w1943 = w1939 | w1942 ;
  assign w1944 = ( w1937 & ~w1939 ) | ( w1937 & w1941 ) | ( ~w1939 & w1941 ) ;
  assign w1945 = ( w1942 & ~w1943 ) | ( w1942 & w1944 ) | ( ~w1943 & w1944 ) ;
  assign w1946 = ( w1935 & w1937 ) | ( w1935 & w1945 ) | ( w1937 & w1945 ) ;
  assign w1947 = ( w1933 & w1935 ) | ( w1933 & w1946 ) | ( w1935 & w1946 ) ;
  assign w1948 = ( w1931 & w1933 ) | ( w1931 & w1947 ) | ( w1933 & w1947 ) ;
  assign w1949 = ( ~w1929 & w1931 ) | ( ~w1929 & w1948 ) | ( w1931 & w1948 ) ;
  assign w1950 = ( w1927 & ~w1929 ) | ( w1927 & w1949 ) | ( ~w1929 & w1949 ) ;
  assign w1951 = ( w1925 & w1927 ) | ( w1925 & w1950 ) | ( w1927 & w1950 ) ;
  assign w1952 = ( w1913 & w1925 ) | ( w1913 & w1951 ) | ( w1925 & w1951 ) ;
  assign w1953 = w1913 ^ w1915 ;
  assign w1954 = ( w1913 & ~w1915 ) | ( w1913 & w1952 ) | ( ~w1915 & w1952 ) ;
  assign w1955 = w1908 ^ w1954 ;
  assign w1956 = w1915 ^ w1955 ;
  assign w1957 = w1923 & w1956 ;
  assign w1958 = ( w1922 & w1923 ) | ( w1922 & ~w1957 ) | ( w1923 & ~w1957 ) ;
  assign w1959 = w285 ^ w1958 ;
  assign w1960 = w679 & w1942 ;
  assign w1961 = ( w536 & w660 ) | ( w536 & w664 ) | ( w660 & w664 ) ;
  assign w1962 = w536 ^ w1961 ;
  assign w1963 = w532 ^ w536 ;
  assign w1964 = w679 & ~w1963 ;
  assign w1965 = w679 & w1963 ;
  assign w1966 = ( ~w532 & w660 ) | ( ~w532 & w664 ) | ( w660 & w664 ) ;
  assign w1967 = ( w660 & w664 ) | ( w660 & ~w1966 ) | ( w664 & ~w1966 ) ;
  assign w1968 = w536 ^ w1967 ;
  assign w1969 = w1942 & w1968 ;
  assign w1970 = w1941 ^ w1967 ;
  assign w1971 = ( w660 & w664 ) | ( w660 & ~w1970 ) | ( w664 & ~w1970 ) ;
  assign w1972 = ( w532 & w1966 ) | ( w532 & ~w1971 ) | ( w1966 & ~w1971 ) ;
  assign w1973 = w1969 ^ w1972 ;
  assign w1974 = ( w532 & w1960 ) | ( w532 & w1973 ) | ( w1960 & w1973 ) ;
  assign w1975 = ~w1960 & w1974 ;
  assign w1976 = w532 & ~w1960 ;
  assign w1977 = w1973 ^ w1976 ;
  assign w1978 = w791 ^ w943 ;
  assign w1979 = w660 ^ w794 ;
  assign w1980 = w1978 & w1979 ;
  assign w1981 = ( w660 & w791 ) | ( w660 & ~w794 ) | ( w791 & ~w794 ) ;
  assign w1982 = ( w791 & w943 ) | ( w791 & w1981 ) | ( w943 & w1981 ) ;
  assign w1983 = w1981 ^ w1982 ;
  assign w1984 = ( w791 & w794 ) | ( w791 & w943 ) | ( w794 & w943 ) ;
  assign w1985 = w794 ^ w1984 ;
  assign w1986 = w1978 & ~w1979 ;
  assign w1987 = ~w1939 & w1983 ;
  assign w1988 = ( w1937 & w1985 ) | ( w1937 & w1987 ) | ( w1985 & w1987 ) ;
  assign w1989 = w1986 | w1988 ;
  assign w1990 = ( w1935 & w1988 ) | ( w1935 & w1989 ) | ( w1988 & w1989 ) ;
  assign w1991 = w1987 | w1990 ;
  assign w1992 = w1935 ^ w1945 ;
  assign w1993 = w1937 ^ w1992 ;
  assign w1994 = w1980 & ~w1993 ;
  assign w1995 = ( w1980 & w1991 ) | ( w1980 & ~w1994 ) | ( w1991 & ~w1994 ) ;
  assign w1996 = w660 ^ w1995 ;
  assign w1997 = w1942 & w1978 ;
  assign w1998 = ( w791 & w794 ) | ( w791 & ~w943 ) | ( w794 & ~w943 ) ;
  assign w1999 = ( w791 & w1942 ) | ( w791 & w1998 ) | ( w1942 & w1998 ) ;
  assign w2000 = ( ~w660 & w791 ) | ( ~w660 & w1998 ) | ( w791 & w1998 ) ;
  assign w2001 = w1999 & ~w2000 ;
  assign w2002 = w660 | w1942 ;
  assign w2003 = w1978 & w2002 ;
  assign w2004 = ( w794 & ~w1942 ) | ( w794 & w2003 ) | ( ~w1942 & w2003 ) ;
  assign w2005 = w1941 ^ w2004 ;
  assign w2006 = w2003 & ~w2005 ;
  assign w2007 = w2001 | w2006 ;
  assign w2008 = ( w791 & ~w794 ) | ( w791 & w943 ) | ( ~w794 & w943 ) ;
  assign w2009 = w794 ^ w2008 ;
  assign w2010 = w1941 & w1978 ;
  assign w2011 = ( w1942 & w2009 ) | ( w1942 & w2010 ) | ( w2009 & w2010 ) ;
  assign w2012 = ( w660 & ~w2007 ) | ( w660 & w2011 ) | ( ~w2007 & w2011 ) ;
  assign w2013 = ~w2007 & w2012 ;
  assign w2014 = ( w660 & w1997 ) | ( w660 & w2013 ) | ( w1997 & w2013 ) ;
  assign w2015 = ~w1997 & w2014 ;
  assign w2016 = w1942 & w1983 ;
  assign w2017 = ( w1941 & w1985 ) | ( w1941 & w2016 ) | ( w1985 & w2016 ) ;
  assign w2018 = w1986 | w2017 ;
  assign w2019 = ( ~w1939 & w2017 ) | ( ~w1939 & w2018 ) | ( w2017 & w2018 ) ;
  assign w2020 = w2016 | w2019 ;
  assign w2021 = w1941 & ~w1942 ;
  assign w2022 = w1939 ^ w2021 ;
  assign w2023 = w1980 & w2022 ;
  assign w2024 = ( w1980 & w2020 ) | ( w1980 & ~w2023 ) | ( w2020 & ~w2023 ) ;
  assign w2025 = w660 ^ w2024 ;
  assign w2026 = w2015 & w2025 ;
  assign w2027 = w1941 & w1983 ;
  assign w2028 = ( ~w1939 & w1985 ) | ( ~w1939 & w2027 ) | ( w1985 & w2027 ) ;
  assign w2029 = w1986 | w2028 ;
  assign w2030 = ( w1937 & w2028 ) | ( w1937 & w2029 ) | ( w2028 & w2029 ) ;
  assign w2031 = w2027 | w2030 ;
  assign w2032 = w1937 ^ w1941 ;
  assign w2033 = w1939 & ~w1941 ;
  assign w2034 = ( w1939 & w1942 ) | ( w1939 & w2033 ) | ( w1942 & w2033 ) ;
  assign w2035 = w2032 ^ w2034 ;
  assign w2036 = w1980 & w2035 ;
  assign w2037 = ( w1980 & w2031 ) | ( w1980 & ~w2036 ) | ( w2031 & ~w2036 ) ;
  assign w2038 = w660 ^ w2037 ;
  assign w2039 = ( w1960 & w2026 ) | ( w1960 & w2038 ) | ( w2026 & w2038 ) ;
  assign w2040 = ( w1977 & w1996 ) | ( w1977 & w2039 ) | ( w1996 & w2039 ) ;
  assign w2041 = w1937 & w1983 ;
  assign w2042 = ( w1935 & w1985 ) | ( w1935 & w2041 ) | ( w1985 & w2041 ) ;
  assign w2043 = w1986 | w2042 ;
  assign w2044 = ( w1933 & w2042 ) | ( w1933 & w2043 ) | ( w2042 & w2043 ) ;
  assign w2045 = w2041 | w2044 ;
  assign w2046 = w1933 ^ w1946 ;
  assign w2047 = w1935 ^ w2046 ;
  assign w2048 = w1980 & ~w2047 ;
  assign w2049 = ( w1980 & w2045 ) | ( w1980 & ~w2048 ) | ( w2045 & ~w2048 ) ;
  assign w2050 = w660 ^ w2049 ;
  assign w2051 = ( w532 & ~w536 ) | ( w532 & w660 ) | ( ~w536 & w660 ) ;
  assign w2052 = ( w660 & w664 ) | ( w660 & w2051 ) | ( w664 & w2051 ) ;
  assign w2053 = w2051 ^ w2052 ;
  assign w2054 = w1941 & w1962 ;
  assign w2055 = ( w1942 & w2053 ) | ( w1942 & w2054 ) | ( w2053 & w2054 ) ;
  assign w2056 = w1964 | w2055 ;
  assign w2057 = ( ~w1939 & w2055 ) | ( ~w1939 & w2056 ) | ( w2055 & w2056 ) ;
  assign w2058 = w2054 | w2057 ;
  assign w2059 = w1965 | w2022 ;
  assign w2060 = ( ~w2022 & w2058 ) | ( ~w2022 & w2059 ) | ( w2058 & w2059 ) ;
  assign w2061 = w532 ^ w2060 ;
  assign w2062 = w1975 & w2061 ;
  assign w2063 = w1975 ^ w2061 ;
  assign w2064 = w2040 ^ w2050 ;
  assign w2065 = w2063 ^ w2064 ;
  assign w2066 = w285 ^ w1067 ;
  assign w2067 = ~w1080 & w2066 ;
  assign w2068 = ( w938 & w943 ) | ( w938 & ~w1067 ) | ( w943 & ~w1067 ) ;
  assign w2069 = ( w285 & w938 ) | ( w285 & w2068 ) | ( w938 & w2068 ) ;
  assign w2070 = w2068 ^ w2069 ;
  assign w2071 = ( w285 & w938 ) | ( w285 & w1067 ) | ( w938 & w1067 ) ;
  assign w2072 = w938 ^ w2071 ;
  assign w2073 = w1927 & w2067 ;
  assign w2074 = ( ~w1929 & w2072 ) | ( ~w1929 & w2073 ) | ( w2072 & w2073 ) ;
  assign w2075 = w2070 | w2074 ;
  assign w2076 = ( w1931 & w2074 ) | ( w1931 & w2075 ) | ( w2074 & w2075 ) ;
  assign w2077 = w2073 | w2076 ;
  assign w2078 = w1927 ^ w1949 ;
  assign w2079 = w1929 ^ w2078 ;
  assign w2080 = w1080 & w2066 ;
  assign w2081 = w2079 & w2080 ;
  assign w2082 = ( w2077 & w2080 ) | ( w2077 & ~w2081 ) | ( w2080 & ~w2081 ) ;
  assign w2083 = w943 ^ w2082 ;
  assign w2084 = ~w1929 & w2067 ;
  assign w2085 = ( w1931 & w2072 ) | ( w1931 & w2084 ) | ( w2072 & w2084 ) ;
  assign w2086 = w2070 | w2085 ;
  assign w2087 = ( w1933 & w2085 ) | ( w1933 & w2086 ) | ( w2085 & w2086 ) ;
  assign w2088 = w2084 | w2087 ;
  assign w2089 = w1929 ^ w1948 ;
  assign w2090 = w1931 ^ w2089 ;
  assign w2091 = w2080 & w2090 ;
  assign w2092 = ( w2080 & w2088 ) | ( w2080 & ~w2091 ) | ( w2088 & ~w2091 ) ;
  assign w2093 = w943 ^ w2092 ;
  assign w2094 = w1996 ^ w2039 ;
  assign w2095 = w1977 ^ w2094 ;
  assign w2096 = w2026 ^ w2038 ;
  assign w2097 = w1960 ^ w2096 ;
  assign w2098 = w1931 & w2067 ;
  assign w2099 = ( w1933 & w2072 ) | ( w1933 & w2098 ) | ( w2072 & w2098 ) ;
  assign w2100 = w2070 | w2099 ;
  assign w2101 = ( w1935 & w2099 ) | ( w1935 & w2100 ) | ( w2099 & w2100 ) ;
  assign w2102 = w2098 | w2101 ;
  assign w2103 = w1931 ^ w1947 ;
  assign w2104 = w1933 ^ w2103 ;
  assign w2105 = w2080 & ~w2104 ;
  assign w2106 = ( w2080 & w2102 ) | ( w2080 & ~w2105 ) | ( w2102 & ~w2105 ) ;
  assign w2107 = w943 ^ w2106 ;
  assign w2108 = w1933 & w2067 ;
  assign w2109 = ( w1935 & w2072 ) | ( w1935 & w2108 ) | ( w2072 & w2108 ) ;
  assign w2110 = w2070 | w2109 ;
  assign w2111 = ( w1937 & w2109 ) | ( w1937 & w2110 ) | ( w2109 & w2110 ) ;
  assign w2112 = w2108 | w2111 ;
  assign w2113 = w2047 & ~w2080 ;
  assign w2114 = ( w2047 & w2112 ) | ( w2047 & ~w2113 ) | ( w2112 & ~w2113 ) ;
  assign w2115 = w943 ^ w2114 ;
  assign w2116 = w2015 ^ w2025 ;
  assign w2117 = w660 & ~w1997 ;
  assign w2118 = w2013 ^ w2117 ;
  assign w2119 = w1935 & w2067 ;
  assign w2120 = ( w1937 & w2072 ) | ( w1937 & w2119 ) | ( w2072 & w2119 ) ;
  assign w2121 = w2070 | w2120 ;
  assign w2122 = ( ~w1939 & w2120 ) | ( ~w1939 & w2121 ) | ( w2120 & w2121 ) ;
  assign w2123 = w2119 | w2122 ;
  assign w2124 = w1993 & ~w2080 ;
  assign w2125 = ( w1993 & w2123 ) | ( w1993 & ~w2124 ) | ( w2123 & ~w2124 ) ;
  assign w2126 = w943 ^ w2125 ;
  assign w2127 = w1942 & w2066 ;
  assign w2128 = ( w285 & w943 ) | ( w285 & w1067 ) | ( w943 & w1067 ) ;
  assign w2129 = w943 & ~w1942 ;
  assign w2130 = ~w1941 & w2129 ;
  assign w2131 = ( w285 & w1067 ) | ( w285 & w2130 ) | ( w1067 & w2130 ) ;
  assign w2132 = ( ~w938 & w943 ) | ( ~w938 & w2131 ) | ( w943 & w2131 ) ;
  assign w2133 = ( w938 & w2129 ) | ( w938 & w2131 ) | ( w2129 & w2131 ) ;
  assign w2134 = ( ~w2128 & w2132 ) | ( ~w2128 & w2133 ) | ( w2132 & w2133 ) ;
  assign w2135 = ~w1939 & w2067 ;
  assign w2136 = ( w1941 & w2072 ) | ( w1941 & w2135 ) | ( w2072 & w2135 ) ;
  assign w2137 = w2070 | w2136 ;
  assign w2138 = ( w1942 & w2136 ) | ( w1942 & w2137 ) | ( w2136 & w2137 ) ;
  assign w2139 = w2135 | w2138 ;
  assign w2140 = w2022 | w2080 ;
  assign w2141 = ( ~w2022 & w2139 ) | ( ~w2022 & w2140 ) | ( w2139 & w2140 ) ;
  assign w2142 = w943 ^ w2141 ;
  assign w2143 = w2134 & w2142 ;
  assign w2144 = w1937 & w2067 ;
  assign w2145 = ( ~w1939 & w2072 ) | ( ~w1939 & w2144 ) | ( w2072 & w2144 ) ;
  assign w2146 = w2070 | w2145 ;
  assign w2147 = ( w1941 & w2145 ) | ( w1941 & w2146 ) | ( w2145 & w2146 ) ;
  assign w2148 = w2144 | w2147 ;
  assign w2149 = w2035 | w2080 ;
  assign w2150 = ( ~w2035 & w2148 ) | ( ~w2035 & w2149 ) | ( w2148 & w2149 ) ;
  assign w2151 = w943 ^ w2150 ;
  assign w2152 = ( w1997 & w2143 ) | ( w1997 & w2151 ) | ( w2143 & w2151 ) ;
  assign w2153 = ( w2118 & w2126 ) | ( w2118 & w2152 ) | ( w2126 & w2152 ) ;
  assign w2154 = ( w2115 & w2116 ) | ( w2115 & w2153 ) | ( w2116 & w2153 ) ;
  assign w2155 = ( w2097 & w2107 ) | ( w2097 & w2154 ) | ( w2107 & w2154 ) ;
  assign w2156 = ( w2093 & w2095 ) | ( w2093 & w2155 ) | ( w2095 & w2155 ) ;
  assign w2157 = ( w2065 & w2083 ) | ( w2065 & w2156 ) | ( w2083 & w2156 ) ;
  assign w2158 = w1935 & w1983 ;
  assign w2159 = ( w1933 & w1985 ) | ( w1933 & w2158 ) | ( w1985 & w2158 ) ;
  assign w2160 = w1986 | w2159 ;
  assign w2161 = ( w1931 & w2159 ) | ( w1931 & w2160 ) | ( w2159 & w2160 ) ;
  assign w2162 = w2158 | w2161 ;
  assign w2163 = ~w1980 & w2104 ;
  assign w2164 = ( w2104 & w2162 ) | ( w2104 & ~w2163 ) | ( w2162 & ~w2163 ) ;
  assign w2165 = w660 ^ w2164 ;
  assign w2166 = ~w1939 & w1962 ;
  assign w2167 = ( w1941 & w2053 ) | ( w1941 & w2166 ) | ( w2053 & w2166 ) ;
  assign w2168 = w1964 | w2167 ;
  assign w2169 = ( w1937 & w2167 ) | ( w1937 & w2168 ) | ( w2167 & w2168 ) ;
  assign w2170 = w2166 | w2169 ;
  assign w2171 = w1965 | w2035 ;
  assign w2172 = ( ~w2035 & w2170 ) | ( ~w2035 & w2171 ) | ( w2170 & w2171 ) ;
  assign w2173 = w532 ^ w2172 ;
  assign w2174 = w532 & w1942 ;
  assign w2175 = ( w2062 & w2173 ) | ( w2062 & w2174 ) | ( w2173 & w2174 ) ;
  assign w2176 = w2062 ^ w2174 ;
  assign w2177 = w2173 ^ w2176 ;
  assign w2178 = ( w2040 & w2050 ) | ( w2040 & w2063 ) | ( w2050 & w2063 ) ;
  assign w2179 = w2165 ^ w2178 ;
  assign w2180 = w2177 ^ w2179 ;
  assign w2181 = w1925 ^ w1950 ;
  assign w2182 = w1927 ^ w2181 ;
  assign w2183 = w1925 & w2067 ;
  assign w2184 = ( w1927 & w2072 ) | ( w1927 & w2183 ) | ( w2072 & w2183 ) ;
  assign w2185 = w2070 | w2184 ;
  assign w2186 = ( ~w1929 & w2184 ) | ( ~w1929 & w2185 ) | ( w2184 & w2185 ) ;
  assign w2187 = w2183 | w2186 ;
  assign w2188 = ~w2080 & w2182 ;
  assign w2189 = ( w2182 & w2187 ) | ( w2182 & ~w2188 ) | ( w2187 & ~w2188 ) ;
  assign w2190 = w943 ^ w2189 ;
  assign w2191 = w2157 ^ w2190 ;
  assign w2192 = w2180 ^ w2191 ;
  assign w2193 = w2083 ^ w2156 ;
  assign w2194 = w2065 ^ w2193 ;
  assign w2195 = w300 & ~w1915 ;
  assign w2196 = ( w1913 & w1917 ) | ( w1913 & w2195 ) | ( w1917 & w2195 ) ;
  assign w2197 = w1911 | w2196 ;
  assign w2198 = ( w1925 & w2196 ) | ( w1925 & w2197 ) | ( w2196 & w2197 ) ;
  assign w2199 = w2195 | w2198 ;
  assign w2200 = w1952 ^ w1953 ;
  assign w2201 = w1923 | w2200 ;
  assign w2202 = ( w2199 & ~w2200 ) | ( w2199 & w2201 ) | ( ~w2200 & w2201 ) ;
  assign w2203 = w285 ^ w2202 ;
  assign w2204 = w2093 ^ w2155 ;
  assign w2205 = w2095 ^ w2204 ;
  assign w2206 = w300 & w1913 ;
  assign w2207 = ( w1917 & w1925 ) | ( w1917 & w2206 ) | ( w1925 & w2206 ) ;
  assign w2208 = w1911 | w2207 ;
  assign w2209 = ( w1927 & w2207 ) | ( w1927 & w2208 ) | ( w2207 & w2208 ) ;
  assign w2210 = w2206 | w2209 ;
  assign w2211 = w1913 ^ w1951 ;
  assign w2212 = w1925 ^ w2211 ;
  assign w2213 = w1923 & ~w2212 ;
  assign w2214 = ( w1923 & w2210 ) | ( w1923 & ~w2213 ) | ( w2210 & ~w2213 ) ;
  assign w2215 = w285 ^ w2214 ;
  assign w2216 = w2107 ^ w2154 ;
  assign w2217 = w2097 ^ w2216 ;
  assign w2218 = w300 & w1925 ;
  assign w2219 = ( w1917 & w1927 ) | ( w1917 & w2218 ) | ( w1927 & w2218 ) ;
  assign w2220 = w1911 | w2219 ;
  assign w2221 = ( ~w1929 & w2219 ) | ( ~w1929 & w2220 ) | ( w2219 & w2220 ) ;
  assign w2222 = w2218 | w2221 ;
  assign w2223 = ~w1923 & w2182 ;
  assign w2224 = ( w2182 & w2222 ) | ( w2182 & ~w2223 ) | ( w2222 & ~w2223 ) ;
  assign w2225 = w285 ^ w2224 ;
  assign w2226 = w2115 ^ w2153 ;
  assign w2227 = w2116 ^ w2226 ;
  assign w2228 = w300 & w1927 ;
  assign w2229 = ( w1917 & ~w1929 ) | ( w1917 & w2228 ) | ( ~w1929 & w2228 ) ;
  assign w2230 = w1911 | w2229 ;
  assign w2231 = ( w1931 & w2229 ) | ( w1931 & w2230 ) | ( w2229 & w2230 ) ;
  assign w2232 = w2228 | w2231 ;
  assign w2233 = w1923 | w2079 ;
  assign w2234 = ( ~w2079 & w2232 ) | ( ~w2079 & w2233 ) | ( w2232 & w2233 ) ;
  assign w2235 = w285 ^ w2234 ;
  assign w2236 = w300 & ~w1929 ;
  assign w2237 = ( w1917 & w1931 ) | ( w1917 & w2236 ) | ( w1931 & w2236 ) ;
  assign w2238 = w1911 | w2237 ;
  assign w2239 = ( w1933 & w2237 ) | ( w1933 & w2238 ) | ( w2237 & w2238 ) ;
  assign w2240 = w2236 | w2239 ;
  assign w2241 = w1923 | w2090 ;
  assign w2242 = ( ~w2090 & w2240 ) | ( ~w2090 & w2241 ) | ( w2240 & w2241 ) ;
  assign w2243 = w285 ^ w2242 ;
  assign w2244 = w2126 ^ w2152 ;
  assign w2245 = w2118 ^ w2244 ;
  assign w2246 = w2143 ^ w2151 ;
  assign w2247 = w1997 ^ w2246 ;
  assign w2248 = w300 & w1931 ;
  assign w2249 = ( w1917 & w1933 ) | ( w1917 & w2248 ) | ( w1933 & w2248 ) ;
  assign w2250 = w1911 | w2249 ;
  assign w2251 = ( w1935 & w2249 ) | ( w1935 & w2250 ) | ( w2249 & w2250 ) ;
  assign w2252 = w2248 | w2251 ;
  assign w2253 = ~w1923 & w2104 ;
  assign w2254 = ( w2104 & w2252 ) | ( w2104 & ~w2253 ) | ( w2252 & ~w2253 ) ;
  assign w2255 = w285 ^ w2254 ;
  assign w2256 = w300 & w1933 ;
  assign w2257 = ( w1917 & w1935 ) | ( w1917 & w2256 ) | ( w1935 & w2256 ) ;
  assign w2258 = w1911 | w2257 ;
  assign w2259 = ( w1937 & w2257 ) | ( w1937 & w2258 ) | ( w2257 & w2258 ) ;
  assign w2260 = w2256 | w2259 ;
  assign w2261 = ~w1923 & w2047 ;
  assign w2262 = ( w2047 & w2260 ) | ( w2047 & ~w2261 ) | ( w2260 & ~w2261 ) ;
  assign w2263 = w285 ^ w2262 ;
  assign w2264 = w2134 ^ w2142 ;
  assign w2265 = w285 & w1067 ;
  assign w2266 = w1942 ^ w2265 ;
  assign w2267 = ( w938 & w2265 ) | ( w938 & w2266 ) | ( w2265 & w2266 ) ;
  assign w2268 = ( w285 & w1067 ) | ( w285 & w1941 ) | ( w1067 & w1941 ) ;
  assign w2269 = w2267 ^ w2268 ;
  assign w2270 = w300 & w1935 ;
  assign w2271 = ( w1917 & w1937 ) | ( w1917 & w2270 ) | ( w1937 & w2270 ) ;
  assign w2272 = w1911 | w2271 ;
  assign w2273 = ( ~w1939 & w2271 ) | ( ~w1939 & w2272 ) | ( w2271 & w2272 ) ;
  assign w2274 = w2270 | w2273 ;
  assign w2275 = ~w1923 & w1993 ;
  assign w2276 = ( w1993 & w2274 ) | ( w1993 & ~w2275 ) | ( w2274 & ~w2275 ) ;
  assign w2277 = w285 ^ w2276 ;
  assign w2278 = ( w285 & w294 ) | ( w285 & w297 ) | ( w294 & w297 ) ;
  assign w2279 = w285 & ~w1942 ;
  assign w2280 = ~w1941 & w2279 ;
  assign w2281 = ( w294 & w297 ) | ( w294 & w2280 ) | ( w297 & w2280 ) ;
  assign w2282 = ( w285 & ~w290 ) | ( w285 & w2281 ) | ( ~w290 & w2281 ) ;
  assign w2283 = ( w290 & w2279 ) | ( w290 & w2281 ) | ( w2279 & w2281 ) ;
  assign w2284 = ( ~w2278 & w2282 ) | ( ~w2278 & w2283 ) | ( w2282 & w2283 ) ;
  assign w2285 = w300 & ~w1939 ;
  assign w2286 = ( w1917 & w1941 ) | ( w1917 & w2285 ) | ( w1941 & w2285 ) ;
  assign w2287 = w1911 | w2286 ;
  assign w2288 = ( w1942 & w2286 ) | ( w1942 & w2287 ) | ( w2286 & w2287 ) ;
  assign w2289 = w2285 | w2288 ;
  assign w2290 = w1923 | w2022 ;
  assign w2291 = ( ~w2022 & w2289 ) | ( ~w2022 & w2290 ) | ( w2289 & w2290 ) ;
  assign w2292 = w285 ^ w2291 ;
  assign w2293 = w2284 & w2292 ;
  assign w2294 = ~w300 & w1937 ;
  assign w2295 = w1911 & w1941 ;
  assign w2296 = ( w1937 & ~w2294 ) | ( w1937 & w2295 ) | ( ~w2294 & w2295 ) ;
  assign w2297 = w1917 | w1939 ;
  assign w2298 = w2035 & ~w2296 ;
  assign w2299 = ( w1923 & w2296 ) | ( w1923 & ~w2298 ) | ( w2296 & ~w2298 ) ;
  assign w2300 = ( ~w1939 & w2297 ) | ( ~w1939 & w2299 ) | ( w2297 & w2299 ) ;
  assign w2301 = w285 ^ w2300 ;
  assign w2302 = ( w2127 & w2293 ) | ( w2127 & w2301 ) | ( w2293 & w2301 ) ;
  assign w2303 = ( w2269 & w2277 ) | ( w2269 & w2302 ) | ( w2277 & w2302 ) ;
  assign w2304 = ( w2263 & w2264 ) | ( w2263 & w2303 ) | ( w2264 & w2303 ) ;
  assign w2305 = ( w2247 & w2255 ) | ( w2247 & w2304 ) | ( w2255 & w2304 ) ;
  assign w2306 = ( w2243 & w2245 ) | ( w2243 & w2305 ) | ( w2245 & w2305 ) ;
  assign w2307 = ( w2227 & w2235 ) | ( w2227 & w2306 ) | ( w2235 & w2306 ) ;
  assign w2308 = ( w2217 & w2225 ) | ( w2217 & w2307 ) | ( w2225 & w2307 ) ;
  assign w2309 = ( w2205 & w2215 ) | ( w2205 & w2308 ) | ( w2215 & w2308 ) ;
  assign w2310 = ( w2194 & w2203 ) | ( w2194 & w2309 ) | ( w2203 & w2309 ) ;
  assign w2311 = w1959 ^ w2310 ;
  assign w2312 = w2192 ^ w2311 ;
  assign w2313 = \pi01 ^ \pi02 ;
  assign w2314 = \pi00 & w2313 ;
  assign w2315 = \pi00 & ~w2313 ;
  assign w2316 = w330 & ~w763 ;
  assign w2317 = ~w492 & w2316 ;
  assign w2318 = ( w437 & ~w492 ) | ( w437 & w1612 ) | ( ~w492 & w1612 ) ;
  assign w2319 = w2317 & ~w2318 ;
  assign w2320 = ( ~w302 & w1706 ) | ( ~w302 & w1794 ) | ( w1706 & w1794 ) ;
  assign w2321 = ~w901 & w2319 ;
  assign w2322 = ( w302 & w511 ) | ( w302 & ~w901 ) | ( w511 & ~w901 ) ;
  assign w2323 = w2321 & ~w2322 ;
  assign w2324 = ~w2320 & w2323 ;
  assign w2325 = w220 | w266 ;
  assign w2326 = ( w220 & ~w244 ) | ( w220 & w2324 ) | ( ~w244 & w2324 ) ;
  assign w2327 = ~w2325 & w2326 ;
  assign w2328 = w305 | w342 ;
  assign w2329 = ( w133 & ~w305 ) | ( w133 & w332 ) | ( ~w305 & w332 ) ;
  assign w2330 = w2328 | w2329 ;
  assign w2331 = w421 | w1525 ;
  assign w2332 = ( w206 & ~w1525 ) | ( w206 & w2330 ) | ( ~w1525 & w2330 ) ;
  assign w2333 = w2331 | w2332 ;
  assign w2334 = ( w234 & w341 ) | ( w234 & ~w374 ) | ( w341 & ~w374 ) ;
  assign w2335 = w221 | w2333 ;
  assign w2336 = ( ~w221 & w374 ) | ( ~w221 & w453 ) | ( w374 & w453 ) ;
  assign w2337 = w2335 | w2336 ;
  assign w2338 = w2334 | w2337 ;
  assign w2339 = w58 | w1526 ;
  assign w2340 = ( ~w58 & w77 ) | ( ~w58 & w2338 ) | ( w77 & w2338 ) ;
  assign w2341 = w2339 | w2340 ;
  assign w2342 = ( w150 & w218 ) | ( w150 & ~w698 ) | ( w218 & ~w698 ) ;
  assign w2343 = w723 | w2341 ;
  assign w2344 = ( w698 & ~w723 ) | ( w698 & w1741 ) | ( ~w723 & w1741 ) ;
  assign w2345 = w2343 | w2344 ;
  assign w2346 = w2342 | w2345 ;
  assign w2347 = ( w173 & w183 ) | ( w173 & ~w228 ) | ( w183 & ~w228 ) ;
  assign w2348 = w141 | w2346 ;
  assign w2349 = ( ~w141 & w228 ) | ( ~w141 & w235 ) | ( w228 & w235 ) ;
  assign w2350 = w2348 | w2349 ;
  assign w2351 = w2347 | w2350 ;
  assign w2352 = w365 | w484 ;
  assign w2353 = ( ~w365 & w452 ) | ( ~w365 & w2351 ) | ( w452 & w2351 ) ;
  assign w2354 = w2352 | w2353 ;
  assign w2355 = w1907 & ~w2354 ;
  assign w2356 = w2327 & w2355 ;
  assign w2357 = w115 | w411 ;
  assign w2358 = w352 | w353 ;
  assign w2359 = w401 | w2358 ;
  assign w2360 = ( ~w401 & w428 ) | ( ~w401 & w1054 ) | ( w428 & w1054 ) ;
  assign w2361 = w2359 | w2360 ;
  assign w2362 = ( ~w320 & w459 ) | ( ~w320 & w509 ) | ( w459 & w509 ) ;
  assign w2363 = w492 | w2361 ;
  assign w2364 = ( w320 & w443 ) | ( w320 & ~w2361 ) | ( w443 & ~w2361 ) ;
  assign w2365 = w2363 | w2364 ;
  assign w2366 = w2362 | w2365 ;
  assign w2367 = ( w126 & ~w2357 ) | ( w126 & w2366 ) | ( ~w2357 & w2366 ) ;
  assign w2368 = w2357 | w2367 ;
  assign w2369 = w2356 ^ w2368 ;
  assign w2370 = \pi02 & ~w26 ;
  assign w2371 = w1907 ^ w2354 ;
  assign w2372 = w2327 ^ w2355 ;
  assign w2373 = w295 | w2372 ;
  assign w2374 = w2370 & w2371 ;
  assign w2375 = ( ~w2372 & w2373 ) | ( ~w2372 & w2374 ) | ( w2373 & w2374 ) ;
  assign w2376 = ( w1908 & ~w1915 ) | ( w1908 & w1954 ) | ( ~w1915 & w1954 ) ;
  assign w2377 = ( w1908 & w2371 ) | ( w1908 & w2376 ) | ( w2371 & w2376 ) ;
  assign w2378 = ( w2371 & ~w2372 ) | ( w2371 & w2377 ) | ( ~w2372 & w2377 ) ;
  assign w2379 = w2369 ^ w2378 ;
  assign w2380 = w2372 ^ w2379 ;
  assign w2381 = ~w2315 & w2369 ;
  assign w2382 = ~w2375 & w2380 ;
  assign w2383 = ( w2314 & w2375 ) | ( w2314 & ~w2382 ) | ( w2375 & ~w2382 ) ;
  assign w2384 = ( w2369 & ~w2381 ) | ( w2369 & w2383 ) | ( ~w2381 & w2383 ) ;
  assign w2385 = w297 ^ w2384 ;
  assign w2386 = w2203 ^ w2309 ;
  assign w2387 = w2194 ^ w2386 ;
  assign w2388 = w2315 & ~w2372 ;
  assign w2389 = ( w295 & w2371 ) | ( w295 & w2388 ) | ( w2371 & w2388 ) ;
  assign w2390 = w2370 | w2389 ;
  assign w2391 = ( w1908 & w2389 ) | ( w1908 & w2390 ) | ( w2389 & w2390 ) ;
  assign w2392 = w2388 | w2391 ;
  assign w2393 = w2372 ^ w2377 ;
  assign w2394 = w2371 ^ w2393 ;
  assign w2395 = w2314 & w2394 ;
  assign w2396 = ( w2314 & w2392 ) | ( w2314 & ~w2395 ) | ( w2392 & ~w2395 ) ;
  assign w2397 = w297 ^ w2396 ;
  assign w2398 = ~w295 & w1908 ;
  assign w2399 = ~w1915 & w2370 ;
  assign w2400 = ( w1908 & ~w2398 ) | ( w1908 & w2399 ) | ( ~w2398 & w2399 ) ;
  assign w2401 = w2371 ^ w2376 ;
  assign w2402 = w1908 ^ w2401 ;
  assign w2403 = ~w2315 & w2371 ;
  assign w2404 = w2400 | w2402 ;
  assign w2405 = ( w2314 & w2400 ) | ( w2314 & w2404 ) | ( w2400 & w2404 ) ;
  assign w2406 = ( w2371 & ~w2403 ) | ( w2371 & w2405 ) | ( ~w2403 & w2405 ) ;
  assign w2407 = w297 ^ w2406 ;
  assign w2408 = w1913 & w2315 ;
  assign w2409 = ( w295 & w1925 ) | ( w295 & w2408 ) | ( w1925 & w2408 ) ;
  assign w2410 = w2370 | w2409 ;
  assign w2411 = ( w1927 & w2409 ) | ( w1927 & w2410 ) | ( w2409 & w2410 ) ;
  assign w2412 = w2408 | w2411 ;
  assign w2413 = w1925 & w2315 ;
  assign w2414 = ( w295 & w1927 ) | ( w295 & w2413 ) | ( w1927 & w2413 ) ;
  assign w2415 = w2370 | w2414 ;
  assign w2416 = ( ~w1929 & w2414 ) | ( ~w1929 & w2415 ) | ( w2414 & w2415 ) ;
  assign w2417 = w2413 | w2416 ;
  assign w2418 = w1927 & w2315 ;
  assign w2419 = ( w295 & ~w1929 ) | ( w295 & w2418 ) | ( ~w1929 & w2418 ) ;
  assign w2420 = w2370 | w2419 ;
  assign w2421 = ( w1931 & w2419 ) | ( w1931 & w2420 ) | ( w2419 & w2420 ) ;
  assign w2422 = w2418 | w2421 ;
  assign w2423 = w1931 & w2315 ;
  assign w2424 = ( w295 & w1933 ) | ( w295 & w2423 ) | ( w1933 & w2423 ) ;
  assign w2425 = w2370 | w2424 ;
  assign w2426 = ( w1935 & w2424 ) | ( w1935 & w2425 ) | ( w2424 & w2425 ) ;
  assign w2427 = w2423 | w2426 ;
  assign w2428 = w1935 & w2315 ;
  assign w2429 = ( w295 & w1937 ) | ( w295 & w2428 ) | ( w1937 & w2428 ) ;
  assign w2430 = w2370 | w2429 ;
  assign w2431 = ( ~w1939 & w2429 ) | ( ~w1939 & w2430 ) | ( w2429 & w2430 ) ;
  assign w2432 = w2428 | w2431 ;
  assign w2433 = ~w1939 & w2315 ;
  assign w2434 = ( w295 & w1941 ) | ( w295 & w2433 ) | ( w1941 & w2433 ) ;
  assign w2435 = w2370 | w2434 ;
  assign w2436 = ( w1942 & w2434 ) | ( w1942 & w2435 ) | ( w2434 & w2435 ) ;
  assign w2437 = w2433 | w2436 ;
  assign w2438 = ~w295 & w1942 ;
  assign w2439 = w1941 & ~w2315 ;
  assign w2440 = ( w297 & ~w1941 ) | ( w297 & w2439 ) | ( ~w1941 & w2439 ) ;
  assign w2441 = ( ~w1942 & w2438 ) | ( ~w1942 & w2440 ) | ( w2438 & w2440 ) ;
  assign w2442 = ~w297 & w2441 ;
  assign w2443 = w1941 ^ w1942 ;
  assign w2444 = ( w2314 & w2442 ) | ( w2314 & w2443 ) | ( w2442 & w2443 ) ;
  assign w2445 = ( w2437 & w2441 ) | ( w2437 & w2444 ) | ( w2441 & w2444 ) ;
  assign w2446 = ( w2441 & w2442 ) | ( w2441 & ~w2445 ) | ( w2442 & ~w2445 ) ;
  assign w2447 = w297 | w2022 ;
  assign w2448 = ( w2022 & ~w2314 ) | ( w2022 & w2446 ) | ( ~w2314 & w2446 ) ;
  assign w2449 = ( w2446 & ~w2447 ) | ( w2446 & w2448 ) | ( ~w2447 & w2448 ) ;
  assign w2450 = \pi00 & w1942 ;
  assign w2451 = w2449 & ~w2450 ;
  assign w2452 = w1937 & ~w2315 ;
  assign w2453 = w1941 & w2370 ;
  assign w2454 = ( w1937 & ~w2452 ) | ( w1937 & w2453 ) | ( ~w2452 & w2453 ) ;
  assign w2455 = w295 | w1939 ;
  assign w2456 = w2035 & w2314 ;
  assign w2457 = ( w2314 & w2454 ) | ( w2314 & ~w2456 ) | ( w2454 & ~w2456 ) ;
  assign w2458 = ( ~w1939 & w2455 ) | ( ~w1939 & w2457 ) | ( w2455 & w2457 ) ;
  assign w2459 = w297 ^ w2458 ;
  assign w2460 = w298 & w1942 ;
  assign w2461 = ( w2451 & w2459 ) | ( w2451 & w2460 ) | ( w2459 & w2460 ) ;
  assign w2462 = w294 & w297 ;
  assign w2463 = w1942 ^ w2462 ;
  assign w2464 = ( w290 & w2462 ) | ( w290 & w2463 ) | ( w2462 & w2463 ) ;
  assign w2465 = ( w294 & w297 ) | ( w294 & w1941 ) | ( w297 & w1941 ) ;
  assign w2466 = w2464 ^ w2465 ;
  assign w2467 = w1993 | w2432 ;
  assign w2468 = ( w2314 & w2432 ) | ( w2314 & w2467 ) | ( w2432 & w2467 ) ;
  assign w2469 = w297 ^ w2468 ;
  assign w2470 = ( w2461 & w2466 ) | ( w2461 & w2469 ) | ( w2466 & w2469 ) ;
  assign w2471 = ~w295 & w1935 ;
  assign w2472 = w1937 & w2370 ;
  assign w2473 = ( w1935 & ~w2471 ) | ( w1935 & w2472 ) | ( ~w2471 & w2472 ) ;
  assign w2474 = w1933 & ~w2315 ;
  assign w2475 = w2047 & ~w2314 ;
  assign w2476 = ( w2047 & w2473 ) | ( w2047 & ~w2475 ) | ( w2473 & ~w2475 ) ;
  assign w2477 = ( w1933 & ~w2474 ) | ( w1933 & w2476 ) | ( ~w2474 & w2476 ) ;
  assign w2478 = w2284 ^ w2292 ;
  assign w2479 = w297 ^ w2477 ;
  assign w2480 = ( w2470 & w2478 ) | ( w2470 & w2479 ) | ( w2478 & w2479 ) ;
  assign w2481 = w2293 ^ w2301 ;
  assign w2482 = w2127 ^ w2481 ;
  assign w2483 = w2104 | w2427 ;
  assign w2484 = ( w2314 & w2427 ) | ( w2314 & w2483 ) | ( w2427 & w2483 ) ;
  assign w2485 = w297 ^ w2484 ;
  assign w2486 = ( w2480 & w2482 ) | ( w2480 & w2485 ) | ( w2482 & w2485 ) ;
  assign w2487 = ~w295 & w1931 ;
  assign w2488 = w1933 & w2370 ;
  assign w2489 = ( w1931 & ~w2487 ) | ( w1931 & w2488 ) | ( ~w2487 & w2488 ) ;
  assign w2490 = w1929 | w2315 ;
  assign w2491 = w2090 | w2314 ;
  assign w2492 = ( ~w2090 & w2489 ) | ( ~w2090 & w2491 ) | ( w2489 & w2491 ) ;
  assign w2493 = ( ~w1929 & w2490 ) | ( ~w1929 & w2492 ) | ( w2490 & w2492 ) ;
  assign w2494 = w297 ^ w2493 ;
  assign w2495 = w2277 ^ w2302 ;
  assign w2496 = w2269 ^ w2495 ;
  assign w2497 = ( w2486 & w2494 ) | ( w2486 & w2496 ) | ( w2494 & w2496 ) ;
  assign w2498 = w2263 ^ w2303 ;
  assign w2499 = w2264 ^ w2498 ;
  assign w2500 = w2079 & ~w2422 ;
  assign w2501 = ( w2314 & w2422 ) | ( w2314 & ~w2500 ) | ( w2422 & ~w2500 ) ;
  assign w2502 = w297 ^ w2501 ;
  assign w2503 = ( w2497 & w2499 ) | ( w2497 & w2502 ) | ( w2499 & w2502 ) ;
  assign w2504 = w2255 ^ w2304 ;
  assign w2505 = w2247 ^ w2504 ;
  assign w2506 = w2182 | w2417 ;
  assign w2507 = ( w2314 & w2417 ) | ( w2314 & w2506 ) | ( w2417 & w2506 ) ;
  assign w2508 = w297 ^ w2507 ;
  assign w2509 = ( w2503 & w2505 ) | ( w2503 & w2508 ) | ( w2505 & w2508 ) ;
  assign w2510 = w2243 ^ w2305 ;
  assign w2511 = w2245 ^ w2510 ;
  assign w2512 = w2212 | w2412 ;
  assign w2513 = ( w2314 & w2412 ) | ( w2314 & w2512 ) | ( w2412 & w2512 ) ;
  assign w2514 = w297 ^ w2513 ;
  assign w2515 = ( w2509 & w2511 ) | ( w2509 & w2514 ) | ( w2511 & w2514 ) ;
  assign w2516 = ~w295 & w1913 ;
  assign w2517 = w1925 & w2370 ;
  assign w2518 = ( w1913 & ~w2516 ) | ( w1913 & w2517 ) | ( ~w2516 & w2517 ) ;
  assign w2519 = w1915 | w2315 ;
  assign w2520 = w2200 & ~w2518 ;
  assign w2521 = ( w2314 & w2518 ) | ( w2314 & ~w2520 ) | ( w2518 & ~w2520 ) ;
  assign w2522 = ( ~w1915 & w2519 ) | ( ~w1915 & w2521 ) | ( w2519 & w2521 ) ;
  assign w2523 = w297 ^ w2522 ;
  assign w2524 = w2235 ^ w2306 ;
  assign w2525 = w2227 ^ w2524 ;
  assign w2526 = ( w2515 & w2523 ) | ( w2515 & w2525 ) | ( w2523 & w2525 ) ;
  assign w2527 = w295 | w1915 ;
  assign w2528 = w1913 & w2370 ;
  assign w2529 = ( ~w1915 & w2527 ) | ( ~w1915 & w2528 ) | ( w2527 & w2528 ) ;
  assign w2530 = w1908 & ~w2315 ;
  assign w2531 = w1956 & ~w2529 ;
  assign w2532 = ( w2314 & w2529 ) | ( w2314 & ~w2531 ) | ( w2529 & ~w2531 ) ;
  assign w2533 = ( w1908 & ~w2530 ) | ( w1908 & w2532 ) | ( ~w2530 & w2532 ) ;
  assign w2534 = w297 ^ w2533 ;
  assign w2535 = w2225 ^ w2307 ;
  assign w2536 = w2217 ^ w2535 ;
  assign w2537 = ( w2526 & w2534 ) | ( w2526 & w2536 ) | ( w2534 & w2536 ) ;
  assign w2538 = w2215 ^ w2308 ;
  assign w2539 = w2205 ^ w2538 ;
  assign w2540 = ( w2407 & w2537 ) | ( w2407 & w2539 ) | ( w2537 & w2539 ) ;
  assign w2541 = ( w2387 & w2397 ) | ( w2387 & w2540 ) | ( w2397 & w2540 ) ;
  assign w2542 = ( w2312 & w2385 ) | ( w2312 & w2541 ) | ( w2385 & w2541 ) ;
  assign w2543 = ( w1959 & w2192 ) | ( w1959 & w2310 ) | ( w2192 & w2310 ) ;
  assign w2544 = w300 & w2371 ;
  assign w2545 = ( w1908 & w1917 ) | ( w1908 & w2544 ) | ( w1917 & w2544 ) ;
  assign w2546 = w1911 | w2545 ;
  assign w2547 = ( ~w1915 & w2545 ) | ( ~w1915 & w2546 ) | ( w2545 & w2546 ) ;
  assign w2548 = w2544 | w2547 ;
  assign w2549 = ~w1923 & w2402 ;
  assign w2550 = ( w2402 & w2548 ) | ( w2402 & ~w2549 ) | ( w2548 & ~w2549 ) ;
  assign w2551 = w285 ^ w2550 ;
  assign w2552 = ( w2157 & w2180 ) | ( w2157 & w2190 ) | ( w2180 & w2190 ) ;
  assign w2553 = ( w2165 & w2177 ) | ( w2165 & w2178 ) | ( w2177 & w2178 ) ;
  assign w2554 = w1933 & w1983 ;
  assign w2555 = ( w1931 & w1985 ) | ( w1931 & w2554 ) | ( w1985 & w2554 ) ;
  assign w2556 = w1986 | w2555 ;
  assign w2557 = ( ~w1929 & w2555 ) | ( ~w1929 & w2556 ) | ( w2555 & w2556 ) ;
  assign w2558 = w2554 | w2557 ;
  assign w2559 = w1980 | w2090 ;
  assign w2560 = ( ~w2090 & w2558 ) | ( ~w2090 & w2559 ) | ( w2558 & w2559 ) ;
  assign w2561 = w660 ^ w2560 ;
  assign w2562 = w1937 & w1962 ;
  assign w2563 = ( ~w1939 & w2053 ) | ( ~w1939 & w2562 ) | ( w2053 & w2562 ) ;
  assign w2564 = w1964 | w2563 ;
  assign w2565 = ( w1935 & w2563 ) | ( w1935 & w2564 ) | ( w2563 & w2564 ) ;
  assign w2566 = w2562 | w2565 ;
  assign w2567 = ( w1965 & w1993 ) | ( w1965 & w2566 ) | ( w1993 & w2566 ) ;
  assign w2568 = w2566 | w2567 ;
  assign w2569 = w532 & ~w1941 ;
  assign w2570 = w2175 ^ w2569 ;
  assign w2571 = w2568 ^ w2570 ;
  assign w2572 = w2553 ^ w2561 ;
  assign w2573 = w2571 ^ w2572 ;
  assign w2574 = w1913 & w2067 ;
  assign w2575 = ( w1925 & w2072 ) | ( w1925 & w2574 ) | ( w2072 & w2574 ) ;
  assign w2576 = w2070 | w2575 ;
  assign w2577 = ( w1927 & w2575 ) | ( w1927 & w2576 ) | ( w2575 & w2576 ) ;
  assign w2578 = w2574 | w2577 ;
  assign w2579 = ~w2080 & w2212 ;
  assign w2580 = ( w2212 & w2578 ) | ( w2212 & ~w2579 ) | ( w2578 & ~w2579 ) ;
  assign w2581 = w943 ^ w2580 ;
  assign w2582 = w2552 ^ w2581 ;
  assign w2583 = w2573 ^ w2582 ;
  assign w2584 = w2543 ^ w2551 ;
  assign w2585 = w2583 ^ w2584 ;
  assign w2586 = ( ~w139 & w420 ) | ( ~w139 & w509 ) | ( w420 & w509 ) ;
  assign w2587 = w492 | w521 ;
  assign w2588 = ( w139 & w353 ) | ( w139 & ~w521 ) | ( w353 & ~w521 ) ;
  assign w2589 = w2587 | w2588 ;
  assign w2590 = w2586 | w2589 ;
  assign w2591 = w227 | w232 ;
  assign w2592 = w410 | w2591 ;
  assign w2593 = ( w188 & ~w410 ) | ( w188 & w2590 ) | ( ~w410 & w2590 ) ;
  assign w2594 = w2592 | w2593 ;
  assign w2595 = w2356 & ~w2368 ;
  assign w2596 = ~w2594 & w2595 ;
  assign w2597 = w2594 ^ w2595 ;
  assign w2598 = ~w295 & w2369 ;
  assign w2599 = w2370 & ~w2372 ;
  assign w2600 = ( w2369 & ~w2598 ) | ( w2369 & w2599 ) | ( ~w2598 & w2599 ) ;
  assign w2601 = ( w2369 & ~w2372 ) | ( w2369 & w2378 ) | ( ~w2372 & w2378 ) ;
  assign w2602 = w2597 ^ w2601 ;
  assign w2603 = w2369 ^ w2602 ;
  assign w2604 = ~w2315 & w2597 ;
  assign w2605 = w2600 | w2603 ;
  assign w2606 = ( w2314 & w2600 ) | ( w2314 & w2605 ) | ( w2600 & w2605 ) ;
  assign w2607 = ( w2597 & ~w2604 ) | ( w2597 & w2606 ) | ( ~w2604 & w2606 ) ;
  assign w2608 = w297 ^ w2607 ;
  assign w2609 = w2542 ^ w2608 ;
  assign w2610 = w2585 ^ w2609 ;
  assign w2611 = w513 | w690 ;
  assign w2612 = w148 | w2611 ;
  assign w2613 = ( w77 & ~w148 ) | ( w77 & w301 ) | ( ~w148 & w301 ) ;
  assign w2614 = w2612 | w2613 ;
  assign w2615 = ( w141 & w183 ) | ( w141 & ~w233 ) | ( w183 & ~w233 ) ;
  assign w2616 = w125 | w2614 ;
  assign w2617 = ( ~w125 & w233 ) | ( ~w125 & w304 ) | ( w233 & w304 ) ;
  assign w2618 = w2616 | w2617 ;
  assign w2619 = w2615 | w2618 ;
  assign w2620 = ( w114 & w128 ) | ( w114 & ~w319 ) | ( w128 & ~w319 ) ;
  assign w2621 = w58 | w2619 ;
  assign w2622 = ( ~w58 & w319 ) | ( ~w58 & w363 ) | ( w319 & w363 ) ;
  assign w2623 = w2621 | w2622 ;
  assign w2624 = w2620 | w2623 ;
  assign w2625 = ( w225 & ~w371 ) | ( w225 & w512 ) | ( ~w371 & w512 ) ;
  assign w2626 = w373 | w1020 ;
  assign w2627 = ( w371 & ~w373 ) | ( w371 & w374 ) | ( ~w373 & w374 ) ;
  assign w2628 = w2626 | w2627 ;
  assign w2629 = w2625 | w2628 ;
  assign w2630 = ( w451 & w478 ) | ( w451 & ~w502 ) | ( w478 & ~w502 ) ;
  assign w2631 = w263 | w2629 ;
  assign w2632 = ( ~w263 & w502 ) | ( ~w263 & w545 ) | ( w502 & w545 ) ;
  assign w2633 = w2631 | w2632 ;
  assign w2634 = w2630 | w2633 ;
  assign w2635 = w223 | w2634 ;
  assign w2636 = w422 | w744 ;
  assign w2637 = ( w303 & ~w744 ) | ( w303 & w2635 ) | ( ~w744 & w2635 ) ;
  assign w2638 = w2636 | w2637 ;
  assign w2639 = ( ~w123 & w905 ) | ( ~w123 & w1833 ) | ( w905 & w1833 ) ;
  assign w2640 = w2624 | w2638 ;
  assign w2641 = ( w123 & w262 ) | ( w123 & ~w2624 ) | ( w262 & ~w2624 ) ;
  assign w2642 = w2640 | w2641 ;
  assign w2643 = w2639 | w2642 ;
  assign w2644 = ( w302 & w333 ) | ( w302 & ~w341 ) | ( w333 & ~w341 ) ;
  assign w2645 = w134 | w2643 ;
  assign w2646 = ( ~w134 & w341 ) | ( ~w134 & w452 ) | ( w341 & w452 ) ;
  assign w2647 = w2645 | w2646 ;
  assign w2648 = w2644 | w2647 ;
  assign w2649 = w2385 ^ w2541 ;
  assign w2650 = w2312 ^ w2649 ;
  assign w2651 = ( w133 & w244 ) | ( w133 & ~w453 ) | ( w244 & ~w453 ) ;
  assign w2652 = w401 | w1673 ;
  assign w2653 = ( ~w401 & w453 ) | ( ~w401 & w544 ) | ( w453 & w544 ) ;
  assign w2654 = w2652 | w2653 ;
  assign w2655 = w2651 | w2654 ;
  assign w2656 = w360 | w510 ;
  assign w2657 = ( ~w360 & w484 ) | ( ~w360 & w2655 ) | ( w484 & w2655 ) ;
  assign w2658 = w2656 | w2657 ;
  assign w2659 = w149 | w347 ;
  assign w2660 = ( w123 & ~w347 ) | ( w123 & w767 ) | ( ~w347 & w767 ) ;
  assign w2661 = w2659 | w2660 ;
  assign w2662 = w374 | w455 ;
  assign w2663 = w301 | w2662 ;
  assign w2664 = ( ~w301 & w364 ) | ( ~w301 & w1811 ) | ( w364 & w1811 ) ;
  assign w2665 = w2663 | w2664 ;
  assign w2666 = ( ~w350 & w2661 ) | ( ~w350 & w2665 ) | ( w2661 & w2665 ) ;
  assign w2667 = w1739 | w2658 ;
  assign w2668 = ( w350 & w421 ) | ( w350 & ~w1739 ) | ( w421 & ~w1739 ) ;
  assign w2669 = w2667 | w2668 ;
  assign w2670 = w2666 | w2669 ;
  assign w2671 = ( w171 & w226 ) | ( w171 & ~w227 ) | ( w226 & ~w227 ) ;
  assign w2672 = w141 | w2670 ;
  assign w2673 = ( ~w141 & w227 ) | ( ~w141 & w322 ) | ( w227 & w322 ) ;
  assign w2674 = w2672 | w2673 ;
  assign w2675 = w2671 | w2674 ;
  assign w2676 = w307 & ~w2675 ;
  assign w2677 = w2397 ^ w2540 ;
  assign w2678 = w2387 ^ w2677 ;
  assign w2679 = ( w2675 & w2676 ) | ( w2675 & w2678 ) | ( w2676 & w2678 ) ;
  assign w2680 = ( ~w348 & w477 ) | ( ~w348 & w2648 ) | ( w477 & w2648 ) ;
  assign w2681 = w348 | w2680 ;
  assign w2682 = ( w2650 & w2679 ) | ( w2650 & w2681 ) | ( w2679 & w2681 ) ;
  assign w2683 = ( w279 & w2610 ) | ( w279 & w2682 ) | ( w2610 & w2682 ) ;
  assign w2684 = ( w244 & w245 ) | ( w244 & ~w354 ) | ( w245 & ~w354 ) ;
  assign w2685 = w94 | w183 ;
  assign w2686 = ( ~w183 & w354 ) | ( ~w183 & w581 ) | ( w354 & w581 ) ;
  assign w2687 = w2685 | w2686 ;
  assign w2688 = w2684 | w2687 ;
  assign w2689 = w451 | w476 ;
  assign w2690 = w215 | w2689 ;
  assign w2691 = ( ~w215 & w319 ) | ( ~w215 & w2688 ) | ( w319 & w2688 ) ;
  assign w2692 = w2690 | w2691 ;
  assign w2693 = ( w192 & w234 ) | ( w192 & ~w355 ) | ( w234 & ~w355 ) ;
  assign w2694 = ~w340 & w1051 ;
  assign w2695 = ( ~w340 & w355 ) | ( ~w340 & w475 ) | ( w355 & w475 ) ;
  assign w2696 = w2694 & ~w2695 ;
  assign w2697 = ~w2693 & w2696 ;
  assign w2698 = ( w174 & ~w230 ) | ( w174 & w1794 ) | ( ~w230 & w1794 ) ;
  assign w2699 = ~w2692 & w2697 ;
  assign w2700 = ( w230 & w322 ) | ( w230 & ~w2692 ) | ( w322 & ~w2692 ) ;
  assign w2701 = w2699 & ~w2700 ;
  assign w2702 = ~w2698 & w2701 ;
  assign w2703 = ( w219 & w226 ) | ( w219 & ~w231 ) | ( w226 & ~w231 ) ;
  assign w2704 = ~w113 & w2702 ;
  assign w2705 = ( ~w113 & w231 ) | ( ~w113 & w546 ) | ( w231 & w546 ) ;
  assign w2706 = w2704 & ~w2705 ;
  assign w2707 = ~w2703 & w2706 ;
  assign w2708 = w2596 ^ w2707 ;
  assign w2709 = ~w295 & w2597 ;
  assign w2710 = w2369 & w2370 ;
  assign w2711 = ( w2597 & ~w2709 ) | ( w2597 & w2710 ) | ( ~w2709 & w2710 ) ;
  assign w2712 = ( w2369 & w2597 ) | ( w2369 & w2601 ) | ( w2597 & w2601 ) ;
  assign w2713 = w2597 ^ w2708 ;
  assign w2714 = w2712 ^ w2713 ;
  assign w2715 = w2315 | w2708 ;
  assign w2716 = ~w2711 & w2714 ;
  assign w2717 = ( w2314 & w2711 ) | ( w2314 & ~w2716 ) | ( w2711 & ~w2716 ) ;
  assign w2718 = ( ~w2708 & w2715 ) | ( ~w2708 & w2717 ) | ( w2715 & w2717 ) ;
  assign w2719 = w297 ^ w2718 ;
  assign w2720 = ( w2543 & w2551 ) | ( w2543 & w2583 ) | ( w2551 & w2583 ) ;
  assign w2721 = ~w1915 & w2067 ;
  assign w2722 = ( w1913 & w2072 ) | ( w1913 & w2721 ) | ( w2072 & w2721 ) ;
  assign w2723 = w2070 | w2722 ;
  assign w2724 = ( w1925 & w2722 ) | ( w1925 & w2723 ) | ( w2722 & w2723 ) ;
  assign w2725 = w2721 | w2724 ;
  assign w2726 = w2080 | w2200 ;
  assign w2727 = ( ~w2200 & w2725 ) | ( ~w2200 & w2726 ) | ( w2725 & w2726 ) ;
  assign w2728 = w943 ^ w2727 ;
  assign w2729 = ( w2553 & w2561 ) | ( w2553 & w2571 ) | ( w2561 & w2571 ) ;
  assign w2730 = w532 & w1941 ;
  assign w2731 = w532 ^ w2568 ;
  assign w2732 = ( w2175 & w2730 ) | ( w2175 & w2731 ) | ( w2730 & w2731 ) ;
  assign w2733 = w1935 & w1962 ;
  assign w2734 = ( w1937 & w2053 ) | ( w1937 & w2733 ) | ( w2053 & w2733 ) ;
  assign w2735 = w1964 | w2734 ;
  assign w2736 = ( w1933 & w2734 ) | ( w1933 & w2735 ) | ( w2734 & w2735 ) ;
  assign w2737 = w2733 | w2736 ;
  assign w2738 = ( w1965 & w2047 ) | ( w1965 & w2737 ) | ( w2047 & w2737 ) ;
  assign w2739 = w2737 | w2738 ;
  assign w2740 = w532 & w1939 ;
  assign w2741 = w2732 ^ w2740 ;
  assign w2742 = w2739 ^ w2741 ;
  assign w2743 = w1931 & w1983 ;
  assign w2744 = ( ~w1929 & w1985 ) | ( ~w1929 & w2743 ) | ( w1985 & w2743 ) ;
  assign w2745 = w1986 | w2744 ;
  assign w2746 = ( w1927 & w2744 ) | ( w1927 & w2745 ) | ( w2744 & w2745 ) ;
  assign w2747 = w2743 | w2746 ;
  assign w2748 = w1980 | w2079 ;
  assign w2749 = ( ~w2079 & w2747 ) | ( ~w2079 & w2748 ) | ( w2747 & w2748 ) ;
  assign w2750 = w660 ^ w2749 ;
  assign w2751 = w2729 ^ w2750 ;
  assign w2752 = w2742 ^ w2751 ;
  assign w2753 = ( w2552 & w2573 ) | ( w2552 & w2581 ) | ( w2573 & w2581 ) ;
  assign w2754 = w2728 ^ w2753 ;
  assign w2755 = w2752 ^ w2754 ;
  assign w2756 = w300 & ~w2372 ;
  assign w2757 = ( w1917 & w2371 ) | ( w1917 & w2756 ) | ( w2371 & w2756 ) ;
  assign w2758 = w1911 | w2757 ;
  assign w2759 = ( w1908 & w2757 ) | ( w1908 & w2758 ) | ( w2757 & w2758 ) ;
  assign w2760 = w2756 | w2759 ;
  assign w2761 = w1923 | w2394 ;
  assign w2762 = ( ~w2394 & w2760 ) | ( ~w2394 & w2761 ) | ( w2760 & w2761 ) ;
  assign w2763 = w285 ^ w2762 ;
  assign w2764 = w2720 ^ w2763 ;
  assign w2765 = w2755 ^ w2764 ;
  assign w2766 = ( w2542 & w2585 ) | ( w2542 & w2608 ) | ( w2585 & w2608 ) ;
  assign w2767 = w2719 ^ w2766 ;
  assign w2768 = w2765 ^ w2767 ;
  assign w2769 = w452 | w545 ;
  assign w2770 = w244 | w2769 ;
  assign w2771 = ( w234 & ~w244 ) | ( w234 & w245 ) | ( ~w244 & w245 ) ;
  assign w2772 = w2770 | w2771 ;
  assign w2773 = ( ~w233 & w1184 ) | ( ~w233 & w2772 ) | ( w1184 & w2772 ) ;
  assign w2774 = w635 | w1682 ;
  assign w2775 = ( w233 & w304 ) | ( w233 & ~w635 ) | ( w304 & ~w635 ) ;
  assign w2776 = w2774 | w2775 ;
  assign w2777 = w2773 | w2776 ;
  assign w2778 = ( w139 & w218 ) | ( w139 & ~w263 ) | ( w218 & ~w263 ) ;
  assign w2779 = w615 | w2777 ;
  assign w2780 = ( w263 & w351 ) | ( w263 & ~w615 ) | ( w351 & ~w615 ) ;
  assign w2781 = w2779 | w2780 ;
  assign w2782 = w2778 | w2781 ;
  assign w2783 = w2683 ^ w2768 ;
  assign w2784 = w2782 ^ w2783 ;
  assign w2785 = w2610 ^ w2682 ;
  assign w2786 = w279 ^ w2785 ;
  assign w2787 = w2784 & w2786 ;
  assign w2788 = w2784 ^ w2786 ;
  assign w2789 = ( w2683 & w2768 ) | ( w2683 & w2782 ) | ( w2768 & w2782 ) ;
  assign w2790 = w242 | w243 ;
  assign w2791 = w707 | w2790 ;
  assign w2792 = ( w463 & ~w707 ) | ( w463 & w1811 ) | ( ~w707 & w1811 ) ;
  assign w2793 = w2791 | w2792 ;
  assign w2794 = w163 | w164 ;
  assign w2795 = w83 | w2794 ;
  assign w2796 = ( ~w83 & w161 ) | ( ~w83 & w2793 ) | ( w161 & w2793 ) ;
  assign w2797 = w2795 | w2796 ;
  assign w2798 = ( w77 & w245 ) | ( w77 & ~w321 ) | ( w245 & ~w321 ) ;
  assign w2799 = ~w769 & w1202 ;
  assign w2800 = ( w321 & w546 ) | ( w321 & w1202 ) | ( w546 & w1202 ) ;
  assign w2801 = w2799 & ~w2800 ;
  assign w2802 = ~w2798 & w2801 ;
  assign w2803 = ( ~w477 & w901 ) | ( ~w477 & w2797 ) | ( w901 & w2797 ) ;
  assign w2804 = ~w1810 & w2802 ;
  assign w2805 = ( w477 & w502 ) | ( w477 & w2802 ) | ( w502 & w2802 ) ;
  assign w2806 = w2804 & ~w2805 ;
  assign w2807 = ~w2803 & w2806 ;
  assign w2808 = w2596 & w2707 ;
  assign w2809 = ( w332 & w371 ) | ( w332 & w2807 ) | ( w371 & w2807 ) ;
  assign w2810 = w2807 & ~w2809 ;
  assign w2811 = w2808 ^ w2810 ;
  assign w2812 = w295 | w2708 ;
  assign w2813 = w2370 & w2597 ;
  assign w2814 = ( ~w2708 & w2812 ) | ( ~w2708 & w2813 ) | ( w2812 & w2813 ) ;
  assign w2815 = ( w2597 & ~w2708 ) | ( w2597 & w2712 ) | ( ~w2708 & w2712 ) ;
  assign w2816 = w2708 ^ w2815 ;
  assign w2817 = w2811 ^ w2816 ;
  assign w2818 = w2315 | w2811 ;
  assign w2819 = w2814 | w2817 ;
  assign w2820 = ( w2314 & w2814 ) | ( w2314 & w2819 ) | ( w2814 & w2819 ) ;
  assign w2821 = ( ~w2811 & w2818 ) | ( ~w2811 & w2820 ) | ( w2818 & w2820 ) ;
  assign w2822 = w297 ^ w2821 ;
  assign w2823 = ( w2720 & w2755 ) | ( w2720 & w2763 ) | ( w2755 & w2763 ) ;
  assign w2824 = w1908 & w2067 ;
  assign w2825 = ( ~w1915 & w2072 ) | ( ~w1915 & w2824 ) | ( w2072 & w2824 ) ;
  assign w2826 = w2070 | w2825 ;
  assign w2827 = ( w1913 & w2825 ) | ( w1913 & w2826 ) | ( w2825 & w2826 ) ;
  assign w2828 = w2824 | w2827 ;
  assign w2829 = w1956 | w2080 ;
  assign w2830 = ( ~w1956 & w2828 ) | ( ~w1956 & w2829 ) | ( w2828 & w2829 ) ;
  assign w2831 = w943 ^ w2830 ;
  assign w2832 = ( w2729 & w2742 ) | ( w2729 & w2750 ) | ( w2742 & w2750 ) ;
  assign w2833 = w532 & ~w1939 ;
  assign w2834 = w532 ^ w2739 ;
  assign w2835 = ( w2732 & w2833 ) | ( w2732 & w2834 ) | ( w2833 & w2834 ) ;
  assign w2836 = w1933 & w1962 ;
  assign w2837 = ( w1935 & w2053 ) | ( w1935 & w2836 ) | ( w2053 & w2836 ) ;
  assign w2838 = w1964 | w2837 ;
  assign w2839 = ( w1931 & w2837 ) | ( w1931 & w2838 ) | ( w2837 & w2838 ) ;
  assign w2840 = w2836 | w2839 ;
  assign w2841 = ( w1965 & w2104 ) | ( w1965 & w2840 ) | ( w2104 & w2840 ) ;
  assign w2842 = w2840 | w2841 ;
  assign w2843 = w532 & ~w1937 ;
  assign w2844 = w2835 ^ w2843 ;
  assign w2845 = w2842 ^ w2844 ;
  assign w2846 = ~w1929 & w1983 ;
  assign w2847 = ( w1927 & w1985 ) | ( w1927 & w2846 ) | ( w1985 & w2846 ) ;
  assign w2848 = w1986 | w2847 ;
  assign w2849 = ( w1925 & w2847 ) | ( w1925 & w2848 ) | ( w2847 & w2848 ) ;
  assign w2850 = w2846 | w2849 ;
  assign w2851 = ~w1980 & w2182 ;
  assign w2852 = ( w2182 & w2850 ) | ( w2182 & ~w2851 ) | ( w2850 & ~w2851 ) ;
  assign w2853 = w660 ^ w2852 ;
  assign w2854 = w2832 ^ w2853 ;
  assign w2855 = w2845 ^ w2854 ;
  assign w2856 = ( w2728 & w2752 ) | ( w2728 & w2753 ) | ( w2752 & w2753 ) ;
  assign w2857 = w2831 ^ w2856 ;
  assign w2858 = w2855 ^ w2857 ;
  assign w2859 = w300 & w2369 ;
  assign w2860 = ( w1917 & ~w2372 ) | ( w1917 & w2859 ) | ( ~w2372 & w2859 ) ;
  assign w2861 = w1911 | w2860 ;
  assign w2862 = ( w2371 & w2860 ) | ( w2371 & w2861 ) | ( w2860 & w2861 ) ;
  assign w2863 = w2859 | w2862 ;
  assign w2864 = w1923 | w2380 ;
  assign w2865 = ( ~w2380 & w2863 ) | ( ~w2380 & w2864 ) | ( w2863 & w2864 ) ;
  assign w2866 = w285 ^ w2865 ;
  assign w2867 = w2823 ^ w2866 ;
  assign w2868 = w2858 ^ w2867 ;
  assign w2869 = ( w2719 & w2765 ) | ( w2719 & w2766 ) | ( w2765 & w2766 ) ;
  assign w2870 = w2822 ^ w2869 ;
  assign w2871 = w2868 ^ w2870 ;
  assign w2872 = w266 | w411 ;
  assign w2873 = ( w126 & ~w266 ) | ( w126 & w365 ) | ( ~w266 & w365 ) ;
  assign w2874 = w2872 | w2873 ;
  assign w2875 = ( w629 & w707 ) | ( w629 & ~w1717 ) | ( w707 & ~w1717 ) ;
  assign w2876 = w257 | w1648 ;
  assign w2877 = ( ~w1648 & w1717 ) | ( ~w1648 & w2874 ) | ( w1717 & w2874 ) ;
  assign w2878 = w2876 | w2877 ;
  assign w2879 = w2875 | w2878 ;
  assign w2880 = ( w149 & ~w172 ) | ( w149 & w2330 ) | ( ~w172 & w2330 ) ;
  assign w2881 = w218 | w2879 ;
  assign w2882 = ( w172 & ~w218 ) | ( w172 & w333 ) | ( ~w218 & w333 ) ;
  assign w2883 = w2881 | w2882 ;
  assign w2884 = w2880 | w2883 ;
  assign w2885 = w83 | w451 ;
  assign w2886 = ( ~w83 & w191 ) | ( ~w83 & w2884 ) | ( w191 & w2884 ) ;
  assign w2887 = w2885 | w2886 ;
  assign w2888 = w2789 ^ w2871 ;
  assign w2889 = w2887 ^ w2888 ;
  assign w2890 = w2787 & w2889 ;
  assign w2891 = w2787 ^ w2889 ;
  assign w2892 = \pi22 ^ \pi23 ;
  assign w2893 = w2788 & w2892 ;
  assign w2894 = w2891 ^ w2893 ;
  assign w2895 = ( w2789 & w2871 ) | ( w2789 & w2887 ) | ( w2871 & w2887 ) ;
  assign w2896 = ( w141 & w236 ) | ( w141 & ~w351 ) | ( w236 & ~w351 ) ;
  assign w2897 = w108 | w128 ;
  assign w2898 = ( ~w128 & w351 ) | ( ~w128 & w412 ) | ( w351 & w412 ) ;
  assign w2899 = w2897 | w2898 ;
  assign w2900 = w2896 | w2899 ;
  assign w2901 = w113 | w2900 ;
  assign w2902 = w263 | w421 ;
  assign w2903 = w2901 | w2902 ;
  assign w2904 = ( w600 & w762 ) | ( w600 & ~w2901 ) | ( w762 & ~w2901 ) ;
  assign w2905 = w2903 | w2904 ;
  assign w2906 = ( w303 & w319 ) | ( w303 & ~w464 ) | ( w319 & ~w464 ) ;
  assign w2907 = w2658 | w2905 ;
  assign w2908 = ( w464 & w511 ) | ( w464 & ~w2905 ) | ( w511 & ~w2905 ) ;
  assign w2909 = w2907 | w2908 ;
  assign w2910 = w2906 | w2909 ;
  assign w2911 = w134 | w513 ;
  assign w2912 = ( ~w134 & w332 ) | ( ~w134 & w2910 ) | ( w332 & w2910 ) ;
  assign w2913 = w2911 | w2912 ;
  assign w2914 = ( w2822 & w2868 ) | ( w2822 & w2869 ) | ( w2868 & w2869 ) ;
  assign w2915 = w2370 | w2708 ;
  assign w2916 = w295 & ~w2811 ;
  assign w2917 = ( ~w2708 & w2915 ) | ( ~w2708 & w2916 ) | ( w2915 & w2916 ) ;
  assign w2918 = ( w2708 & w2811 ) | ( w2708 & ~w2815 ) | ( w2811 & ~w2815 ) ;
  assign w2919 = w2811 | w2918 ;
  assign w2920 = w2314 | w2917 ;
  assign w2921 = w2811 ^ w2918 ;
  assign w2922 = ( w2917 & w2920 ) | ( w2917 & w2921 ) | ( w2920 & w2921 ) ;
  assign w2923 = w297 ^ w2922 ;
  assign w2924 = ( w2823 & w2858 ) | ( w2823 & w2866 ) | ( w2858 & w2866 ) ;
  assign w2925 = w2067 & w2371 ;
  assign w2926 = ( w1908 & w2072 ) | ( w1908 & w2925 ) | ( w2072 & w2925 ) ;
  assign w2927 = w2070 | w2926 ;
  assign w2928 = ( ~w1915 & w2926 ) | ( ~w1915 & w2927 ) | ( w2926 & w2927 ) ;
  assign w2929 = w2925 | w2928 ;
  assign w2930 = ~w2080 & w2402 ;
  assign w2931 = ( w2402 & w2929 ) | ( w2402 & ~w2930 ) | ( w2929 & ~w2930 ) ;
  assign w2932 = w943 ^ w2931 ;
  assign w2933 = ( w2832 & w2845 ) | ( w2832 & w2853 ) | ( w2845 & w2853 ) ;
  assign w2934 = w532 & w1937 ;
  assign w2935 = w532 ^ w2842 ;
  assign w2936 = ( w2835 & w2934 ) | ( w2835 & w2935 ) | ( w2934 & w2935 ) ;
  assign w2937 = w1931 & w1962 ;
  assign w2938 = ( w1933 & w2053 ) | ( w1933 & w2937 ) | ( w2053 & w2937 ) ;
  assign w2939 = w1964 | w2938 ;
  assign w2940 = ( ~w1929 & w2938 ) | ( ~w1929 & w2939 ) | ( w2938 & w2939 ) ;
  assign w2941 = w2937 | w2940 ;
  assign w2942 = ( w1965 & ~w2090 ) | ( w1965 & w2941 ) | ( ~w2090 & w2941 ) ;
  assign w2943 = w2941 | w2942 ;
  assign w2944 = w532 & ~w1935 ;
  assign w2945 = w2936 ^ w2944 ;
  assign w2946 = w2943 ^ w2945 ;
  assign w2947 = w1927 & w1983 ;
  assign w2948 = ( w1925 & w1985 ) | ( w1925 & w2947 ) | ( w1985 & w2947 ) ;
  assign w2949 = w1986 | w2948 ;
  assign w2950 = ( w1913 & w2948 ) | ( w1913 & w2949 ) | ( w2948 & w2949 ) ;
  assign w2951 = w2947 | w2950 ;
  assign w2952 = ~w1980 & w2212 ;
  assign w2953 = ( w2212 & w2951 ) | ( w2212 & ~w2952 ) | ( w2951 & ~w2952 ) ;
  assign w2954 = w660 ^ w2953 ;
  assign w2955 = w2933 ^ w2954 ;
  assign w2956 = w2946 ^ w2955 ;
  assign w2957 = ( w2831 & w2855 ) | ( w2831 & w2856 ) | ( w2855 & w2856 ) ;
  assign w2958 = w2932 ^ w2957 ;
  assign w2959 = w2956 ^ w2958 ;
  assign w2960 = w300 & w2597 ;
  assign w2961 = ( w1917 & w2369 ) | ( w1917 & w2960 ) | ( w2369 & w2960 ) ;
  assign w2962 = w1911 | w2961 ;
  assign w2963 = ( ~w2372 & w2961 ) | ( ~w2372 & w2962 ) | ( w2961 & w2962 ) ;
  assign w2964 = w2960 | w2963 ;
  assign w2965 = ~w1923 & w2603 ;
  assign w2966 = ( w2603 & w2964 ) | ( w2603 & ~w2965 ) | ( w2964 & ~w2965 ) ;
  assign w2967 = w285 ^ w2966 ;
  assign w2968 = w2924 ^ w2967 ;
  assign w2969 = w2959 ^ w2968 ;
  assign w2970 = w2914 ^ w2969 ;
  assign w2971 = w2923 ^ w2970 ;
  assign w2972 = ( w2895 & w2913 ) | ( w2895 & w2971 ) | ( w2913 & w2971 ) ;
  assign w2973 = w2895 ^ w2971 ;
  assign w2974 = w2913 ^ w2973 ;
  assign w2975 = w2890 & w2974 ;
  assign w2976 = w2890 ^ w2974 ;
  assign w2977 = w2788 | w2891 ;
  assign w2978 = w2892 & w2977 ;
  assign w2979 = w2976 ^ w2978 ;
  assign w2980 = ( w401 & w868 ) | ( w401 & ~w1717 ) | ( w868 & ~w1717 ) ;
  assign w2981 = w1194 | w1558 ;
  assign w2982 = ( ~w1558 & w1717 ) | ( ~w1558 & w2614 ) | ( w1717 & w2614 ) ;
  assign w2983 = w2981 | w2982 ;
  assign w2984 = w2980 | w2983 ;
  assign w2985 = ( w172 & ~w322 ) | ( w172 & w359 ) | ( ~w322 & w359 ) ;
  assign w2986 = w689 | w2984 ;
  assign w2987 = ( w322 & w374 ) | ( w322 & ~w689 ) | ( w374 & ~w689 ) ;
  assign w2988 = w2986 | w2987 ;
  assign w2989 = w2985 | w2988 ;
  assign w2990 = w71 | w266 ;
  assign w2991 = ( ~w71 & w245 ) | ( ~w71 & w2989 ) | ( w245 & w2989 ) ;
  assign w2992 = w2990 | w2991 ;
  assign w2993 = ( w2914 & w2923 ) | ( w2914 & w2969 ) | ( w2923 & w2969 ) ;
  assign w2994 = ( w2924 & w2959 ) | ( w2924 & w2967 ) | ( w2959 & w2967 ) ;
  assign w2995 = w2370 & ~w2811 ;
  assign w2996 = w2314 | w2995 ;
  assign w2997 = ( ~w2919 & w2995 ) | ( ~w2919 & w2996 ) | ( w2995 & w2996 ) ;
  assign w2998 = w297 ^ w2997 ;
  assign w2999 = w2067 & ~w2372 ;
  assign w3000 = ( w2072 & w2371 ) | ( w2072 & w2999 ) | ( w2371 & w2999 ) ;
  assign w3001 = w2070 | w3000 ;
  assign w3002 = ( w1908 & w3000 ) | ( w1908 & w3001 ) | ( w3000 & w3001 ) ;
  assign w3003 = w2999 | w3002 ;
  assign w3004 = w2080 | w2394 ;
  assign w3005 = ( ~w2394 & w3003 ) | ( ~w2394 & w3004 ) | ( w3003 & w3004 ) ;
  assign w3006 = w943 ^ w3005 ;
  assign w3007 = ( w2933 & w2946 ) | ( w2933 & w2954 ) | ( w2946 & w2954 ) ;
  assign w3008 = w532 & w1935 ;
  assign w3009 = w532 ^ w2943 ;
  assign w3010 = ( w2936 & w3008 ) | ( w2936 & w3009 ) | ( w3008 & w3009 ) ;
  assign w3011 = ~w1929 & w1962 ;
  assign w3012 = ( w1931 & w2053 ) | ( w1931 & w3011 ) | ( w2053 & w3011 ) ;
  assign w3013 = w1964 | w3012 ;
  assign w3014 = ( w1927 & w3012 ) | ( w1927 & w3013 ) | ( w3012 & w3013 ) ;
  assign w3015 = w3011 | w3014 ;
  assign w3016 = ( w1965 & ~w2079 ) | ( w1965 & w3015 ) | ( ~w2079 & w3015 ) ;
  assign w3017 = w3015 | w3016 ;
  assign w3018 = w532 & ~w1933 ;
  assign w3019 = w3010 ^ w3018 ;
  assign w3020 = w3017 ^ w3019 ;
  assign w3021 = w1925 & w1983 ;
  assign w3022 = ( w1913 & w1985 ) | ( w1913 & w3021 ) | ( w1985 & w3021 ) ;
  assign w3023 = w1986 | w3022 ;
  assign w3024 = ( ~w1915 & w3022 ) | ( ~w1915 & w3023 ) | ( w3022 & w3023 ) ;
  assign w3025 = w3021 | w3024 ;
  assign w3026 = w1980 | w2200 ;
  assign w3027 = ( ~w2200 & w3025 ) | ( ~w2200 & w3026 ) | ( w3025 & w3026 ) ;
  assign w3028 = w660 ^ w3027 ;
  assign w3029 = w3007 ^ w3028 ;
  assign w3030 = w3020 ^ w3029 ;
  assign w3031 = ( w2932 & w2956 ) | ( w2932 & w2957 ) | ( w2956 & w2957 ) ;
  assign w3032 = w3006 ^ w3031 ;
  assign w3033 = w3030 ^ w3032 ;
  assign w3034 = w300 & ~w2708 ;
  assign w3035 = ( w1917 & w2597 ) | ( w1917 & w3034 ) | ( w2597 & w3034 ) ;
  assign w3036 = w1911 | w3035 ;
  assign w3037 = ( w2369 & w3035 ) | ( w2369 & w3036 ) | ( w3035 & w3036 ) ;
  assign w3038 = w3034 | w3037 ;
  assign w3039 = w1923 | w2714 ;
  assign w3040 = ( ~w2714 & w3038 ) | ( ~w2714 & w3039 ) | ( w3038 & w3039 ) ;
  assign w3041 = w285 ^ w3040 ;
  assign w3042 = w2998 ^ w3041 ;
  assign w3043 = w3033 ^ w3042 ;
  assign w3044 = w2993 ^ w3043 ;
  assign w3045 = w2994 ^ w3044 ;
  assign w3046 = w2972 ^ w3045 ;
  assign w3047 = w2992 ^ w3046 ;
  assign w3048 = w2975 & w3047 ;
  assign w3049 = w2975 ^ w3047 ;
  assign w3050 = w2976 | w2977 ;
  assign w3051 = w2892 & w3050 ;
  assign w3052 = w3049 ^ w3051 ;
  assign w3053 = ( w2972 & w2992 ) | ( w2972 & w3045 ) | ( w2992 & w3045 ) ;
  assign w3054 = w341 | w351 ;
  assign w3055 = w83 | w3054 ;
  assign w3056 = ( ~w83 & w141 ) | ( ~w83 & w306 ) | ( w141 & w306 ) ;
  assign w3057 = w3055 | w3056 ;
  assign w3058 = ( ~w636 & w900 ) | ( ~w636 & w3057 ) | ( w900 & w3057 ) ;
  assign w3059 = w706 | w1843 ;
  assign w3060 = ( w636 & w1794 ) | ( w636 & ~w1843 ) | ( w1794 & ~w1843 ) ;
  assign w3061 = w3059 | w3060 ;
  assign w3062 = w3058 | w3061 ;
  assign w3063 = w175 | w581 ;
  assign w3064 = ( ~w175 & w197 ) | ( ~w175 & w3062 ) | ( w197 & w3062 ) ;
  assign w3065 = w3063 | w3064 ;
  assign w3066 = ( w2993 & w2994 ) | ( w2993 & w3043 ) | ( w2994 & w3043 ) ;
  assign w3067 = ( w2998 & w3033 ) | ( w2998 & w3041 ) | ( w3033 & w3041 ) ;
  assign w3068 = ( w3006 & w3030 ) | ( w3006 & w3031 ) | ( w3030 & w3031 ) ;
  assign w3069 = ( w3007 & w3020 ) | ( w3007 & w3028 ) | ( w3020 & w3028 ) ;
  assign w3070 = w1927 & w1962 ;
  assign w3071 = ( ~w1929 & w2053 ) | ( ~w1929 & w3070 ) | ( w2053 & w3070 ) ;
  assign w3072 = w1964 | w3071 ;
  assign w3073 = ( w1925 & w3071 ) | ( w1925 & w3072 ) | ( w3071 & w3072 ) ;
  assign w3074 = w3070 | w3073 ;
  assign w3075 = ~w1965 & w2182 ;
  assign w3076 = ( w2182 & w3074 ) | ( w2182 & ~w3075 ) | ( w3074 & ~w3075 ) ;
  assign w3077 = w532 ^ w3076 ;
  assign w3078 = w532 & w1931 ;
  assign w3079 = w297 ^ w3078 ;
  assign w3080 = w3077 ^ w3079 ;
  assign w3081 = w532 & w1933 ;
  assign w3082 = w532 ^ w3017 ;
  assign w3083 = ( w3010 & w3081 ) | ( w3010 & w3082 ) | ( w3081 & w3082 ) ;
  assign w3084 = w1913 & w1983 ;
  assign w3085 = ( ~w1915 & w1985 ) | ( ~w1915 & w3084 ) | ( w1985 & w3084 ) ;
  assign w3086 = w1986 | w3085 ;
  assign w3087 = ( w1908 & w3085 ) | ( w1908 & w3086 ) | ( w3085 & w3086 ) ;
  assign w3088 = w3084 | w3087 ;
  assign w3089 = w1956 | w1980 ;
  assign w3090 = ( ~w1956 & w3088 ) | ( ~w1956 & w3089 ) | ( w3088 & w3089 ) ;
  assign w3091 = w660 ^ w3090 ;
  assign w3092 = w3080 ^ w3091 ;
  assign w3093 = w3083 ^ w3092 ;
  assign w3094 = w2067 & w2369 ;
  assign w3095 = ( w2072 & ~w2372 ) | ( w2072 & w3094 ) | ( ~w2372 & w3094 ) ;
  assign w3096 = w2070 | w3095 ;
  assign w3097 = ( w2371 & w3095 ) | ( w2371 & w3096 ) | ( w3095 & w3096 ) ;
  assign w3098 = w3094 | w3097 ;
  assign w3099 = w2080 | w2380 ;
  assign w3100 = ( ~w2380 & w3098 ) | ( ~w2380 & w3099 ) | ( w3098 & w3099 ) ;
  assign w3101 = w943 ^ w3100 ;
  assign w3102 = w3069 ^ w3101 ;
  assign w3103 = w3093 ^ w3102 ;
  assign w3104 = w300 & ~w2811 ;
  assign w3105 = ( w1917 & ~w2708 ) | ( w1917 & w3104 ) | ( ~w2708 & w3104 ) ;
  assign w3106 = w1911 | w3105 ;
  assign w3107 = ( w2597 & w3105 ) | ( w2597 & w3106 ) | ( w3105 & w3106 ) ;
  assign w3108 = w3104 | w3107 ;
  assign w3109 = ~w1923 & w2817 ;
  assign w3110 = ( w2817 & w3108 ) | ( w2817 & ~w3109 ) | ( w3108 & ~w3109 ) ;
  assign w3111 = w285 ^ w3110 ;
  assign w3112 = w3068 ^ w3111 ;
  assign w3113 = w3103 ^ w3112 ;
  assign w3114 = w3066 ^ w3067 ;
  assign w3115 = w3113 ^ w3114 ;
  assign w3116 = w3053 ^ w3115 ;
  assign w3117 = w3065 ^ w3116 ;
  assign w3118 = w3048 & w3117 ;
  assign w3119 = w3048 ^ w3117 ;
  assign w3120 = w3049 | w3050 ;
  assign w3121 = w2892 & w3120 ;
  assign w3122 = w3119 ^ w3121 ;
  assign w3123 = ( w3053 & w3065 ) | ( w3053 & w3115 ) | ( w3065 & w3115 ) ;
  assign w3124 = ( w322 & ~w363 ) | ( w322 & w479 ) | ( ~w363 & w479 ) ;
  assign w3125 = w363 | w3124 ;
  assign w3126 = w172 | w3125 ;
  assign w3127 = ( w94 & w189 ) | ( w94 & ~w3125 ) | ( w189 & ~w3125 ) ;
  assign w3128 = w3126 | w3127 ;
  assign w3129 = ( w320 & ~w1688 ) | ( w320 & w3128 ) | ( ~w1688 & w3128 ) ;
  assign w3130 = w2341 | w2797 ;
  assign w3131 = ( w1688 & ~w2797 ) | ( w1688 & w2874 ) | ( ~w2797 & w2874 ) ;
  assign w3132 = w3130 | w3131 ;
  assign w3133 = w3129 | w3132 ;
  assign w3134 = ( w175 & w244 ) | ( w175 & ~w304 ) | ( w244 & ~w304 ) ;
  assign w3135 = w373 | w3133 ;
  assign w3136 = ( w304 & ~w373 ) | ( w304 & w422 ) | ( ~w373 & w422 ) ;
  assign w3137 = w3135 | w3136 ;
  assign w3138 = w3134 | w3137 ;
  assign w3139 = ( w3066 & w3067 ) | ( w3066 & w3113 ) | ( w3067 & w3113 ) ;
  assign w3140 = ( w3068 & w3103 ) | ( w3068 & w3111 ) | ( w3103 & w3111 ) ;
  assign w3141 = ( w3069 & w3093 ) | ( w3069 & w3101 ) | ( w3093 & w3101 ) ;
  assign w3142 = w2067 & w2597 ;
  assign w3143 = ( w2072 & w2369 ) | ( w2072 & w3142 ) | ( w2369 & w3142 ) ;
  assign w3144 = w2070 | w3143 ;
  assign w3145 = ( ~w2372 & w3143 ) | ( ~w2372 & w3144 ) | ( w3143 & w3144 ) ;
  assign w3146 = w3142 | w3145 ;
  assign w3147 = ~w2080 & w2603 ;
  assign w3148 = ( w2603 & w3146 ) | ( w2603 & ~w3147 ) | ( w3146 & ~w3147 ) ;
  assign w3149 = w943 ^ w3148 ;
  assign w3150 = ( w3080 & w3083 ) | ( w3080 & w3091 ) | ( w3083 & w3091 ) ;
  assign w3151 = ( w297 & w3077 ) | ( w297 & w3078 ) | ( w3077 & w3078 ) ;
  assign w3152 = w532 & ~w1929 ;
  assign w3153 = w297 ^ w3152 ;
  assign w3154 = w3151 ^ w3153 ;
  assign w3155 = w1925 & w1962 ;
  assign w3156 = ( w1927 & w2053 ) | ( w1927 & w3155 ) | ( w2053 & w3155 ) ;
  assign w3157 = w1964 | w3156 ;
  assign w3158 = ( w1913 & w3156 ) | ( w1913 & w3157 ) | ( w3156 & w3157 ) ;
  assign w3159 = w3155 | w3158 ;
  assign w3160 = ~w1965 & w2212 ;
  assign w3161 = ( w2212 & w3159 ) | ( w2212 & ~w3160 ) | ( w3159 & ~w3160 ) ;
  assign w3162 = w532 ^ w3161 ;
  assign w3163 = ~w1915 & w1983 ;
  assign w3164 = ( w1908 & w1985 ) | ( w1908 & w3163 ) | ( w1985 & w3163 ) ;
  assign w3165 = w1986 | w3164 ;
  assign w3166 = ( w2371 & w3164 ) | ( w2371 & w3165 ) | ( w3164 & w3165 ) ;
  assign w3167 = w3163 | w3166 ;
  assign w3168 = ~w1980 & w2402 ;
  assign w3169 = ( w2402 & w3167 ) | ( w2402 & ~w3168 ) | ( w3167 & ~w3168 ) ;
  assign w3170 = w660 ^ w3169 ;
  assign w3171 = w3154 ^ w3170 ;
  assign w3172 = w3162 ^ w3171 ;
  assign w3173 = w3149 ^ w3172 ;
  assign w3174 = w3150 ^ w3173 ;
  assign w3175 = w1917 & ~w2811 ;
  assign w3176 = ( w1911 & ~w2708 ) | ( w1911 & w3175 ) | ( ~w2708 & w3175 ) ;
  assign w3177 = ( w2708 & w2815 ) | ( w2708 & ~w3176 ) | ( w2815 & ~w3176 ) ;
  assign w3178 = ( w1923 & w2811 ) | ( w1923 & ~w2815 ) | ( w2811 & ~w2815 ) ;
  assign w3179 = ( w3175 & w3177 ) | ( w3175 & w3178 ) | ( w3177 & w3178 ) ;
  assign w3180 = w2708 & w2811 ;
  assign w3181 = ( w3176 & w3179 ) | ( w3176 & ~w3180 ) | ( w3179 & ~w3180 ) ;
  assign w3182 = w285 ^ w3141 ;
  assign w3183 = w3174 ^ w3182 ;
  assign w3184 = w3181 ^ w3183 ;
  assign w3185 = w3139 ^ w3140 ;
  assign w3186 = w3184 ^ w3185 ;
  assign w3187 = w3123 ^ w3186 ;
  assign w3188 = w3138 ^ w3187 ;
  assign w3189 = w3118 & w3188 ;
  assign w3190 = w3118 ^ w3188 ;
  assign w3191 = w3119 | w3120 ;
  assign w3192 = w2892 & w3191 ;
  assign w3193 = w3190 ^ w3192 ;
  assign w3194 = ( w3123 & w3138 ) | ( w3123 & w3186 ) | ( w3138 & w3186 ) ;
  assign w3195 = ( w77 & w126 ) | ( w77 & ~w321 ) | ( w126 & ~w321 ) ;
  assign w3196 = w578 | w1797 ;
  assign w3197 = ( w321 & w342 ) | ( w321 & ~w578 ) | ( w342 & ~w578 ) ;
  assign w3198 = w3196 | w3197 ;
  assign w3199 = w3195 | w3198 ;
  assign w3200 = ( w373 & w901 ) | ( w373 & ~w1717 ) | ( w901 & ~w1717 ) ;
  assign w3201 = w150 | w3199 ;
  assign w3202 = ( ~w150 & w361 ) | ( ~w150 & w1717 ) | ( w361 & w1717 ) ;
  assign w3203 = w3201 | w3202 ;
  assign w3204 = w3200 | w3203 ;
  assign w3205 = ( w895 & w1837 ) | ( w895 & ~w2357 ) | ( w1837 & ~w2357 ) ;
  assign w3206 = w261 | w3204 ;
  assign w3207 = ( w343 & w2357 ) | ( w343 & ~w3204 ) | ( w2357 & ~w3204 ) ;
  assign w3208 = w3206 | w3207 ;
  assign w3209 = w3205 | w3208 ;
  assign w3210 = ( w141 & w164 ) | ( w141 & ~w169 ) | ( w164 & ~w169 ) ;
  assign w3211 = w139 | w3209 ;
  assign w3212 = ( ~w139 & w169 ) | ( ~w139 & w453 ) | ( w169 & w453 ) ;
  assign w3213 = w3211 | w3212 ;
  assign w3214 = w3210 | w3213 ;
  assign w3215 = ( w3139 & w3140 ) | ( w3139 & w3184 ) | ( w3140 & w3184 ) ;
  assign w3216 = w285 ^ w3181 ;
  assign w3217 = ( w3141 & w3174 ) | ( w3141 & w3216 ) | ( w3174 & w3216 ) ;
  assign w3218 = ( w3149 & w3150 ) | ( w3149 & w3172 ) | ( w3150 & w3172 ) ;
  assign w3219 = w1911 & ~w2811 ;
  assign w3220 = w1923 | w3219 ;
  assign w3221 = ( ~w2919 & w3219 ) | ( ~w2919 & w3220 ) | ( w3219 & w3220 ) ;
  assign w3222 = w285 ^ w3221 ;
  assign w3223 = w2067 & ~w2708 ;
  assign w3224 = ( w2072 & w2597 ) | ( w2072 & w3223 ) | ( w2597 & w3223 ) ;
  assign w3225 = w2070 | w3224 ;
  assign w3226 = ( w2369 & w3224 ) | ( w2369 & w3225 ) | ( w3224 & w3225 ) ;
  assign w3227 = w3223 | w3226 ;
  assign w3228 = w2080 | w2714 ;
  assign w3229 = ( ~w2714 & w3227 ) | ( ~w2714 & w3228 ) | ( w3227 & w3228 ) ;
  assign w3230 = w943 ^ w3229 ;
  assign w3231 = ( w3154 & w3162 ) | ( w3154 & w3170 ) | ( w3162 & w3170 ) ;
  assign w3232 = ( w297 & w3151 ) | ( w297 & w3152 ) | ( w3151 & w3152 ) ;
  assign w3233 = w532 & w1927 ;
  assign w3234 = w297 ^ w3233 ;
  assign w3235 = w3232 ^ w3234 ;
  assign w3236 = w1913 & w1962 ;
  assign w3237 = ( w1925 & w2053 ) | ( w1925 & w3236 ) | ( w2053 & w3236 ) ;
  assign w3238 = w1964 | w3237 ;
  assign w3239 = ( ~w1915 & w3237 ) | ( ~w1915 & w3238 ) | ( w3237 & w3238 ) ;
  assign w3240 = w3236 | w3239 ;
  assign w3241 = w1965 | w2200 ;
  assign w3242 = ( ~w2200 & w3240 ) | ( ~w2200 & w3241 ) | ( w3240 & w3241 ) ;
  assign w3243 = w532 ^ w3242 ;
  assign w3244 = w1908 & w1983 ;
  assign w3245 = ( w1985 & w2371 ) | ( w1985 & w3244 ) | ( w2371 & w3244 ) ;
  assign w3246 = w1986 | w3245 ;
  assign w3247 = ( ~w2372 & w3245 ) | ( ~w2372 & w3246 ) | ( w3245 & w3246 ) ;
  assign w3248 = w3244 | w3247 ;
  assign w3249 = w1980 | w2394 ;
  assign w3250 = ( ~w2394 & w3248 ) | ( ~w2394 & w3249 ) | ( w3248 & w3249 ) ;
  assign w3251 = w660 ^ w3250 ;
  assign w3252 = w3235 ^ w3251 ;
  assign w3253 = w3243 ^ w3252 ;
  assign w3254 = w3230 ^ w3253 ;
  assign w3255 = w3231 ^ w3254 ;
  assign w3256 = w3222 ^ w3255 ;
  assign w3257 = w3218 ^ w3256 ;
  assign w3258 = w3215 ^ w3257 ;
  assign w3259 = w3217 ^ w3258 ;
  assign w3260 = w3194 ^ w3259 ;
  assign w3261 = w3214 ^ w3260 ;
  assign w3262 = w3189 & w3261 ;
  assign w3263 = w3189 ^ w3261 ;
  assign w3264 = w3190 | w3191 ;
  assign w3265 = w2892 & w3264 ;
  assign w3266 = w3263 ^ w3265 ;
  assign w3267 = ( w3194 & w3214 ) | ( w3194 & w3259 ) | ( w3214 & w3259 ) ;
  assign w3268 = ( w3218 & w3222 ) | ( w3218 & w3255 ) | ( w3222 & w3255 ) ;
  assign w3269 = ( w3230 & w3231 ) | ( w3230 & w3253 ) | ( w3231 & w3253 ) ;
  assign w3270 = w2067 & ~w2811 ;
  assign w3271 = ( w2072 & ~w2708 ) | ( w2072 & w3270 ) | ( ~w2708 & w3270 ) ;
  assign w3272 = w2070 | w3271 ;
  assign w3273 = ( w2597 & w3271 ) | ( w2597 & w3272 ) | ( w3271 & w3272 ) ;
  assign w3274 = w3270 | w3273 ;
  assign w3275 = ~w2080 & w2817 ;
  assign w3276 = ( w2817 & w3274 ) | ( w2817 & ~w3275 ) | ( w3274 & ~w3275 ) ;
  assign w3277 = w943 ^ w3276 ;
  assign w3278 = ( w3235 & w3243 ) | ( w3235 & w3251 ) | ( w3243 & w3251 ) ;
  assign w3279 = ( w297 & w3232 ) | ( w297 & w3233 ) | ( w3232 & w3233 ) ;
  assign w3280 = ~w1915 & w1962 ;
  assign w3281 = ( w1913 & w2053 ) | ( w1913 & w3280 ) | ( w2053 & w3280 ) ;
  assign w3282 = w1964 | w3281 ;
  assign w3283 = ( w1908 & w3281 ) | ( w1908 & w3282 ) | ( w3281 & w3282 ) ;
  assign w3284 = w3280 | w3283 ;
  assign w3285 = w1956 | w1965 ;
  assign w3286 = ( ~w1956 & w3284 ) | ( ~w1956 & w3285 ) | ( w3284 & w3285 ) ;
  assign w3287 = w532 ^ w3286 ;
  assign w3288 = w3279 ^ w3287 ;
  assign w3289 = w285 ^ w3288 ;
  assign w3290 = w297 ^ w3289 ;
  assign w3291 = w532 & w1925 ;
  assign w3292 = w3290 ^ w3291 ;
  assign w3293 = w1983 & w2371 ;
  assign w3294 = ( w1985 & ~w2372 ) | ( w1985 & w3293 ) | ( ~w2372 & w3293 ) ;
  assign w3295 = w1986 | w3294 ;
  assign w3296 = ( w2369 & w3294 ) | ( w2369 & w3295 ) | ( w3294 & w3295 ) ;
  assign w3297 = w3293 | w3296 ;
  assign w3298 = w1980 | w2380 ;
  assign w3299 = ( ~w2380 & w3297 ) | ( ~w2380 & w3298 ) | ( w3297 & w3298 ) ;
  assign w3300 = w660 ^ w3299 ;
  assign w3301 = w3278 ^ w3300 ;
  assign w3302 = w3292 ^ w3301 ;
  assign w3303 = w3269 ^ w3277 ;
  assign w3304 = w3302 ^ w3303 ;
  assign w3305 = ( w3215 & w3217 ) | ( w3215 & w3257 ) | ( w3217 & w3257 ) ;
  assign w3306 = w3268 ^ w3305 ;
  assign w3307 = w3304 ^ w3306 ;
  assign w3308 = w333 | w3125 ;
  assign w3309 = ( w125 & w1651 ) | ( w125 & ~w3125 ) | ( w1651 & ~w3125 ) ;
  assign w3310 = w3308 | w3309 ;
  assign w3311 = ( w108 & ~w123 ) | ( w108 & w763 ) | ( ~w123 & w763 ) ;
  assign w3312 = w3204 | w3310 ;
  assign w3313 = ( w123 & w197 ) | ( w123 & ~w3204 ) | ( w197 & ~w3204 ) ;
  assign w3314 = w3312 | w3313 ;
  assign w3315 = w3311 | w3314 ;
  assign w3316 = ( w226 & w353 ) | ( w226 & ~w451 ) | ( w353 & ~w451 ) ;
  assign w3317 = w163 | w3315 ;
  assign w3318 = ( ~w163 & w451 ) | ( ~w163 & w502 ) | ( w451 & w502 ) ;
  assign w3319 = w3317 | w3318 ;
  assign w3320 = w3316 | w3319 ;
  assign w3321 = w3267 ^ w3307 ;
  assign w3322 = w3320 ^ w3321 ;
  assign w3323 = w3262 & w3322 ;
  assign w3324 = w3262 ^ w3322 ;
  assign w3325 = w3263 | w3264 ;
  assign w3326 = w2892 & w3325 ;
  assign w3327 = w3324 ^ w3326 ;
  assign w3328 = ( w3267 & w3307 ) | ( w3267 & w3320 ) | ( w3307 & w3320 ) ;
  assign w3329 = w227 | w229 ;
  assign w3330 = w601 | w3329 ;
  assign w3331 = ( w160 & ~w601 ) | ( w160 & w1541 ) | ( ~w601 & w1541 ) ;
  assign w3332 = w3330 | w3331 ;
  assign w3333 = ( w162 & w219 ) | ( w162 & ~w233 ) | ( w219 & ~w233 ) ;
  assign w3334 = w71 | w3332 ;
  assign w3335 = ( ~w71 & w233 ) | ( ~w71 & w452 ) | ( w233 & w452 ) ;
  assign w3336 = w3334 | w3335 ;
  assign w3337 = w3333 | w3336 ;
  assign w3338 = w364 | w453 ;
  assign w3339 = w1719 | w3338 ;
  assign w3340 = ( w164 & w904 ) | ( w164 & ~w1719 ) | ( w904 & ~w1719 ) ;
  assign w3341 = w3339 | w3340 ;
  assign w3342 = ( w215 & ~w265 ) | ( w215 & w3341 ) | ( ~w265 & w3341 ) ;
  assign w3343 = w2638 | w3337 ;
  assign w3344 = ( w265 & w412 ) | ( w265 & ~w3337 ) | ( w412 & ~w3337 ) ;
  assign w3345 = w3343 | w3344 ;
  assign w3346 = w3342 | w3345 ;
  assign w3347 = w365 | w476 ;
  assign w3348 = w232 | w3347 ;
  assign w3349 = ( ~w232 & w332 ) | ( ~w232 & w3346 ) | ( w332 & w3346 ) ;
  assign w3350 = w3348 | w3349 ;
  assign w3351 = ( w3268 & w3304 ) | ( w3268 & w3305 ) | ( w3304 & w3305 ) ;
  assign w3352 = ( w3269 & w3277 ) | ( w3269 & w3302 ) | ( w3277 & w3302 ) ;
  assign w3353 = w2072 & ~w2811 ;
  assign w3354 = ( w2070 & ~w2708 ) | ( w2070 & w3353 ) | ( ~w2708 & w3353 ) ;
  assign w3355 = ( w2708 & w2815 ) | ( w2708 & ~w3354 ) | ( w2815 & ~w3354 ) ;
  assign w3356 = ( w2080 & w2811 ) | ( w2080 & ~w2815 ) | ( w2811 & ~w2815 ) ;
  assign w3357 = ( w3353 & w3355 ) | ( w3353 & w3356 ) | ( w3355 & w3356 ) ;
  assign w3358 = ( ~w3180 & w3354 ) | ( ~w3180 & w3357 ) | ( w3354 & w3357 ) ;
  assign w3359 = ( w3278 & w3292 ) | ( w3278 & w3300 ) | ( w3292 & w3300 ) ;
  assign w3360 = w285 ^ w297 ;
  assign w3361 = w3291 ^ w3360 ;
  assign w3362 = ( w3279 & w3287 ) | ( w3279 & w3361 ) | ( w3287 & w3361 ) ;
  assign w3363 = w1908 & w1962 ;
  assign w3364 = ( ~w1915 & w2053 ) | ( ~w1915 & w3363 ) | ( w2053 & w3363 ) ;
  assign w3365 = w1964 | w3364 ;
  assign w3366 = ( w2371 & w3364 ) | ( w2371 & w3365 ) | ( w3364 & w3365 ) ;
  assign w3367 = w3363 | w3366 ;
  assign w3368 = ~w1965 & w2402 ;
  assign w3369 = ( w2402 & w3367 ) | ( w2402 & ~w3368 ) | ( w3367 & ~w3368 ) ;
  assign w3370 = w532 ^ w3369 ;
  assign w3371 = w532 & w1913 ;
  assign w3372 = w3370 ^ w3371 ;
  assign w3373 = ( w285 & w297 ) | ( w285 & ~w3291 ) | ( w297 & ~w3291 ) ;
  assign w3374 = w3372 ^ w3373 ;
  assign w3375 = w1983 & ~w2372 ;
  assign w3376 = ( w1985 & w2369 ) | ( w1985 & w3375 ) | ( w2369 & w3375 ) ;
  assign w3377 = w1986 | w3376 ;
  assign w3378 = ( w2597 & w3376 ) | ( w2597 & w3377 ) | ( w3376 & w3377 ) ;
  assign w3379 = w3375 | w3378 ;
  assign w3380 = ~w1980 & w2603 ;
  assign w3381 = ( w2603 & w3379 ) | ( w2603 & ~w3380 ) | ( w3379 & ~w3380 ) ;
  assign w3382 = w660 ^ w3381 ;
  assign w3383 = w3374 ^ w3382 ;
  assign w3384 = w3362 ^ w3383 ;
  assign w3385 = w943 ^ w3359 ;
  assign w3386 = w3358 ^ w3385 ;
  assign w3387 = w3384 ^ w3386 ;
  assign w3388 = w3351 ^ w3352 ;
  assign w3389 = w3387 ^ w3388 ;
  assign w3390 = w3328 ^ w3389 ;
  assign w3391 = w3350 ^ w3390 ;
  assign w3392 = w3323 & w3391 ;
  assign w3393 = w3323 ^ w3391 ;
  assign w3394 = w3324 | w3325 ;
  assign w3395 = w2892 & w3394 ;
  assign w3396 = w3393 ^ w3395 ;
  assign w3397 = ( w3328 & w3350 ) | ( w3328 & w3389 ) | ( w3350 & w3389 ) ;
  assign w3398 = ( w712 & w763 ) | ( w712 & ~w2330 ) | ( w763 & ~w2330 ) ;
  assign w3399 = w210 | w1810 ;
  assign w3400 = ( ~w210 & w2330 ) | ( ~w210 & w2357 ) | ( w2330 & w2357 ) ;
  assign w3401 = w3399 | w3400 ;
  assign w3402 = w3398 | w3401 ;
  assign w3403 = ( w233 & w242 ) | ( w233 & ~w333 ) | ( w242 & ~w333 ) ;
  assign w3404 = w114 | w3402 ;
  assign w3405 = ( ~w114 & w333 ) | ( ~w114 & w343 ) | ( w333 & w343 ) ;
  assign w3406 = w3404 | w3405 ;
  assign w3407 = w3403 | w3406 ;
  assign w3408 = ( ~w224 & w360 ) | ( ~w224 & w3407 ) | ( w360 & w3407 ) ;
  assign w3409 = w224 | w3408 ;
  assign w3410 = w943 ^ w3358 ;
  assign w3411 = ( w3359 & w3384 ) | ( w3359 & w3410 ) | ( w3384 & w3410 ) ;
  assign w3412 = ( ~w3370 & w3371 ) | ( ~w3370 & w3373 ) | ( w3371 & w3373 ) ;
  assign w3413 = w1962 & w2371 ;
  assign w3414 = ( w1908 & w2053 ) | ( w1908 & w3413 ) | ( w2053 & w3413 ) ;
  assign w3415 = w1964 | w3414 ;
  assign w3416 = ( ~w2372 & w3414 ) | ( ~w2372 & w3415 ) | ( w3414 & w3415 ) ;
  assign w3417 = w3413 | w3416 ;
  assign w3418 = w1965 | w2394 ;
  assign w3419 = ( ~w2394 & w3417 ) | ( ~w2394 & w3418 ) | ( w3417 & w3418 ) ;
  assign w3420 = w532 ^ w3419 ;
  assign w3421 = w532 & ~w1953 ;
  assign w3422 = w3420 ^ w3421 ;
  assign w3423 = w1983 & w2369 ;
  assign w3424 = ( w1985 & w2597 ) | ( w1985 & w3423 ) | ( w2597 & w3423 ) ;
  assign w3425 = w1986 | w3424 ;
  assign w3426 = ( ~w2708 & w3424 ) | ( ~w2708 & w3425 ) | ( w3424 & w3425 ) ;
  assign w3427 = w3423 | w3426 ;
  assign w3428 = w1980 | w2714 ;
  assign w3429 = ( ~w2714 & w3427 ) | ( ~w2714 & w3428 ) | ( w3427 & w3428 ) ;
  assign w3430 = w660 ^ w3429 ;
  assign w3431 = w3422 ^ w3430 ;
  assign w3432 = w3412 ^ w3431 ;
  assign w3433 = ( w3362 & w3374 ) | ( w3362 & w3382 ) | ( w3374 & w3382 ) ;
  assign w3434 = w2070 & ~w2811 ;
  assign w3435 = w2080 | w3434 ;
  assign w3436 = ( ~w2919 & w3434 ) | ( ~w2919 & w3435 ) | ( w3434 & w3435 ) ;
  assign w3437 = w943 ^ w3436 ;
  assign w3438 = w3432 ^ w3437 ;
  assign w3439 = w3433 ^ w3438 ;
  assign w3440 = ( w3351 & w3352 ) | ( w3351 & w3387 ) | ( w3352 & w3387 ) ;
  assign w3441 = w3439 ^ w3440 ;
  assign w3442 = w3411 ^ w3441 ;
  assign w3443 = w3397 ^ w3442 ;
  assign w3444 = w3409 ^ w3443 ;
  assign w3445 = w3392 & w3444 ;
  assign w3446 = w3392 ^ w3444 ;
  assign w3447 = w3393 | w3394 ;
  assign w3448 = w2892 & w3447 ;
  assign w3449 = w3446 ^ w3448 ;
  assign w3450 = ( w3397 & w3409 ) | ( w3397 & w3442 ) | ( w3409 & w3442 ) ;
  assign w3451 = w267 | w512 ;
  assign w3452 = w483 | w3451 ;
  assign w3453 = ( w218 & ~w483 ) | ( w218 & w645 ) | ( ~w483 & w645 ) ;
  assign w3454 = w3452 | w3453 ;
  assign w3455 = ( w901 & ~w2357 ) | ( w901 & w2624 ) | ( ~w2357 & w2624 ) ;
  assign w3456 = w986 | w3454 ;
  assign w3457 = ( w171 & ~w986 ) | ( w171 & w2357 ) | ( ~w986 & w2357 ) ;
  assign w3458 = w3456 | w3457 ;
  assign w3459 = w3455 | w3458 ;
  assign w3460 = w192 | w321 ;
  assign w3461 = ( ~w192 & w318 ) | ( ~w192 & w3459 ) | ( w318 & w3459 ) ;
  assign w3462 = w3460 | w3461 ;
  assign w3463 = ( w3411 & w3439 ) | ( w3411 & w3440 ) | ( w3439 & w3440 ) ;
  assign w3464 = ( w3432 & w3433 ) | ( w3432 & w3437 ) | ( w3433 & w3437 ) ;
  assign w3465 = w532 ^ w3420 ;
  assign w3466 = ( w1913 & ~w1915 ) | ( w1913 & w3465 ) | ( ~w1915 & w3465 ) ;
  assign w3467 = ( ~w1913 & w3420 ) | ( ~w1913 & w3466 ) | ( w3420 & w3466 ) ;
  assign w3468 = ( ~w943 & w1908 ) | ( ~w943 & w1913 ) | ( w1908 & w1913 ) ;
  assign w3469 = w532 & w3468 ;
  assign w3470 = w1962 & ~w2372 ;
  assign w3471 = ( w2053 & w2371 ) | ( w2053 & w3470 ) | ( w2371 & w3470 ) ;
  assign w3472 = w1964 | w3471 ;
  assign w3473 = ( w2369 & w3471 ) | ( w2369 & w3472 ) | ( w3471 & w3472 ) ;
  assign w3474 = w3470 | w3473 ;
  assign w3475 = w1965 | w2380 ;
  assign w3476 = ( ~w2380 & w3474 ) | ( ~w2380 & w3475 ) | ( w3474 & w3475 ) ;
  assign w3477 = w532 ^ w3476 ;
  assign w3478 = w1908 ^ w1913 ;
  assign w3479 = w532 & w3478 ;
  assign w3480 = w3467 ^ w3477 ;
  assign w3481 = w943 ^ w3480 ;
  assign w3482 = w3479 ^ w3481 ;
  assign w3483 = ( w3412 & w3422 ) | ( w3412 & ~w3430 ) | ( w3422 & ~w3430 ) ;
  assign w3484 = w1983 & w2597 ;
  assign w3485 = ( w1985 & ~w2708 ) | ( w1985 & w3484 ) | ( ~w2708 & w3484 ) ;
  assign w3486 = w1986 | w3485 ;
  assign w3487 = ( ~w2811 & w3485 ) | ( ~w2811 & w3486 ) | ( w3485 & w3486 ) ;
  assign w3488 = w3484 | w3487 ;
  assign w3489 = ~w1980 & w2817 ;
  assign w3490 = ( w2817 & w3488 ) | ( w2817 & ~w3489 ) | ( w3488 & ~w3489 ) ;
  assign w3491 = w660 ^ w3490 ;
  assign w3492 = w3483 ^ w3491 ;
  assign w3493 = w3482 ^ w3492 ;
  assign w3494 = w3463 ^ w3464 ;
  assign w3495 = w3493 ^ w3494 ;
  assign w3496 = w3450 ^ w3495 ;
  assign w3497 = w3462 ^ w3496 ;
  assign w3498 = w3445 & w3497 ;
  assign w3499 = w3445 ^ w3497 ;
  assign w3500 = w3446 | w3447 ;
  assign w3501 = w2892 & w3500 ;
  assign w3502 = w3499 ^ w3501 ;
  assign w3503 = ( w3450 & w3462 ) | ( w3450 & w3495 ) | ( w3462 & w3495 ) ;
  assign w3504 = w477 | w894 ;
  assign w3505 = ( w171 & w506 ) | ( w171 & ~w894 ) | ( w506 & ~w894 ) ;
  assign w3506 = w3504 | w3505 ;
  assign w3507 = w342 | w3506 ;
  assign w3508 = w459 | w3507 ;
  assign w3509 = ( ~w459 & w628 ) | ( ~w459 & w2692 ) | ( w628 & w2692 ) ;
  assign w3510 = w3508 | w3509 ;
  assign w3511 = ( w3463 & w3464 ) | ( w3463 & w3493 ) | ( w3464 & w3493 ) ;
  assign w3512 = ( w3482 & w3483 ) | ( w3482 & ~w3491 ) | ( w3483 & ~w3491 ) ;
  assign w3513 = w943 ^ w3479 ;
  assign w3514 = ( w3467 & w3477 ) | ( w3467 & ~w3513 ) | ( w3477 & ~w3513 ) ;
  assign w3515 = w532 & w2371 ;
  assign w3516 = w1962 & w2369 ;
  assign w3517 = ( w2053 & ~w2372 ) | ( w2053 & w3516 ) | ( ~w2372 & w3516 ) ;
  assign w3518 = w1964 | w3517 ;
  assign w3519 = ( w2597 & w3517 ) | ( w2597 & w3518 ) | ( w3517 & w3518 ) ;
  assign w3520 = w3516 | w3519 ;
  assign w3521 = ~w1965 & w2603 ;
  assign w3522 = ( w2603 & w3520 ) | ( w2603 & ~w3521 ) | ( w3520 & ~w3521 ) ;
  assign w3523 = w532 ^ w3522 ;
  assign w3524 = w3515 ^ w3523 ;
  assign w3525 = w3469 ^ w3524 ;
  assign w3526 = w1985 & ~w2811 ;
  assign w3527 = ( w1983 & ~w2708 ) | ( w1983 & w3526 ) | ( ~w2708 & w3526 ) ;
  assign w3528 = ( w2708 & w2815 ) | ( w2708 & ~w3527 ) | ( w2815 & ~w3527 ) ;
  assign w3529 = ( w1980 & w2811 ) | ( w1980 & ~w2815 ) | ( w2811 & ~w2815 ) ;
  assign w3530 = ( w3526 & w3528 ) | ( w3526 & w3529 ) | ( w3528 & w3529 ) ;
  assign w3531 = ( ~w3180 & w3527 ) | ( ~w3180 & w3530 ) | ( w3527 & w3530 ) ;
  assign w3532 = w660 ^ w3514 ;
  assign w3533 = w3525 ^ w3532 ;
  assign w3534 = w3531 ^ w3533 ;
  assign w3535 = w3511 ^ w3512 ;
  assign w3536 = w3534 ^ w3535 ;
  assign w3537 = w3503 ^ w3536 ;
  assign w3538 = w3510 ^ w3537 ;
  assign w3539 = w3498 & w3538 ;
  assign w3540 = w3498 ^ w3538 ;
  assign w3541 = w3499 | w3500 ;
  assign w3542 = w2892 & w3541 ;
  assign w3543 = w3540 ^ w3542 ;
  assign w3544 = ( w3503 & w3510 ) | ( w3503 & w3536 ) | ( w3510 & w3536 ) ;
  assign w3545 = w242 | w341 ;
  assign w3546 = w183 | w3545 ;
  assign w3547 = ( w174 & ~w183 ) | ( w174 & w215 ) | ( ~w183 & w215 ) ;
  assign w3548 = w3546 | w3547 ;
  assign w3549 = ( ~w197 & w868 ) | ( ~w197 & w3548 ) | ( w868 & w3548 ) ;
  assign w3550 = w1621 | w2901 ;
  assign w3551 = ( w197 & w244 ) | ( w197 & ~w2901 ) | ( w244 & ~w2901 ) ;
  assign w3552 = w3550 | w3551 ;
  assign w3553 = w3549 | w3552 ;
  assign w3554 = w125 | w219 ;
  assign w3555 = w384 | w3554 ;
  assign w3556 = ( w115 & ~w384 ) | ( w115 & w3553 ) | ( ~w384 & w3553 ) ;
  assign w3557 = w3555 | w3556 ;
  assign w3558 = ( ~w3511 & w3512 ) | ( ~w3511 & w3534 ) | ( w3512 & w3534 ) ;
  assign w3559 = w660 ^ w3531 ;
  assign w3560 = ( w3514 & ~w3525 ) | ( w3514 & w3559 ) | ( ~w3525 & w3559 ) ;
  assign w3561 = w1983 & ~w2811 ;
  assign w3562 = w1980 | w3561 ;
  assign w3563 = ( ~w2919 & w3561 ) | ( ~w2919 & w3562 ) | ( w3561 & w3562 ) ;
  assign w3564 = w660 ^ w3563 ;
  assign w3565 = w1962 & w2597 ;
  assign w3566 = ( w2053 & w2369 ) | ( w2053 & w3565 ) | ( w2369 & w3565 ) ;
  assign w3567 = w1964 | w3566 ;
  assign w3568 = ( ~w2708 & w3566 ) | ( ~w2708 & w3567 ) | ( w3566 & w3567 ) ;
  assign w3569 = w3565 | w3568 ;
  assign w3570 = w1965 | w2714 ;
  assign w3571 = ( ~w2714 & w3569 ) | ( ~w2714 & w3570 ) | ( w3569 & w3570 ) ;
  assign w3572 = w532 ^ w3571 ;
  assign w3573 = ( w3469 & ~w3515 ) | ( w3469 & w3523 ) | ( ~w3515 & w3523 ) ;
  assign w3574 = w532 & ~w2372 ;
  assign w3575 = ( w3515 & w3573 ) | ( w3515 & ~w3574 ) | ( w3573 & ~w3574 ) ;
  assign w3576 = w3573 ^ w3574 ;
  assign w3577 = w3515 ^ w3576 ;
  assign w3578 = w3564 ^ w3572 ;
  assign w3579 = w3577 ^ w3578 ;
  assign w3580 = w3558 ^ w3579 ;
  assign w3581 = w3560 ^ w3580 ;
  assign w3582 = w3544 ^ w3581 ;
  assign w3583 = w3557 ^ w3582 ;
  assign w3584 = w3539 & w3583 ;
  assign w3585 = w3539 ^ w3583 ;
  assign w3586 = w3540 | w3541 ;
  assign w3587 = w2892 & w3586 ;
  assign w3588 = w3585 ^ w3587 ;
  assign w3589 = ( w3544 & w3557 ) | ( w3544 & w3581 ) | ( w3557 & w3581 ) ;
  assign w3590 = w364 | w400 ;
  assign w3591 = w197 | w3590 ;
  assign w3592 = ( w83 & ~w197 ) | ( w83 & w263 ) | ( ~w197 & w263 ) ;
  assign w3593 = w3591 | w3592 ;
  assign w3594 = ( w150 & w905 ) | ( w150 & ~w2874 ) | ( w905 & ~w2874 ) ;
  assign w3595 = w317 | w1537 ;
  assign w3596 = ( ~w1537 & w2874 ) | ( ~w1537 & w3593 ) | ( w2874 & w3593 ) ;
  assign w3597 = w3595 | w3596 ;
  assign w3598 = w3594 | w3597 ;
  assign w3599 = ( w164 & w202 ) | ( w164 & ~w265 ) | ( w202 & ~w265 ) ;
  assign w3600 = w2658 | w3598 ;
  assign w3601 = ( w265 & w349 ) | ( w265 & ~w3598 ) | ( w349 & ~w3598 ) ;
  assign w3602 = w3600 | w3601 ;
  assign w3603 = w3599 | w3602 ;
  assign w3604 = w128 | w477 ;
  assign w3605 = ( ~w128 & w355 ) | ( ~w128 & w3603 ) | ( w355 & w3603 ) ;
  assign w3606 = w3604 | w3605 ;
  assign w3607 = ( w3558 & ~w3560 ) | ( w3558 & w3579 ) | ( ~w3560 & w3579 ) ;
  assign w3608 = w1962 & ~w2708 ;
  assign w3609 = ( w2053 & w2597 ) | ( w2053 & w3608 ) | ( w2597 & w3608 ) ;
  assign w3610 = w1964 | w3609 ;
  assign w3611 = ( ~w2811 & w3609 ) | ( ~w2811 & w3610 ) | ( w3609 & w3610 ) ;
  assign w3612 = w3608 | w3611 ;
  assign w3613 = ~w1965 & w2817 ;
  assign w3614 = ( w2817 & w3612 ) | ( w2817 & ~w3613 ) | ( w3612 & ~w3613 ) ;
  assign w3615 = w532 ^ w3614 ;
  assign w3616 = w2369 ^ w2372 ;
  assign w3617 = w532 & ~w3616 ;
  assign w3618 = w3575 ^ w3615 ;
  assign w3619 = w660 ^ w3618 ;
  assign w3620 = w3617 ^ w3619 ;
  assign w3621 = ( w3564 & w3572 ) | ( w3564 & ~w3577 ) | ( w3572 & ~w3577 ) ;
  assign w3622 = w3607 ^ w3620 ;
  assign w3623 = w3621 ^ w3622 ;
  assign w3624 = ( w3589 & w3606 ) | ( w3589 & w3623 ) | ( w3606 & w3623 ) ;
  assign w3625 = w3589 ^ w3623 ;
  assign w3626 = w3606 ^ w3625 ;
  assign w3627 = w3584 & w3626 ;
  assign w3628 = w3584 ^ w3626 ;
  assign w3629 = w3585 | w3586 ;
  assign w3630 = w2892 & w3629 ;
  assign w3631 = w3628 ^ w3630 ;
  assign w3632 = ( ~w197 & w480 ) | ( ~w197 & w1811 ) | ( w480 & w1811 ) ;
  assign w3633 = w892 | w1552 ;
  assign w3634 = ( w197 & w244 ) | ( w197 & ~w892 ) | ( w244 & ~w892 ) ;
  assign w3635 = w3633 | w3634 ;
  assign w3636 = w3632 | w3635 ;
  assign w3637 = ( ~w124 & w908 ) | ( ~w124 & w2357 ) | ( w908 & w2357 ) ;
  assign w3638 = w1182 | w3636 ;
  assign w3639 = ( w124 & w173 ) | ( w124 & ~w1182 ) | ( w173 & ~w1182 ) ;
  assign w3640 = w3638 | w3639 ;
  assign w3641 = w3637 | w3640 ;
  assign w3642 = ( w342 & w349 ) | ( w342 & ~w374 ) | ( w349 & ~w374 ) ;
  assign w3643 = w105 | w3641 ;
  assign w3644 = ( ~w105 & w374 ) | ( ~w105 & w513 ) | ( w374 & w513 ) ;
  assign w3645 = w3643 | w3644 ;
  assign w3646 = w3642 | w3645 ;
  assign w3647 = ( w3607 & w3620 ) | ( w3607 & ~w3621 ) | ( w3620 & ~w3621 ) ;
  assign w3648 = w660 ^ w3617 ;
  assign w3649 = ( w3575 & w3615 ) | ( w3575 & ~w3648 ) | ( w3615 & ~w3648 ) ;
  assign w3650 = w1962 & ~w2811 ;
  assign w3651 = ( w2708 & w2811 ) | ( w2708 & w2815 ) | ( w2811 & w2815 ) ;
  assign w3652 = ( w1965 & w2708 ) | ( w1965 & w3651 ) | ( w2708 & w3651 ) ;
  assign w3653 = w2053 | w2708 ;
  assign w3654 = ( ~w2708 & w3652 ) | ( ~w2708 & w3653 ) | ( w3652 & w3653 ) ;
  assign w3655 = w2708 & w3651 ;
  assign w3656 = ( w3650 & w3654 ) | ( w3650 & ~w3655 ) | ( w3654 & ~w3655 ) ;
  assign w3657 = ( w660 & ~w2369 ) | ( w660 & w2372 ) | ( ~w2369 & w2372 ) ;
  assign w3658 = w2597 ^ w3657 ;
  assign w3659 = w532 & w3658 ;
  assign w3660 = w3656 ^ w3659 ;
  assign w3661 = w3647 ^ w3649 ;
  assign w3662 = w3660 ^ w3661 ;
  assign w3663 = w3624 ^ w3662 ;
  assign w3664 = w3646 ^ w3663 ;
  assign w3665 = w3627 & w3664 ;
  assign w3666 = w3627 ^ w3664 ;
  assign w3667 = w3628 | w3629 ;
  assign w3668 = w2892 & w3667 ;
  assign w3669 = w3666 ^ w3668 ;
  assign w3670 = ( w3624 & w3646 ) | ( w3624 & w3662 ) | ( w3646 & w3662 ) ;
  assign w3671 = w262 | w343 ;
  assign w3672 = ( ~w262 & w334 ) | ( ~w262 & w1033 ) | ( w334 & w1033 ) ;
  assign w3673 = w3671 | w3672 ;
  assign w3674 = ( w350 & ~w895 ) | ( w350 & w998 ) | ( ~w895 & w998 ) ;
  assign w3675 = w1750 | w3673 ;
  assign w3676 = ( w895 & ~w1750 ) | ( w895 & w3548 ) | ( ~w1750 & w3548 ) ;
  assign w3677 = w3675 | w3676 ;
  assign w3678 = w3674 | w3677 ;
  assign w3679 = ( w225 & w234 ) | ( w225 & ~w360 ) | ( w234 & ~w360 ) ;
  assign w3680 = w105 | w3678 ;
  assign w3681 = ( ~w105 & w360 ) | ( ~w105 & w513 ) | ( w360 & w513 ) ;
  assign w3682 = w3680 | w3681 ;
  assign w3683 = w3679 | w3682 ;
  assign w3684 = w690 | w3683 ;
  assign w3685 = w2053 & ~w2811 ;
  assign w3686 = w1965 | w3685 ;
  assign w3687 = ( ~w2919 & w3685 ) | ( ~w2919 & w3686 ) | ( w3685 & w3686 ) ;
  assign w3688 = w532 ^ w3687 ;
  assign w3689 = ( w2597 & w3656 ) | ( w2597 & ~w3657 ) | ( w3656 & ~w3657 ) ;
  assign w3690 = w532 ^ w3656 ;
  assign w3691 = ( ~w2597 & w3689 ) | ( ~w2597 & w3690 ) | ( w3689 & w3690 ) ;
  assign w3692 = ( w3647 & ~w3649 ) | ( w3647 & w3660 ) | ( ~w3649 & w3660 ) ;
  assign w3693 = w532 & ~w2713 ;
  assign w3694 = w3688 ^ w3691 ;
  assign w3695 = w3692 ^ w3694 ;
  assign w3696 = w3693 ^ w3695 ;
  assign w3697 = ( w3670 & w3684 ) | ( w3670 & w3696 ) | ( w3684 & w3696 ) ;
  assign w3698 = w3670 ^ w3696 ;
  assign w3699 = w3684 ^ w3698 ;
  assign w3700 = w3665 & w3699 ;
  assign w3701 = w3665 ^ w3699 ;
  assign w3702 = w3666 | w3667 ;
  assign w3703 = w2892 & w3702 ;
  assign w3704 = w3701 ^ w3703 ;
  assign w3705 = ( ~w173 & w1623 ) | ( ~w173 & w3593 ) | ( w1623 & w3593 ) ;
  assign w3706 = w241 | w1684 ;
  assign w3707 = ( w173 & ~w241 ) | ( w173 & w510 ) | ( ~w241 & w510 ) ;
  assign w3708 = w3706 | w3707 ;
  assign w3709 = w3705 | w3708 ;
  assign w3710 = ( w216 & ~w453 ) | ( w216 & w482 ) | ( ~w453 & w482 ) ;
  assign w3711 = w2661 | w3709 ;
  assign w3712 = ( w453 & w484 ) | ( w453 & ~w2661 ) | ( w484 & ~w2661 ) ;
  assign w3713 = w3711 | w3712 ;
  assign w3714 = w3710 | w3713 ;
  assign w3715 = ( ~w2597 & w2708 ) | ( ~w2597 & w3692 ) | ( w2708 & w3692 ) ;
  assign w3716 = w532 ^ w3692 ;
  assign w3717 = ( ~w2597 & w2708 ) | ( ~w2597 & w3716 ) | ( w2708 & w3716 ) ;
  assign w3718 = ( w3692 & ~w3715 ) | ( w3692 & w3717 ) | ( ~w3715 & w3717 ) ;
  assign w3719 = ( w3688 & w3691 ) | ( w3688 & w3718 ) | ( w3691 & w3718 ) ;
  assign w3720 = ( w2597 & w3692 ) | ( w2597 & w3718 ) | ( w3692 & w3718 ) ;
  assign w3721 = w3719 ^ w3720 ;
  assign w3722 = w2597 ^ w2811 ;
  assign w3723 = w532 & w3722 ;
  assign w3724 = w3721 ^ w3723 ;
  assign w3725 = ( w3697 & w3714 ) | ( w3697 & w3724 ) | ( w3714 & w3724 ) ;
  assign w3726 = w3697 ^ w3724 ;
  assign w3727 = w3714 ^ w3726 ;
  assign w3728 = w3700 & w3727 ;
  assign w3729 = w3700 ^ w3727 ;
  assign w3730 = w3701 | w3702 ;
  assign w3731 = w2892 & w3730 ;
  assign w3732 = w3729 ^ w3731 ;
  assign w3733 = ( w150 & w222 ) | ( w150 & ~w307 ) | ( w222 & ~w307 ) ;
  assign w3734 = w140 | w147 ;
  assign w3735 = ( ~w147 & w307 ) | ( ~w147 & w411 ) | ( w307 & w411 ) ;
  assign w3736 = w3734 | w3735 ;
  assign w3737 = w3733 | w3736 ;
  assign w3738 = ( ~w267 & w823 ) | ( ~w267 & w3737 ) | ( w823 & w3737 ) ;
  assign w3739 = w267 | w3738 ;
  assign w3740 = ( ~w125 & w905 ) | ( ~w125 & w3739 ) | ( w905 & w3739 ) ;
  assign w3741 = w563 | w2341 ;
  assign w3742 = ( w125 & w215 ) | ( w125 & ~w563 ) | ( w215 & ~w563 ) ;
  assign w3743 = w3741 | w3742 ;
  assign w3744 = w3740 | w3743 ;
  assign w3745 = w223 | w372 ;
  assign w3746 = ( ~w223 & w302 ) | ( ~w223 & w3744 ) | ( w302 & w3744 ) ;
  assign w3747 = w3745 | w3746 ;
  assign w3748 = w3725 & w3747 ;
  assign w3749 = w3725 ^ w3747 ;
  assign w3750 = w3728 ^ w3749 ;
  assign w3751 = w3729 | w3730 ;
  assign w3752 = w2892 & w3751 ;
  assign w3753 = w3750 ^ w3752 ;
  assign w3754 = w3728 & w3749 ;
  assign w3755 = w1041 | w1529 ;
  assign w3756 = ( w580 & w600 ) | ( w580 & ~w1041 ) | ( w600 & ~w1041 ) ;
  assign w3757 = w3755 | w3756 ;
  assign w3758 = ( ~w173 & w911 ) | ( ~w173 & w991 ) | ( w911 & w991 ) ;
  assign w3759 = w2635 | w3757 ;
  assign w3760 = ( w173 & w235 ) | ( w173 & ~w3757 ) | ( w235 & ~w3757 ) ;
  assign w3761 = w3759 | w3760 ;
  assign w3762 = w3758 | w3761 ;
  assign w3763 = w215 | w361 ;
  assign w3764 = ( ~w215 & w245 ) | ( ~w215 & w3762 ) | ( w245 & w3762 ) ;
  assign w3765 = w3763 | w3764 ;
  assign w3766 = w3748 & w3765 ;
  assign w3767 = w3748 | w3765 ;
  assign w3768 = w3754 & w3767 ;
  assign w3769 = w3754 ^ w3767 ;
  assign w3770 = ( w3766 & w3767 ) | ( w3766 & ~w3769 ) | ( w3767 & ~w3769 ) ;
  assign w3771 = ( w3754 & w3769 ) | ( w3754 & ~w3770 ) | ( w3769 & ~w3770 ) ;
  assign w3772 = w3750 | w3751 ;
  assign w3773 = w2892 & w3772 ;
  assign w3774 = w3771 ^ w3773 ;
  assign w3775 = w375 | w3125 ;
  assign w3776 = w860 | w3775 ;
  assign w3777 = ( ~w860 & w1893 ) | ( ~w860 & w3673 ) | ( w1893 & w3673 ) ;
  assign w3778 = w3776 | w3777 ;
  assign w3779 = ( w133 & w146 ) | ( w133 & ~w216 ) | ( w146 & ~w216 ) ;
  assign w3780 = w126 | w3778 ;
  assign w3781 = ( ~w126 & w216 ) | ( ~w126 & w452 ) | ( w216 & w452 ) ;
  assign w3782 = w3780 | w3781 ;
  assign w3783 = w3779 | w3782 ;
  assign w3784 = ( ~w214 & w303 ) | ( ~w214 & w3783 ) | ( w303 & w3783 ) ;
  assign w3785 = w214 | w3784 ;
  assign w3786 = w3766 & w3785 ;
  assign w3787 = w3766 ^ w3785 ;
  assign w3788 = w3768 & w3787 ;
  assign w3789 = w3768 ^ w3787 ;
  assign w3790 = w3771 | w3772 ;
  assign w3791 = w2892 & w3790 ;
  assign w3792 = w3789 ^ w3791 ;
  assign w3793 = w305 | w464 ;
  assign w3794 = w509 | w3793 ;
  assign w3795 = ( w189 & ~w509 ) | ( w189 & w925 ) | ( ~w509 & w925 ) ;
  assign w3796 = w3794 | w3795 ;
  assign w3797 = ( w197 & ~w235 ) | ( w197 & w373 ) | ( ~w235 & w373 ) ;
  assign w3798 = w3337 | w3796 ;
  assign w3799 = ( w235 & w318 ) | ( w235 & ~w3337 ) | ( w318 & ~w3337 ) ;
  assign w3800 = w3798 | w3799 ;
  assign w3801 = w3797 | w3800 ;
  assign w3802 = w226 | w546 ;
  assign w3803 = w220 | w3802 ;
  assign w3804 = ( ~w220 & w221 ) | ( ~w220 & w3801 ) | ( w221 & w3801 ) ;
  assign w3805 = w3803 | w3804 ;
  assign w3806 = w3786 & w3805 ;
  assign w3807 = w3786 | w3805 ;
  assign w3808 = w3788 & w3807 ;
  assign w3809 = w3788 ^ w3807 ;
  assign w3810 = ( w3806 & w3807 ) | ( w3806 & ~w3809 ) | ( w3807 & ~w3809 ) ;
  assign w3811 = ( w3788 & w3809 ) | ( w3788 & ~w3810 ) | ( w3809 & ~w3810 ) ;
  assign w3812 = w3789 | w3790 ;
  assign w3813 = w2892 & w3812 ;
  assign w3814 = w3811 ^ w3813 ;
  assign w3815 = ( w139 & ~w349 ) | ( w139 & w509 ) | ( ~w349 & w509 ) ;
  assign w3816 = w450 | w496 ;
  assign w3817 = ( w349 & w353 ) | ( w349 & ~w496 ) | ( w353 & ~w496 ) ;
  assign w3818 = w3816 | w3817 ;
  assign w3819 = w3815 | w3818 ;
  assign w3820 = w364 | w3819 ;
  assign w3821 = w3806 & w3820 ;
  assign w3822 = w3806 ^ w3820 ;
  assign w3823 = w3808 & w3822 ;
  assign w3824 = w3808 ^ w3822 ;
  assign w3825 = w3811 | w3812 ;
  assign w3826 = w2892 & w3825 ;
  assign w3827 = w3824 ^ w3826 ;
  assign w3828 = w450 | w524 ;
  assign w3829 = w3821 & w3828 ;
  assign w3830 = ( w3821 & w3823 ) | ( w3821 & w3828 ) | ( w3823 & w3828 ) ;
  assign w3831 = w3823 & w3830 ;
  assign w3832 = w3821 | w3823 ;
  assign w3833 = w3821 ^ w3823 ;
  assign w3834 = ( w3828 & w3832 ) | ( w3828 & ~w3833 ) | ( w3832 & ~w3833 ) ;
  assign w3835 = w3832 ^ w3834 ;
  assign w3836 = w3824 | w3825 ;
  assign w3837 = w2892 & w3836 ;
  assign w3838 = w3835 ^ w3837 ;
  assign w3839 = w3835 | w3836 ;
  assign w3840 = w2892 & w3839 ;
  assign w3841 = w3831 ^ w3840 ;
  assign w3842 = w3829 ^ w3841 ;
  assign w3843 = \pi22 & ~w3842 ;
  assign w3844 = ( w45 & ~w3842 ) | ( w45 & w3843 ) | ( ~w3842 & w3843 ) ;
  assign w3845 = ( ~w3829 & w3831 ) | ( ~w3829 & w3839 ) | ( w3831 & w3839 ) ;
  assign w3846 = w3829 ^ w3845 ;
  assign w3847 = \pi23 & ~w45 ;
  assign w3848 = ~\pi22 & w3847 ;
  assign w3849 = ( w2892 & w3846 ) | ( w2892 & w3848 ) | ( w3846 & w3848 ) ;
  assign \po00 = w2788 ;
  assign \po01 = w2894 ;
  assign \po02 = w2979 ;
  assign \po03 = w3052 ;
  assign \po04 = w3122 ;
  assign \po05 = w3193 ;
  assign \po06 = w3266 ;
  assign \po07 = w3327 ;
  assign \po08 = w3396 ;
  assign \po09 = w3449 ;
  assign \po10 = w3502 ;
  assign \po11 = w3543 ;
  assign \po12 = w3588 ;
  assign \po13 = w3631 ;
  assign \po14 = w3669 ;
  assign \po15 = w3704 ;
  assign \po16 = w3732 ;
  assign \po17 = w3753 ;
  assign \po18 = w3774 ;
  assign \po19 = w3792 ;
  assign \po20 = w3814 ;
  assign \po21 = w3827 ;
  assign \po22 = w3838 ;
  assign \po23 = ~w3844 ;
  assign \po24 = w3849 ;
endmodule
