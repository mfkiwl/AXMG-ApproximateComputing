module div( \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 );
  input \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 ;
  output \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 ;
  wire zero , w129 , w130 , w131 , w132 , w133 , w134 , w135 , w136 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w146 , w147 , w148 , w149 , w150 , w151 , w152 , w153 , w154 , w155 , w156 , w157 , w158 , w159 , w160 , w161 , w162 , w163 , w164 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w174 , w175 , w176 , w177 , w178 , w179 , w180 , w181 , w182 , w183 , w184 , w185 , w186 , w187 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w203 , w204 , w205 , w206 , w207 , w208 , w209 , w210 , w211 , w212 , w213 , w214 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w224 , w225 , w226 , w227 , w228 , w229 , w230 , w231 , w232 , w233 , w234 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w250 , w251 , w252 , w253 , w254 , w255 , w256 , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 , w2495 , w2496 , w2497 , w2498 , w2499 , w2500 , w2501 , w2502 , w2503 , w2504 , w2505 , w2506 , w2507 , w2508 , w2509 , w2510 , w2511 , w2512 , w2513 , w2514 , w2515 , w2516 , w2517 , w2518 , w2519 , w2520 , w2521 , w2522 , w2523 , w2524 , w2525 , w2526 , w2527 , w2528 , w2529 , w2530 , w2531 , w2532 , w2533 , w2534 , w2535 , w2536 , w2537 , w2538 , w2539 , w2540 , w2541 , w2542 , w2543 , w2544 , w2545 , w2546 , w2547 , w2548 , w2549 , w2550 , w2551 , w2552 , w2553 , w2554 , w2555 , w2556 , w2557 , w2558 , w2559 , w2560 , w2561 , w2562 , w2563 , w2564 , w2565 , w2566 , w2567 , w2568 , w2569 , w2570 , w2571 , w2572 , w2573 , w2574 , w2575 , w2576 , w2577 , w2578 , w2579 , w2580 , w2581 , w2582 , w2583 , w2584 , w2585 , w2586 , w2587 , w2588 , w2589 , w2590 , w2591 , w2592 , w2593 , w2594 , w2595 , w2596 , w2597 , w2598 , w2599 , w2600 , w2601 , w2602 , w2603 , w2604 , w2605 , w2606 , w2607 , w2608 , w2609 , w2610 , w2611 , w2612 , w2613 , w2614 , w2615 , w2616 , w2617 , w2618 , w2619 , w2620 , w2621 , w2622 , w2623 , w2624 , w2625 , w2626 , w2627 , w2628 , w2629 , w2630 , w2631 , w2632 , w2633 , w2634 , w2635 , w2636 , w2637 , w2638 , w2639 , w2640 , w2641 , w2642 , w2643 , w2644 , w2645 , w2646 , w2647 , w2648 , w2649 , w2650 , w2651 , w2652 , w2653 , w2654 , w2655 , w2656 , w2657 , w2658 , w2659 , w2660 , w2661 , w2662 , w2663 , w2664 , w2665 , w2666 , w2667 , w2668 , w2669 , w2670 , w2671 , w2672 , w2673 , w2674 , w2675 , w2676 , w2677 , w2678 , w2679 , w2680 , w2681 , w2682 , w2683 , w2684 , w2685 , w2686 , w2687 , w2688 , w2689 , w2690 , w2691 , w2692 , w2693 , w2694 , w2695 , w2696 , w2697 , w2698 , w2699 , w2700 , w2701 , w2702 , w2703 , w2704 , w2705 , w2706 , w2707 , w2708 , w2709 , w2710 , w2711 , w2712 , w2713 , w2714 , w2715 , w2716 , w2717 , w2718 , w2719 , w2720 , w2721 , w2722 , w2723 , w2724 , w2725 , w2726 , w2727 , w2728 , w2729 , w2730 , w2731 , w2732 , w2733 , w2734 , w2735 , w2736 , w2737 , w2738 , w2739 , w2740 , w2741 , w2742 , w2743 , w2744 , w2745 , w2746 , w2747 , w2748 , w2749 , w2750 , w2751 , w2752 , w2753 , w2754 , w2755 , w2756 , w2757 , w2758 , w2759 , w2760 , w2761 , w2762 , w2763 , w2764 , w2765 , w2766 , w2767 , w2768 , w2769 , w2770 , w2771 , w2772 , w2773 , w2774 , w2775 , w2776 , w2777 , w2778 , w2779 , w2780 , w2781 , w2782 , w2783 , w2784 , w2785 , w2786 , w2787 , w2788 , w2789 , w2790 , w2791 , w2792 , w2793 , w2794 , w2795 , w2796 , w2797 , w2798 , w2799 , w2800 , w2801 , w2802 , w2803 , w2804 , w2805 , w2806 , w2807 , w2808 , w2809 , w2810 , w2811 , w2812 , w2813 , w2814 , w2815 , w2816 , w2817 , w2818 , w2819 , w2820 , w2821 , w2822 , w2823 , w2824 , w2825 , w2826 , w2827 , w2828 , w2829 , w2830 , w2831 , w2832 , w2833 , w2834 , w2835 , w2836 , w2837 , w2838 , w2839 , w2840 , w2841 , w2842 , w2843 , w2844 , w2845 , w2846 , w2847 , w2848 , w2849 , w2850 , w2851 , w2852 , w2853 , w2854 , w2855 , w2856 , w2857 , w2858 , w2859 , w2860 , w2861 , w2862 , w2863 , w2864 , w2865 , w2866 , w2867 , w2868 , w2869 , w2870 , w2871 , w2872 , w2873 , w2874 , w2875 , w2876 , w2877 , w2878 , w2879 , w2880 , w2881 , w2882 , w2883 , w2884 , w2885 , w2886 , w2887 , w2888 , w2889 , w2890 , w2891 , w2892 , w2893 , w2894 , w2895 , w2896 , w2897 , w2898 , w2899 , w2900 , w2901 , w2902 , w2903 , w2904 , w2905 , w2906 , w2907 , w2908 , w2909 , w2910 , w2911 , w2912 , w2913 , w2914 , w2915 , w2916 , w2917 , w2918 , w2919 , w2920 , w2921 , w2922 , w2923 , w2924 , w2925 , w2926 , w2927 , w2928 , w2929 , w2930 , w2931 , w2932 , w2933 , w2934 , w2935 , w2936 , w2937 , w2938 , w2939 , w2940 , w2941 , w2942 , w2943 , w2944 , w2945 , w2946 , w2947 , w2948 , w2949 , w2950 , w2951 , w2952 , w2953 , w2954 , w2955 , w2956 , w2957 , w2958 , w2959 , w2960 , w2961 , w2962 , w2963 , w2964 , w2965 , w2966 , w2967 , w2968 , w2969 , w2970 , w2971 , w2972 , w2973 , w2974 , w2975 , w2976 , w2977 , w2978 , w2979 , w2980 , w2981 , w2982 , w2983 , w2984 , w2985 , w2986 , w2987 , w2988 , w2989 , w2990 , w2991 , w2992 , w2993 , w2994 , w2995 , w2996 , w2997 , w2998 , w2999 , w3000 , w3001 , w3002 , w3003 , w3004 , w3005 , w3006 , w3007 , w3008 , w3009 , w3010 , w3011 , w3012 , w3013 , w3014 , w3015 , w3016 , w3017 , w3018 , w3019 , w3020 , w3021 , w3022 , w3023 , w3024 , w3025 , w3026 , w3027 , w3028 , w3029 , w3030 , w3031 , w3032 , w3033 , w3034 , w3035 , w3036 , w3037 , w3038 , w3039 , w3040 , w3041 , w3042 , w3043 , w3044 , w3045 , w3046 , w3047 , w3048 , w3049 , w3050 , w3051 , w3052 , w3053 , w3054 , w3055 , w3056 , w3057 , w3058 , w3059 , w3060 , w3061 , w3062 , w3063 , w3064 , w3065 , w3066 , w3067 , w3068 , w3069 , w3070 , w3071 , w3072 , w3073 , w3074 , w3075 , w3076 , w3077 , w3078 , w3079 , w3080 , w3081 , w3082 , w3083 , w3084 , w3085 , w3086 , w3087 , w3088 , w3089 , w3090 , w3091 , w3092 , w3093 , w3094 , w3095 , w3096 , w3097 , w3098 , w3099 , w3100 , w3101 , w3102 , w3103 , w3104 , w3105 , w3106 , w3107 , w3108 , w3109 , w3110 , w3111 , w3112 , w3113 , w3114 , w3115 , w3116 , w3117 , w3118 , w3119 , w3120 , w3121 , w3122 , w3123 , w3124 , w3125 , w3126 , w3127 , w3128 , w3129 , w3130 , w3131 , w3132 , w3133 , w3134 , w3135 , w3136 , w3137 , w3138 , w3139 , w3140 , w3141 , w3142 , w3143 , w3144 , w3145 , w3146 , w3147 , w3148 , w3149 , w3150 , w3151 , w3152 , w3153 , w3154 , w3155 , w3156 , w3157 , w3158 , w3159 , w3160 , w3161 , w3162 , w3163 , w3164 , w3165 , w3166 , w3167 , w3168 , w3169 , w3170 , w3171 , w3172 , w3173 , w3174 , w3175 , w3176 , w3177 , w3178 , w3179 , w3180 , w3181 , w3182 , w3183 , w3184 , w3185 , w3186 , w3187 , w3188 , w3189 , w3190 , w3191 , w3192 , w3193 , w3194 , w3195 , w3196 , w3197 , w3198 , w3199 , w3200 , w3201 , w3202 , w3203 , w3204 , w3205 , w3206 , w3207 , w3208 , w3209 , w3210 , w3211 , w3212 , w3213 , w3214 , w3215 , w3216 , w3217 , w3218 , w3219 , w3220 , w3221 , w3222 , w3223 , w3224 , w3225 , w3226 , w3227 , w3228 , w3229 , w3230 , w3231 , w3232 , w3233 , w3234 , w3235 , w3236 , w3237 , w3238 , w3239 , w3240 , w3241 , w3242 , w3243 , w3244 , w3245 , w3246 , w3247 , w3248 , w3249 , w3250 , w3251 , w3252 , w3253 , w3254 , w3255 , w3256 , w3257 , w3258 , w3259 , w3260 , w3261 , w3262 , w3263 , w3264 , w3265 , w3266 , w3267 , w3268 , w3269 , w3270 , w3271 , w3272 , w3273 , w3274 , w3275 , w3276 , w3277 , w3278 , w3279 , w3280 , w3281 , w3282 , w3283 , w3284 , w3285 , w3286 , w3287 , w3288 , w3289 , w3290 , w3291 , w3292 , w3293 , w3294 , w3295 , w3296 , w3297 , w3298 , w3299 , w3300 , w3301 , w3302 , w3303 , w3304 , w3305 , w3306 , w3307 , w3308 , w3309 , w3310 , w3311 , w3312 , w3313 , w3314 , w3315 , w3316 , w3317 , w3318 , w3319 , w3320 , w3321 , w3322 , w3323 , w3324 , w3325 , w3326 , w3327 , w3328 , w3329 , w3330 , w3331 , w3332 , w3333 , w3334 , w3335 , w3336 , w3337 , w3338 , w3339 , w3340 , w3341 , w3342 , w3343 , w3344 , w3345 , w3346 , w3347 , w3348 , w3349 , w3350 , w3351 , w3352 , w3353 , w3354 , w3355 , w3356 , w3357 , w3358 , w3359 , w3360 , w3361 , w3362 , w3363 , w3364 , w3365 , w3366 , w3367 , w3368 , w3369 , w3370 , w3371 , w3372 , w3373 , w3374 , w3375 , w3376 , w3377 , w3378 , w3379 , w3380 , w3381 , w3382 , w3383 , w3384 , w3385 , w3386 , w3387 , w3388 , w3389 , w3390 , w3391 , w3392 , w3393 , w3394 , w3395 , w3396 , w3397 , w3398 , w3399 , w3400 , w3401 , w3402 , w3403 , w3404 , w3405 , w3406 , w3407 , w3408 , w3409 , w3410 , w3411 , w3412 , w3413 , w3414 , w3415 , w3416 , w3417 , w3418 , w3419 , w3420 , w3421 , w3422 , w3423 , w3424 , w3425 , w3426 , w3427 , w3428 , w3429 , w3430 , w3431 , w3432 , w3433 , w3434 , w3435 , w3436 , w3437 , w3438 , w3439 , w3440 , w3441 , w3442 , w3443 , w3444 , w3445 , w3446 , w3447 , w3448 , w3449 , w3450 , w3451 , w3452 , w3453 , w3454 , w3455 , w3456 , w3457 , w3458 , w3459 , w3460 , w3461 , w3462 , w3463 , w3464 , w3465 , w3466 , w3467 , w3468 , w3469 , w3470 , w3471 , w3472 , w3473 , w3474 , w3475 , w3476 , w3477 , w3478 , w3479 , w3480 , w3481 , w3482 , w3483 , w3484 , w3485 , w3486 , w3487 , w3488 , w3489 , w3490 , w3491 , w3492 , w3493 , w3494 , w3495 , w3496 , w3497 , w3498 , w3499 , w3500 , w3501 , w3502 , w3503 , w3504 , w3505 , w3506 , w3507 , w3508 , w3509 , w3510 , w3511 , w3512 , w3513 , w3514 , w3515 , w3516 , w3517 , w3518 , w3519 , w3520 , w3521 , w3522 , w3523 , w3524 , w3525 , w3526 , w3527 , w3528 , w3529 , w3530 , w3531 , w3532 , w3533 , w3534 , w3535 , w3536 , w3537 , w3538 , w3539 , w3540 , w3541 , w3542 , w3543 , w3544 , w3545 , w3546 , w3547 , w3548 , w3549 , w3550 , w3551 , w3552 , w3553 , w3554 , w3555 , w3556 , w3557 , w3558 , w3559 , w3560 , w3561 , w3562 , w3563 , w3564 , w3565 , w3566 , w3567 , w3568 , w3569 , w3570 , w3571 , w3572 , w3573 , w3574 , w3575 , w3576 , w3577 , w3578 , w3579 , w3580 , w3581 , w3582 , w3583 , w3584 , w3585 , w3586 , w3587 , w3588 , w3589 , w3590 , w3591 , w3592 , w3593 , w3594 , w3595 , w3596 , w3597 , w3598 , w3599 , w3600 , w3601 , w3602 , w3603 , w3604 , w3605 , w3606 , w3607 , w3608 , w3609 , w3610 , w3611 , w3612 , w3613 , w3614 , w3615 , w3616 , w3617 , w3618 , w3619 , w3620 , w3621 , w3622 , w3623 , w3624 , w3625 , w3626 , w3627 , w3628 , w3629 , w3630 , w3631 , w3632 , w3633 , w3634 , w3635 , w3636 , w3637 , w3638 , w3639 , w3640 , w3641 , w3642 , w3643 , w3644 , w3645 , w3646 , w3647 , w3648 , w3649 , w3650 , w3651 , w3652 , w3653 , w3654 , w3655 , w3656 , w3657 , w3658 , w3659 , w3660 , w3661 , w3662 , w3663 , w3664 , w3665 , w3666 , w3667 , w3668 , w3669 , w3670 , w3671 , w3672 , w3673 , w3674 , w3675 , w3676 , w3677 , w3678 , w3679 , w3680 , w3681 , w3682 , w3683 , w3684 , w3685 , w3686 , w3687 , w3688 , w3689 , w3690 , w3691 , w3692 , w3693 , w3694 , w3695 , w3696 , w3697 , w3698 , w3699 , w3700 , w3701 , w3702 , w3703 , w3704 , w3705 , w3706 , w3707 , w3708 , w3709 , w3710 , w3711 , w3712 , w3713 , w3714 , w3715 , w3716 , w3717 , w3718 , w3719 , w3720 , w3721 , w3722 , w3723 , w3724 , w3725 , w3726 , w3727 , w3728 , w3729 , w3730 , w3731 , w3732 , w3733 , w3734 , w3735 , w3736 , w3737 , w3738 , w3739 , w3740 , w3741 , w3742 , w3743 , w3744 , w3745 , w3746 , w3747 , w3748 , w3749 , w3750 , w3751 , w3752 , w3753 , w3754 , w3755 , w3756 , w3757 , w3758 , w3759 , w3760 , w3761 , w3762 , w3763 , w3764 , w3765 , w3766 , w3767 , w3768 , w3769 , w3770 , w3771 , w3772 , w3773 , w3774 , w3775 , w3776 , w3777 , w3778 , w3779 , w3780 , w3781 , w3782 , w3783 , w3784 , w3785 , w3786 , w3787 , w3788 , w3789 , w3790 , w3791 , w3792 , w3793 , w3794 , w3795 , w3796 , w3797 , w3798 , w3799 , w3800 , w3801 , w3802 , w3803 , w3804 , w3805 , w3806 , w3807 , w3808 , w3809 , w3810 , w3811 , w3812 , w3813 , w3814 , w3815 , w3816 , w3817 , w3818 , w3819 , w3820 , w3821 , w3822 , w3823 , w3824 , w3825 , w3826 , w3827 , w3828 , w3829 , w3830 , w3831 , w3832 , w3833 , w3834 , w3835 , w3836 , w3837 , w3838 , w3839 , w3840 , w3841 , w3842 , w3843 , w3844 , w3845 , w3846 , w3847 , w3848 , w3849 , w3850 , w3851 , w3852 , w3853 , w3854 , w3855 , w3856 , w3857 , w3858 , w3859 , w3860 , w3861 , w3862 , w3863 , w3864 , w3865 , w3866 , w3867 , w3868 , w3869 , w3870 , w3871 , w3872 , w3873 , w3874 , w3875 , w3876 , w3877 , w3878 , w3879 , w3880 , w3881 , w3882 , w3883 , w3884 , w3885 , w3886 , w3887 , w3888 , w3889 , w3890 , w3891 , w3892 , w3893 , w3894 , w3895 , w3896 , w3897 , w3898 , w3899 , w3900 , w3901 , w3902 , w3903 , w3904 , w3905 , w3906 , w3907 , w3908 , w3909 , w3910 , w3911 , w3912 , w3913 , w3914 , w3915 , w3916 , w3917 , w3918 , w3919 , w3920 , w3921 , w3922 , w3923 , w3924 , w3925 , w3926 , w3927 , w3928 , w3929 , w3930 , w3931 , w3932 , w3933 , w3934 , w3935 , w3936 , w3937 , w3938 , w3939 , w3940 , w3941 , w3942 , w3943 , w3944 , w3945 , w3946 , w3947 , w3948 , w3949 , w3950 , w3951 , w3952 , w3953 , w3954 , w3955 , w3956 , w3957 , w3958 , w3959 , w3960 , w3961 , w3962 , w3963 , w3964 , w3965 , w3966 , w3967 , w3968 , w3969 , w3970 , w3971 , w3972 , w3973 , w3974 , w3975 , w3976 , w3977 , w3978 , w3979 , w3980 , w3981 , w3982 , w3983 , w3984 , w3985 , w3986 , w3987 , w3988 , w3989 , w3990 , w3991 , w3992 , w3993 , w3994 , w3995 , w3996 , w3997 , w3998 , w3999 , w4000 , w4001 , w4002 , w4003 , w4004 , w4005 , w4006 , w4007 , w4008 , w4009 , w4010 , w4011 , w4012 , w4013 , w4014 , w4015 , w4016 , w4017 , w4018 , w4019 , w4020 , w4021 , w4022 , w4023 , w4024 , w4025 , w4026 , w4027 , w4028 , w4029 , w4030 , w4031 , w4032 , w4033 , w4034 , w4035 , w4036 , w4037 , w4038 , w4039 , w4040 , w4041 , w4042 , w4043 , w4044 , w4045 , w4046 , w4047 , w4048 , w4049 , w4050 , w4051 , w4052 , w4053 , w4054 , w4055 , w4056 , w4057 , w4058 , w4059 , w4060 , w4061 , w4062 , w4063 , w4064 , w4065 , w4066 , w4067 , w4068 , w4069 , w4070 , w4071 , w4072 , w4073 , w4074 , w4075 , w4076 , w4077 , w4078 , w4079 , w4080 , w4081 , w4082 , w4083 , w4084 , w4085 , w4086 , w4087 , w4088 , w4089 , w4090 , w4091 , w4092 , w4093 , w4094 , w4095 , w4096 , w4097 , w4098 , w4099 , w4100 , w4101 , w4102 , w4103 , w4104 , w4105 , w4106 , w4107 , w4108 , w4109 , w4110 , w4111 , w4112 , w4113 , w4114 , w4115 , w4116 , w4117 , w4118 , w4119 , w4120 , w4121 , w4122 , w4123 , w4124 , w4125 , w4126 , w4127 , w4128 , w4129 , w4130 , w4131 , w4132 , w4133 , w4134 , w4135 , w4136 , w4137 , w4138 , w4139 , w4140 , w4141 , w4142 , w4143 , w4144 , w4145 , w4146 , w4147 , w4148 , w4149 , w4150 , w4151 , w4152 , w4153 , w4154 , w4155 , w4156 , w4157 , w4158 , w4159 , w4160 , w4161 , w4162 , w4163 , w4164 , w4165 , w4166 , w4167 , w4168 , w4169 , w4170 , w4171 , w4172 , w4173 , w4174 , w4175 , w4176 , w4177 , w4178 , w4179 , w4180 , w4181 , w4182 , w4183 , w4184 , w4185 , w4186 , w4187 , w4188 , w4189 , w4190 , w4191 , w4192 , w4193 , w4194 , w4195 , w4196 , w4197 , w4198 , w4199 , w4200 , w4201 , w4202 , w4203 , w4204 , w4205 , w4206 , w4207 , w4208 , w4209 , w4210 , w4211 , w4212 , w4213 , w4214 , w4215 , w4216 , w4217 , w4218 , w4219 , w4220 , w4221 , w4222 , w4223 , w4224 , w4225 , w4226 , w4227 , w4228 , w4229 , w4230 , w4231 , w4232 , w4233 , w4234 , w4235 , w4236 , w4237 , w4238 , w4239 , w4240 , w4241 , w4242 , w4243 , w4244 , w4245 , w4246 , w4247 , w4248 , w4249 , w4250 , w4251 , w4252 , w4253 , w4254 , w4255 , w4256 , w4257 , w4258 , w4259 , w4260 , w4261 , w4262 , w4263 , w4264 , w4265 , w4266 , w4267 , w4268 , w4269 , w4270 , w4271 , w4272 , w4273 , w4274 , w4275 , w4276 , w4277 , w4278 , w4279 , w4280 , w4281 , w4282 , w4283 , w4284 , w4285 , w4286 , w4287 , w4288 , w4289 , w4290 , w4291 , w4292 , w4293 , w4294 , w4295 , w4296 , w4297 , w4298 , w4299 , w4300 , w4301 , w4302 , w4303 , w4304 , w4305 , w4306 , w4307 , w4308 , w4309 , w4310 , w4311 , w4312 , w4313 , w4314 , w4315 , w4316 , w4317 , w4318 , w4319 , w4320 , w4321 , w4322 , w4323 , w4324 , w4325 , w4326 , w4327 , w4328 , w4329 , w4330 , w4331 , w4332 , w4333 , w4334 , w4335 , w4336 , w4337 , w4338 , w4339 , w4340 , w4341 , w4342 , w4343 , w4344 , w4345 , w4346 , w4347 , w4348 , w4349 , w4350 , w4351 , w4352 , w4353 , w4354 , w4355 , w4356 , w4357 , w4358 , w4359 , w4360 , w4361 , w4362 , w4363 , w4364 , w4365 , w4366 , w4367 , w4368 , w4369 , w4370 , w4371 , w4372 , w4373 , w4374 , w4375 , w4376 , w4377 , w4378 , w4379 , w4380 , w4381 , w4382 , w4383 , w4384 , w4385 , w4386 , w4387 , w4388 , w4389 , w4390 , w4391 , w4392 , w4393 , w4394 , w4395 , w4396 , w4397 , w4398 , w4399 , w4400 , w4401 , w4402 , w4403 , w4404 , w4405 , w4406 , w4407 , w4408 , w4409 , w4410 , w4411 , w4412 , w4413 , w4414 , w4415 , w4416 , w4417 , w4418 , w4419 , w4420 , w4421 , w4422 , w4423 , w4424 , w4425 , w4426 , w4427 , w4428 , w4429 , w4430 , w4431 , w4432 , w4433 , w4434 , w4435 , w4436 , w4437 , w4438 , w4439 , w4440 , w4441 , w4442 , w4443 , w4444 , w4445 , w4446 , w4447 , w4448 , w4449 , w4450 , w4451 , w4452 , w4453 , w4454 , w4455 , w4456 , w4457 , w4458 , w4459 , w4460 , w4461 , w4462 , w4463 , w4464 , w4465 , w4466 , w4467 , w4468 , w4469 , w4470 , w4471 , w4472 , w4473 , w4474 , w4475 , w4476 , w4477 , w4478 , w4479 , w4480 , w4481 , w4482 , w4483 , w4484 , w4485 , w4486 , w4487 , w4488 , w4489 , w4490 , w4491 , w4492 , w4493 , w4494 , w4495 , w4496 , w4497 , w4498 , w4499 , w4500 , w4501 , w4502 , w4503 , w4504 , w4505 , w4506 , w4507 , w4508 , w4509 , w4510 , w4511 , w4512 , w4513 , w4514 , w4515 , w4516 , w4517 , w4518 , w4519 , w4520 , w4521 , w4522 , w4523 , w4524 , w4525 , w4526 , w4527 , w4528 , w4529 , w4530 , w4531 , w4532 , w4533 , w4534 , w4535 , w4536 , w4537 , w4538 , w4539 , w4540 , w4541 , w4542 , w4543 , w4544 , w4545 , w4546 , w4547 , w4548 , w4549 , w4550 , w4551 , w4552 , w4553 , w4554 , w4555 , w4556 , w4557 , w4558 , w4559 , w4560 , w4561 , w4562 , w4563 , w4564 , w4565 , w4566 , w4567 , w4568 , w4569 , w4570 , w4571 , w4572 , w4573 , w4574 , w4575 , w4576 , w4577 , w4578 , w4579 , w4580 , w4581 , w4582 , w4583 , w4584 , w4585 , w4586 , w4587 , w4588 , w4589 , w4590 , w4591 , w4592 , w4593 , w4594 , w4595 , w4596 , w4597 , w4598 , w4599 , w4600 , w4601 , w4602 , w4603 , w4604 , w4605 , w4606 , w4607 , w4608 , w4609 , w4610 , w4611 , w4612 , w4613 , w4614 , w4615 , w4616 , w4617 , w4618 , w4619 , w4620 , w4621 , w4622 , w4623 , w4624 , w4625 , w4626 , w4627 , w4628 , w4629 , w4630 , w4631 , w4632 , w4633 , w4634 , w4635 , w4636 , w4637 , w4638 , w4639 , w4640 , w4641 , w4642 , w4643 , w4644 , w4645 , w4646 , w4647 , w4648 , w4649 , w4650 , w4651 , w4652 , w4653 , w4654 , w4655 , w4656 , w4657 , w4658 , w4659 , w4660 , w4661 , w4662 , w4663 , w4664 , w4665 , w4666 , w4667 , w4668 , w4669 , w4670 , w4671 , w4672 , w4673 , w4674 , w4675 , w4676 , w4677 , w4678 , w4679 , w4680 , w4681 , w4682 , w4683 , w4684 , w4685 , w4686 , w4687 , w4688 , w4689 , w4690 , w4691 , w4692 , w4693 , w4694 , w4695 , w4696 , w4697 , w4698 , w4699 , w4700 , w4701 , w4702 , w4703 , w4704 , w4705 , w4706 , w4707 , w4708 , w4709 , w4710 , w4711 , w4712 , w4713 , w4714 , w4715 , w4716 , w4717 , w4718 , w4719 , w4720 , w4721 , w4722 , w4723 , w4724 , w4725 , w4726 , w4727 , w4728 , w4729 , w4730 , w4731 , w4732 , w4733 , w4734 , w4735 , w4736 , w4737 , w4738 , w4739 , w4740 , w4741 , w4742 , w4743 , w4744 , w4745 , w4746 , w4747 , w4748 , w4749 , w4750 , w4751 , w4752 , w4753 , w4754 , w4755 , w4756 , w4757 , w4758 , w4759 , w4760 , w4761 , w4762 , w4763 , w4764 , w4765 , w4766 , w4767 , w4768 , w4769 , w4770 , w4771 , w4772 , w4773 , w4774 , w4775 , w4776 , w4777 , w4778 , w4779 , w4780 , w4781 , w4782 , w4783 , w4784 , w4785 , w4786 , w4787 , w4788 , w4789 , w4790 , w4791 , w4792 , w4793 , w4794 , w4795 , w4796 , w4797 , w4798 , w4799 , w4800 , w4801 , w4802 , w4803 , w4804 , w4805 , w4806 , w4807 , w4808 , w4809 , w4810 , w4811 , w4812 , w4813 , w4814 , w4815 , w4816 , w4817 , w4818 , w4819 , w4820 , w4821 , w4822 , w4823 , w4824 , w4825 , w4826 , w4827 , w4828 , w4829 , w4830 , w4831 , w4832 , w4833 , w4834 , w4835 , w4836 , w4837 , w4838 , w4839 , w4840 , w4841 , w4842 , w4843 , w4844 , w4845 , w4846 , w4847 , w4848 , w4849 , w4850 , w4851 , w4852 , w4853 , w4854 , w4855 , w4856 , w4857 , w4858 , w4859 , w4860 , w4861 , w4862 , w4863 , w4864 , w4865 , w4866 , w4867 , w4868 , w4869 , w4870 , w4871 , w4872 , w4873 , w4874 , w4875 , w4876 , w4877 , w4878 , w4879 , w4880 , w4881 , w4882 , w4883 , w4884 , w4885 , w4886 , w4887 , w4888 , w4889 , w4890 , w4891 , w4892 , w4893 , w4894 , w4895 , w4896 , w4897 , w4898 , w4899 , w4900 , w4901 , w4902 , w4903 , w4904 , w4905 , w4906 , w4907 , w4908 , w4909 , w4910 , w4911 , w4912 , w4913 , w4914 , w4915 , w4916 , w4917 , w4918 , w4919 , w4920 , w4921 , w4922 , w4923 , w4924 , w4925 , w4926 , w4927 , w4928 , w4929 , w4930 , w4931 , w4932 , w4933 , w4934 , w4935 , w4936 , w4937 , w4938 , w4939 , w4940 , w4941 , w4942 , w4943 , w4944 , w4945 , w4946 , w4947 , w4948 , w4949 , w4950 , w4951 , w4952 , w4953 , w4954 , w4955 , w4956 , w4957 , w4958 , w4959 , w4960 , w4961 , w4962 , w4963 , w4964 , w4965 , w4966 , w4967 , w4968 , w4969 , w4970 , w4971 , w4972 , w4973 , w4974 , w4975 , w4976 , w4977 , w4978 , w4979 , w4980 , w4981 , w4982 , w4983 , w4984 , w4985 , w4986 , w4987 , w4988 , w4989 , w4990 , w4991 , w4992 , w4993 , w4994 , w4995 , w4996 , w4997 , w4998 , w4999 , w5000 , w5001 , w5002 , w5003 , w5004 , w5005 , w5006 , w5007 , w5008 , w5009 , w5010 , w5011 , w5012 , w5013 , w5014 , w5015 , w5016 , w5017 , w5018 , w5019 , w5020 , w5021 , w5022 , w5023 , w5024 , w5025 , w5026 , w5027 , w5028 , w5029 , w5030 , w5031 , w5032 , w5033 , w5034 , w5035 , w5036 , w5037 , w5038 , w5039 , w5040 , w5041 , w5042 , w5043 , w5044 , w5045 , w5046 , w5047 , w5048 , w5049 , w5050 , w5051 , w5052 , w5053 , w5054 , w5055 , w5056 , w5057 , w5058 , w5059 , w5060 , w5061 , w5062 , w5063 , w5064 , w5065 , w5066 , w5067 , w5068 , w5069 , w5070 , w5071 , w5072 , w5073 , w5074 , w5075 , w5076 , w5077 , w5078 , w5079 , w5080 , w5081 , w5082 , w5083 , w5084 , w5085 , w5086 , w5087 , w5088 , w5089 , w5090 , w5091 , w5092 , w5093 , w5094 , w5095 , w5096 , w5097 , w5098 , w5099 , w5100 , w5101 , w5102 , w5103 , w5104 , w5105 , w5106 , w5107 , w5108 , w5109 , w5110 , w5111 , w5112 , w5113 , w5114 , w5115 , w5116 , w5117 , w5118 , w5119 , w5120 , w5121 , w5122 , w5123 , w5124 , w5125 , w5126 , w5127 , w5128 , w5129 , w5130 , w5131 , w5132 , w5133 , w5134 , w5135 , w5136 , w5137 , w5138 , w5139 , w5140 , w5141 , w5142 , w5143 , w5144 , w5145 , w5146 , w5147 , w5148 , w5149 , w5150 , w5151 , w5152 , w5153 , w5154 , w5155 , w5156 , w5157 , w5158 , w5159 , w5160 , w5161 , w5162 , w5163 , w5164 , w5165 , w5166 , w5167 , w5168 , w5169 , w5170 , w5171 , w5172 , w5173 , w5174 , w5175 , w5176 , w5177 , w5178 , w5179 , w5180 , w5181 , w5182 , w5183 , w5184 , w5185 , w5186 , w5187 , w5188 , w5189 , w5190 , w5191 , w5192 , w5193 , w5194 , w5195 , w5196 , w5197 , w5198 , w5199 , w5200 , w5201 , w5202 , w5203 , w5204 , w5205 , w5206 , w5207 , w5208 , w5209 , w5210 , w5211 , w5212 , w5213 , w5214 , w5215 , w5216 , w5217 , w5218 , w5219 , w5220 , w5221 , w5222 , w5223 , w5224 , w5225 , w5226 , w5227 , w5228 , w5229 , w5230 , w5231 , w5232 , w5233 , w5234 , w5235 , w5236 , w5237 , w5238 , w5239 , w5240 , w5241 , w5242 , w5243 , w5244 , w5245 , w5246 , w5247 , w5248 , w5249 , w5250 , w5251 , w5252 , w5253 , w5254 , w5255 , w5256 , w5257 , w5258 , w5259 , w5260 , w5261 , w5262 , w5263 , w5264 , w5265 , w5266 , w5267 , w5268 , w5269 , w5270 , w5271 , w5272 , w5273 , w5274 , w5275 , w5276 , w5277 , w5278 , w5279 , w5280 , w5281 , w5282 , w5283 , w5284 , w5285 , w5286 , w5287 , w5288 , w5289 , w5290 , w5291 , w5292 , w5293 , w5294 , w5295 , w5296 , w5297 , w5298 , w5299 , w5300 , w5301 , w5302 , w5303 , w5304 , w5305 , w5306 , w5307 , w5308 , w5309 , w5310 , w5311 , w5312 , w5313 , w5314 , w5315 , w5316 , w5317 , w5318 , w5319 , w5320 , w5321 , w5322 , w5323 , w5324 , w5325 , w5326 , w5327 , w5328 , w5329 , w5330 , w5331 , w5332 , w5333 , w5334 , w5335 , w5336 , w5337 , w5338 , w5339 , w5340 , w5341 , w5342 , w5343 , w5344 , w5345 , w5346 , w5347 , w5348 , w5349 , w5350 , w5351 , w5352 , w5353 , w5354 , w5355 , w5356 , w5357 , w5358 , w5359 , w5360 , w5361 , w5362 , w5363 , w5364 , w5365 , w5366 , w5367 , w5368 , w5369 , w5370 , w5371 , w5372 , w5373 , w5374 , w5375 , w5376 , w5377 , w5378 , w5379 , w5380 , w5381 , w5382 , w5383 , w5384 , w5385 , w5386 , w5387 , w5388 , w5389 , w5390 , w5391 , w5392 , w5393 , w5394 , w5395 , w5396 , w5397 , w5398 , w5399 , w5400 , w5401 , w5402 , w5403 , w5404 , w5405 , w5406 , w5407 , w5408 , w5409 , w5410 , w5411 , w5412 , w5413 , w5414 , w5415 , w5416 , w5417 , w5418 , w5419 , w5420 , w5421 , w5422 , w5423 , w5424 , w5425 , w5426 , w5427 , w5428 , w5429 , w5430 , w5431 , w5432 , w5433 , w5434 , w5435 , w5436 , w5437 , w5438 , w5439 , w5440 , w5441 , w5442 , w5443 , w5444 , w5445 , w5446 , w5447 , w5448 , w5449 , w5450 , w5451 , w5452 , w5453 , w5454 , w5455 , w5456 , w5457 , w5458 , w5459 , w5460 , w5461 , w5462 , w5463 , w5464 , w5465 , w5466 , w5467 , w5468 , w5469 , w5470 , w5471 , w5472 , w5473 , w5474 , w5475 , w5476 , w5477 , w5478 , w5479 , w5480 , w5481 , w5482 , w5483 , w5484 , w5485 , w5486 , w5487 , w5488 , w5489 , w5490 , w5491 , w5492 , w5493 , w5494 , w5495 , w5496 , w5497 , w5498 , w5499 , w5500 , w5501 , w5502 , w5503 , w5504 , w5505 , w5506 , w5507 , w5508 , w5509 , w5510 , w5511 , w5512 , w5513 , w5514 , w5515 , w5516 , w5517 , w5518 , w5519 , w5520 , w5521 , w5522 , w5523 , w5524 , w5525 , w5526 , w5527 , w5528 , w5529 , w5530 , w5531 , w5532 , w5533 , w5534 , w5535 , w5536 , w5537 , w5538 , w5539 , w5540 , w5541 , w5542 , w5543 , w5544 , w5545 , w5546 , w5547 , w5548 , w5549 , w5550 , w5551 , w5552 , w5553 , w5554 , w5555 , w5556 , w5557 , w5558 , w5559 , w5560 , w5561 , w5562 , w5563 , w5564 , w5565 , w5566 , w5567 , w5568 , w5569 , w5570 , w5571 , w5572 , w5573 , w5574 , w5575 , w5576 , w5577 , w5578 , w5579 , w5580 , w5581 , w5582 , w5583 , w5584 , w5585 , w5586 , w5587 , w5588 , w5589 , w5590 , w5591 , w5592 , w5593 , w5594 , w5595 , w5596 , w5597 , w5598 , w5599 , w5600 , w5601 , w5602 , w5603 , w5604 , w5605 , w5606 , w5607 , w5608 , w5609 , w5610 , w5611 , w5612 , w5613 , w5614 , w5615 , w5616 , w5617 , w5618 , w5619 , w5620 , w5621 , w5622 , w5623 , w5624 , w5625 , w5626 , w5627 , w5628 , w5629 , w5630 , w5631 , w5632 , w5633 , w5634 , w5635 , w5636 , w5637 , w5638 , w5639 , w5640 , w5641 , w5642 , w5643 , w5644 , w5645 , w5646 , w5647 , w5648 , w5649 , w5650 , w5651 , w5652 , w5653 , w5654 , w5655 , w5656 , w5657 , w5658 , w5659 , w5660 , w5661 , w5662 , w5663 , w5664 , w5665 , w5666 , w5667 , w5668 , w5669 , w5670 , w5671 , w5672 , w5673 , w5674 , w5675 , w5676 , w5677 , w5678 , w5679 , w5680 , w5681 , w5682 , w5683 , w5684 , w5685 , w5686 , w5687 , w5688 , w5689 , w5690 , w5691 , w5692 , w5693 , w5694 , w5695 , w5696 , w5697 , w5698 , w5699 , w5700 , w5701 , w5702 , w5703 , w5704 , w5705 , w5706 , w5707 , w5708 , w5709 , w5710 , w5711 , w5712 , w5713 , w5714 , w5715 , w5716 , w5717 , w5718 , w5719 , w5720 , w5721 , w5722 , w5723 , w5724 , w5725 , w5726 , w5727 , w5728 , w5729 , w5730 , w5731 , w5732 , w5733 , w5734 , w5735 , w5736 , w5737 , w5738 , w5739 , w5740 , w5741 , w5742 , w5743 , w5744 , w5745 , w5746 , w5747 , w5748 , w5749 , w5750 , w5751 , w5752 , w5753 , w5754 , w5755 , w5756 , w5757 , w5758 , w5759 , w5760 , w5761 , w5762 , w5763 , w5764 , w5765 , w5766 , w5767 , w5768 , w5769 , w5770 , w5771 , w5772 , w5773 , w5774 , w5775 , w5776 , w5777 , w5778 , w5779 , w5780 , w5781 , w5782 , w5783 , w5784 , w5785 , w5786 , w5787 , w5788 , w5789 , w5790 , w5791 , w5792 , w5793 , w5794 , w5795 , w5796 , w5797 , w5798 , w5799 , w5800 , w5801 , w5802 , w5803 , w5804 , w5805 , w5806 , w5807 , w5808 , w5809 , w5810 , w5811 , w5812 , w5813 , w5814 , w5815 , w5816 , w5817 , w5818 , w5819 , w5820 , w5821 , w5822 , w5823 , w5824 , w5825 , w5826 , w5827 , w5828 , w5829 , w5830 , w5831 , w5832 , w5833 , w5834 , w5835 , w5836 , w5837 , w5838 , w5839 , w5840 , w5841 , w5842 , w5843 , w5844 , w5845 , w5846 , w5847 , w5848 , w5849 , w5850 , w5851 , w5852 , w5853 , w5854 , w5855 , w5856 , w5857 , w5858 , w5859 , w5860 , w5861 , w5862 , w5863 , w5864 , w5865 , w5866 , w5867 , w5868 , w5869 , w5870 , w5871 , w5872 , w5873 , w5874 , w5875 , w5876 , w5877 , w5878 , w5879 , w5880 , w5881 , w5882 , w5883 , w5884 , w5885 , w5886 , w5887 , w5888 , w5889 , w5890 , w5891 , w5892 , w5893 , w5894 , w5895 , w5896 , w5897 , w5898 , w5899 , w5900 , w5901 , w5902 , w5903 , w5904 , w5905 , w5906 , w5907 , w5908 , w5909 , w5910 , w5911 , w5912 , w5913 , w5914 , w5915 , w5916 , w5917 , w5918 , w5919 , w5920 , w5921 , w5922 , w5923 , w5924 , w5925 , w5926 , w5927 , w5928 , w5929 , w5930 , w5931 , w5932 , w5933 , w5934 , w5935 , w5936 , w5937 , w5938 , w5939 , w5940 , w5941 , w5942 , w5943 , w5944 , w5945 , w5946 , w5947 , w5948 , w5949 , w5950 , w5951 , w5952 , w5953 , w5954 , w5955 , w5956 , w5957 , w5958 , w5959 , w5960 , w5961 , w5962 , w5963 , w5964 , w5965 , w5966 , w5967 , w5968 , w5969 , w5970 , w5971 , w5972 , w5973 , w5974 , w5975 , w5976 , w5977 , w5978 , w5979 , w5980 , w5981 , w5982 , w5983 , w5984 , w5985 , w5986 , w5987 , w5988 , w5989 , w5990 , w5991 , w5992 , w5993 , w5994 , w5995 , w5996 , w5997 , w5998 , w5999 , w6000 , w6001 , w6002 , w6003 , w6004 , w6005 , w6006 , w6007 , w6008 , w6009 , w6010 , w6011 , w6012 , w6013 , w6014 , w6015 , w6016 , w6017 , w6018 , w6019 , w6020 , w6021 , w6022 , w6023 , w6024 , w6025 , w6026 , w6027 , w6028 , w6029 , w6030 , w6031 , w6032 , w6033 , w6034 , w6035 , w6036 , w6037 , w6038 , w6039 , w6040 , w6041 , w6042 , w6043 , w6044 , w6045 , w6046 , w6047 , w6048 , w6049 , w6050 , w6051 , w6052 , w6053 , w6054 , w6055 , w6056 , w6057 , w6058 , w6059 , w6060 , w6061 , w6062 , w6063 , w6064 , w6065 , w6066 , w6067 , w6068 , w6069 , w6070 , w6071 , w6072 , w6073 , w6074 , w6075 , w6076 , w6077 , w6078 , w6079 , w6080 , w6081 , w6082 , w6083 , w6084 , w6085 , w6086 , w6087 , w6088 , w6089 , w6090 , w6091 , w6092 , w6093 , w6094 , w6095 , w6096 , w6097 , w6098 , w6099 , w6100 , w6101 , w6102 , w6103 , w6104 , w6105 , w6106 , w6107 , w6108 , w6109 , w6110 , w6111 , w6112 , w6113 , w6114 , w6115 , w6116 , w6117 , w6118 , w6119 , w6120 , w6121 , w6122 , w6123 , w6124 , w6125 , w6126 , w6127 , w6128 , w6129 , w6130 , w6131 , w6132 , w6133 , w6134 , w6135 , w6136 , w6137 , w6138 , w6139 , w6140 , w6141 , w6142 , w6143 , w6144 , w6145 , w6146 , w6147 , w6148 , w6149 , w6150 , w6151 , w6152 , w6153 , w6154 , w6155 , w6156 , w6157 , w6158 , w6159 , w6160 , w6161 , w6162 , w6163 , w6164 , w6165 , w6166 , w6167 , w6168 , w6169 , w6170 , w6171 , w6172 , w6173 , w6174 , w6175 , w6176 , w6177 , w6178 , w6179 , w6180 , w6181 , w6182 , w6183 , w6184 , w6185 , w6186 , w6187 , w6188 , w6189 , w6190 , w6191 , w6192 , w6193 , w6194 , w6195 , w6196 , w6197 , w6198 , w6199 , w6200 , w6201 , w6202 , w6203 , w6204 , w6205 , w6206 , w6207 , w6208 , w6209 , w6210 , w6211 , w6212 , w6213 , w6214 , w6215 , w6216 , w6217 , w6218 , w6219 , w6220 , w6221 , w6222 , w6223 , w6224 , w6225 , w6226 , w6227 , w6228 , w6229 , w6230 , w6231 , w6232 , w6233 , w6234 , w6235 , w6236 , w6237 , w6238 , w6239 , w6240 , w6241 , w6242 , w6243 , w6244 , w6245 , w6246 , w6247 , w6248 , w6249 , w6250 , w6251 , w6252 , w6253 , w6254 , w6255 , w6256 , w6257 , w6258 , w6259 , w6260 , w6261 , w6262 , w6263 , w6264 , w6265 , w6266 , w6267 , w6268 , w6269 , w6270 , w6271 , w6272 , w6273 , w6274 , w6275 , w6276 , w6277 , w6278 , w6279 , w6280 , w6281 , w6282 , w6283 , w6284 , w6285 , w6286 , w6287 , w6288 , w6289 , w6290 , w6291 , w6292 , w6293 , w6294 , w6295 , w6296 , w6297 , w6298 , w6299 , w6300 , w6301 , w6302 , w6303 , w6304 , w6305 , w6306 , w6307 , w6308 , w6309 , w6310 , w6311 , w6312 , w6313 , w6314 , w6315 , w6316 , w6317 , w6318 , w6319 , w6320 , w6321 , w6322 , w6323 , w6324 , w6325 , w6326 , w6327 , w6328 , w6329 , w6330 , w6331 , w6332 , w6333 , w6334 , w6335 , w6336 , w6337 , w6338 , w6339 , w6340 , w6341 , w6342 , w6343 , w6344 , w6345 , w6346 , w6347 , w6348 , w6349 , w6350 , w6351 , w6352 , w6353 , w6354 , w6355 , w6356 , w6357 , w6358 , w6359 , w6360 , w6361 , w6362 , w6363 , w6364 , w6365 , w6366 , w6367 , w6368 , w6369 , w6370 , w6371 , w6372 , w6373 , w6374 , w6375 , w6376 , w6377 , w6378 , w6379 , w6380 , w6381 , w6382 , w6383 , w6384 , w6385 , w6386 , w6387 , w6388 , w6389 , w6390 , w6391 , w6392 , w6393 , w6394 , w6395 , w6396 , w6397 , w6398 , w6399 , w6400 , w6401 , w6402 , w6403 , w6404 , w6405 , w6406 , w6407 , w6408 , w6409 , w6410 , w6411 , w6412 , w6413 , w6414 , w6415 , w6416 , w6417 , w6418 , w6419 , w6420 , w6421 , w6422 , w6423 , w6424 , w6425 , w6426 , w6427 , w6428 , w6429 , w6430 , w6431 , w6432 , w6433 , w6434 , w6435 , w6436 , w6437 , w6438 , w6439 , w6440 , w6441 , w6442 , w6443 , w6444 , w6445 , w6446 , w6447 , w6448 , w6449 , w6450 , w6451 , w6452 , w6453 , w6454 , w6455 , w6456 , w6457 , w6458 , w6459 , w6460 , w6461 , w6462 , w6463 , w6464 , w6465 , w6466 , w6467 , w6468 , w6469 , w6470 , w6471 , w6472 , w6473 , w6474 , w6475 , w6476 , w6477 , w6478 , w6479 , w6480 , w6481 , w6482 , w6483 , w6484 , w6485 , w6486 , w6487 , w6488 , w6489 , w6490 , w6491 , w6492 , w6493 , w6494 , w6495 , w6496 , w6497 , w6498 , w6499 , w6500 , w6501 , w6502 , w6503 , w6504 , w6505 , w6506 , w6507 , w6508 , w6509 , w6510 , w6511 , w6512 , w6513 , w6514 , w6515 , w6516 , w6517 , w6518 , w6519 , w6520 , w6521 , w6522 , w6523 , w6524 , w6525 , w6526 , w6527 , w6528 , w6529 , w6530 , w6531 , w6532 , w6533 , w6534 , w6535 , w6536 , w6537 , w6538 , w6539 , w6540 , w6541 , w6542 , w6543 , w6544 , w6545 , w6546 , w6547 , w6548 , w6549 , w6550 , w6551 , w6552 , w6553 , w6554 , w6555 , w6556 , w6557 , w6558 , w6559 , w6560 , w6561 , w6562 , w6563 , w6564 , w6565 , w6566 , w6567 , w6568 , w6569 , w6570 , w6571 , w6572 , w6573 , w6574 , w6575 , w6576 , w6577 , w6578 , w6579 , w6580 , w6581 , w6582 , w6583 , w6584 , w6585 , w6586 , w6587 , w6588 , w6589 , w6590 , w6591 , w6592 , w6593 , w6594 , w6595 , w6596 , w6597 , w6598 , w6599 , w6600 , w6601 , w6602 , w6603 , w6604 , w6605 , w6606 , w6607 , w6608 , w6609 , w6610 , w6611 , w6612 , w6613 , w6614 , w6615 , w6616 , w6617 , w6618 , w6619 , w6620 , w6621 , w6622 , w6623 , w6624 , w6625 , w6626 , w6627 , w6628 , w6629 , w6630 , w6631 , w6632 , w6633 , w6634 , w6635 , w6636 , w6637 , w6638 , w6639 , w6640 , w6641 , w6642 , w6643 , w6644 , w6645 , w6646 , w6647 , w6648 , w6649 , w6650 , w6651 , w6652 , w6653 , w6654 , w6655 , w6656 , w6657 , w6658 , w6659 , w6660 , w6661 , w6662 , w6663 , w6664 , w6665 , w6666 , w6667 , w6668 , w6669 , w6670 , w6671 , w6672 , w6673 , w6674 , w6675 , w6676 , w6677 , w6678 , w6679 , w6680 , w6681 , w6682 , w6683 , w6684 , w6685 , w6686 , w6687 , w6688 , w6689 , w6690 , w6691 , w6692 , w6693 , w6694 , w6695 , w6696 , w6697 , w6698 , w6699 , w6700 , w6701 , w6702 , w6703 , w6704 , w6705 , w6706 , w6707 , w6708 , w6709 , w6710 , w6711 , w6712 , w6713 , w6714 , w6715 , w6716 , w6717 , w6718 , w6719 , w6720 , w6721 , w6722 , w6723 , w6724 , w6725 , w6726 , w6727 , w6728 , w6729 , w6730 , w6731 , w6732 , w6733 , w6734 , w6735 , w6736 , w6737 , w6738 , w6739 , w6740 , w6741 , w6742 , w6743 , w6744 , w6745 , w6746 , w6747 , w6748 , w6749 , w6750 , w6751 , w6752 , w6753 , w6754 , w6755 , w6756 , w6757 , w6758 , w6759 , w6760 , w6761 , w6762 , w6763 , w6764 , w6765 , w6766 , w6767 , w6768 , w6769 , w6770 , w6771 , w6772 , w6773 , w6774 , w6775 , w6776 , w6777 , w6778 , w6779 , w6780 , w6781 , w6782 , w6783 , w6784 , w6785 , w6786 , w6787 , w6788 , w6789 , w6790 , w6791 , w6792 , w6793 , w6794 , w6795 , w6796 , w6797 , w6798 , w6799 , w6800 , w6801 , w6802 , w6803 , w6804 , w6805 , w6806 , w6807 , w6808 , w6809 , w6810 , w6811 , w6812 , w6813 , w6814 , w6815 , w6816 , w6817 , w6818 , w6819 , w6820 , w6821 , w6822 , w6823 , w6824 , w6825 , w6826 , w6827 , w6828 , w6829 , w6830 , w6831 , w6832 , w6833 , w6834 , w6835 , w6836 , w6837 , w6838 , w6839 , w6840 , w6841 , w6842 , w6843 , w6844 , w6845 , w6846 , w6847 , w6848 , w6849 , w6850 , w6851 , w6852 , w6853 , w6854 , w6855 , w6856 , w6857 , w6858 , w6859 , w6860 , w6861 , w6862 , w6863 , w6864 , w6865 , w6866 , w6867 , w6868 , w6869 , w6870 , w6871 , w6872 , w6873 , w6874 , w6875 , w6876 , w6877 , w6878 , w6879 , w6880 , w6881 , w6882 , w6883 , w6884 , w6885 , w6886 , w6887 , w6888 , w6889 , w6890 , w6891 , w6892 , w6893 , w6894 , w6895 , w6896 , w6897 , w6898 , w6899 , w6900 , w6901 , w6902 , w6903 , w6904 , w6905 , w6906 , w6907 , w6908 , w6909 , w6910 , w6911 , w6912 , w6913 , w6914 , w6915 , w6916 , w6917 , w6918 , w6919 , w6920 , w6921 , w6922 , w6923 , w6924 , w6925 , w6926 , w6927 , w6928 , w6929 , w6930 , w6931 , w6932 , w6933 , w6934 , w6935 , w6936 , w6937 , w6938 , w6939 , w6940 , w6941 , w6942 , w6943 , w6944 , w6945 , w6946 , w6947 , w6948 , w6949 , w6950 , w6951 , w6952 , w6953 , w6954 , w6955 , w6956 , w6957 , w6958 , w6959 , w6960 , w6961 , w6962 , w6963 , w6964 , w6965 , w6966 , w6967 , w6968 , w6969 , w6970 , w6971 , w6972 , w6973 , w6974 , w6975 , w6976 , w6977 , w6978 , w6979 , w6980 , w6981 , w6982 , w6983 , w6984 , w6985 , w6986 , w6987 , w6988 , w6989 , w6990 , w6991 , w6992 , w6993 , w6994 , w6995 , w6996 , w6997 , w6998 , w6999 , w7000 , w7001 , w7002 , w7003 , w7004 , w7005 , w7006 , w7007 , w7008 , w7009 , w7010 , w7011 , w7012 , w7013 , w7014 , w7015 , w7016 , w7017 , w7018 , w7019 , w7020 , w7021 , w7022 , w7023 , w7024 , w7025 , w7026 , w7027 , w7028 , w7029 , w7030 , w7031 , w7032 , w7033 , w7034 , w7035 , w7036 , w7037 , w7038 , w7039 , w7040 , w7041 , w7042 , w7043 , w7044 , w7045 , w7046 , w7047 , w7048 , w7049 , w7050 , w7051 , w7052 , w7053 , w7054 , w7055 , w7056 , w7057 , w7058 , w7059 , w7060 , w7061 , w7062 , w7063 , w7064 , w7065 , w7066 , w7067 , w7068 , w7069 , w7070 , w7071 , w7072 , w7073 , w7074 , w7075 , w7076 , w7077 , w7078 , w7079 , w7080 , w7081 , w7082 , w7083 , w7084 , w7085 , w7086 , w7087 , w7088 , w7089 , w7090 , w7091 , w7092 , w7093 , w7094 , w7095 , w7096 , w7097 , w7098 , w7099 , w7100 , w7101 , w7102 , w7103 , w7104 , w7105 , w7106 , w7107 , w7108 , w7109 , w7110 , w7111 , w7112 , w7113 , w7114 , w7115 , w7116 , w7117 , w7118 , w7119 , w7120 , w7121 , w7122 , w7123 , w7124 , w7125 , w7126 , w7127 , w7128 , w7129 , w7130 , w7131 , w7132 , w7133 , w7134 , w7135 , w7136 , w7137 , w7138 , w7139 , w7140 , w7141 , w7142 , w7143 , w7144 , w7145 , w7146 , w7147 , w7148 , w7149 , w7150 , w7151 , w7152 , w7153 , w7154 , w7155 , w7156 , w7157 , w7158 , w7159 , w7160 , w7161 , w7162 , w7163 , w7164 , w7165 , w7166 , w7167 , w7168 , w7169 , w7170 , w7171 , w7172 , w7173 , w7174 , w7175 , w7176 , w7177 , w7178 , w7179 , w7180 , w7181 , w7182 , w7183 , w7184 , w7185 , w7186 , w7187 , w7188 , w7189 , w7190 , w7191 , w7192 , w7193 , w7194 , w7195 , w7196 , w7197 , w7198 , w7199 , w7200 , w7201 , w7202 , w7203 , w7204 , w7205 , w7206 , w7207 , w7208 , w7209 , w7210 , w7211 , w7212 , w7213 , w7214 , w7215 , w7216 , w7217 , w7218 , w7219 , w7220 , w7221 , w7222 , w7223 , w7224 , w7225 , w7226 , w7227 , w7228 , w7229 , w7230 , w7231 , w7232 , w7233 , w7234 , w7235 , w7236 , w7237 , w7238 , w7239 , w7240 , w7241 , w7242 , w7243 , w7244 , w7245 , w7246 , w7247 , w7248 , w7249 , w7250 , w7251 , w7252 , w7253 , w7254 , w7255 , w7256 , w7257 , w7258 , w7259 , w7260 , w7261 , w7262 , w7263 , w7264 , w7265 , w7266 , w7267 , w7268 , w7269 , w7270 , w7271 , w7272 , w7273 , w7274 , w7275 , w7276 , w7277 , w7278 , w7279 , w7280 , w7281 , w7282 , w7283 , w7284 , w7285 , w7286 , w7287 , w7288 , w7289 , w7290 , w7291 , w7292 , w7293 , w7294 , w7295 , w7296 , w7297 , w7298 , w7299 , w7300 , w7301 , w7302 , w7303 , w7304 , w7305 , w7306 , w7307 , w7308 , w7309 , w7310 , w7311 , w7312 , w7313 , w7314 , w7315 , w7316 , w7317 , w7318 , w7319 , w7320 , w7321 , w7322 , w7323 , w7324 , w7325 , w7326 , w7327 , w7328 , w7329 , w7330 , w7331 , w7332 , w7333 , w7334 , w7335 , w7336 , w7337 , w7338 , w7339 , w7340 , w7341 , w7342 , w7343 , w7344 , w7345 , w7346 , w7347 , w7348 , w7349 , w7350 , w7351 , w7352 , w7353 , w7354 , w7355 , w7356 , w7357 , w7358 , w7359 , w7360 , w7361 , w7362 , w7363 , w7364 , w7365 , w7366 , w7367 , w7368 , w7369 , w7370 , w7371 , w7372 , w7373 , w7374 , w7375 , w7376 , w7377 , w7378 , w7379 , w7380 , w7381 , w7382 , w7383 , w7384 , w7385 , w7386 , w7387 , w7388 , w7389 , w7390 , w7391 , w7392 , w7393 , w7394 , w7395 , w7396 , w7397 , w7398 , w7399 , w7400 , w7401 , w7402 , w7403 , w7404 , w7405 , w7406 , w7407 , w7408 , w7409 , w7410 , w7411 , w7412 , w7413 , w7414 , w7415 , w7416 , w7417 , w7418 , w7419 , w7420 , w7421 , w7422 , w7423 , w7424 , w7425 , w7426 , w7427 , w7428 , w7429 , w7430 , w7431 , w7432 , w7433 , w7434 , w7435 , w7436 , w7437 , w7438 , w7439 , w7440 , w7441 , w7442 , w7443 , w7444 , w7445 , w7446 , w7447 , w7448 , w7449 , w7450 , w7451 , w7452 , w7453 , w7454 , w7455 , w7456 , w7457 , w7458 , w7459 , w7460 , w7461 , w7462 , w7463 , w7464 , w7465 , w7466 , w7467 , w7468 , w7469 , w7470 , w7471 , w7472 , w7473 , w7474 , w7475 , w7476 , w7477 , w7478 , w7479 , w7480 , w7481 , w7482 , w7483 , w7484 , w7485 , w7486 , w7487 , w7488 , w7489 , w7490 , w7491 , w7492 , w7493 , w7494 , w7495 , w7496 , w7497 , w7498 , w7499 , w7500 , w7501 , w7502 , w7503 , w7504 , w7505 , w7506 , w7507 , w7508 , w7509 , w7510 , w7511 , w7512 , w7513 , w7514 , w7515 , w7516 , w7517 , w7518 , w7519 , w7520 , w7521 , w7522 , w7523 , w7524 , w7525 , w7526 , w7527 , w7528 , w7529 , w7530 , w7531 , w7532 , w7533 , w7534 , w7535 , w7536 , w7537 , w7538 , w7539 , w7540 , w7541 , w7542 , w7543 , w7544 , w7545 , w7546 , w7547 , w7548 , w7549 , w7550 , w7551 , w7552 , w7553 , w7554 , w7555 , w7556 , w7557 , w7558 , w7559 , w7560 , w7561 , w7562 , w7563 , w7564 , w7565 , w7566 , w7567 , w7568 , w7569 , w7570 , w7571 , w7572 , w7573 , w7574 , w7575 , w7576 , w7577 , w7578 , w7579 , w7580 , w7581 , w7582 , w7583 , w7584 , w7585 , w7586 , w7587 , w7588 , w7589 , w7590 , w7591 , w7592 , w7593 , w7594 , w7595 , w7596 , w7597 , w7598 , w7599 , w7600 , w7601 , w7602 , w7603 , w7604 , w7605 , w7606 , w7607 , w7608 , w7609 , w7610 , w7611 , w7612 , w7613 , w7614 , w7615 , w7616 , w7617 , w7618 , w7619 , w7620 , w7621 , w7622 , w7623 , w7624 , w7625 , w7626 , w7627 , w7628 , w7629 , w7630 , w7631 , w7632 , w7633 , w7634 , w7635 , w7636 , w7637 , w7638 , w7639 , w7640 , w7641 , w7642 , w7643 , w7644 , w7645 , w7646 , w7647 , w7648 , w7649 , w7650 , w7651 , w7652 , w7653 , w7654 , w7655 , w7656 , w7657 , w7658 , w7659 , w7660 , w7661 , w7662 , w7663 , w7664 , w7665 , w7666 , w7667 , w7668 , w7669 , w7670 , w7671 , w7672 , w7673 , w7674 , w7675 , w7676 , w7677 , w7678 , w7679 , w7680 , w7681 , w7682 , w7683 , w7684 , w7685 , w7686 , w7687 , w7688 , w7689 , w7690 , w7691 , w7692 , w7693 , w7694 , w7695 , w7696 , w7697 , w7698 , w7699 , w7700 , w7701 , w7702 , w7703 , w7704 , w7705 , w7706 , w7707 , w7708 , w7709 , w7710 , w7711 , w7712 , w7713 , w7714 , w7715 , w7716 , w7717 , w7718 , w7719 , w7720 , w7721 , w7722 , w7723 , w7724 , w7725 , w7726 , w7727 , w7728 , w7729 , w7730 , w7731 , w7732 , w7733 , w7734 , w7735 , w7736 , w7737 , w7738 , w7739 , w7740 , w7741 , w7742 , w7743 , w7744 , w7745 , w7746 , w7747 , w7748 , w7749 , w7750 , w7751 , w7752 , w7753 , w7754 , w7755 , w7756 , w7757 , w7758 , w7759 , w7760 , w7761 , w7762 , w7763 , w7764 , w7765 , w7766 , w7767 , w7768 , w7769 , w7770 , w7771 , w7772 , w7773 , w7774 , w7775 , w7776 , w7777 , w7778 , w7779 , w7780 , w7781 , w7782 , w7783 , w7784 , w7785 , w7786 , w7787 , w7788 , w7789 , w7790 , w7791 , w7792 , w7793 , w7794 , w7795 , w7796 , w7797 , w7798 , w7799 , w7800 , w7801 , w7802 , w7803 , w7804 , w7805 , w7806 , w7807 , w7808 , w7809 , w7810 , w7811 , w7812 , w7813 , w7814 , w7815 , w7816 , w7817 , w7818 , w7819 , w7820 , w7821 , w7822 , w7823 , w7824 , w7825 , w7826 , w7827 , w7828 , w7829 , w7830 , w7831 , w7832 , w7833 , w7834 , w7835 , w7836 , w7837 , w7838 , w7839 , w7840 , w7841 , w7842 , w7843 , w7844 , w7845 , w7846 , w7847 , w7848 , w7849 , w7850 , w7851 , w7852 , w7853 , w7854 , w7855 , w7856 , w7857 , w7858 , w7859 , w7860 , w7861 , w7862 , w7863 , w7864 , w7865 , w7866 , w7867 , w7868 , w7869 , w7870 , w7871 , w7872 , w7873 , w7874 , w7875 , w7876 , w7877 , w7878 , w7879 , w7880 , w7881 , w7882 , w7883 , w7884 , w7885 , w7886 , w7887 , w7888 , w7889 , w7890 , w7891 , w7892 , w7893 , w7894 , w7895 , w7896 , w7897 , w7898 , w7899 , w7900 , w7901 , w7902 , w7903 , w7904 , w7905 , w7906 , w7907 , w7908 , w7909 , w7910 , w7911 , w7912 , w7913 , w7914 , w7915 , w7916 , w7917 , w7918 , w7919 , w7920 , w7921 , w7922 , w7923 , w7924 , w7925 , w7926 , w7927 , w7928 , w7929 , w7930 , w7931 , w7932 , w7933 , w7934 , w7935 , w7936 , w7937 , w7938 , w7939 , w7940 , w7941 , w7942 , w7943 , w7944 , w7945 , w7946 , w7947 , w7948 , w7949 , w7950 , w7951 , w7952 , w7953 , w7954 , w7955 , w7956 , w7957 , w7958 , w7959 , w7960 , w7961 , w7962 , w7963 , w7964 , w7965 , w7966 , w7967 , w7968 , w7969 , w7970 , w7971 , w7972 , w7973 , w7974 , w7975 , w7976 , w7977 , w7978 , w7979 , w7980 , w7981 , w7982 , w7983 , w7984 , w7985 , w7986 , w7987 , w7988 , w7989 , w7990 , w7991 , w7992 , w7993 , w7994 , w7995 , w7996 , w7997 , w7998 , w7999 , w8000 , w8001 , w8002 , w8003 , w8004 , w8005 , w8006 , w8007 , w8008 , w8009 , w8010 , w8011 , w8012 , w8013 , w8014 , w8015 , w8016 , w8017 , w8018 , w8019 , w8020 , w8021 , w8022 , w8023 , w8024 , w8025 , w8026 , w8027 , w8028 , w8029 , w8030 , w8031 , w8032 , w8033 , w8034 , w8035 , w8036 , w8037 , w8038 , w8039 , w8040 , w8041 , w8042 , w8043 , w8044 , w8045 , w8046 , w8047 , w8048 , w8049 , w8050 , w8051 , w8052 , w8053 , w8054 , w8055 , w8056 , w8057 , w8058 , w8059 , w8060 , w8061 , w8062 , w8063 , w8064 , w8065 , w8066 , w8067 , w8068 , w8069 , w8070 , w8071 , w8072 , w8073 , w8074 , w8075 , w8076 , w8077 , w8078 , w8079 , w8080 , w8081 , w8082 , w8083 , w8084 , w8085 , w8086 , w8087 , w8088 , w8089 , w8090 , w8091 , w8092 , w8093 , w8094 , w8095 , w8096 , w8097 , w8098 , w8099 , w8100 , w8101 , w8102 , w8103 , w8104 , w8105 , w8106 , w8107 , w8108 , w8109 , w8110 , w8111 , w8112 , w8113 , w8114 , w8115 , w8116 , w8117 , w8118 , w8119 , w8120 , w8121 , w8122 , w8123 , w8124 , w8125 , w8126 , w8127 , w8128 , w8129 , w8130 , w8131 , w8132 , w8133 , w8134 , w8135 , w8136 , w8137 , w8138 , w8139 , w8140 , w8141 , w8142 , w8143 , w8144 , w8145 , w8146 , w8147 , w8148 , w8149 , w8150 , w8151 , w8152 , w8153 , w8154 , w8155 , w8156 , w8157 , w8158 , w8159 , w8160 , w8161 , w8162 , w8163 , w8164 , w8165 , w8166 , w8167 , w8168 , w8169 , w8170 , w8171 , w8172 , w8173 , w8174 , w8175 , w8176 , w8177 , w8178 , w8179 , w8180 , w8181 , w8182 , w8183 , w8184 , w8185 , w8186 , w8187 , w8188 , w8189 , w8190 , w8191 , w8192 , w8193 , w8194 , w8195 , w8196 , w8197 , w8198 , w8199 , w8200 , w8201 , w8202 , w8203 , w8204 , w8205 , w8206 , w8207 , w8208 , w8209 , w8210 , w8211 , w8212 , w8213 , w8214 , w8215 , w8216 , w8217 , w8218 , w8219 , w8220 , w8221 , w8222 , w8223 , w8224 , w8225 , w8226 , w8227 , w8228 , w8229 , w8230 , w8231 , w8232 , w8233 , w8234 , w8235 , w8236 , w8237 , w8238 , w8239 , w8240 , w8241 , w8242 , w8243 , w8244 , w8245 , w8246 , w8247 , w8248 , w8249 , w8250 , w8251 , w8252 , w8253 , w8254 , w8255 , w8256 , w8257 , w8258 , w8259 , w8260 , w8261 , w8262 , w8263 , w8264 , w8265 , w8266 , w8267 , w8268 , w8269 , w8270 , w8271 , w8272 , w8273 , w8274 , w8275 , w8276 , w8277 , w8278 , w8279 , w8280 , w8281 , w8282 , w8283 , w8284 , w8285 , w8286 , w8287 , w8288 , w8289 , w8290 , w8291 , w8292 , w8293 , w8294 , w8295 , w8296 , w8297 , w8298 , w8299 , w8300 , w8301 , w8302 , w8303 , w8304 , w8305 , w8306 , w8307 , w8308 , w8309 , w8310 , w8311 , w8312 , w8313 , w8314 , w8315 , w8316 , w8317 , w8318 , w8319 , w8320 , w8321 , w8322 , w8323 , w8324 , w8325 , w8326 , w8327 , w8328 , w8329 , w8330 , w8331 , w8332 , w8333 , w8334 , w8335 , w8336 , w8337 , w8338 , w8339 , w8340 , w8341 , w8342 , w8343 , w8344 , w8345 , w8346 , w8347 , w8348 , w8349 , w8350 , w8351 , w8352 , w8353 , w8354 , w8355 , w8356 , w8357 , w8358 , w8359 , w8360 , w8361 , w8362 , w8363 , w8364 , w8365 , w8366 , w8367 , w8368 , w8369 , w8370 , w8371 , w8372 , w8373 , w8374 , w8375 , w8376 , w8377 , w8378 , w8379 , w8380 , w8381 , w8382 , w8383 , w8384 , w8385 , w8386 , w8387 , w8388 , w8389 , w8390 , w8391 , w8392 , w8393 , w8394 , w8395 , w8396 , w8397 , w8398 , w8399 , w8400 , w8401 , w8402 , w8403 , w8404 , w8405 , w8406 , w8407 , w8408 , w8409 , w8410 , w8411 , w8412 , w8413 , w8414 , w8415 , w8416 , w8417 , w8418 , w8419 , w8420 , w8421 , w8422 , w8423 , w8424 , w8425 , w8426 , w8427 , w8428 , w8429 , w8430 , w8431 , w8432 , w8433 , w8434 , w8435 , w8436 , w8437 , w8438 , w8439 , w8440 , w8441 , w8442 , w8443 , w8444 , w8445 , w8446 , w8447 , w8448 , w8449 , w8450 , w8451 , w8452 , w8453 , w8454 , w8455 , w8456 , w8457 , w8458 , w8459 , w8460 , w8461 , w8462 , w8463 , w8464 , w8465 , w8466 , w8467 , w8468 , w8469 , w8470 , w8471 , w8472 , w8473 , w8474 , w8475 , w8476 , w8477 , w8478 , w8479 , w8480 , w8481 , w8482 , w8483 , w8484 , w8485 , w8486 , w8487 , w8488 , w8489 , w8490 , w8491 , w8492 , w8493 , w8494 , w8495 , w8496 , w8497 , w8498 , w8499 , w8500 , w8501 , w8502 , w8503 , w8504 , w8505 , w8506 , w8507 , w8508 , w8509 , w8510 , w8511 , w8512 , w8513 , w8514 , w8515 , w8516 , w8517 , w8518 , w8519 , w8520 , w8521 , w8522 , w8523 , w8524 , w8525 , w8526 , w8527 , w8528 , w8529 , w8530 , w8531 , w8532 , w8533 , w8534 , w8535 , w8536 , w8537 , w8538 , w8539 , w8540 , w8541 , w8542 , w8543 , w8544 , w8545 , w8546 , w8547 , w8548 , w8549 , w8550 , w8551 , w8552 , w8553 , w8554 , w8555 , w8556 , w8557 , w8558 , w8559 , w8560 , w8561 , w8562 , w8563 , w8564 , w8565 , w8566 , w8567 , w8568 , w8569 , w8570 , w8571 , w8572 , w8573 , w8574 , w8575 , w8576 , w8577 , w8578 , w8579 , w8580 , w8581 , w8582 , w8583 , w8584 , w8585 , w8586 , w8587 , w8588 , w8589 , w8590 , w8591 , w8592 , w8593 , w8594 , w8595 , w8596 , w8597 , w8598 , w8599 , w8600 , w8601 , w8602 , w8603 , w8604 , w8605 , w8606 , w8607 , w8608 , w8609 , w8610 , w8611 , w8612 , w8613 , w8614 , w8615 , w8616 , w8617 , w8618 , w8619 , w8620 , w8621 , w8622 , w8623 , w8624 , w8625 , w8626 , w8627 , w8628 , w8629 , w8630 , w8631 , w8632 , w8633 , w8634 , w8635 , w8636 , w8637 , w8638 , w8639 , w8640 , w8641 , w8642 , w8643 , w8644 , w8645 , w8646 , w8647 , w8648 , w8649 , w8650 , w8651 , w8652 , w8653 , w8654 , w8655 , w8656 , w8657 , w8658 , w8659 , w8660 , w8661 , w8662 , w8663 , w8664 , w8665 , w8666 , w8667 , w8668 , w8669 , w8670 , w8671 , w8672 , w8673 , w8674 , w8675 , w8676 , w8677 , w8678 , w8679 , w8680 , w8681 , w8682 , w8683 , w8684 , w8685 , w8686 , w8687 , w8688 , w8689 , w8690 , w8691 , w8692 , w8693 , w8694 , w8695 , w8696 , w8697 , w8698 , w8699 , w8700 , w8701 , w8702 , w8703 , w8704 , w8705 , w8706 , w8707 , w8708 , w8709 , w8710 , w8711 , w8712 , w8713 , w8714 , w8715 , w8716 , w8717 , w8718 , w8719 , w8720 , w8721 , w8722 , w8723 , w8724 , w8725 , w8726 , w8727 , w8728 , w8729 , w8730 , w8731 , w8732 , w8733 , w8734 , w8735 , w8736 , w8737 , w8738 , w8739 , w8740 , w8741 , w8742 , w8743 , w8744 , w8745 , w8746 , w8747 , w8748 , w8749 , w8750 , w8751 , w8752 , w8753 , w8754 , w8755 , w8756 , w8757 , w8758 , w8759 , w8760 , w8761 , w8762 , w8763 , w8764 , w8765 , w8766 , w8767 , w8768 , w8769 , w8770 , w8771 , w8772 , w8773 , w8774 , w8775 , w8776 , w8777 , w8778 , w8779 , w8780 , w8781 , w8782 , w8783 , w8784 , w8785 , w8786 , w8787 , w8788 , w8789 , w8790 , w8791 , w8792 , w8793 , w8794 , w8795 , w8796 , w8797 , w8798 , w8799 , w8800 , w8801 , w8802 , w8803 , w8804 , w8805 , w8806 , w8807 , w8808 , w8809 , w8810 , w8811 , w8812 , w8813 , w8814 , w8815 , w8816 , w8817 , w8818 , w8819 , w8820 , w8821 , w8822 , w8823 , w8824 , w8825 , w8826 , w8827 , w8828 , w8829 , w8830 , w8831 , w8832 , w8833 , w8834 , w8835 , w8836 , w8837 , w8838 , w8839 , w8840 , w8841 , w8842 , w8843 , w8844 , w8845 , w8846 , w8847 , w8848 , w8849 , w8850 , w8851 , w8852 , w8853 , w8854 , w8855 , w8856 , w8857 , w8858 , w8859 , w8860 , w8861 , w8862 , w8863 , w8864 , w8865 , w8866 , w8867 , w8868 , w8869 , w8870 , w8871 , w8872 , w8873 , w8874 , w8875 , w8876 , w8877 , w8878 , w8879 , w8880 , w8881 , w8882 , w8883 , w8884 , w8885 , w8886 , w8887 , w8888 , w8889 , w8890 , w8891 , w8892 , w8893 , w8894 , w8895 , w8896 , w8897 , w8898 , w8899 , w8900 , w8901 , w8902 , w8903 , w8904 , w8905 , w8906 , w8907 , w8908 , w8909 , w8910 , w8911 , w8912 , w8913 , w8914 , w8915 , w8916 , w8917 , w8918 , w8919 , w8920 , w8921 , w8922 , w8923 , w8924 , w8925 , w8926 , w8927 , w8928 , w8929 , w8930 , w8931 , w8932 , w8933 , w8934 , w8935 , w8936 , w8937 , w8938 , w8939 , w8940 , w8941 , w8942 , w8943 , w8944 , w8945 , w8946 , w8947 , w8948 , w8949 , w8950 , w8951 , w8952 , w8953 , w8954 , w8955 , w8956 , w8957 , w8958 , w8959 , w8960 , w8961 , w8962 , w8963 , w8964 , w8965 , w8966 , w8967 , w8968 , w8969 , w8970 , w8971 , w8972 , w8973 , w8974 , w8975 , w8976 , w8977 , w8978 , w8979 , w8980 , w8981 , w8982 , w8983 , w8984 , w8985 , w8986 , w8987 , w8988 , w8989 , w8990 , w8991 , w8992 , w8993 , w8994 , w8995 , w8996 , w8997 , w8998 , w8999 , w9000 , w9001 , w9002 , w9003 , w9004 , w9005 , w9006 , w9007 , w9008 , w9009 , w9010 , w9011 , w9012 , w9013 , w9014 , w9015 , w9016 , w9017 , w9018 , w9019 , w9020 , w9021 , w9022 , w9023 , w9024 , w9025 , w9026 , w9027 , w9028 , w9029 , w9030 , w9031 , w9032 , w9033 , w9034 , w9035 , w9036 , w9037 , w9038 , w9039 , w9040 , w9041 , w9042 , w9043 , w9044 , w9045 , w9046 , w9047 , w9048 , w9049 , w9050 , w9051 , w9052 , w9053 , w9054 , w9055 , w9056 , w9057 , w9058 , w9059 , w9060 , w9061 , w9062 , w9063 , w9064 , w9065 , w9066 , w9067 , w9068 , w9069 , w9070 , w9071 , w9072 , w9073 , w9074 , w9075 , w9076 , w9077 , w9078 , w9079 , w9080 , w9081 , w9082 , w9083 , w9084 , w9085 , w9086 , w9087 , w9088 , w9089 , w9090 , w9091 , w9092 , w9093 , w9094 , w9095 , w9096 , w9097 , w9098 , w9099 , w9100 , w9101 , w9102 , w9103 , w9104 , w9105 , w9106 , w9107 , w9108 , w9109 , w9110 , w9111 , w9112 , w9113 , w9114 , w9115 , w9116 , w9117 , w9118 , w9119 , w9120 , w9121 , w9122 , w9123 , w9124 , w9125 , w9126 , w9127 , w9128 , w9129 , w9130 , w9131 , w9132 , w9133 , w9134 , w9135 , w9136 , w9137 , w9138 , w9139 , w9140 , w9141 , w9142 , w9143 , w9144 , w9145 , w9146 , w9147 , w9148 , w9149 , w9150 , w9151 , w9152 , w9153 , w9154 , w9155 , w9156 , w9157 , w9158 , w9159 , w9160 , w9161 , w9162 , w9163 , w9164 , w9165 , w9166 , w9167 , w9168 , w9169 , w9170 , w9171 , w9172 , w9173 , w9174 , w9175 , w9176 , w9177 , w9178 , w9179 , w9180 , w9181 , w9182 , w9183 , w9184 , w9185 , w9186 , w9187 , w9188 , w9189 , w9190 , w9191 , w9192 , w9193 , w9194 , w9195 , w9196 , w9197 , w9198 , w9199 , w9200 , w9201 , w9202 , w9203 , w9204 , w9205 , w9206 , w9207 , w9208 , w9209 , w9210 , w9211 , w9212 , w9213 , w9214 , w9215 , w9216 , w9217 , w9218 , w9219 , w9220 , w9221 , w9222 , w9223 , w9224 , w9225 , w9226 , w9227 , w9228 , w9229 , w9230 , w9231 , w9232 , w9233 , w9234 , w9235 , w9236 , w9237 , w9238 , w9239 , w9240 , w9241 , w9242 , w9243 , w9244 , w9245 , w9246 , w9247 , w9248 , w9249 , w9250 , w9251 , w9252 , w9253 , w9254 , w9255 , w9256 , w9257 , w9258 , w9259 , w9260 , w9261 , w9262 , w9263 , w9264 , w9265 , w9266 , w9267 , w9268 , w9269 , w9270 , w9271 , w9272 , w9273 , w9274 , w9275 , w9276 , w9277 , w9278 , w9279 , w9280 , w9281 , w9282 , w9283 , w9284 , w9285 , w9286 , w9287 , w9288 , w9289 , w9290 , w9291 , w9292 , w9293 , w9294 , w9295 , w9296 , w9297 , w9298 , w9299 , w9300 , w9301 , w9302 , w9303 , w9304 , w9305 , w9306 , w9307 , w9308 , w9309 , w9310 , w9311 , w9312 , w9313 , w9314 , w9315 , w9316 , w9317 , w9318 , w9319 , w9320 , w9321 , w9322 , w9323 , w9324 , w9325 , w9326 , w9327 , w9328 , w9329 , w9330 , w9331 , w9332 , w9333 , w9334 , w9335 , w9336 , w9337 , w9338 , w9339 , w9340 , w9341 , w9342 , w9343 , w9344 , w9345 , w9346 , w9347 , w9348 , w9349 , w9350 , w9351 , w9352 , w9353 , w9354 , w9355 , w9356 , w9357 , w9358 , w9359 , w9360 , w9361 , w9362 , w9363 , w9364 , w9365 , w9366 , w9367 , w9368 , w9369 , w9370 , w9371 , w9372 , w9373 , w9374 , w9375 , w9376 , w9377 , w9378 , w9379 , w9380 , w9381 , w9382 , w9383 , w9384 , w9385 , w9386 , w9387 , w9388 , w9389 , w9390 , w9391 , w9392 , w9393 , w9394 , w9395 , w9396 , w9397 , w9398 , w9399 , w9400 , w9401 , w9402 , w9403 , w9404 , w9405 , w9406 , w9407 , w9408 , w9409 , w9410 , w9411 , w9412 , w9413 , w9414 , w9415 , w9416 , w9417 , w9418 , w9419 , w9420 , w9421 , w9422 , w9423 , w9424 , w9425 , w9426 , w9427 , w9428 , w9429 , w9430 , w9431 , w9432 , w9433 , w9434 , w9435 , w9436 , w9437 , w9438 , w9439 , w9440 , w9441 , w9442 , w9443 , w9444 , w9445 , w9446 , w9447 , w9448 , w9449 , w9450 , w9451 , w9452 , w9453 , w9454 , w9455 , w9456 , w9457 , w9458 , w9459 , w9460 , w9461 , w9462 , w9463 , w9464 , w9465 , w9466 , w9467 , w9468 , w9469 , w9470 , w9471 , w9472 , w9473 , w9474 , w9475 , w9476 , w9477 , w9478 , w9479 , w9480 , w9481 , w9482 , w9483 , w9484 , w9485 , w9486 , w9487 , w9488 , w9489 , w9490 , w9491 , w9492 , w9493 , w9494 , w9495 , w9496 , w9497 , w9498 , w9499 , w9500 , w9501 , w9502 , w9503 , w9504 , w9505 , w9506 , w9507 , w9508 , w9509 , w9510 , w9511 , w9512 , w9513 , w9514 , w9515 , w9516 , w9517 , w9518 , w9519 , w9520 , w9521 , w9522 , w9523 , w9524 , w9525 , w9526 , w9527 , w9528 , w9529 , w9530 , w9531 , w9532 , w9533 , w9534 , w9535 , w9536 , w9537 , w9538 , w9539 , w9540 , w9541 , w9542 , w9543 , w9544 , w9545 , w9546 , w9547 , w9548 , w9549 , w9550 , w9551 , w9552 , w9553 , w9554 , w9555 , w9556 , w9557 , w9558 , w9559 , w9560 , w9561 , w9562 , w9563 , w9564 , w9565 , w9566 , w9567 , w9568 , w9569 , w9570 , w9571 , w9572 , w9573 , w9574 , w9575 , w9576 , w9577 , w9578 , w9579 , w9580 , w9581 , w9582 , w9583 , w9584 , w9585 , w9586 , w9587 , w9588 , w9589 , w9590 , w9591 , w9592 , w9593 , w9594 , w9595 , w9596 , w9597 , w9598 , w9599 , w9600 , w9601 , w9602 , w9603 , w9604 , w9605 , w9606 , w9607 , w9608 , w9609 , w9610 , w9611 , w9612 , w9613 , w9614 , w9615 , w9616 , w9617 , w9618 , w9619 , w9620 , w9621 , w9622 , w9623 , w9624 , w9625 , w9626 , w9627 , w9628 , w9629 , w9630 , w9631 , w9632 , w9633 , w9634 , w9635 , w9636 , w9637 , w9638 , w9639 , w9640 , w9641 , w9642 , w9643 , w9644 , w9645 , w9646 , w9647 , w9648 , w9649 , w9650 , w9651 , w9652 , w9653 , w9654 , w9655 , w9656 , w9657 , w9658 , w9659 , w9660 , w9661 , w9662 , w9663 , w9664 , w9665 , w9666 , w9667 , w9668 , w9669 , w9670 , w9671 , w9672 , w9673 , w9674 , w9675 , w9676 , w9677 , w9678 , w9679 , w9680 , w9681 , w9682 , w9683 , w9684 , w9685 , w9686 , w9687 , w9688 , w9689 , w9690 , w9691 , w9692 , w9693 , w9694 , w9695 , w9696 , w9697 , w9698 , w9699 , w9700 , w9701 , w9702 , w9703 , w9704 , w9705 , w9706 , w9707 , w9708 , w9709 , w9710 , w9711 , w9712 , w9713 , w9714 , w9715 , w9716 , w9717 , w9718 , w9719 , w9720 , w9721 , w9722 , w9723 , w9724 , w9725 , w9726 , w9727 , w9728 , w9729 , w9730 , w9731 , w9732 , w9733 , w9734 , w9735 , w9736 , w9737 , w9738 , w9739 , w9740 , w9741 , w9742 , w9743 , w9744 , w9745 , w9746 , w9747 , w9748 , w9749 , w9750 , w9751 , w9752 , w9753 , w9754 , w9755 , w9756 , w9757 , w9758 , w9759 , w9760 , w9761 , w9762 , w9763 , w9764 , w9765 , w9766 , w9767 , w9768 , w9769 , w9770 , w9771 , w9772 , w9773 , w9774 , w9775 , w9776 , w9777 , w9778 , w9779 , w9780 , w9781 , w9782 , w9783 , w9784 , w9785 , w9786 , w9787 , w9788 , w9789 , w9790 , w9791 , w9792 , w9793 , w9794 , w9795 , w9796 , w9797 , w9798 , w9799 , w9800 , w9801 , w9802 , w9803 , w9804 , w9805 , w9806 , w9807 , w9808 , w9809 , w9810 , w9811 , w9812 , w9813 , w9814 , w9815 , w9816 , w9817 , w9818 , w9819 , w9820 , w9821 , w9822 , w9823 , w9824 , w9825 , w9826 , w9827 , w9828 , w9829 , w9830 , w9831 , w9832 , w9833 , w9834 , w9835 , w9836 , w9837 , w9838 , w9839 , w9840 , w9841 , w9842 , w9843 , w9844 , w9845 , w9846 , w9847 , w9848 , w9849 , w9850 , w9851 , w9852 , w9853 , w9854 , w9855 , w9856 , w9857 , w9858 , w9859 , w9860 , w9861 , w9862 , w9863 , w9864 , w9865 , w9866 , w9867 , w9868 , w9869 , w9870 , w9871 , w9872 , w9873 , w9874 , w9875 , w9876 , w9877 , w9878 , w9879 , w9880 , w9881 , w9882 , w9883 , w9884 , w9885 , w9886 , w9887 , w9888 , w9889 , w9890 , w9891 , w9892 , w9893 , w9894 , w9895 , w9896 , w9897 , w9898 , w9899 , w9900 , w9901 , w9902 , w9903 , w9904 , w9905 , w9906 , w9907 , w9908 , w9909 , w9910 , w9911 , w9912 , w9913 , w9914 , w9915 , w9916 , w9917 , w9918 , w9919 , w9920 , w9921 , w9922 , w9923 , w9924 , w9925 , w9926 , w9927 , w9928 , w9929 , w9930 , w9931 , w9932 , w9933 , w9934 , w9935 , w9936 , w9937 , w9938 , w9939 , w9940 , w9941 , w9942 , w9943 , w9944 , w9945 , w9946 , w9947 , w9948 , w9949 , w9950 , w9951 , w9952 , w9953 , w9954 , w9955 , w9956 , w9957 , w9958 , w9959 , w9960 , w9961 , w9962 , w9963 , w9964 , w9965 , w9966 , w9967 , w9968 , w9969 , w9970 , w9971 , w9972 , w9973 , w9974 , w9975 , w9976 , w9977 , w9978 , w9979 , w9980 , w9981 , w9982 , w9983 , w9984 , w9985 , w9986 , w9987 , w9988 , w9989 , w9990 , w9991 , w9992 , w9993 , w9994 , w9995 , w9996 , w9997 , w9998 , w9999 , w10000 , w10001 , w10002 , w10003 , w10004 , w10005 , w10006 , w10007 , w10008 , w10009 , w10010 , w10011 , w10012 , w10013 , w10014 , w10015 , w10016 , w10017 , w10018 , w10019 , w10020 , w10021 , w10022 , w10023 , w10024 , w10025 , w10026 , w10027 , w10028 , w10029 , w10030 , w10031 , w10032 , w10033 , w10034 , w10035 , w10036 , w10037 , w10038 , w10039 , w10040 , w10041 , w10042 , w10043 , w10044 , w10045 , w10046 , w10047 , w10048 , w10049 , w10050 , w10051 , w10052 , w10053 , w10054 , w10055 , w10056 , w10057 , w10058 , w10059 , w10060 , w10061 , w10062 , w10063 , w10064 , w10065 , w10066 , w10067 , w10068 , w10069 , w10070 , w10071 , w10072 , w10073 , w10074 , w10075 , w10076 , w10077 , w10078 , w10079 , w10080 , w10081 , w10082 , w10083 , w10084 , w10085 , w10086 , w10087 , w10088 , w10089 , w10090 , w10091 , w10092 , w10093 , w10094 , w10095 , w10096 , w10097 , w10098 , w10099 , w10100 , w10101 , w10102 , w10103 , w10104 , w10105 , w10106 , w10107 , w10108 , w10109 , w10110 , w10111 , w10112 , w10113 , w10114 , w10115 , w10116 , w10117 , w10118 , w10119 , w10120 , w10121 , w10122 , w10123 , w10124 , w10125 , w10126 , w10127 , w10128 , w10129 , w10130 , w10131 , w10132 , w10133 , w10134 , w10135 , w10136 , w10137 , w10138 , w10139 , w10140 , w10141 , w10142 , w10143 , w10144 , w10145 , w10146 , w10147 , w10148 , w10149 , w10150 , w10151 , w10152 , w10153 , w10154 , w10155 , w10156 , w10157 , w10158 , w10159 , w10160 , w10161 , w10162 , w10163 , w10164 , w10165 , w10166 , w10167 , w10168 , w10169 , w10170 , w10171 , w10172 , w10173 , w10174 , w10175 , w10176 , w10177 , w10178 , w10179 , w10180 , w10181 , w10182 , w10183 , w10184 , w10185 , w10186 , w10187 , w10188 , w10189 , w10190 , w10191 , w10192 , w10193 , w10194 , w10195 , w10196 , w10197 , w10198 , w10199 , w10200 , w10201 , w10202 , w10203 , w10204 , w10205 , w10206 , w10207 , w10208 , w10209 , w10210 , w10211 , w10212 , w10213 , w10214 , w10215 , w10216 , w10217 , w10218 , w10219 , w10220 , w10221 , w10222 , w10223 , w10224 , w10225 , w10226 , w10227 , w10228 , w10229 , w10230 , w10231 , w10232 , w10233 , w10234 , w10235 , w10236 , w10237 , w10238 , w10239 , w10240 , w10241 , w10242 , w10243 , w10244 , w10245 , w10246 , w10247 , w10248 , w10249 , w10250 , w10251 , w10252 , w10253 , w10254 , w10255 , w10256 , w10257 , w10258 , w10259 , w10260 , w10261 , w10262 , w10263 , w10264 , w10265 , w10266 , w10267 , w10268 , w10269 , w10270 , w10271 , w10272 , w10273 , w10274 , w10275 , w10276 , w10277 , w10278 , w10279 , w10280 , w10281 , w10282 , w10283 , w10284 , w10285 , w10286 , w10287 , w10288 , w10289 , w10290 , w10291 , w10292 , w10293 , w10294 , w10295 , w10296 , w10297 , w10298 , w10299 , w10300 , w10301 , w10302 , w10303 , w10304 , w10305 , w10306 , w10307 , w10308 , w10309 , w10310 , w10311 , w10312 , w10313 , w10314 , w10315 , w10316 , w10317 , w10318 , w10319 , w10320 , w10321 , w10322 , w10323 , w10324 , w10325 , w10326 , w10327 , w10328 , w10329 , w10330 , w10331 , w10332 , w10333 , w10334 , w10335 , w10336 , w10337 , w10338 , w10339 , w10340 , w10341 , w10342 , w10343 , w10344 , w10345 , w10346 , w10347 , w10348 , w10349 , w10350 , w10351 , w10352 , w10353 , w10354 , w10355 , w10356 , w10357 , w10358 , w10359 , w10360 , w10361 , w10362 , w10363 , w10364 , w10365 , w10366 , w10367 , w10368 , w10369 , w10370 , w10371 , w10372 , w10373 , w10374 , w10375 , w10376 , w10377 , w10378 , w10379 , w10380 , w10381 , w10382 , w10383 , w10384 , w10385 , w10386 , w10387 , w10388 , w10389 , w10390 , w10391 , w10392 , w10393 , w10394 , w10395 , w10396 , w10397 , w10398 , w10399 , w10400 , w10401 , w10402 , w10403 , w10404 , w10405 , w10406 , w10407 , w10408 , w10409 , w10410 , w10411 , w10412 , w10413 , w10414 , w10415 , w10416 , w10417 , w10418 , w10419 , w10420 , w10421 , w10422 , w10423 , w10424 , w10425 , w10426 , w10427 , w10428 , w10429 , w10430 , w10431 , w10432 , w10433 , w10434 , w10435 , w10436 , w10437 , w10438 , w10439 , w10440 , w10441 , w10442 , w10443 , w10444 , w10445 , w10446 , w10447 , w10448 , w10449 , w10450 , w10451 , w10452 , w10453 , w10454 , w10455 , w10456 , w10457 , w10458 , w10459 , w10460 , w10461 , w10462 , w10463 , w10464 , w10465 , w10466 , w10467 , w10468 , w10469 , w10470 , w10471 , w10472 , w10473 , w10474 , w10475 , w10476 , w10477 , w10478 , w10479 , w10480 , w10481 , w10482 , w10483 , w10484 , w10485 , w10486 , w10487 , w10488 , w10489 , w10490 , w10491 , w10492 , w10493 , w10494 , w10495 , w10496 , w10497 , w10498 , w10499 , w10500 , w10501 , w10502 , w10503 , w10504 , w10505 , w10506 , w10507 , w10508 , w10509 , w10510 , w10511 , w10512 , w10513 , w10514 , w10515 , w10516 , w10517 , w10518 , w10519 , w10520 , w10521 , w10522 , w10523 , w10524 , w10525 , w10526 , w10527 , w10528 , w10529 , w10530 , w10531 , w10532 , w10533 , w10534 , w10535 , w10536 , w10537 , w10538 , w10539 , w10540 , w10541 , w10542 , w10543 , w10544 , w10545 , w10546 , w10547 , w10548 , w10549 , w10550 , w10551 , w10552 , w10553 , w10554 , w10555 , w10556 , w10557 , w10558 , w10559 , w10560 , w10561 , w10562 , w10563 , w10564 , w10565 , w10566 , w10567 , w10568 , w10569 , w10570 , w10571 , w10572 , w10573 , w10574 , w10575 , w10576 , w10577 , w10578 , w10579 , w10580 , w10581 , w10582 , w10583 , w10584 , w10585 , w10586 , w10587 , w10588 , w10589 , w10590 , w10591 , w10592 , w10593 , w10594 , w10595 , w10596 , w10597 , w10598 , w10599 , w10600 , w10601 , w10602 , w10603 , w10604 , w10605 , w10606 , w10607 , w10608 , w10609 , w10610 , w10611 , w10612 , w10613 , w10614 , w10615 , w10616 , w10617 , w10618 , w10619 , w10620 , w10621 , w10622 , w10623 , w10624 , w10625 , w10626 , w10627 , w10628 , w10629 , w10630 , w10631 , w10632 , w10633 , w10634 , w10635 , w10636 , w10637 , w10638 , w10639 , w10640 , w10641 , w10642 , w10643 , w10644 , w10645 , w10646 , w10647 , w10648 , w10649 , w10650 , w10651 , w10652 , w10653 , w10654 , w10655 , w10656 , w10657 , w10658 , w10659 , w10660 , w10661 , w10662 , w10663 , w10664 , w10665 , w10666 , w10667 , w10668 , w10669 , w10670 , w10671 , w10672 , w10673 , w10674 , w10675 , w10676 , w10677 , w10678 , w10679 , w10680 , w10681 , w10682 , w10683 , w10684 , w10685 , w10686 , w10687 , w10688 , w10689 , w10690 , w10691 , w10692 , w10693 , w10694 , w10695 , w10696 , w10697 , w10698 , w10699 , w10700 , w10701 , w10702 , w10703 , w10704 , w10705 , w10706 , w10707 , w10708 , w10709 , w10710 , w10711 , w10712 , w10713 , w10714 , w10715 , w10716 , w10717 , w10718 , w10719 , w10720 , w10721 , w10722 , w10723 , w10724 , w10725 , w10726 , w10727 , w10728 , w10729 , w10730 , w10731 , w10732 , w10733 , w10734 , w10735 , w10736 , w10737 , w10738 , w10739 , w10740 , w10741 , w10742 , w10743 , w10744 , w10745 , w10746 , w10747 , w10748 , w10749 , w10750 , w10751 , w10752 , w10753 , w10754 , w10755 , w10756 , w10757 , w10758 , w10759 , w10760 , w10761 , w10762 , w10763 , w10764 , w10765 , w10766 , w10767 , w10768 , w10769 , w10770 , w10771 , w10772 , w10773 , w10774 , w10775 , w10776 , w10777 , w10778 , w10779 , w10780 , w10781 , w10782 , w10783 , w10784 , w10785 , w10786 , w10787 , w10788 , w10789 , w10790 , w10791 , w10792 , w10793 , w10794 , w10795 , w10796 , w10797 , w10798 , w10799 , w10800 , w10801 , w10802 , w10803 , w10804 , w10805 , w10806 , w10807 , w10808 , w10809 , w10810 , w10811 , w10812 , w10813 , w10814 , w10815 , w10816 , w10817 , w10818 , w10819 , w10820 , w10821 , w10822 , w10823 , w10824 , w10825 , w10826 , w10827 , w10828 , w10829 , w10830 , w10831 , w10832 , w10833 , w10834 , w10835 , w10836 , w10837 , w10838 , w10839 , w10840 , w10841 , w10842 , w10843 , w10844 , w10845 , w10846 , w10847 , w10848 , w10849 , w10850 , w10851 , w10852 , w10853 , w10854 , w10855 , w10856 , w10857 , w10858 , w10859 , w10860 , w10861 , w10862 , w10863 , w10864 , w10865 , w10866 , w10867 , w10868 , w10869 , w10870 , w10871 , w10872 , w10873 , w10874 , w10875 , w10876 , w10877 , w10878 , w10879 , w10880 , w10881 , w10882 , w10883 , w10884 , w10885 , w10886 , w10887 , w10888 , w10889 , w10890 , w10891 , w10892 , w10893 , w10894 , w10895 , w10896 , w10897 , w10898 , w10899 , w10900 , w10901 , w10902 , w10903 , w10904 , w10905 , w10906 , w10907 , w10908 , w10909 , w10910 , w10911 , w10912 , w10913 , w10914 , w10915 , w10916 , w10917 , w10918 , w10919 , w10920 , w10921 , w10922 , w10923 , w10924 , w10925 , w10926 , w10927 , w10928 , w10929 , w10930 , w10931 , w10932 , w10933 , w10934 , w10935 , w10936 , w10937 , w10938 , w10939 , w10940 , w10941 , w10942 , w10943 , w10944 , w10945 , w10946 , w10947 , w10948 , w10949 , w10950 , w10951 , w10952 , w10953 , w10954 , w10955 , w10956 , w10957 , w10958 , w10959 , w10960 , w10961 , w10962 , w10963 , w10964 , w10965 , w10966 , w10967 , w10968 , w10969 , w10970 , w10971 , w10972 , w10973 , w10974 , w10975 , w10976 , w10977 , w10978 , w10979 , w10980 , w10981 , w10982 , w10983 , w10984 , w10985 , w10986 , w10987 , w10988 , w10989 , w10990 , w10991 , w10992 , w10993 , w10994 , w10995 , w10996 , w10997 , w10998 , w10999 , w11000 , w11001 , w11002 , w11003 , w11004 , w11005 , w11006 , w11007 , w11008 , w11009 , w11010 , w11011 , w11012 , w11013 , w11014 , w11015 , w11016 , w11017 , w11018 , w11019 , w11020 , w11021 , w11022 , w11023 , w11024 , w11025 , w11026 , w11027 , w11028 , w11029 , w11030 , w11031 , w11032 , w11033 , w11034 , w11035 , w11036 , w11037 , w11038 , w11039 , w11040 , w11041 , w11042 , w11043 , w11044 , w11045 , w11046 , w11047 , w11048 , w11049 , w11050 , w11051 , w11052 , w11053 , w11054 , w11055 , w11056 , w11057 , w11058 , w11059 , w11060 , w11061 , w11062 , w11063 , w11064 , w11065 , w11066 , w11067 , w11068 , w11069 , w11070 , w11071 , w11072 , w11073 , w11074 , w11075 , w11076 , w11077 , w11078 , w11079 , w11080 , w11081 , w11082 , w11083 , w11084 , w11085 , w11086 , w11087 , w11088 , w11089 , w11090 , w11091 , w11092 , w11093 , w11094 , w11095 , w11096 , w11097 , w11098 , w11099 , w11100 , w11101 , w11102 , w11103 , w11104 , w11105 , w11106 , w11107 , w11108 , w11109 , w11110 , w11111 , w11112 , w11113 , w11114 , w11115 , w11116 , w11117 , w11118 , w11119 , w11120 , w11121 , w11122 , w11123 , w11124 , w11125 , w11126 , w11127 , w11128 , w11129 , w11130 , w11131 , w11132 , w11133 , w11134 , w11135 , w11136 , w11137 , w11138 , w11139 , w11140 , w11141 , w11142 , w11143 , w11144 , w11145 , w11146 , w11147 , w11148 , w11149 , w11150 , w11151 , w11152 , w11153 , w11154 , w11155 , w11156 , w11157 , w11158 , w11159 , w11160 , w11161 , w11162 , w11163 , w11164 , w11165 , w11166 , w11167 , w11168 , w11169 , w11170 , w11171 , w11172 , w11173 , w11174 , w11175 , w11176 , w11177 , w11178 , w11179 , w11180 , w11181 , w11182 , w11183 , w11184 , w11185 , w11186 , w11187 , w11188 , w11189 , w11190 , w11191 , w11192 , w11193 , w11194 , w11195 , w11196 , w11197 , w11198 , w11199 , w11200 , w11201 , w11202 , w11203 , w11204 , w11205 , w11206 , w11207 , w11208 , w11209 , w11210 , w11211 , w11212 , w11213 , w11214 , w11215 , w11216 , w11217 , w11218 , w11219 , w11220 , w11221 , w11222 , w11223 , w11224 , w11225 , w11226 , w11227 , w11228 , w11229 , w11230 , w11231 , w11232 , w11233 , w11234 , w11235 , w11236 , w11237 , w11238 , w11239 , w11240 , w11241 , w11242 , w11243 , w11244 , w11245 , w11246 , w11247 , w11248 , w11249 , w11250 , w11251 , w11252 , w11253 , w11254 , w11255 , w11256 , w11257 , w11258 , w11259 , w11260 , w11261 , w11262 , w11263 , w11264 , w11265 , w11266 , w11267 , w11268 , w11269 , w11270 , w11271 , w11272 , w11273 , w11274 , w11275 , w11276 , w11277 , w11278 , w11279 , w11280 , w11281 , w11282 , w11283 , w11284 , w11285 , w11286 , w11287 , w11288 , w11289 , w11290 , w11291 , w11292 , w11293 , w11294 , w11295 , w11296 , w11297 , w11298 , w11299 , w11300 , w11301 , w11302 , w11303 , w11304 , w11305 , w11306 , w11307 , w11308 , w11309 , w11310 , w11311 , w11312 , w11313 , w11314 , w11315 , w11316 , w11317 , w11318 , w11319 , w11320 , w11321 , w11322 , w11323 , w11324 , w11325 , w11326 , w11327 , w11328 , w11329 , w11330 , w11331 , w11332 , w11333 , w11334 , w11335 , w11336 , w11337 , w11338 , w11339 , w11340 , w11341 , w11342 , w11343 , w11344 , w11345 , w11346 , w11347 , w11348 , w11349 , w11350 , w11351 , w11352 , w11353 , w11354 , w11355 , w11356 , w11357 , w11358 , w11359 , w11360 , w11361 , w11362 , w11363 , w11364 , w11365 , w11366 , w11367 , w11368 , w11369 , w11370 , w11371 , w11372 , w11373 , w11374 , w11375 , w11376 , w11377 , w11378 , w11379 , w11380 , w11381 , w11382 , w11383 , w11384 , w11385 , w11386 , w11387 , w11388 , w11389 , w11390 , w11391 , w11392 , w11393 , w11394 , w11395 , w11396 , w11397 , w11398 , w11399 , w11400 , w11401 , w11402 , w11403 , w11404 , w11405 , w11406 , w11407 , w11408 , w11409 , w11410 , w11411 , w11412 , w11413 , w11414 , w11415 , w11416 , w11417 , w11418 , w11419 , w11420 , w11421 , w11422 , w11423 , w11424 , w11425 , w11426 , w11427 , w11428 , w11429 , w11430 , w11431 , w11432 , w11433 , w11434 , w11435 , w11436 , w11437 , w11438 , w11439 , w11440 , w11441 , w11442 , w11443 , w11444 , w11445 , w11446 , w11447 , w11448 , w11449 , w11450 , w11451 , w11452 , w11453 , w11454 , w11455 , w11456 , w11457 , w11458 , w11459 , w11460 , w11461 , w11462 , w11463 , w11464 , w11465 , w11466 , w11467 , w11468 , w11469 , w11470 , w11471 , w11472 , w11473 , w11474 , w11475 , w11476 , w11477 , w11478 , w11479 , w11480 , w11481 , w11482 , w11483 , w11484 , w11485 , w11486 , w11487 , w11488 , w11489 , w11490 , w11491 , w11492 , w11493 , w11494 , w11495 , w11496 , w11497 , w11498 , w11499 , w11500 , w11501 , w11502 , w11503 , w11504 , w11505 , w11506 , w11507 , w11508 , w11509 , w11510 , w11511 , w11512 , w11513 , w11514 , w11515 , w11516 , w11517 , w11518 , w11519 , w11520 , w11521 , w11522 , w11523 , w11524 , w11525 , w11526 , w11527 , w11528 , w11529 , w11530 , w11531 , w11532 , w11533 , w11534 , w11535 , w11536 , w11537 , w11538 , w11539 , w11540 , w11541 , w11542 , w11543 , w11544 , w11545 , w11546 , w11547 , w11548 , w11549 , w11550 , w11551 , w11552 , w11553 , w11554 , w11555 , w11556 , w11557 , w11558 , w11559 , w11560 , w11561 , w11562 , w11563 , w11564 , w11565 , w11566 , w11567 , w11568 , w11569 , w11570 , w11571 , w11572 , w11573 , w11574 , w11575 , w11576 , w11577 , w11578 , w11579 , w11580 , w11581 , w11582 , w11583 , w11584 , w11585 , w11586 , w11587 , w11588 , w11589 , w11590 , w11591 , w11592 , w11593 , w11594 , w11595 , w11596 , w11597 , w11598 , w11599 , w11600 , w11601 , w11602 , w11603 , w11604 , w11605 , w11606 , w11607 , w11608 , w11609 , w11610 , w11611 , w11612 , w11613 , w11614 , w11615 , w11616 , w11617 , w11618 , w11619 , w11620 , w11621 , w11622 , w11623 , w11624 , w11625 , w11626 , w11627 , w11628 , w11629 , w11630 , w11631 , w11632 , w11633 , w11634 , w11635 , w11636 , w11637 , w11638 , w11639 , w11640 , w11641 , w11642 , w11643 , w11644 , w11645 , w11646 , w11647 , w11648 , w11649 , w11650 , w11651 , w11652 , w11653 , w11654 , w11655 , w11656 , w11657 , w11658 , w11659 , w11660 , w11661 , w11662 , w11663 , w11664 , w11665 , w11666 , w11667 , w11668 , w11669 , w11670 , w11671 , w11672 , w11673 , w11674 , w11675 , w11676 , w11677 , w11678 , w11679 , w11680 , w11681 , w11682 , w11683 , w11684 , w11685 , w11686 , w11687 , w11688 , w11689 , w11690 , w11691 , w11692 , w11693 , w11694 , w11695 , w11696 , w11697 , w11698 , w11699 , w11700 , w11701 , w11702 , w11703 , w11704 , w11705 , w11706 , w11707 , w11708 , w11709 , w11710 , w11711 , w11712 , w11713 , w11714 , w11715 , w11716 , w11717 , w11718 , w11719 , w11720 , w11721 , w11722 , w11723 , w11724 , w11725 , w11726 , w11727 , w11728 , w11729 , w11730 , w11731 , w11732 , w11733 , w11734 , w11735 , w11736 , w11737 , w11738 , w11739 , w11740 , w11741 , w11742 , w11743 , w11744 , w11745 , w11746 , w11747 , w11748 , w11749 , w11750 , w11751 , w11752 , w11753 , w11754 , w11755 , w11756 , w11757 , w11758 , w11759 , w11760 , w11761 , w11762 , w11763 , w11764 , w11765 , w11766 , w11767 , w11768 , w11769 , w11770 , w11771 , w11772 , w11773 , w11774 , w11775 , w11776 , w11777 , w11778 , w11779 , w11780 , w11781 , w11782 , w11783 , w11784 , w11785 , w11786 , w11787 , w11788 , w11789 , w11790 , w11791 , w11792 , w11793 , w11794 , w11795 , w11796 , w11797 , w11798 , w11799 , w11800 , w11801 , w11802 , w11803 , w11804 , w11805 , w11806 , w11807 , w11808 , w11809 , w11810 , w11811 , w11812 , w11813 , w11814 , w11815 , w11816 , w11817 , w11818 , w11819 , w11820 , w11821 , w11822 , w11823 , w11824 , w11825 , w11826 , w11827 , w11828 , w11829 , w11830 , w11831 , w11832 , w11833 , w11834 , w11835 , w11836 , w11837 , w11838 , w11839 , w11840 , w11841 , w11842 , w11843 , w11844 , w11845 , w11846 , w11847 , w11848 , w11849 , w11850 , w11851 , w11852 , w11853 , w11854 , w11855 , w11856 , w11857 , w11858 , w11859 , w11860 , w11861 , w11862 , w11863 , w11864 , w11865 , w11866 , w11867 , w11868 , w11869 , w11870 , w11871 , w11872 , w11873 , w11874 , w11875 , w11876 , w11877 , w11878 , w11879 , w11880 , w11881 , w11882 , w11883 , w11884 , w11885 , w11886 , w11887 , w11888 , w11889 , w11890 , w11891 , w11892 , w11893 , w11894 , w11895 , w11896 , w11897 , w11898 , w11899 , w11900 , w11901 , w11902 , w11903 , w11904 , w11905 , w11906 , w11907 , w11908 , w11909 , w11910 , w11911 , w11912 , w11913 , w11914 , w11915 , w11916 , w11917 , w11918 , w11919 , w11920 , w11921 , w11922 , w11923 , w11924 , w11925 , w11926 , w11927 , w11928 , w11929 , w11930 , w11931 , w11932 , w11933 , w11934 , w11935 , w11936 , w11937 , w11938 , w11939 , w11940 , w11941 , w11942 , w11943 , w11944 , w11945 , w11946 , w11947 , w11948 , w11949 , w11950 , w11951 , w11952 , w11953 , w11954 , w11955 , w11956 , w11957 , w11958 , w11959 , w11960 , w11961 , w11962 , w11963 , w11964 , w11965 , w11966 , w11967 , w11968 , w11969 , w11970 , w11971 , w11972 , w11973 , w11974 , w11975 , w11976 , w11977 , w11978 , w11979 , w11980 , w11981 , w11982 , w11983 , w11984 , w11985 , w11986 , w11987 , w11988 , w11989 , w11990 , w11991 , w11992 , w11993 , w11994 , w11995 , w11996 , w11997 , w11998 , w11999 , w12000 , w12001 , w12002 , w12003 , w12004 , w12005 , w12006 , w12007 , w12008 , w12009 , w12010 , w12011 , w12012 , w12013 , w12014 , w12015 , w12016 , w12017 , w12018 , w12019 , w12020 , w12021 , w12022 , w12023 , w12024 , w12025 , w12026 , w12027 , w12028 , w12029 , w12030 , w12031 , w12032 , w12033 , w12034 , w12035 , w12036 , w12037 , w12038 , w12039 , w12040 , w12041 , w12042 , w12043 , w12044 , w12045 , w12046 , w12047 , w12048 , w12049 , w12050 , w12051 , w12052 , w12053 , w12054 , w12055 , w12056 , w12057 , w12058 , w12059 , w12060 , w12061 , w12062 , w12063 , w12064 , w12065 , w12066 , w12067 , w12068 , w12069 , w12070 , w12071 , w12072 , w12073 , w12074 , w12075 , w12076 , w12077 , w12078 , w12079 , w12080 , w12081 , w12082 , w12083 , w12084 , w12085 , w12086 , w12087 , w12088 , w12089 , w12090 , w12091 , w12092 , w12093 , w12094 , w12095 , w12096 , w12097 , w12098 , w12099 , w12100 , w12101 , w12102 , w12103 , w12104 , w12105 , w12106 , w12107 , w12108 , w12109 , w12110 , w12111 , w12112 , w12113 , w12114 , w12115 , w12116 , w12117 , w12118 , w12119 , w12120 , w12121 , w12122 , w12123 , w12124 , w12125 , w12126 , w12127 , w12128 , w12129 , w12130 , w12131 , w12132 , w12133 , w12134 , w12135 , w12136 , w12137 , w12138 , w12139 , w12140 , w12141 , w12142 , w12143 , w12144 , w12145 , w12146 , w12147 , w12148 , w12149 , w12150 , w12151 , w12152 , w12153 , w12154 , w12155 , w12156 , w12157 , w12158 , w12159 , w12160 , w12161 , w12162 , w12163 , w12164 , w12165 , w12166 , w12167 , w12168 , w12169 , w12170 , w12171 , w12172 , w12173 , w12174 , w12175 , w12176 , w12177 , w12178 , w12179 , w12180 , w12181 , w12182 , w12183 , w12184 , w12185 , w12186 , w12187 , w12188 , w12189 , w12190 , w12191 , w12192 , w12193 , w12194 , w12195 , w12196 , w12197 , w12198 , w12199 , w12200 , w12201 , w12202 , w12203 , w12204 , w12205 , w12206 , w12207 , w12208 , w12209 , w12210 , w12211 , w12212 , w12213 , w12214 , w12215 , w12216 , w12217 , w12218 , w12219 , w12220 , w12221 , w12222 , w12223 , w12224 , w12225 , w12226 , w12227 , w12228 , w12229 , w12230 , w12231 , w12232 , w12233 , w12234 , w12235 , w12236 , w12237 , w12238 , w12239 , w12240 , w12241 , w12242 , w12243 , w12244 , w12245 , w12246 , w12247 , w12248 , w12249 , w12250 , w12251 , w12252 , w12253 , w12254 , w12255 , w12256 , w12257 , w12258 , w12259 , w12260 , w12261 , w12262 , w12263 , w12264 , w12265 , w12266 , w12267 , w12268 , w12269 , w12270 , w12271 , w12272 , w12273 , w12274 , w12275 , w12276 , w12277 , w12278 , w12279 , w12280 , w12281 , w12282 , w12283 , w12284 , w12285 , w12286 , w12287 , w12288 , w12289 , w12290 , w12291 , w12292 , w12293 , w12294 , w12295 , w12296 , w12297 , w12298 , w12299 , w12300 , w12301 , w12302 , w12303 , w12304 , w12305 , w12306 , w12307 , w12308 , w12309 , w12310 , w12311 , w12312 , w12313 , w12314 , w12315 , w12316 , w12317 , w12318 , w12319 , w12320 , w12321 , w12322 , w12323 , w12324 , w12325 , w12326 , w12327 , w12328 , w12329 , w12330 , w12331 , w12332 , w12333 , w12334 , w12335 , w12336 , w12337 , w12338 , w12339 , w12340 , w12341 , w12342 , w12343 , w12344 , w12345 , w12346 , w12347 , w12348 , w12349 , w12350 , w12351 , w12352 , w12353 , w12354 , w12355 , w12356 , w12357 , w12358 , w12359 , w12360 , w12361 , w12362 , w12363 , w12364 , w12365 , w12366 , w12367 , w12368 , w12369 , w12370 , w12371 , w12372 , w12373 , w12374 , w12375 , w12376 , w12377 , w12378 , w12379 , w12380 , w12381 , w12382 , w12383 , w12384 , w12385 , w12386 , w12387 , w12388 , w12389 , w12390 , w12391 , w12392 , w12393 , w12394 , w12395 , w12396 , w12397 , w12398 , w12399 , w12400 , w12401 , w12402 , w12403 , w12404 , w12405 , w12406 , w12407 , w12408 , w12409 , w12410 , w12411 , w12412 , w12413 , w12414 , w12415 , w12416 , w12417 , w12418 , w12419 , w12420 , w12421 , w12422 , w12423 , w12424 , w12425 , w12426 , w12427 , w12428 , w12429 , w12430 , w12431 , w12432 , w12433 , w12434 , w12435 , w12436 , w12437 , w12438 , w12439 , w12440 , w12441 , w12442 , w12443 , w12444 , w12445 , w12446 , w12447 , w12448 , w12449 , w12450 , w12451 , w12452 , w12453 , w12454 , w12455 , w12456 , w12457 , w12458 , w12459 , w12460 , w12461 , w12462 , w12463 , w12464 , w12465 , w12466 , w12467 , w12468 , w12469 , w12470 , w12471 , w12472 , w12473 , w12474 , w12475 , w12476 , w12477 , w12478 , w12479 , w12480 , w12481 , w12482 , w12483 , w12484 , w12485 , w12486 , w12487 , w12488 , w12489 , w12490 , w12491 , w12492 , w12493 , w12494 , w12495 , w12496 , w12497 , w12498 , w12499 , w12500 , w12501 , w12502 , w12503 , w12504 , w12505 , w12506 , w12507 , w12508 , w12509 , w12510 , w12511 , w12512 , w12513 , w12514 , w12515 , w12516 , w12517 , w12518 , w12519 , w12520 , w12521 , w12522 , w12523 , w12524 , w12525 , w12526 , w12527 , w12528 , w12529 , w12530 , w12531 , w12532 , w12533 , w12534 , w12535 , w12536 , w12537 , w12538 , w12539 , w12540 , w12541 , w12542 , w12543 , w12544 , w12545 , w12546 , w12547 , w12548 , w12549 , w12550 , w12551 , w12552 , w12553 , w12554 , w12555 , w12556 , w12557 , w12558 , w12559 , w12560 , w12561 , w12562 , w12563 , w12564 , w12565 , w12566 , w12567 , w12568 , w12569 , w12570 , w12571 , w12572 , w12573 , w12574 , w12575 , w12576 , w12577 , w12578 , w12579 , w12580 , w12581 , w12582 , w12583 , w12584 , w12585 , w12586 , w12587 , w12588 , w12589 , w12590 , w12591 , w12592 , w12593 , w12594 , w12595 , w12596 , w12597 , w12598 , w12599 , w12600 , w12601 , w12602 , w12603 , w12604 , w12605 , w12606 , w12607 , w12608 , w12609 , w12610 , w12611 , w12612 , w12613 , w12614 , w12615 , w12616 , w12617 , w12618 , w12619 , w12620 , w12621 , w12622 , w12623 , w12624 , w12625 , w12626 , w12627 , w12628 , w12629 , w12630 , w12631 , w12632 , w12633 , w12634 , w12635 , w12636 , w12637 , w12638 , w12639 , w12640 , w12641 , w12642 , w12643 , w12644 , w12645 , w12646 , w12647 , w12648 , w12649 , w12650 , w12651 , w12652 , w12653 , w12654 , w12655 , w12656 , w12657 , w12658 , w12659 , w12660 , w12661 , w12662 , w12663 , w12664 , w12665 , w12666 , w12667 , w12668 , w12669 , w12670 , w12671 , w12672 , w12673 , w12674 , w12675 , w12676 , w12677 , w12678 , w12679 , w12680 , w12681 , w12682 , w12683 , w12684 , w12685 , w12686 , w12687 , w12688 , w12689 , w12690 , w12691 , w12692 , w12693 , w12694 , w12695 , w12696 , w12697 , w12698 , w12699 , w12700 , w12701 , w12702 , w12703 , w12704 , w12705 , w12706 , w12707 , w12708 , w12709 , w12710 , w12711 , w12712 , w12713 , w12714 , w12715 , w12716 , w12717 , w12718 , w12719 , w12720 , w12721 , w12722 , w12723 , w12724 , w12725 , w12726 , w12727 , w12728 , w12729 , w12730 , w12731 , w12732 , w12733 , w12734 , w12735 , w12736 , w12737 , w12738 , w12739 , w12740 , w12741 , w12742 , w12743 , w12744 , w12745 , w12746 , w12747 , w12748 , w12749 , w12750 , w12751 , w12752 , w12753 , w12754 , w12755 , w12756 , w12757 , w12758 , w12759 , w12760 , w12761 , w12762 , w12763 , w12764 , w12765 , w12766 , w12767 , w12768 , w12769 , w12770 , w12771 , w12772 , w12773 , w12774 , w12775 , w12776 , w12777 , w12778 , w12779 , w12780 , w12781 , w12782 , w12783 , w12784 , w12785 , w12786 , w12787 , w12788 , w12789 , w12790 , w12791 , w12792 , w12793 , w12794 , w12795 , w12796 , w12797 , w12798 , w12799 , w12800 , w12801 , w12802 , w12803 , w12804 , w12805 , w12806 , w12807 , w12808 , w12809 , w12810 , w12811 , w12812 , w12813 , w12814 , w12815 , w12816 , w12817 , w12818 , w12819 , w12820 , w12821 , w12822 , w12823 , w12824 , w12825 , w12826 , w12827 , w12828 , w12829 , w12830 , w12831 , w12832 , w12833 , w12834 , w12835 , w12836 , w12837 , w12838 , w12839 , w12840 , w12841 , w12842 , w12843 , w12844 , w12845 , w12846 , w12847 , w12848 , w12849 , w12850 , w12851 , w12852 , w12853 , w12854 , w12855 , w12856 , w12857 , w12858 , w12859 , w12860 , w12861 , w12862 , w12863 , w12864 , w12865 , w12866 , w12867 , w12868 , w12869 , w12870 , w12871 , w12872 , w12873 , w12874 , w12875 , w12876 , w12877 , w12878 , w12879 , w12880 , w12881 , w12882 , w12883 , w12884 , w12885 , w12886 , w12887 , w12888 , w12889 , w12890 , w12891 , w12892 , w12893 , w12894 , w12895 , w12896 , w12897 , w12898 , w12899 , w12900 , w12901 , w12902 , w12903 , w12904 , w12905 , w12906 , w12907 , w12908 , w12909 , w12910 , w12911 , w12912 , w12913 , w12914 , w12915 , w12916 , w12917 , w12918 , w12919 , w12920 , w12921 , w12922 , w12923 , w12924 , w12925 , w12926 , w12927 , w12928 , w12929 , w12930 , w12931 , w12932 , w12933 , w12934 , w12935 , w12936 , w12937 , w12938 , w12939 , w12940 , w12941 , w12942 , w12943 , w12944 , w12945 , w12946 , w12947 , w12948 , w12949 , w12950 , w12951 , w12952 , w12953 , w12954 , w12955 , w12956 , w12957 , w12958 , w12959 , w12960 , w12961 , w12962 , w12963 , w12964 , w12965 , w12966 , w12967 , w12968 , w12969 , w12970 , w12971 , w12972 , w12973 , w12974 , w12975 , w12976 , w12977 , w12978 , w12979 , w12980 , w12981 , w12982 , w12983 , w12984 , w12985 , w12986 , w12987 , w12988 , w12989 , w12990 , w12991 , w12992 , w12993 , w12994 , w12995 , w12996 , w12997 , w12998 , w12999 , w13000 , w13001 , w13002 , w13003 , w13004 , w13005 , w13006 , w13007 , w13008 , w13009 , w13010 , w13011 , w13012 , w13013 , w13014 , w13015 , w13016 , w13017 , w13018 , w13019 , w13020 , w13021 , w13022 , w13023 , w13024 , w13025 , w13026 , w13027 , w13028 , w13029 , w13030 , w13031 , w13032 , w13033 , w13034 , w13035 , w13036 , w13037 , w13038 , w13039 , w13040 , w13041 , w13042 , w13043 , w13044 , w13045 , w13046 , w13047 , w13048 , w13049 , w13050 , w13051 , w13052 , w13053 , w13054 , w13055 , w13056 , w13057 , w13058 , w13059 , w13060 , w13061 , w13062 , w13063 , w13064 , w13065 , w13066 , w13067 , w13068 , w13069 , w13070 , w13071 , w13072 , w13073 , w13074 , w13075 , w13076 , w13077 , w13078 , w13079 , w13080 , w13081 , w13082 , w13083 , w13084 , w13085 , w13086 , w13087 , w13088 , w13089 , w13090 , w13091 , w13092 , w13093 , w13094 , w13095 , w13096 , w13097 , w13098 , w13099 , w13100 , w13101 , w13102 , w13103 , w13104 , w13105 , w13106 , w13107 , w13108 , w13109 , w13110 , w13111 , w13112 , w13113 , w13114 , w13115 , w13116 , w13117 , w13118 , w13119 , w13120 , w13121 , w13122 , w13123 , w13124 , w13125 , w13126 , w13127 , w13128 , w13129 , w13130 , w13131 , w13132 , w13133 , w13134 , w13135 , w13136 , w13137 , w13138 , w13139 , w13140 , w13141 , w13142 , w13143 , w13144 , w13145 , w13146 , w13147 , w13148 , w13149 , w13150 , w13151 , w13152 , w13153 , w13154 , w13155 , w13156 , w13157 , w13158 , w13159 , w13160 , w13161 , w13162 , w13163 , w13164 , w13165 , w13166 , w13167 , w13168 , w13169 , w13170 , w13171 , w13172 , w13173 , w13174 , w13175 , w13176 , w13177 , w13178 , w13179 , w13180 , w13181 , w13182 , w13183 , w13184 , w13185 , w13186 , w13187 , w13188 , w13189 , w13190 , w13191 , w13192 , w13193 , w13194 , w13195 , w13196 , w13197 , w13198 , w13199 , w13200 , w13201 , w13202 , w13203 , w13204 , w13205 , w13206 , w13207 , w13208 , w13209 , w13210 , w13211 , w13212 , w13213 , w13214 , w13215 , w13216 , w13217 , w13218 , w13219 , w13220 , w13221 , w13222 , w13223 , w13224 , w13225 , w13226 , w13227 , w13228 , w13229 , w13230 , w13231 , w13232 , w13233 , w13234 , w13235 , w13236 , w13237 , w13238 , w13239 , w13240 , w13241 , w13242 , w13243 , w13244 , w13245 , w13246 , w13247 , w13248 , w13249 , w13250 , w13251 , w13252 , w13253 , w13254 , w13255 , w13256 , w13257 , w13258 , w13259 , w13260 , w13261 , w13262 , w13263 , w13264 , w13265 , w13266 , w13267 , w13268 , w13269 , w13270 , w13271 , w13272 , w13273 , w13274 , w13275 , w13276 , w13277 , w13278 , w13279 , w13280 , w13281 , w13282 , w13283 , w13284 , w13285 , w13286 , w13287 , w13288 , w13289 , w13290 , w13291 , w13292 , w13293 , w13294 , w13295 , w13296 , w13297 , w13298 , w13299 , w13300 , w13301 , w13302 , w13303 , w13304 , w13305 , w13306 , w13307 , w13308 , w13309 , w13310 , w13311 , w13312 , w13313 , w13314 , w13315 , w13316 , w13317 , w13318 , w13319 , w13320 , w13321 , w13322 , w13323 , w13324 , w13325 , w13326 , w13327 , w13328 , w13329 , w13330 , w13331 , w13332 , w13333 , w13334 , w13335 , w13336 , w13337 , w13338 , w13339 , w13340 , w13341 , w13342 , w13343 , w13344 , w13345 , w13346 , w13347 , w13348 , w13349 , w13350 , w13351 , w13352 , w13353 , w13354 , w13355 , w13356 , w13357 , w13358 , w13359 , w13360 , w13361 , w13362 , w13363 , w13364 , w13365 , w13366 , w13367 , w13368 , w13369 , w13370 , w13371 , w13372 , w13373 , w13374 , w13375 , w13376 , w13377 , w13378 , w13379 , w13380 , w13381 , w13382 , w13383 , w13384 , w13385 , w13386 , w13387 , w13388 , w13389 , w13390 , w13391 , w13392 , w13393 , w13394 , w13395 , w13396 , w13397 , w13398 , w13399 , w13400 , w13401 , w13402 , w13403 , w13404 , w13405 , w13406 , w13407 , w13408 , w13409 , w13410 , w13411 , w13412 , w13413 , w13414 , w13415 , w13416 , w13417 , w13418 , w13419 , w13420 , w13421 , w13422 , w13423 , w13424 , w13425 , w13426 , w13427 , w13428 , w13429 , w13430 , w13431 , w13432 , w13433 , w13434 , w13435 , w13436 , w13437 , w13438 , w13439 , w13440 , w13441 , w13442 , w13443 , w13444 , w13445 , w13446 , w13447 , w13448 , w13449 , w13450 , w13451 , w13452 , w13453 , w13454 , w13455 , w13456 , w13457 , w13458 , w13459 , w13460 , w13461 , w13462 , w13463 , w13464 , w13465 , w13466 , w13467 , w13468 , w13469 , w13470 , w13471 , w13472 , w13473 , w13474 , w13475 , w13476 , w13477 , w13478 , w13479 , w13480 , w13481 , w13482 , w13483 , w13484 , w13485 , w13486 , w13487 , w13488 , w13489 , w13490 , w13491 , w13492 , w13493 , w13494 , w13495 , w13496 , w13497 , w13498 , w13499 , w13500 , w13501 , w13502 , w13503 , w13504 , w13505 , w13506 , w13507 , w13508 , w13509 , w13510 , w13511 , w13512 , w13513 , w13514 , w13515 , w13516 , w13517 , w13518 , w13519 , w13520 , w13521 , w13522 , w13523 , w13524 , w13525 , w13526 , w13527 , w13528 , w13529 , w13530 , w13531 , w13532 , w13533 , w13534 , w13535 , w13536 , w13537 , w13538 , w13539 , w13540 , w13541 , w13542 , w13543 , w13544 , w13545 , w13546 , w13547 , w13548 , w13549 , w13550 , w13551 , w13552 , w13553 , w13554 , w13555 , w13556 , w13557 , w13558 , w13559 , w13560 , w13561 , w13562 , w13563 , w13564 , w13565 , w13566 , w13567 , w13568 , w13569 , w13570 , w13571 , w13572 , w13573 , w13574 , w13575 , w13576 , w13577 , w13578 , w13579 , w13580 , w13581 , w13582 , w13583 , w13584 , w13585 , w13586 , w13587 , w13588 , w13589 , w13590 , w13591 , w13592 , w13593 , w13594 , w13595 , w13596 , w13597 , w13598 , w13599 , w13600 , w13601 , w13602 , w13603 , w13604 , w13605 , w13606 , w13607 , w13608 , w13609 , w13610 , w13611 , w13612 , w13613 , w13614 , w13615 , w13616 , w13617 , w13618 , w13619 , w13620 , w13621 , w13622 , w13623 , w13624 , w13625 , w13626 , w13627 , w13628 , w13629 , w13630 , w13631 , w13632 , w13633 , w13634 , w13635 , w13636 , w13637 , w13638 , w13639 , w13640 , w13641 , w13642 , w13643 , w13644 , w13645 , w13646 , w13647 , w13648 , w13649 , w13650 , w13651 , w13652 , w13653 , w13654 , w13655 , w13656 , w13657 , w13658 , w13659 , w13660 , w13661 , w13662 , w13663 , w13664 , w13665 , w13666 , w13667 , w13668 , w13669 , w13670 , w13671 , w13672 , w13673 , w13674 , w13675 , w13676 , w13677 , w13678 , w13679 , w13680 , w13681 , w13682 , w13683 , w13684 , w13685 , w13686 , w13687 , w13688 , w13689 , w13690 , w13691 , w13692 , w13693 , w13694 , w13695 , w13696 , w13697 , w13698 , w13699 , w13700 , w13701 , w13702 , w13703 , w13704 , w13705 , w13706 , w13707 , w13708 , w13709 , w13710 , w13711 , w13712 , w13713 , w13714 , w13715 , w13716 , w13717 , w13718 , w13719 , w13720 , w13721 , w13722 , w13723 , w13724 , w13725 , w13726 , w13727 , w13728 , w13729 , w13730 , w13731 , w13732 , w13733 , w13734 , w13735 , w13736 , w13737 , w13738 , w13739 , w13740 , w13741 , w13742 , w13743 , w13744 , w13745 , w13746 , w13747 , w13748 , w13749 , w13750 , w13751 , w13752 , w13753 , w13754 , w13755 , w13756 , w13757 , w13758 , w13759 , w13760 , w13761 , w13762 , w13763 , w13764 , w13765 , w13766 , w13767 , w13768 , w13769 , w13770 , w13771 , w13772 , w13773 , w13774 , w13775 , w13776 , w13777 , w13778 , w13779 , w13780 , w13781 , w13782 , w13783 , w13784 , w13785 , w13786 , w13787 , w13788 , w13789 , w13790 , w13791 , w13792 , w13793 , w13794 , w13795 , w13796 , w13797 , w13798 , w13799 , w13800 , w13801 , w13802 , w13803 , w13804 , w13805 , w13806 , w13807 , w13808 , w13809 , w13810 , w13811 , w13812 , w13813 , w13814 , w13815 , w13816 , w13817 , w13818 , w13819 , w13820 , w13821 , w13822 , w13823 , w13824 , w13825 , w13826 , w13827 , w13828 , w13829 , w13830 , w13831 , w13832 , w13833 , w13834 , w13835 , w13836 , w13837 , w13838 , w13839 , w13840 , w13841 , w13842 , w13843 , w13844 , w13845 , w13846 , w13847 , w13848 , w13849 , w13850 , w13851 , w13852 , w13853 , w13854 , w13855 , w13856 , w13857 , w13858 , w13859 , w13860 , w13861 , w13862 , w13863 , w13864 , w13865 , w13866 , w13867 , w13868 , w13869 , w13870 , w13871 , w13872 , w13873 , w13874 , w13875 , w13876 , w13877 , w13878 , w13879 , w13880 , w13881 , w13882 , w13883 , w13884 , w13885 , w13886 , w13887 , w13888 , w13889 , w13890 , w13891 , w13892 , w13893 , w13894 , w13895 , w13896 , w13897 , w13898 , w13899 , w13900 , w13901 , w13902 , w13903 , w13904 , w13905 , w13906 , w13907 , w13908 , w13909 , w13910 , w13911 , w13912 , w13913 , w13914 , w13915 , w13916 , w13917 , w13918 , w13919 , w13920 , w13921 , w13922 , w13923 , w13924 , w13925 , w13926 , w13927 , w13928 , w13929 , w13930 , w13931 , w13932 , w13933 , w13934 , w13935 , w13936 , w13937 , w13938 , w13939 , w13940 , w13941 , w13942 , w13943 , w13944 , w13945 , w13946 , w13947 , w13948 , w13949 , w13950 , w13951 , w13952 , w13953 , w13954 , w13955 , w13956 , w13957 , w13958 , w13959 , w13960 , w13961 , w13962 , w13963 , w13964 , w13965 , w13966 , w13967 , w13968 , w13969 , w13970 , w13971 , w13972 , w13973 , w13974 , w13975 , w13976 , w13977 , w13978 , w13979 , w13980 , w13981 , w13982 , w13983 , w13984 , w13985 , w13986 , w13987 , w13988 , w13989 , w13990 , w13991 , w13992 , w13993 , w13994 , w13995 , w13996 , w13997 , w13998 , w13999 , w14000 , w14001 , w14002 , w14003 , w14004 , w14005 , w14006 , w14007 , w14008 , w14009 , w14010 , w14011 , w14012 , w14013 , w14014 , w14015 , w14016 , w14017 , w14018 , w14019 , w14020 , w14021 , w14022 , w14023 , w14024 , w14025 , w14026 , w14027 , w14028 , w14029 , w14030 , w14031 , w14032 , w14033 , w14034 , w14035 , w14036 , w14037 , w14038 , w14039 , w14040 , w14041 , w14042 , w14043 , w14044 , w14045 , w14046 , w14047 , w14048 , w14049 , w14050 , w14051 , w14052 , w14053 , w14054 , w14055 , w14056 , w14057 , w14058 , w14059 , w14060 , w14061 , w14062 , w14063 , w14064 , w14065 , w14066 , w14067 , w14068 , w14069 , w14070 , w14071 , w14072 , w14073 , w14074 , w14075 , w14076 , w14077 , w14078 , w14079 , w14080 , w14081 , w14082 , w14083 , w14084 , w14085 , w14086 , w14087 , w14088 , w14089 , w14090 , w14091 , w14092 , w14093 , w14094 , w14095 , w14096 , w14097 , w14098 , w14099 , w14100 , w14101 , w14102 , w14103 , w14104 , w14105 , w14106 , w14107 , w14108 , w14109 , w14110 , w14111 , w14112 , w14113 , w14114 , w14115 , w14116 , w14117 , w14118 , w14119 , w14120 , w14121 , w14122 , w14123 , w14124 , w14125 , w14126 , w14127 , w14128 , w14129 , w14130 , w14131 , w14132 , w14133 , w14134 , w14135 , w14136 , w14137 , w14138 , w14139 , w14140 , w14141 , w14142 , w14143 , w14144 , w14145 , w14146 , w14147 , w14148 , w14149 , w14150 , w14151 , w14152 , w14153 , w14154 , w14155 , w14156 , w14157 , w14158 , w14159 , w14160 , w14161 , w14162 , w14163 , w14164 , w14165 , w14166 , w14167 , w14168 , w14169 , w14170 , w14171 , w14172 , w14173 , w14174 , w14175 , w14176 , w14177 , w14178 , w14179 , w14180 , w14181 , w14182 , w14183 , w14184 , w14185 , w14186 , w14187 , w14188 , w14189 , w14190 , w14191 , w14192 , w14193 , w14194 , w14195 , w14196 , w14197 , w14198 , w14199 , w14200 , w14201 , w14202 , w14203 , w14204 , w14205 , w14206 , w14207 , w14208 , w14209 , w14210 , w14211 , w14212 , w14213 , w14214 , w14215 , w14216 , w14217 , w14218 , w14219 , w14220 , w14221 , w14222 , w14223 , w14224 , w14225 , w14226 , w14227 , w14228 , w14229 , w14230 , w14231 , w14232 , w14233 , w14234 , w14235 , w14236 , w14237 , w14238 , w14239 , w14240 , w14241 , w14242 , w14243 , w14244 , w14245 , w14246 , w14247 , w14248 , w14249 , w14250 , w14251 , w14252 , w14253 , w14254 , w14255 , w14256 , w14257 , w14258 , w14259 , w14260 , w14261 , w14262 , w14263 , w14264 , w14265 , w14266 , w14267 , w14268 , w14269 , w14270 , w14271 , w14272 , w14273 , w14274 , w14275 , w14276 , w14277 , w14278 , w14279 , w14280 , w14281 , w14282 , w14283 , w14284 , w14285 , w14286 , w14287 , w14288 , w14289 , w14290 , w14291 , w14292 , w14293 , w14294 , w14295 , w14296 , w14297 , w14298 , w14299 , w14300 , w14301 , w14302 , w14303 , w14304 , w14305 , w14306 , w14307 , w14308 , w14309 , w14310 , w14311 , w14312 , w14313 , w14314 , w14315 , w14316 , w14317 , w14318 , w14319 , w14320 , w14321 , w14322 , w14323 , w14324 , w14325 , w14326 , w14327 , w14328 , w14329 , w14330 , w14331 , w14332 , w14333 , w14334 , w14335 , w14336 , w14337 , w14338 , w14339 , w14340 , w14341 , w14342 , w14343 , w14344 , w14345 , w14346 , w14347 , w14348 , w14349 , w14350 , w14351 , w14352 , w14353 , w14354 , w14355 , w14356 , w14357 , w14358 , w14359 , w14360 , w14361 , w14362 , w14363 , w14364 , w14365 , w14366 , w14367 , w14368 , w14369 , w14370 , w14371 , w14372 , w14373 , w14374 , w14375 , w14376 , w14377 , w14378 , w14379 , w14380 , w14381 , w14382 , w14383 , w14384 , w14385 , w14386 , w14387 , w14388 , w14389 , w14390 , w14391 , w14392 , w14393 , w14394 , w14395 , w14396 , w14397 , w14398 , w14399 , w14400 , w14401 , w14402 , w14403 , w14404 , w14405 , w14406 , w14407 , w14408 , w14409 , w14410 , w14411 , w14412 , w14413 , w14414 , w14415 , w14416 , w14417 , w14418 , w14419 , w14420 , w14421 , w14422 , w14423 , w14424 , w14425 , w14426 , w14427 , w14428 , w14429 , w14430 , w14431 , w14432 , w14433 , w14434 , w14435 , w14436 , w14437 , w14438 , w14439 , w14440 , w14441 , w14442 , w14443 , w14444 , w14445 , w14446 , w14447 , w14448 , w14449 , w14450 , w14451 , w14452 , w14453 , w14454 , w14455 , w14456 , w14457 , w14458 , w14459 , w14460 , w14461 , w14462 , w14463 , w14464 , w14465 , w14466 , w14467 , w14468 , w14469 , w14470 , w14471 , w14472 , w14473 , w14474 , w14475 , w14476 , w14477 , w14478 , w14479 , w14480 , w14481 , w14482 , w14483 , w14484 , w14485 , w14486 , w14487 , w14488 , w14489 , w14490 , w14491 , w14492 , w14493 , w14494 , w14495 , w14496 , w14497 , w14498 , w14499 , w14500 , w14501 , w14502 , w14503 , w14504 , w14505 , w14506 , w14507 , w14508 , w14509 , w14510 , w14511 , w14512 , w14513 , w14514 , w14515 , w14516 , w14517 , w14518 , w14519 , w14520 , w14521 , w14522 , w14523 , w14524 , w14525 , w14526 , w14527 , w14528 , w14529 , w14530 , w14531 , w14532 , w14533 , w14534 , w14535 , w14536 , w14537 , w14538 , w14539 , w14540 , w14541 , w14542 , w14543 , w14544 , w14545 , w14546 , w14547 , w14548 , w14549 , w14550 , w14551 , w14552 , w14553 , w14554 , w14555 , w14556 , w14557 , w14558 , w14559 , w14560 , w14561 , w14562 , w14563 , w14564 , w14565 , w14566 , w14567 , w14568 , w14569 , w14570 , w14571 , w14572 , w14573 , w14574 , w14575 , w14576 , w14577 , w14578 , w14579 , w14580 , w14581 , w14582 , w14583 , w14584 , w14585 , w14586 , w14587 , w14588 , w14589 , w14590 , w14591 , w14592 , w14593 , w14594 , w14595 , w14596 , w14597 , w14598 , w14599 , w14600 , w14601 , w14602 , w14603 , w14604 , w14605 , w14606 , w14607 , w14608 , w14609 , w14610 , w14611 , w14612 , w14613 , w14614 , w14615 , w14616 , w14617 , w14618 , w14619 , w14620 , w14621 , w14622 , w14623 , w14624 , w14625 , w14626 , w14627 , w14628 , w14629 , w14630 , w14631 , w14632 , w14633 , w14634 , w14635 , w14636 , w14637 , w14638 , w14639 , w14640 , w14641 , w14642 , w14643 , w14644 , w14645 , w14646 , w14647 , w14648 , w14649 , w14650 , w14651 , w14652 , w14653 , w14654 , w14655 , w14656 , w14657 , w14658 , w14659 , w14660 , w14661 , w14662 , w14663 , w14664 , w14665 , w14666 , w14667 , w14668 , w14669 , w14670 , w14671 , w14672 , w14673 , w14674 , w14675 , w14676 , w14677 , w14678 , w14679 , w14680 , w14681 , w14682 , w14683 , w14684 , w14685 , w14686 , w14687 , w14688 , w14689 , w14690 , w14691 , w14692 , w14693 , w14694 , w14695 , w14696 , w14697 , w14698 , w14699 , w14700 , w14701 , w14702 , w14703 , w14704 , w14705 , w14706 , w14707 , w14708 , w14709 , w14710 , w14711 , w14712 , w14713 , w14714 , w14715 , w14716 , w14717 , w14718 , w14719 , w14720 , w14721 , w14722 , w14723 , w14724 , w14725 , w14726 , w14727 , w14728 , w14729 , w14730 , w14731 , w14732 , w14733 , w14734 , w14735 , w14736 , w14737 , w14738 , w14739 , w14740 , w14741 , w14742 , w14743 , w14744 , w14745 , w14746 , w14747 , w14748 , w14749 , w14750 , w14751 , w14752 , w14753 , w14754 , w14755 , w14756 , w14757 , w14758 , w14759 , w14760 , w14761 , w14762 , w14763 , w14764 , w14765 , w14766 , w14767 , w14768 , w14769 , w14770 , w14771 , w14772 , w14773 , w14774 , w14775 , w14776 , w14777 , w14778 , w14779 , w14780 , w14781 , w14782 , w14783 , w14784 , w14785 , w14786 , w14787 , w14788 , w14789 , w14790 , w14791 , w14792 , w14793 , w14794 , w14795 , w14796 , w14797 , w14798 , w14799 , w14800 , w14801 , w14802 , w14803 , w14804 , w14805 , w14806 , w14807 , w14808 , w14809 , w14810 , w14811 , w14812 , w14813 , w14814 , w14815 , w14816 , w14817 , w14818 , w14819 , w14820 , w14821 , w14822 , w14823 , w14824 , w14825 , w14826 , w14827 , w14828 , w14829 , w14830 , w14831 , w14832 , w14833 , w14834 , w14835 , w14836 , w14837 , w14838 , w14839 , w14840 , w14841 , w14842 , w14843 , w14844 , w14845 , w14846 , w14847 , w14848 , w14849 , w14850 , w14851 , w14852 , w14853 , w14854 , w14855 , w14856 , w14857 , w14858 , w14859 , w14860 , w14861 , w14862 , w14863 , w14864 , w14865 , w14866 , w14867 , w14868 , w14869 , w14870 , w14871 , w14872 , w14873 , w14874 , w14875 , w14876 , w14877 , w14878 , w14879 , w14880 , w14881 , w14882 , w14883 , w14884 , w14885 , w14886 , w14887 , w14888 , w14889 , w14890 , w14891 , w14892 , w14893 , w14894 , w14895 , w14896 , w14897 , w14898 , w14899 , w14900 , w14901 , w14902 , w14903 , w14904 , w14905 , w14906 , w14907 , w14908 , w14909 , w14910 , w14911 , w14912 , w14913 , w14914 , w14915 , w14916 , w14917 , w14918 , w14919 , w14920 , w14921 , w14922 , w14923 , w14924 , w14925 , w14926 , w14927 , w14928 , w14929 , w14930 , w14931 , w14932 , w14933 , w14934 , w14935 , w14936 , w14937 , w14938 , w14939 , w14940 , w14941 , w14942 , w14943 , w14944 , w14945 , w14946 , w14947 , w14948 , w14949 , w14950 , w14951 , w14952 , w14953 , w14954 , w14955 , w14956 , w14957 , w14958 , w14959 , w14960 , w14961 , w14962 , w14963 , w14964 , w14965 , w14966 , w14967 , w14968 , w14969 , w14970 , w14971 , w14972 , w14973 , w14974 , w14975 , w14976 , w14977 , w14978 , w14979 , w14980 , w14981 , w14982 , w14983 , w14984 , w14985 , w14986 , w14987 , w14988 , w14989 , w14990 , w14991 , w14992 , w14993 , w14994 , w14995 , w14996 , w14997 , w14998 , w14999 , w15000 , w15001 , w15002 , w15003 , w15004 , w15005 , w15006 , w15007 , w15008 , w15009 , w15010 , w15011 , w15012 , w15013 , w15014 , w15015 , w15016 , w15017 , w15018 , w15019 , w15020 , w15021 , w15022 , w15023 , w15024 , w15025 , w15026 , w15027 , w15028 , w15029 , w15030 , w15031 , w15032 , w15033 , w15034 , w15035 , w15036 , w15037 , w15038 , w15039 , w15040 , w15041 , w15042 , w15043 , w15044 , w15045 , w15046 , w15047 , w15048 , w15049 , w15050 , w15051 , w15052 , w15053 , w15054 , w15055 , w15056 , w15057 , w15058 , w15059 , w15060 , w15061 , w15062 , w15063 , w15064 , w15065 , w15066 , w15067 , w15068 , w15069 , w15070 , w15071 , w15072 , w15073 , w15074 , w15075 , w15076 , w15077 , w15078 , w15079 , w15080 , w15081 , w15082 , w15083 , w15084 , w15085 , w15086 , w15087 , w15088 , w15089 , w15090 , w15091 , w15092 , w15093 , w15094 , w15095 , w15096 , w15097 , w15098 , w15099 , w15100 , w15101 , w15102 , w15103 , w15104 , w15105 , w15106 , w15107 , w15108 , w15109 , w15110 , w15111 , w15112 , w15113 , w15114 , w15115 , w15116 , w15117 , w15118 , w15119 , w15120 , w15121 , w15122 , w15123 , w15124 , w15125 , w15126 , w15127 , w15128 , w15129 , w15130 , w15131 , w15132 , w15133 , w15134 , w15135 , w15136 , w15137 , w15138 , w15139 , w15140 , w15141 , w15142 , w15143 , w15144 , w15145 , w15146 , w15147 , w15148 , w15149 , w15150 , w15151 , w15152 , w15153 , w15154 , w15155 , w15156 , w15157 , w15158 , w15159 , w15160 , w15161 , w15162 , w15163 , w15164 , w15165 , w15166 , w15167 , w15168 , w15169 , w15170 , w15171 , w15172 , w15173 , w15174 , w15175 , w15176 , w15177 , w15178 , w15179 , w15180 , w15181 , w15182 , w15183 , w15184 , w15185 , w15186 , w15187 , w15188 , w15189 , w15190 , w15191 , w15192 , w15193 , w15194 , w15195 , w15196 , w15197 , w15198 , w15199 , w15200 , w15201 , w15202 , w15203 , w15204 , w15205 , w15206 , w15207 , w15208 , w15209 , w15210 , w15211 , w15212 , w15213 , w15214 , w15215 , w15216 , w15217 , w15218 , w15219 , w15220 , w15221 , w15222 , w15223 , w15224 , w15225 , w15226 , w15227 , w15228 , w15229 , w15230 , w15231 , w15232 , w15233 , w15234 , w15235 , w15236 , w15237 , w15238 , w15239 , w15240 , w15241 , w15242 , w15243 , w15244 , w15245 , w15246 , w15247 , w15248 , w15249 , w15250 , w15251 , w15252 , w15253 , w15254 , w15255 , w15256 , w15257 , w15258 , w15259 , w15260 , w15261 , w15262 , w15263 , w15264 , w15265 , w15266 , w15267 , w15268 , w15269 , w15270 , w15271 , w15272 , w15273 , w15274 , w15275 , w15276 , w15277 , w15278 , w15279 , w15280 , w15281 , w15282 , w15283 , w15284 , w15285 , w15286 , w15287 , w15288 , w15289 , w15290 , w15291 , w15292 , w15293 , w15294 , w15295 , w15296 , w15297 , w15298 , w15299 , w15300 , w15301 , w15302 , w15303 , w15304 , w15305 , w15306 , w15307 , w15308 , w15309 , w15310 , w15311 , w15312 , w15313 , w15314 , w15315 , w15316 , w15317 , w15318 , w15319 , w15320 , w15321 , w15322 , w15323 , w15324 , w15325 , w15326 , w15327 , w15328 , w15329 , w15330 , w15331 , w15332 , w15333 , w15334 , w15335 , w15336 , w15337 , w15338 , w15339 , w15340 , w15341 , w15342 , w15343 , w15344 , w15345 , w15346 , w15347 , w15348 , w15349 , w15350 , w15351 , w15352 , w15353 , w15354 , w15355 , w15356 , w15357 , w15358 , w15359 , w15360 , w15361 , w15362 , w15363 , w15364 , w15365 , w15366 , w15367 , w15368 , w15369 , w15370 , w15371 , w15372 , w15373 , w15374 , w15375 , w15376 , w15377 , w15378 , w15379 , w15380 , w15381 , w15382 , w15383 , w15384 , w15385 , w15386 , w15387 , w15388 , w15389 , w15390 , w15391 , w15392 , w15393 , w15394 , w15395 , w15396 , w15397 , w15398 , w15399 , w15400 , w15401 , w15402 , w15403 , w15404 , w15405 , w15406 , w15407 , w15408 , w15409 , w15410 , w15411 , w15412 , w15413 , w15414 , w15415 , w15416 , w15417 , w15418 , w15419 , w15420 , w15421 , w15422 , w15423 , w15424 , w15425 , w15426 , w15427 , w15428 , w15429 , w15430 , w15431 , w15432 , w15433 , w15434 , w15435 , w15436 , w15437 , w15438 , w15439 , w15440 , w15441 , w15442 , w15443 , w15444 , w15445 , w15446 , w15447 , w15448 , w15449 , w15450 , w15451 , w15452 , w15453 , w15454 , w15455 , w15456 , w15457 , w15458 , w15459 , w15460 , w15461 , w15462 , w15463 , w15464 , w15465 , w15466 , w15467 , w15468 , w15469 , w15470 , w15471 , w15472 , w15473 , w15474 , w15475 , w15476 , w15477 , w15478 , w15479 , w15480 , w15481 , w15482 , w15483 , w15484 , w15485 , w15486 , w15487 , w15488 , w15489 , w15490 , w15491 , w15492 , w15493 , w15494 , w15495 , w15496 , w15497 , w15498 , w15499 , w15500 , w15501 , w15502 , w15503 , w15504 , w15505 , w15506 , w15507 , w15508 , w15509 , w15510 , w15511 , w15512 , w15513 , w15514 , w15515 , w15516 , w15517 , w15518 , w15519 , w15520 , w15521 , w15522 , w15523 , w15524 , w15525 , w15526 , w15527 , w15528 , w15529 , w15530 , w15531 , w15532 , w15533 , w15534 , w15535 , w15536 , w15537 , w15538 , w15539 , w15540 , w15541 , w15542 , w15543 , w15544 , w15545 , w15546 , w15547 , w15548 , w15549 , w15550 , w15551 , w15552 , w15553 , w15554 , w15555 , w15556 , w15557 , w15558 , w15559 , w15560 , w15561 , w15562 , w15563 , w15564 , w15565 , w15566 , w15567 , w15568 , w15569 , w15570 , w15571 , w15572 , w15573 , w15574 , w15575 , w15576 , w15577 , w15578 , w15579 , w15580 , w15581 , w15582 , w15583 , w15584 , w15585 , w15586 , w15587 , w15588 , w15589 , w15590 , w15591 , w15592 , w15593 , w15594 , w15595 , w15596 , w15597 , w15598 , w15599 , w15600 , w15601 , w15602 , w15603 , w15604 , w15605 , w15606 , w15607 , w15608 , w15609 , w15610 , w15611 , w15612 , w15613 , w15614 , w15615 , w15616 , w15617 , w15618 , w15619 , w15620 , w15621 , w15622 , w15623 , w15624 , w15625 , w15626 , w15627 , w15628 , w15629 , w15630 , w15631 , w15632 , w15633 , w15634 , w15635 , w15636 , w15637 , w15638 , w15639 , w15640 , w15641 , w15642 , w15643 , w15644 , w15645 , w15646 , w15647 , w15648 , w15649 , w15650 , w15651 , w15652 , w15653 , w15654 , w15655 , w15656 , w15657 , w15658 , w15659 , w15660 , w15661 , w15662 , w15663 , w15664 , w15665 , w15666 , w15667 , w15668 , w15669 , w15670 , w15671 , w15672 , w15673 , w15674 , w15675 , w15676 , w15677 , w15678 , w15679 , w15680 , w15681 , w15682 , w15683 , w15684 , w15685 , w15686 , w15687 , w15688 , w15689 , w15690 , w15691 , w15692 , w15693 , w15694 , w15695 , w15696 , w15697 , w15698 , w15699 , w15700 , w15701 , w15702 , w15703 , w15704 , w15705 , w15706 , w15707 , w15708 , w15709 , w15710 , w15711 , w15712 , w15713 , w15714 , w15715 , w15716 , w15717 , w15718 , w15719 , w15720 , w15721 , w15722 , w15723 , w15724 , w15725 , w15726 , w15727 , w15728 , w15729 , w15730 , w15731 , w15732 , w15733 , w15734 , w15735 , w15736 , w15737 , w15738 , w15739 , w15740 , w15741 , w15742 , w15743 , w15744 , w15745 , w15746 , w15747 , w15748 , w15749 , w15750 , w15751 , w15752 , w15753 , w15754 , w15755 , w15756 , w15757 , w15758 , w15759 , w15760 , w15761 , w15762 , w15763 , w15764 , w15765 , w15766 , w15767 , w15768 , w15769 , w15770 , w15771 , w15772 , w15773 , w15774 , w15775 , w15776 , w15777 , w15778 , w15779 , w15780 , w15781 , w15782 , w15783 , w15784 , w15785 , w15786 , w15787 , w15788 , w15789 , w15790 , w15791 , w15792 , w15793 , w15794 , w15795 , w15796 , w15797 , w15798 , w15799 , w15800 , w15801 , w15802 , w15803 , w15804 , w15805 , w15806 , w15807 , w15808 , w15809 , w15810 , w15811 , w15812 , w15813 , w15814 , w15815 , w15816 , w15817 , w15818 , w15819 , w15820 , w15821 , w15822 , w15823 , w15824 , w15825 , w15826 , w15827 , w15828 , w15829 , w15830 , w15831 , w15832 , w15833 , w15834 , w15835 , w15836 , w15837 , w15838 , w15839 , w15840 , w15841 , w15842 , w15843 , w15844 , w15845 , w15846 , w15847 , w15848 , w15849 , w15850 , w15851 , w15852 , w15853 , w15854 , w15855 , w15856 , w15857 , w15858 , w15859 , w15860 , w15861 , w15862 , w15863 , w15864 , w15865 , w15866 , w15867 , w15868 , w15869 , w15870 , w15871 , w15872 , w15873 , w15874 , w15875 , w15876 , w15877 , w15878 , w15879 , w15880 , w15881 , w15882 , w15883 , w15884 , w15885 , w15886 , w15887 , w15888 , w15889 , w15890 , w15891 , w15892 , w15893 , w15894 , w15895 , w15896 , w15897 , w15898 , w15899 , w15900 , w15901 , w15902 , w15903 , w15904 , w15905 , w15906 , w15907 , w15908 , w15909 , w15910 , w15911 , w15912 , w15913 , w15914 , w15915 , w15916 , w15917 , w15918 , w15919 , w15920 , w15921 , w15922 , w15923 , w15924 , w15925 , w15926 , w15927 , w15928 , w15929 , w15930 , w15931 , w15932 , w15933 , w15934 , w15935 , w15936 , w15937 , w15938 , w15939 , w15940 , w15941 , w15942 , w15943 , w15944 , w15945 , w15946 , w15947 , w15948 , w15949 , w15950 , w15951 , w15952 , w15953 , w15954 , w15955 , w15956 , w15957 , w15958 , w15959 , w15960 , w15961 , w15962 , w15963 , w15964 , w15965 , w15966 , w15967 , w15968 , w15969 , w15970 , w15971 , w15972 , w15973 , w15974 , w15975 , w15976 , w15977 , w15978 , w15979 , w15980 , w15981 , w15982 , w15983 , w15984 , w15985 , w15986 , w15987 , w15988 , w15989 , w15990 , w15991 , w15992 , w15993 , w15994 , w15995 , w15996 , w15997 , w15998 , w15999 , w16000 , w16001 , w16002 , w16003 , w16004 , w16005 , w16006 , w16007 , w16008 , w16009 , w16010 , w16011 , w16012 , w16013 , w16014 , w16015 , w16016 , w16017 , w16018 , w16019 , w16020 , w16021 , w16022 , w16023 , w16024 , w16025 , w16026 , w16027 , w16028 , w16029 , w16030 , w16031 , w16032 , w16033 , w16034 , w16035 , w16036 , w16037 , w16038 , w16039 , w16040 , w16041 , w16042 , w16043 , w16044 , w16045 , w16046 , w16047 , w16048 , w16049 , w16050 , w16051 , w16052 , w16053 , w16054 , w16055 , w16056 , w16057 , w16058 , w16059 , w16060 , w16061 , w16062 , w16063 , w16064 , w16065 , w16066 , w16067 , w16068 , w16069 , w16070 , w16071 , w16072 , w16073 , w16074 , w16075 , w16076 , w16077 , w16078 , w16079 , w16080 , w16081 , w16082 , w16083 , w16084 , w16085 , w16086 , w16087 , w16088 , w16089 , w16090 , w16091 , w16092 , w16093 , w16094 , w16095 , w16096 , w16097 , w16098 , w16099 , w16100 , w16101 , w16102 , w16103 , w16104 , w16105 , w16106 , w16107 , w16108 , w16109 , w16110 , w16111 , w16112 , w16113 , w16114 , w16115 , w16116 , w16117 , w16118 , w16119 , w16120 , w16121 , w16122 , w16123 , w16124 , w16125 , w16126 , w16127 , w16128 , w16129 , w16130 , w16131 , w16132 , w16133 , w16134 , w16135 , w16136 , w16137 , w16138 , w16139 , w16140 , w16141 , w16142 , w16143 , w16144 , w16145 , w16146 , w16147 , w16148 , w16149 , w16150 , w16151 , w16152 , w16153 , w16154 , w16155 , w16156 , w16157 , w16158 , w16159 , w16160 , w16161 , w16162 , w16163 , w16164 , w16165 , w16166 , w16167 , w16168 , w16169 , w16170 , w16171 , w16172 , w16173 , w16174 , w16175 , w16176 , w16177 , w16178 , w16179 , w16180 , w16181 , w16182 , w16183 , w16184 , w16185 , w16186 , w16187 , w16188 , w16189 , w16190 , w16191 , w16192 , w16193 , w16194 , w16195 , w16196 , w16197 , w16198 , w16199 , w16200 , w16201 , w16202 , w16203 , w16204 , w16205 , w16206 , w16207 , w16208 , w16209 , w16210 , w16211 , w16212 , w16213 , w16214 , w16215 , w16216 , w16217 , w16218 , w16219 , w16220 , w16221 , w16222 , w16223 , w16224 , w16225 , w16226 , w16227 , w16228 , w16229 , w16230 , w16231 , w16232 , w16233 , w16234 , w16235 , w16236 , w16237 , w16238 , w16239 , w16240 , w16241 , w16242 , w16243 , w16244 , w16245 , w16246 , w16247 , w16248 , w16249 , w16250 , w16251 , w16252 , w16253 , w16254 , w16255 , w16256 , w16257 , w16258 , w16259 , w16260 , w16261 , w16262 , w16263 , w16264 , w16265 , w16266 , w16267 , w16268 , w16269 , w16270 , w16271 , w16272 , w16273 , w16274 , w16275 , w16276 , w16277 , w16278 , w16279 , w16280 , w16281 , w16282 , w16283 , w16284 , w16285 , w16286 , w16287 , w16288 , w16289 , w16290 , w16291 , w16292 , w16293 , w16294 , w16295 , w16296 , w16297 , w16298 , w16299 , w16300 , w16301 , w16302 , w16303 , w16304 , w16305 , w16306 , w16307 , w16308 , w16309 , w16310 , w16311 , w16312 , w16313 , w16314 , w16315 , w16316 , w16317 , w16318 , w16319 , w16320 , w16321 , w16322 , w16323 , w16324 , w16325 , w16326 , w16327 , w16328 , w16329 , w16330 , w16331 , w16332 , w16333 , w16334 , w16335 , w16336 , w16337 , w16338 , w16339 , w16340 , w16341 , w16342 , w16343 , w16344 , w16345 , w16346 , w16347 , w16348 , w16349 , w16350 , w16351 , w16352 , w16353 , w16354 , w16355 , w16356 , w16357 , w16358 , w16359 , w16360 , w16361 , w16362 , w16363 , w16364 , w16365 , w16366 , w16367 , w16368 , w16369 , w16370 , w16371 , w16372 , w16373 , w16374 , w16375 , w16376 , w16377 , w16378 , w16379 , w16380 , w16381 , w16382 , w16383 , w16384 , w16385 , w16386 , w16387 , w16388 , w16389 , w16390 , w16391 , w16392 , w16393 , w16394 , w16395 , w16396 , w16397 , w16398 , w16399 , w16400 , w16401 , w16402 , w16403 , w16404 , w16405 , w16406 , w16407 , w16408 , w16409 , w16410 , w16411 , w16412 , w16413 , w16414 , w16415 , w16416 , w16417 , w16418 , w16419 , w16420 , w16421 , w16422 , w16423 , w16424 , w16425 , w16426 , w16427 , w16428 , w16429 , w16430 , w16431 , w16432 , w16433 , w16434 , w16435 , w16436 , w16437 , w16438 , w16439 , w16440 , w16441 , w16442 , w16443 , w16444 , w16445 , w16446 , w16447 , w16448 , w16449 , w16450 , w16451 , w16452 , w16453 , w16454 , w16455 , w16456 , w16457 , w16458 , w16459 , w16460 , w16461 , w16462 , w16463 , w16464 , w16465 , w16466 , w16467 , w16468 , w16469 , w16470 , w16471 , w16472 , w16473 , w16474 , w16475 , w16476 , w16477 , w16478 , w16479 , w16480 , w16481 , w16482 , w16483 , w16484 , w16485 , w16486 , w16487 , w16488 , w16489 , w16490 , w16491 , w16492 , w16493 , w16494 , w16495 , w16496 , w16497 , w16498 , w16499 , w16500 , w16501 , w16502 , w16503 , w16504 , w16505 , w16506 , w16507 , w16508 , w16509 , w16510 , w16511 , w16512 , w16513 , w16514 , w16515 , w16516 , w16517 , w16518 , w16519 , w16520 , w16521 , w16522 , w16523 , w16524 , w16525 , w16526 , w16527 , w16528 , w16529 , w16530 , w16531 , w16532 , w16533 , w16534 , w16535 , w16536 , w16537 , w16538 , w16539 , w16540 , w16541 , w16542 , w16543 , w16544 , w16545 , w16546 , w16547 , w16548 , w16549 , w16550 , w16551 , w16552 , w16553 , w16554 , w16555 , w16556 , w16557 , w16558 , w16559 , w16560 , w16561 , w16562 , w16563 , w16564 , w16565 , w16566 , w16567 , w16568 , w16569 , w16570 , w16571 , w16572 , w16573 , w16574 , w16575 , w16576 , w16577 , w16578 , w16579 , w16580 , w16581 , w16582 , w16583 , w16584 , w16585 , w16586 , w16587 , w16588 , w16589 , w16590 , w16591 , w16592 , w16593 , w16594 , w16595 , w16596 , w16597 , w16598 , w16599 , w16600 , w16601 , w16602 , w16603 , w16604 , w16605 , w16606 , w16607 , w16608 , w16609 , w16610 , w16611 , w16612 , w16613 , w16614 , w16615 , w16616 , w16617 , w16618 , w16619 , w16620 , w16621 , w16622 , w16623 , w16624 , w16625 , w16626 , w16627 , w16628 , w16629 , w16630 , w16631 , w16632 , w16633 , w16634 , w16635 , w16636 , w16637 , w16638 , w16639 , w16640 , w16641 , w16642 , w16643 , w16644 , w16645 , w16646 , w16647 , w16648 , w16649 , w16650 , w16651 , w16652 , w16653 , w16654 , w16655 , w16656 , w16657 , w16658 , w16659 , w16660 , w16661 , w16662 , w16663 , w16664 , w16665 , w16666 , w16667 , w16668 , w16669 , w16670 , w16671 , w16672 , w16673 , w16674 , w16675 , w16676 , w16677 , w16678 , w16679 , w16680 , w16681 , w16682 , w16683 , w16684 , w16685 , w16686 , w16687 , w16688 , w16689 , w16690 , w16691 , w16692 , w16693 , w16694 , w16695 , w16696 , w16697 , w16698 , w16699 , w16700 , w16701 , w16702 , w16703 , w16704 , w16705 , w16706 , w16707 , w16708 , w16709 , w16710 , w16711 , w16712 , w16713 , w16714 , w16715 , w16716 , w16717 , w16718 , w16719 , w16720 , w16721 , w16722 , w16723 , w16724 , w16725 , w16726 , w16727 , w16728 , w16729 , w16730 , w16731 , w16732 , w16733 , w16734 , w16735 , w16736 , w16737 , w16738 , w16739 , w16740 , w16741 , w16742 , w16743 , w16744 , w16745 , w16746 , w16747 , w16748 , w16749 , w16750 , w16751 , w16752 , w16753 , w16754 , w16755 , w16756 , w16757 , w16758 , w16759 , w16760 , w16761 , w16762 , w16763 , w16764 , w16765 , w16766 , w16767 , w16768 , w16769 , w16770 , w16771 , w16772 , w16773 , w16774 , w16775 , w16776 , w16777 , w16778 , w16779 , w16780 , w16781 , w16782 , w16783 , w16784 , w16785 , w16786 , w16787 , w16788 , w16789 , w16790 , w16791 , w16792 , w16793 , w16794 , w16795 , w16796 , w16797 , w16798 , w16799 , w16800 , w16801 , w16802 , w16803 , w16804 , w16805 , w16806 , w16807 , w16808 , w16809 , w16810 , w16811 , w16812 , w16813 , w16814 , w16815 , w16816 , w16817 , w16818 , w16819 , w16820 , w16821 , w16822 , w16823 , w16824 , w16825 , w16826 , w16827 , w16828 , w16829 , w16830 , w16831 , w16832 , w16833 , w16834 , w16835 , w16836 , w16837 , w16838 , w16839 , w16840 , w16841 , w16842 , w16843 , w16844 , w16845 , w16846 , w16847 , w16848 , w16849 , w16850 , w16851 , w16852 , w16853 , w16854 , w16855 , w16856 , w16857 , w16858 , w16859 , w16860 , w16861 , w16862 , w16863 , w16864 , w16865 , w16866 , w16867 , w16868 , w16869 , w16870 , w16871 , w16872 , w16873 , w16874 , w16875 , w16876 , w16877 , w16878 , w16879 , w16880 , w16881 , w16882 , w16883 , w16884 , w16885 , w16886 , w16887 , w16888 , w16889 , w16890 , w16891 , w16892 , w16893 , w16894 , w16895 , w16896 , w16897 , w16898 , w16899 , w16900 , w16901 , w16902 , w16903 , w16904 , w16905 , w16906 , w16907 , w16908 , w16909 , w16910 , w16911 , w16912 , w16913 , w16914 , w16915 , w16916 , w16917 , w16918 , w16919 , w16920 , w16921 , w16922 , w16923 , w16924 , w16925 , w16926 , w16927 , w16928 , w16929 , w16930 , w16931 , w16932 , w16933 , w16934 , w16935 , w16936 , w16937 , w16938 , w16939 , w16940 , w16941 , w16942 , w16943 , w16944 , w16945 , w16946 , w16947 , w16948 , w16949 , w16950 , w16951 , w16952 , w16953 , w16954 , w16955 , w16956 , w16957 , w16958 , w16959 , w16960 , w16961 , w16962 , w16963 , w16964 , w16965 , w16966 , w16967 , w16968 , w16969 , w16970 , w16971 , w16972 , w16973 , w16974 , w16975 , w16976 , w16977 , w16978 , w16979 , w16980 , w16981 , w16982 , w16983 , w16984 , w16985 , w16986 , w16987 , w16988 , w16989 , w16990 , w16991 , w16992 , w16993 , w16994 , w16995 , w16996 , w16997 , w16998 , w16999 , w17000 , w17001 , w17002 , w17003 , w17004 , w17005 , w17006 , w17007 , w17008 , w17009 , w17010 , w17011 , w17012 , w17013 , w17014 , w17015 , w17016 , w17017 , w17018 , w17019 , w17020 , w17021 , w17022 , w17023 , w17024 , w17025 , w17026 , w17027 , w17028 , w17029 , w17030 , w17031 , w17032 , w17033 , w17034 , w17035 , w17036 , w17037 , w17038 , w17039 , w17040 , w17041 , w17042 , w17043 , w17044 , w17045 , w17046 , w17047 , w17048 , w17049 , w17050 , w17051 , w17052 , w17053 , w17054 , w17055 , w17056 , w17057 , w17058 , w17059 , w17060 , w17061 , w17062 , w17063 , w17064 , w17065 , w17066 , w17067 , w17068 , w17069 , w17070 , w17071 , w17072 , w17073 , w17074 , w17075 , w17076 , w17077 , w17078 , w17079 , w17080 , w17081 , w17082 , w17083 , w17084 , w17085 , w17086 , w17087 , w17088 , w17089 , w17090 , w17091 , w17092 , w17093 , w17094 , w17095 , w17096 , w17097 , w17098 , w17099 , w17100 , w17101 , w17102 , w17103 , w17104 , w17105 , w17106 , w17107 , w17108 , w17109 , w17110 , w17111 , w17112 , w17113 , w17114 , w17115 , w17116 , w17117 , w17118 , w17119 , w17120 , w17121 , w17122 , w17123 , w17124 , w17125 , w17126 , w17127 , w17128 , w17129 , w17130 , w17131 , w17132 , w17133 , w17134 , w17135 , w17136 , w17137 , w17138 , w17139 , w17140 , w17141 , w17142 , w17143 , w17144 , w17145 , w17146 , w17147 , w17148 , w17149 , w17150 , w17151 , w17152 , w17153 , w17154 , w17155 , w17156 , w17157 , w17158 , w17159 , w17160 , w17161 , w17162 , w17163 , w17164 , w17165 , w17166 , w17167 , w17168 , w17169 , w17170 , w17171 , w17172 , w17173 , w17174 , w17175 , w17176 , w17177 , w17178 , w17179 , w17180 , w17181 , w17182 , w17183 , w17184 , w17185 , w17186 , w17187 , w17188 , w17189 , w17190 , w17191 , w17192 , w17193 , w17194 , w17195 , w17196 , w17197 , w17198 , w17199 , w17200 , w17201 , w17202 , w17203 , w17204 , w17205 , w17206 , w17207 , w17208 , w17209 , w17210 , w17211 , w17212 , w17213 , w17214 , w17215 , w17216 , w17217 , w17218 , w17219 , w17220 , w17221 , w17222 , w17223 , w17224 , w17225 , w17226 , w17227 , w17228 , w17229 , w17230 , w17231 , w17232 , w17233 , w17234 , w17235 , w17236 , w17237 , w17238 , w17239 , w17240 , w17241 , w17242 , w17243 , w17244 , w17245 , w17246 , w17247 , w17248 , w17249 , w17250 , w17251 , w17252 , w17253 , w17254 , w17255 , w17256 , w17257 , w17258 , w17259 , w17260 , w17261 , w17262 , w17263 , w17264 , w17265 , w17266 , w17267 , w17268 , w17269 , w17270 , w17271 , w17272 , w17273 , w17274 , w17275 , w17276 , w17277 , w17278 , w17279 , w17280 , w17281 , w17282 , w17283 , w17284 , w17285 , w17286 , w17287 , w17288 , w17289 , w17290 , w17291 , w17292 , w17293 , w17294 , w17295 , w17296 , w17297 , w17298 , w17299 , w17300 , w17301 , w17302 , w17303 , w17304 , w17305 , w17306 , w17307 , w17308 , w17309 , w17310 , w17311 , w17312 , w17313 , w17314 , w17315 , w17316 , w17317 , w17318 , w17319 , w17320 , w17321 , w17322 , w17323 , w17324 , w17325 , w17326 , w17327 , w17328 , w17329 , w17330 , w17331 , w17332 , w17333 , w17334 , w17335 , w17336 , w17337 , w17338 , w17339 , w17340 , w17341 , w17342 , w17343 , w17344 , w17345 , w17346 , w17347 , w17348 , w17349 , w17350 , w17351 , w17352 , w17353 , w17354 , w17355 , w17356 , w17357 , w17358 , w17359 , w17360 , w17361 , w17362 , w17363 , w17364 , w17365 , w17366 , w17367 , w17368 , w17369 , w17370 , w17371 , w17372 , w17373 , w17374 , w17375 , w17376 , w17377 , w17378 , w17379 , w17380 , w17381 , w17382 , w17383 , w17384 , w17385 , w17386 , w17387 , w17388 , w17389 , w17390 , w17391 , w17392 , w17393 , w17394 , w17395 , w17396 , w17397 , w17398 , w17399 , w17400 , w17401 , w17402 , w17403 , w17404 , w17405 , w17406 , w17407 , w17408 , w17409 , w17410 , w17411 , w17412 , w17413 , w17414 , w17415 , w17416 , w17417 , w17418 , w17419 , w17420 , w17421 , w17422 , w17423 , w17424 , w17425 , w17426 , w17427 , w17428 , w17429 , w17430 , w17431 , w17432 , w17433 , w17434 , w17435 , w17436 , w17437 , w17438 , w17439 , w17440 , w17441 , w17442 , w17443 , w17444 , w17445 , w17446 , w17447 , w17448 , w17449 , w17450 , w17451 , w17452 , w17453 , w17454 , w17455 , w17456 , w17457 , w17458 , w17459 , w17460 , w17461 , w17462 , w17463 , w17464 , w17465 , w17466 , w17467 , w17468 , w17469 , w17470 , w17471 , w17472 , w17473 , w17474 , w17475 , w17476 , w17477 , w17478 , w17479 , w17480 , w17481 , w17482 , w17483 , w17484 , w17485 , w17486 , w17487 , w17488 , w17489 , w17490 , w17491 , w17492 , w17493 , w17494 , w17495 , w17496 , w17497 , w17498 , w17499 , w17500 , w17501 , w17502 , w17503 , w17504 , w17505 , w17506 , w17507 , w17508 , w17509 , w17510 , w17511 , w17512 , w17513 , w17514 , w17515 , w17516 , w17517 , w17518 , w17519 , w17520 , w17521 , w17522 , w17523 , w17524 , w17525 , w17526 , w17527 , w17528 , w17529 , w17530 , w17531 , w17532 , w17533 , w17534 , w17535 , w17536 , w17537 , w17538 , w17539 , w17540 , w17541 , w17542 , w17543 , w17544 , w17545 , w17546 , w17547 , w17548 , w17549 , w17550 , w17551 , w17552 , w17553 , w17554 , w17555 , w17556 , w17557 , w17558 , w17559 , w17560 , w17561 , w17562 , w17563 , w17564 , w17565 , w17566 , w17567 , w17568 , w17569 , w17570 , w17571 , w17572 , w17573 , w17574 , w17575 , w17576 , w17577 , w17578 , w17579 , w17580 , w17581 , w17582 , w17583 , w17584 , w17585 , w17586 , w17587 , w17588 , w17589 , w17590 , w17591 , w17592 , w17593 , w17594 , w17595 , w17596 , w17597 , w17598 , w17599 , w17600 , w17601 , w17602 , w17603 , w17604 , w17605 , w17606 , w17607 , w17608 , w17609 , w17610 , w17611 , w17612 , w17613 , w17614 , w17615 , w17616 , w17617 , w17618 , w17619 , w17620 , w17621 , w17622 , w17623 , w17624 , w17625 , w17626 , w17627 , w17628 , w17629 , w17630 , w17631 , w17632 , w17633 , w17634 , w17635 , w17636 , w17637 , w17638 , w17639 , w17640 , w17641 , w17642 , w17643 , w17644 , w17645 , w17646 , w17647 , w17648 , w17649 , w17650 , w17651 , w17652 , w17653 , w17654 , w17655 , w17656 , w17657 , w17658 , w17659 , w17660 , w17661 , w17662 , w17663 , w17664 , w17665 , w17666 , w17667 , w17668 , w17669 , w17670 , w17671 , w17672 , w17673 , w17674 , w17675 , w17676 , w17677 , w17678 , w17679 , w17680 , w17681 , w17682 , w17683 , w17684 , w17685 , w17686 , w17687 , w17688 , w17689 , w17690 , w17691 , w17692 , w17693 , w17694 , w17695 , w17696 , w17697 , w17698 , w17699 , w17700 , w17701 , w17702 , w17703 , w17704 , w17705 , w17706 , w17707 , w17708 , w17709 , w17710 , w17711 , w17712 , w17713 , w17714 , w17715 , w17716 , w17717 , w17718 , w17719 , w17720 , w17721 , w17722 , w17723 , w17724 , w17725 , w17726 , w17727 , w17728 , w17729 , w17730 , w17731 , w17732 , w17733 , w17734 , w17735 , w17736 , w17737 , w17738 , w17739 , w17740 , w17741 , w17742 , w17743 , w17744 , w17745 , w17746 , w17747 , w17748 , w17749 , w17750 , w17751 , w17752 , w17753 , w17754 , w17755 , w17756 , w17757 , w17758 , w17759 , w17760 , w17761 , w17762 , w17763 , w17764 , w17765 , w17766 , w17767 , w17768 , w17769 , w17770 , w17771 , w17772 , w17773 , w17774 , w17775 , w17776 , w17777 , w17778 , w17779 , w17780 , w17781 , w17782 , w17783 , w17784 , w17785 , w17786 , w17787 , w17788 , w17789 , w17790 , w17791 , w17792 , w17793 , w17794 , w17795 , w17796 , w17797 , w17798 , w17799 , w17800 , w17801 , w17802 , w17803 , w17804 , w17805 , w17806 , w17807 , w17808 , w17809 , w17810 , w17811 , w17812 , w17813 , w17814 , w17815 , w17816 , w17817 , w17818 , w17819 , w17820 , w17821 , w17822 , w17823 , w17824 , w17825 , w17826 , w17827 , w17828 , w17829 , w17830 , w17831 , w17832 , w17833 , w17834 , w17835 , w17836 , w17837 , w17838 , w17839 , w17840 , w17841 , w17842 , w17843 , w17844 , w17845 , w17846 , w17847 , w17848 , w17849 , w17850 , w17851 , w17852 , w17853 , w17854 , w17855 , w17856 , w17857 , w17858 , w17859 , w17860 , w17861 , w17862 , w17863 , w17864 , w17865 , w17866 , w17867 , w17868 , w17869 , w17870 , w17871 , w17872 , w17873 , w17874 , w17875 , w17876 , w17877 , w17878 , w17879 , w17880 , w17881 , w17882 , w17883 , w17884 , w17885 , w17886 , w17887 , w17888 , w17889 , w17890 , w17891 , w17892 , w17893 , w17894 , w17895 , w17896 , w17897 , w17898 , w17899 , w17900 , w17901 , w17902 , w17903 , w17904 , w17905 , w17906 , w17907 , w17908 , w17909 , w17910 , w17911 , w17912 , w17913 , w17914 , w17915 , w17916 , w17917 , w17918 , w17919 , w17920 , w17921 , w17922 , w17923 , w17924 , w17925 , w17926 , w17927 , w17928 , w17929 , w17930 , w17931 , w17932 , w17933 , w17934 , w17935 , w17936 , w17937 , w17938 , w17939 , w17940 , w17941 , w17942 , w17943 , w17944 , w17945 , w17946 , w17947 , w17948 , w17949 , w17950 , w17951 , w17952 , w17953 , w17954 , w17955 , w17956 , w17957 , w17958 , w17959 , w17960 , w17961 , w17962 , w17963 , w17964 , w17965 , w17966 , w17967 , w17968 , w17969 , w17970 , w17971 , w17972 , w17973 , w17974 , w17975 , w17976 , w17977 , w17978 , w17979 , w17980 , w17981 , w17982 , w17983 , w17984 , w17985 , w17986 , w17987 , w17988 , w17989 , w17990 , w17991 , w17992 , w17993 , w17994 , w17995 , w17996 , w17997 , w17998 , w17999 , w18000 , w18001 , w18002 , w18003 , w18004 , w18005 , w18006 , w18007 , w18008 , w18009 , w18010 , w18011 , w18012 , w18013 , w18014 , w18015 , w18016 , w18017 , w18018 , w18019 , w18020 , w18021 , w18022 , w18023 , w18024 , w18025 , w18026 , w18027 , w18028 , w18029 , w18030 , w18031 , w18032 , w18033 , w18034 , w18035 , w18036 , w18037 , w18038 , w18039 , w18040 , w18041 , w18042 , w18043 , w18044 , w18045 , w18046 , w18047 , w18048 , w18049 , w18050 , w18051 , w18052 , w18053 , w18054 , w18055 , w18056 , w18057 , w18058 , w18059 , w18060 , w18061 , w18062 , w18063 , w18064 , w18065 , w18066 , w18067 , w18068 , w18069 , w18070 , w18071 , w18072 , w18073 , w18074 , w18075 , w18076 , w18077 , w18078 , w18079 , w18080 , w18081 , w18082 , w18083 , w18084 , w18085 , w18086 , w18087 , w18088 , w18089 , w18090 , w18091 , w18092 , w18093 , w18094 , w18095 , w18096 , w18097 , w18098 , w18099 , w18100 , w18101 , w18102 , w18103 , w18104 , w18105 , w18106 , w18107 , w18108 , w18109 , w18110 , w18111 , w18112 , w18113 , w18114 , w18115 , w18116 , w18117 , w18118 , w18119 , w18120 , w18121 , w18122 , w18123 , w18124 , w18125 , w18126 , w18127 , w18128 , w18129 , w18130 , w18131 , w18132 , w18133 , w18134 , w18135 , w18136 , w18137 , w18138 , w18139 , w18140 , w18141 , w18142 , w18143 , w18144 , w18145 , w18146 , w18147 , w18148 , w18149 , w18150 , w18151 , w18152 , w18153 , w18154 , w18155 , w18156 , w18157 , w18158 , w18159 , w18160 , w18161 , w18162 , w18163 , w18164 , w18165 , w18166 , w18167 , w18168 , w18169 , w18170 , w18171 , w18172 , w18173 , w18174 , w18175 , w18176 , w18177 , w18178 , w18179 , w18180 , w18181 , w18182 , w18183 , w18184 , w18185 , w18186 , w18187 , w18188 , w18189 , w18190 , w18191 , w18192 , w18193 , w18194 , w18195 , w18196 , w18197 , w18198 , w18199 , w18200 , w18201 , w18202 , w18203 , w18204 , w18205 , w18206 , w18207 , w18208 , w18209 , w18210 , w18211 , w18212 , w18213 , w18214 , w18215 , w18216 , w18217 , w18218 , w18219 , w18220 , w18221 , w18222 , w18223 , w18224 , w18225 , w18226 , w18227 , w18228 , w18229 , w18230 , w18231 , w18232 , w18233 , w18234 , w18235 , w18236 , w18237 , w18238 , w18239 , w18240 , w18241 , w18242 , w18243 , w18244 , w18245 , w18246 , w18247 , w18248 , w18249 , w18250 , w18251 , w18252 , w18253 , w18254 , w18255 , w18256 , w18257 , w18258 , w18259 , w18260 , w18261 , w18262 , w18263 , w18264 , w18265 , w18266 , w18267 , w18268 , w18269 , w18270 , w18271 , w18272 , w18273 , w18274 , w18275 , w18276 , w18277 , w18278 , w18279 , w18280 , w18281 , w18282 , w18283 , w18284 , w18285 , w18286 , w18287 , w18288 , w18289 , w18290 , w18291 , w18292 , w18293 , w18294 , w18295 , w18296 , w18297 , w18298 , w18299 , w18300 , w18301 , w18302 , w18303 , w18304 , w18305 , w18306 , w18307 , w18308 , w18309 , w18310 , w18311 , w18312 , w18313 , w18314 , w18315 , w18316 , w18317 , w18318 , w18319 , w18320 , w18321 , w18322 , w18323 , w18324 , w18325 , w18326 , w18327 , w18328 , w18329 , w18330 , w18331 , w18332 , w18333 , w18334 , w18335 , w18336 , w18337 , w18338 , w18339 , w18340 , w18341 , w18342 , w18343 , w18344 , w18345 , w18346 , w18347 , w18348 , w18349 , w18350 , w18351 , w18352 , w18353 , w18354 , w18355 , w18356 , w18357 , w18358 , w18359 , w18360 , w18361 , w18362 , w18363 , w18364 , w18365 , w18366 , w18367 , w18368 , w18369 , w18370 , w18371 , w18372 , w18373 , w18374 , w18375 , w18376 , w18377 , w18378 , w18379 , w18380 , w18381 , w18382 , w18383 , w18384 , w18385 , w18386 , w18387 , w18388 , w18389 , w18390 , w18391 , w18392 , w18393 , w18394 , w18395 , w18396 , w18397 , w18398 , w18399 , w18400 , w18401 , w18402 , w18403 , w18404 , w18405 , w18406 , w18407 , w18408 , w18409 , w18410 , w18411 , w18412 , w18413 , w18414 , w18415 , w18416 , w18417 , w18418 , w18419 , w18420 , w18421 , w18422 , w18423 , w18424 , w18425 , w18426 , w18427 , w18428 , w18429 , w18430 , w18431 , w18432 , w18433 , w18434 , w18435 , w18436 , w18437 , w18438 , w18439 , w18440 , w18441 , w18442 , w18443 , w18444 , w18445 , w18446 , w18447 , w18448 , w18449 , w18450 , w18451 , w18452 , w18453 , w18454 , w18455 , w18456 , w18457 , w18458 , w18459 , w18460 , w18461 , w18462 , w18463 , w18464 , w18465 , w18466 , w18467 , w18468 , w18469 , w18470 , w18471 , w18472 , w18473 , w18474 , w18475 , w18476 , w18477 , w18478 , w18479 , w18480 , w18481 , w18482 , w18483 , w18484 , w18485 , w18486 , w18487 , w18488 , w18489 , w18490 , w18491 , w18492 , w18493 , w18494 , w18495 , w18496 , w18497 , w18498 , w18499 , w18500 , w18501 , w18502 , w18503 , w18504 , w18505 , w18506 , w18507 , w18508 , w18509 , w18510 , w18511 , w18512 , w18513 , w18514 , w18515 , w18516 , w18517 , w18518 , w18519 , w18520 , w18521 , w18522 , w18523 , w18524 , w18525 , w18526 , w18527 , w18528 , w18529 , w18530 , w18531 , w18532 , w18533 , w18534 , w18535 , w18536 , w18537 , w18538 , w18539 , w18540 , w18541 , w18542 , w18543 , w18544 , w18545 , w18546 , w18547 , w18548 , w18549 , w18550 , w18551 , w18552 , w18553 , w18554 , w18555 , w18556 , w18557 , w18558 , w18559 , w18560 , w18561 , w18562 , w18563 , w18564 , w18565 , w18566 , w18567 , w18568 , w18569 , w18570 , w18571 , w18572 , w18573 , w18574 , w18575 , w18576 , w18577 , w18578 , w18579 , w18580 , w18581 , w18582 , w18583 , w18584 , w18585 , w18586 , w18587 , w18588 , w18589 , w18590 , w18591 , w18592 , w18593 , w18594 , w18595 , w18596 , w18597 , w18598 , w18599 , w18600 , w18601 , w18602 , w18603 , w18604 , w18605 , w18606 , w18607 , w18608 , w18609 , w18610 , w18611 , w18612 , w18613 , w18614 , w18615 , w18616 , w18617 , w18618 , w18619 , w18620 , w18621 , w18622 , w18623 , w18624 , w18625 , w18626 , w18627 , w18628 , w18629 , w18630 , w18631 , w18632 , w18633 , w18634 , w18635 , w18636 , w18637 , w18638 , w18639 , w18640 , w18641 , w18642 , w18643 , w18644 , w18645 , w18646 , w18647 , w18648 , w18649 , w18650 , w18651 , w18652 , w18653 , w18654 , w18655 , w18656 , w18657 , w18658 , w18659 , w18660 , w18661 , w18662 , w18663 , w18664 , w18665 , w18666 , w18667 , w18668 , w18669 , w18670 , w18671 , w18672 , w18673 , w18674 , w18675 , w18676 , w18677 , w18678 , w18679 , w18680 , w18681 , w18682 , w18683 , w18684 , w18685 , w18686 , w18687 , w18688 , w18689 , w18690 , w18691 , w18692 , w18693 , w18694 , w18695 , w18696 , w18697 , w18698 , w18699 , w18700 , w18701 , w18702 , w18703 , w18704 , w18705 , w18706 , w18707 , w18708 , w18709 , w18710 , w18711 , w18712 , w18713 , w18714 , w18715 , w18716 , w18717 , w18718 , w18719 , w18720 , w18721 , w18722 , w18723 , w18724 , w18725 , w18726 , w18727 , w18728 , w18729 , w18730 , w18731 , w18732 , w18733 , w18734 , w18735 , w18736 , w18737 , w18738 , w18739 , w18740 , w18741 , w18742 , w18743 , w18744 , w18745 , w18746 , w18747 , w18748 , w18749 , w18750 , w18751 , w18752 , w18753 , w18754 , w18755 , w18756 , w18757 , w18758 , w18759 , w18760 , w18761 , w18762 , w18763 , w18764 , w18765 , w18766 , w18767 , w18768 , w18769 , w18770 , w18771 , w18772 , w18773 , w18774 , w18775 , w18776 , w18777 , w18778 , w18779 , w18780 , w18781 , w18782 , w18783 , w18784 , w18785 , w18786 , w18787 , w18788 , w18789 , w18790 , w18791 , w18792 , w18793 , w18794 , w18795 , w18796 , w18797 , w18798 , w18799 , w18800 , w18801 , w18802 , w18803 , w18804 , w18805 , w18806 , w18807 , w18808 , w18809 , w18810 , w18811 , w18812 , w18813 , w18814 , w18815 , w18816 , w18817 , w18818 , w18819 , w18820 , w18821 , w18822 , w18823 , w18824 , w18825 , w18826 , w18827 , w18828 , w18829 , w18830 , w18831 , w18832 , w18833 , w18834 , w18835 , w18836 , w18837 , w18838 , w18839 , w18840 , w18841 , w18842 , w18843 , w18844 , w18845 , w18846 , w18847 , w18848 , w18849 , w18850 , w18851 , w18852 , w18853 , w18854 , w18855 , w18856 , w18857 , w18858 , w18859 , w18860 , w18861 , w18862 , w18863 , w18864 , w18865 , w18866 , w18867 , w18868 , w18869 , w18870 , w18871 , w18872 , w18873 , w18874 , w18875 , w18876 , w18877 , w18878 , w18879 , w18880 , w18881 , w18882 , w18883 , w18884 , w18885 , w18886 , w18887 , w18888 , w18889 , w18890 , w18891 , w18892 , w18893 , w18894 , w18895 , w18896 , w18897 , w18898 , w18899 , w18900 , w18901 , w18902 , w18903 , w18904 , w18905 , w18906 , w18907 , w18908 , w18909 , w18910 , w18911 , w18912 , w18913 , w18914 , w18915 , w18916 , w18917 , w18918 , w18919 , w18920 , w18921 , w18922 , w18923 , w18924 , w18925 , w18926 , w18927 , w18928 , w18929 , w18930 , w18931 , w18932 , w18933 , w18934 , w18935 , w18936 , w18937 , w18938 , w18939 , w18940 , w18941 , w18942 , w18943 , w18944 , w18945 , w18946 , w18947 , w18948 , w18949 , w18950 , w18951 , w18952 , w18953 , w18954 , w18955 , w18956 , w18957 , w18958 , w18959 , w18960 , w18961 , w18962 , w18963 , w18964 , w18965 , w18966 , w18967 , w18968 , w18969 , w18970 , w18971 , w18972 , w18973 , w18974 , w18975 , w18976 , w18977 , w18978 , w18979 , w18980 , w18981 , w18982 , w18983 , w18984 , w18985 , w18986 , w18987 , w18988 , w18989 , w18990 , w18991 , w18992 , w18993 , w18994 , w18995 , w18996 , w18997 , w18998 , w18999 , w19000 , w19001 , w19002 , w19003 , w19004 , w19005 , w19006 , w19007 , w19008 , w19009 , w19010 , w19011 , w19012 , w19013 , w19014 , w19015 , w19016 , w19017 , w19018 , w19019 , w19020 , w19021 , w19022 , w19023 , w19024 , w19025 , w19026 , w19027 , w19028 , w19029 , w19030 , w19031 , w19032 , w19033 , w19034 , w19035 , w19036 , w19037 , w19038 , w19039 , w19040 , w19041 , w19042 , w19043 , w19044 , w19045 , w19046 , w19047 , w19048 , w19049 , w19050 , w19051 , w19052 , w19053 , w19054 , w19055 , w19056 , w19057 , w19058 , w19059 , w19060 , w19061 , w19062 , w19063 , w19064 , w19065 , w19066 , w19067 , w19068 , w19069 , w19070 , w19071 , w19072 , w19073 , w19074 , w19075 , w19076 , w19077 , w19078 , w19079 , w19080 , w19081 , w19082 , w19083 , w19084 , w19085 , w19086 , w19087 , w19088 , w19089 , w19090 , w19091 , w19092 , w19093 , w19094 , w19095 , w19096 , w19097 , w19098 , w19099 , w19100 , w19101 , w19102 , w19103 , w19104 , w19105 , w19106 , w19107 , w19108 , w19109 , w19110 , w19111 , w19112 , w19113 , w19114 , w19115 , w19116 , w19117 , w19118 , w19119 , w19120 , w19121 , w19122 , w19123 , w19124 , w19125 , w19126 , w19127 , w19128 , w19129 , w19130 , w19131 , w19132 , w19133 , w19134 , w19135 , w19136 , w19137 , w19138 , w19139 , w19140 , w19141 , w19142 , w19143 , w19144 , w19145 , w19146 , w19147 , w19148 , w19149 , w19150 , w19151 , w19152 , w19153 , w19154 , w19155 , w19156 , w19157 , w19158 , w19159 , w19160 , w19161 , w19162 , w19163 , w19164 , w19165 , w19166 , w19167 , w19168 , w19169 , w19170 , w19171 , w19172 , w19173 , w19174 , w19175 , w19176 , w19177 , w19178 , w19179 , w19180 , w19181 , w19182 , w19183 , w19184 , w19185 , w19186 , w19187 , w19188 , w19189 , w19190 , w19191 , w19192 , w19193 , w19194 , w19195 , w19196 , w19197 , w19198 , w19199 , w19200 , w19201 , w19202 , w19203 , w19204 , w19205 , w19206 , w19207 , w19208 , w19209 , w19210 , w19211 , w19212 , w19213 , w19214 , w19215 , w19216 , w19217 , w19218 , w19219 , w19220 , w19221 , w19222 , w19223 , w19224 , w19225 , w19226 , w19227 , w19228 , w19229 , w19230 , w19231 , w19232 , w19233 , w19234 , w19235 , w19236 , w19237 , w19238 , w19239 , w19240 , w19241 , w19242 , w19243 , w19244 , w19245 , w19246 , w19247 , w19248 , w19249 , w19250 , w19251 , w19252 , w19253 , w19254 , w19255 , w19256 , w19257 , w19258 , w19259 , w19260 , w19261 , w19262 , w19263 , w19264 , w19265 , w19266 , w19267 , w19268 , w19269 , w19270 , w19271 , w19272 , w19273 , w19274 , w19275 , w19276 , w19277 , w19278 , w19279 , w19280 , w19281 , w19282 , w19283 , w19284 , w19285 , w19286 , w19287 , w19288 , w19289 , w19290 , w19291 , w19292 , w19293 , w19294 , w19295 , w19296 , w19297 , w19298 , w19299 , w19300 , w19301 , w19302 , w19303 , w19304 , w19305 , w19306 , w19307 , w19308 , w19309 , w19310 , w19311 , w19312 , w19313 , w19314 , w19315 , w19316 , w19317 , w19318 , w19319 , w19320 , w19321 , w19322 , w19323 , w19324 , w19325 , w19326 , w19327 , w19328 , w19329 , w19330 , w19331 , w19332 , w19333 , w19334 , w19335 , w19336 , w19337 , w19338 , w19339 , w19340 , w19341 , w19342 , w19343 , w19344 , w19345 , w19346 , w19347 , w19348 , w19349 , w19350 , w19351 , w19352 , w19353 , w19354 , w19355 , w19356 , w19357 , w19358 , w19359 , w19360 , w19361 , w19362 , w19363 , w19364 , w19365 , w19366 , w19367 , w19368 , w19369 , w19370 , w19371 , w19372 , w19373 , w19374 , w19375 , w19376 , w19377 , w19378 , w19379 , w19380 , w19381 , w19382 , w19383 , w19384 , w19385 , w19386 , w19387 , w19388 , w19389 , w19390 , w19391 , w19392 , w19393 , w19394 , w19395 , w19396 , w19397 , w19398 , w19399 , w19400 , w19401 , w19402 , w19403 , w19404 , w19405 , w19406 , w19407 , w19408 , w19409 , w19410 , w19411 , w19412 , w19413 , w19414 , w19415 , w19416 , w19417 , w19418 , w19419 , w19420 , w19421 , w19422 , w19423 , w19424 , w19425 , w19426 , w19427 , w19428 , w19429 , w19430 , w19431 , w19432 , w19433 , w19434 , w19435 , w19436 , w19437 , w19438 , w19439 , w19440 , w19441 , w19442 , w19443 , w19444 , w19445 , w19446 , w19447 , w19448 , w19449 , w19450 , w19451 , w19452 , w19453 , w19454 , w19455 , w19456 , w19457 , w19458 , w19459 , w19460 , w19461 , w19462 , w19463 , w19464 , w19465 , w19466 , w19467 , w19468 , w19469 , w19470 , w19471 , w19472 , w19473 , w19474 , w19475 , w19476 , w19477 , w19478 , w19479 , w19480 , w19481 , w19482 , w19483 , w19484 , w19485 , w19486 , w19487 , w19488 , w19489 , w19490 , w19491 , w19492 , w19493 , w19494 , w19495 , w19496 , w19497 , w19498 , w19499 , w19500 , w19501 , w19502 , w19503 , w19504 , w19505 , w19506 , w19507 , w19508 , w19509 , w19510 , w19511 , w19512 , w19513 , w19514 , w19515 , w19516 , w19517 , w19518 , w19519 , w19520 , w19521 , w19522 , w19523 , w19524 , w19525 , w19526 , w19527 , w19528 , w19529 , w19530 , w19531 , w19532 , w19533 , w19534 , w19535 , w19536 , w19537 , w19538 , w19539 , w19540 , w19541 , w19542 , w19543 , w19544 , w19545 , w19546 , w19547 , w19548 , w19549 , w19550 , w19551 , w19552 , w19553 , w19554 , w19555 , w19556 , w19557 , w19558 , w19559 , w19560 , w19561 , w19562 , w19563 , w19564 , w19565 , w19566 , w19567 , w19568 , w19569 , w19570 , w19571 , w19572 , w19573 , w19574 , w19575 , w19576 , w19577 , w19578 , w19579 , w19580 , w19581 , w19582 , w19583 , w19584 , w19585 , w19586 , w19587 , w19588 , w19589 , w19590 , w19591 , w19592 , w19593 , w19594 , w19595 , w19596 , w19597 , w19598 , w19599 , w19600 , w19601 , w19602 , w19603 , w19604 , w19605 , w19606 , w19607 , w19608 , w19609 , w19610 , w19611 , w19612 , w19613 , w19614 , w19615 , w19616 , w19617 , w19618 , w19619 , w19620 , w19621 , w19622 , w19623 , w19624 , w19625 , w19626 , w19627 , w19628 , w19629 , w19630 , w19631 , w19632 , w19633 , w19634 , w19635 , w19636 , w19637 , w19638 , w19639 , w19640 , w19641 , w19642 , w19643 , w19644 , w19645 , w19646 , w19647 , w19648 , w19649 , w19650 , w19651 , w19652 , w19653 , w19654 , w19655 , w19656 , w19657 , w19658 , w19659 , w19660 , w19661 , w19662 , w19663 , w19664 , w19665 , w19666 , w19667 , w19668 , w19669 , w19670 , w19671 , w19672 , w19673 , w19674 , w19675 , w19676 , w19677 , w19678 , w19679 , w19680 , w19681 , w19682 , w19683 , w19684 , w19685 , w19686 , w19687 , w19688 , w19689 , w19690 , w19691 , w19692 , w19693 , w19694 , w19695 , w19696 , w19697 , w19698 , w19699 , w19700 , w19701 , w19702 , w19703 , w19704 , w19705 , w19706 , w19707 , w19708 , w19709 , w19710 , w19711 , w19712 , w19713 , w19714 , w19715 , w19716 , w19717 , w19718 , w19719 , w19720 , w19721 , w19722 , w19723 , w19724 , w19725 , w19726 , w19727 , w19728 , w19729 , w19730 , w19731 , w19732 , w19733 , w19734 , w19735 , w19736 , w19737 , w19738 , w19739 , w19740 , w19741 , w19742 , w19743 , w19744 , w19745 , w19746 , w19747 , w19748 , w19749 , w19750 , w19751 , w19752 , w19753 , w19754 , w19755 , w19756 , w19757 , w19758 , w19759 , w19760 , w19761 , w19762 , w19763 , w19764 , w19765 , w19766 , w19767 , w19768 , w19769 , w19770 , w19771 , w19772 , w19773 , w19774 , w19775 , w19776 , w19777 , w19778 , w19779 , w19780 , w19781 , w19782 , w19783 , w19784 , w19785 , w19786 , w19787 , w19788 , w19789 , w19790 , w19791 , w19792 , w19793 , w19794 , w19795 , w19796 , w19797 , w19798 , w19799 , w19800 , w19801 , w19802 , w19803 , w19804 , w19805 , w19806 , w19807 , w19808 , w19809 , w19810 , w19811 , w19812 , w19813 , w19814 , w19815 , w19816 , w19817 , w19818 , w19819 , w19820 , w19821 , w19822 , w19823 , w19824 , w19825 , w19826 , w19827 , w19828 , w19829 , w19830 , w19831 , w19832 , w19833 , w19834 , w19835 , w19836 , w19837 , w19838 , w19839 , w19840 , w19841 , w19842 , w19843 , w19844 , w19845 , w19846 , w19847 , w19848 , w19849 , w19850 , w19851 , w19852 , w19853 , w19854 , w19855 , w19856 , w19857 , w19858 , w19859 , w19860 , w19861 , w19862 , w19863 , w19864 , w19865 , w19866 , w19867 , w19868 , w19869 , w19870 , w19871 , w19872 , w19873 , w19874 , w19875 , w19876 , w19877 , w19878 , w19879 , w19880 , w19881 , w19882 , w19883 , w19884 , w19885 , w19886 , w19887 , w19888 , w19889 , w19890 , w19891 , w19892 , w19893 , w19894 , w19895 , w19896 , w19897 , w19898 , w19899 , w19900 , w19901 , w19902 , w19903 , w19904 , w19905 , w19906 , w19907 , w19908 , w19909 , w19910 , w19911 , w19912 , w19913 , w19914 , w19915 , w19916 , w19917 , w19918 , w19919 , w19920 , w19921 , w19922 , w19923 , w19924 , w19925 , w19926 , w19927 , w19928 , w19929 , w19930 , w19931 , w19932 , w19933 , w19934 , w19935 , w19936 , w19937 , w19938 , w19939 , w19940 , w19941 , w19942 , w19943 , w19944 , w19945 , w19946 , w19947 , w19948 , w19949 , w19950 , w19951 , w19952 , w19953 , w19954 , w19955 , w19956 , w19957 , w19958 , w19959 , w19960 , w19961 , w19962 , w19963 , w19964 , w19965 , w19966 , w19967 , w19968 , w19969 , w19970 , w19971 , w19972 , w19973 , w19974 , w19975 , w19976 , w19977 , w19978 , w19979 , w19980 , w19981 , w19982 , w19983 , w19984 , w19985 , w19986 , w19987 , w19988 , w19989 , w19990 , w19991 , w19992 , w19993 , w19994 , w19995 , w19996 , w19997 , w19998 , w19999 , w20000 , w20001 , w20002 , w20003 , w20004 , w20005 , w20006 , w20007 , w20008 , w20009 , w20010 , w20011 , w20012 , w20013 , w20014 , w20015 , w20016 , w20017 , w20018 , w20019 , w20020 , w20021 , w20022 , w20023 , w20024 , w20025 , w20026 , w20027 , w20028 , w20029 , w20030 , w20031 , w20032 , w20033 , w20034 , w20035 , w20036 , w20037 , w20038 , w20039 , w20040 , w20041 , w20042 , w20043 , w20044 , w20045 , w20046 , w20047 , w20048 , w20049 , w20050 , w20051 , w20052 , w20053 , w20054 , w20055 , w20056 , w20057 , w20058 , w20059 , w20060 , w20061 , w20062 , w20063 , w20064 , w20065 , w20066 , w20067 , w20068 , w20069 , w20070 , w20071 , w20072 , w20073 , w20074 , w20075 , w20076 , w20077 , w20078 , w20079 , w20080 , w20081 , w20082 , w20083 , w20084 , w20085 , w20086 , w20087 , w20088 , w20089 , w20090 , w20091 , w20092 , w20093 , w20094 , w20095 , w20096 , w20097 , w20098 , w20099 , w20100 , w20101 , w20102 , w20103 , w20104 , w20105 , w20106 , w20107 , w20108 , w20109 , w20110 , w20111 , w20112 , w20113 , w20114 , w20115 , w20116 , w20117 , w20118 , w20119 , w20120 , w20121 , w20122 , w20123 , w20124 , w20125 , w20126 , w20127 , w20128 , w20129 , w20130 , w20131 , w20132 , w20133 , w20134 , w20135 , w20136 , w20137 , w20138 , w20139 , w20140 , w20141 , w20142 , w20143 , w20144 , w20145 , w20146 , w20147 , w20148 , w20149 , w20150 , w20151 , w20152 , w20153 , w20154 , w20155 , w20156 , w20157 , w20158 , w20159 , w20160 , w20161 , w20162 , w20163 , w20164 , w20165 , w20166 , w20167 , w20168 , w20169 , w20170 , w20171 , w20172 , w20173 , w20174 , w20175 , w20176 , w20177 , w20178 , w20179 , w20180 , w20181 , w20182 , w20183 , w20184 , w20185 , w20186 , w20187 , w20188 , w20189 , w20190 , w20191 , w20192 , w20193 , w20194 , w20195 , w20196 , w20197 , w20198 , w20199 , w20200 , w20201 , w20202 , w20203 , w20204 , w20205 , w20206 , w20207 , w20208 , w20209 , w20210 , w20211 , w20212 , w20213 , w20214 , w20215 , w20216 , w20217 , w20218 , w20219 , w20220 , w20221 , w20222 , w20223 , w20224 , w20225 , w20226 , w20227 , w20228 , w20229 , w20230 , w20231 , w20232 , w20233 , w20234 , w20235 , w20236 , w20237 , w20238 , w20239 , w20240 , w20241 , w20242 , w20243 , w20244 , w20245 , w20246 , w20247 , w20248 , w20249 , w20250 , w20251 , w20252 , w20253 , w20254 , w20255 , w20256 , w20257 , w20258 , w20259 , w20260 , w20261 , w20262 , w20263 , w20264 , w20265 , w20266 , w20267 , w20268 , w20269 , w20270 , w20271 , w20272 , w20273 , w20274 , w20275 , w20276 , w20277 , w20278 , w20279 , w20280 , w20281 , w20282 , w20283 , w20284 , w20285 , w20286 , w20287 , w20288 , w20289 , w20290 , w20291 , w20292 , w20293 , w20294 , w20295 , w20296 , w20297 , w20298 , w20299 , w20300 , w20301 , w20302 , w20303 , w20304 , w20305 , w20306 , w20307 , w20308 , w20309 , w20310 , w20311 , w20312 , w20313 , w20314 , w20315 , w20316 , w20317 , w20318 , w20319 , w20320 , w20321 , w20322 , w20323 , w20324 , w20325 , w20326 , w20327 , w20328 , w20329 , w20330 , w20331 , w20332 , w20333 , w20334 , w20335 , w20336 , w20337 , w20338 , w20339 , w20340 , w20341 , w20342 , w20343 , w20344 , w20345 , w20346 , w20347 , w20348 , w20349 , w20350 , w20351 , w20352 , w20353 , w20354 , w20355 , w20356 , w20357 , w20358 , w20359 , w20360 , w20361 , w20362 , w20363 , w20364 , w20365 , w20366 , w20367 , w20368 , w20369 , w20370 , w20371 , w20372 , w20373 , w20374 , w20375 , w20376 , w20377 , w20378 , w20379 , w20380 , w20381 , w20382 , w20383 , w20384 , w20385 , w20386 , w20387 , w20388 , w20389 , w20390 , w20391 , w20392 , w20393 , w20394 , w20395 , w20396 , w20397 , w20398 , w20399 , w20400 , w20401 , w20402 , w20403 , w20404 , w20405 , w20406 , w20407 , w20408 , w20409 , w20410 , w20411 , w20412 , w20413 , w20414 , w20415 , w20416 , w20417 , w20418 , w20419 , w20420 , w20421 , w20422 , w20423 , w20424 , w20425 , w20426 , w20427 , w20428 , w20429 , w20430 , w20431 , w20432 , w20433 , w20434 , w20435 , w20436 , w20437 , w20438 , w20439 , w20440 , w20441 , w20442 , w20443 , w20444 , w20445 , w20446 , w20447 , w20448 , w20449 , w20450 , w20451 , w20452 , w20453 , w20454 , w20455 , w20456 , w20457 , w20458 , w20459 , w20460 , w20461 , w20462 , w20463 , w20464 , w20465 , w20466 , w20467 , w20468 , w20469 , w20470 , w20471 , w20472 , w20473 , w20474 , w20475 , w20476 , w20477 , w20478 , w20479 , w20480 , w20481 , w20482 , w20483 , w20484 , w20485 , w20486 , w20487 , w20488 , w20489 , w20490 , w20491 , w20492 , w20493 , w20494 , w20495 , w20496 , w20497 , w20498 , w20499 , w20500 , w20501 , w20502 , w20503 , w20504 , w20505 , w20506 , w20507 , w20508 , w20509 , w20510 , w20511 , w20512 , w20513 , w20514 , w20515 , w20516 , w20517 , w20518 , w20519 , w20520 , w20521 , w20522 , w20523 , w20524 , w20525 , w20526 , w20527 , w20528 , w20529 , w20530 , w20531 , w20532 , w20533 , w20534 , w20535 , w20536 , w20537 , w20538 , w20539 , w20540 , w20541 , w20542 , w20543 , w20544 , w20545 , w20546 , w20547 , w20548 , w20549 , w20550 , w20551 , w20552 , w20553 , w20554 , w20555 , w20556 , w20557 , w20558 , w20559 , w20560 , w20561 , w20562 , w20563 , w20564 , w20565 , w20566 , w20567 , w20568 , w20569 , w20570 , w20571 , w20572 , w20573 , w20574 , w20575 , w20576 , w20577 , w20578 , w20579 , w20580 , w20581 , w20582 , w20583 , w20584 , w20585 , w20586 , w20587 , w20588 , w20589 , w20590 , w20591 , w20592 , w20593 , w20594 , w20595 , w20596 , w20597 , w20598 , w20599 , w20600 , w20601 , w20602 , w20603 , w20604 , w20605 , w20606 , w20607 , w20608 , w20609 , w20610 , w20611 , w20612 , w20613 , w20614 , w20615 , w20616 , w20617 , w20618 , w20619 , w20620 , w20621 , w20622 , w20623 , w20624 , w20625 , w20626 , w20627 , w20628 , w20629 , w20630 , w20631 , w20632 , w20633 , w20634 , w20635 , w20636 , w20637 , w20638 , w20639 , w20640 , w20641 , w20642 , w20643 , w20644 , w20645 , w20646 , w20647 , w20648 , w20649 , w20650 , w20651 , w20652 , w20653 , w20654 , w20655 , w20656 , w20657 , w20658 , w20659 , w20660 , w20661 , w20662 , w20663 , w20664 , w20665 , w20666 , w20667 , w20668 , w20669 , w20670 , w20671 , w20672 , w20673 , w20674 , w20675 , w20676 , w20677 , w20678 , w20679 , w20680 , w20681 , w20682 , w20683 , w20684 , w20685 , w20686 , w20687 , w20688 , w20689 , w20690 , w20691 , w20692 , w20693 , w20694 , w20695 , w20696 , w20697 , w20698 , w20699 , w20700 , w20701 , w20702 , w20703 , w20704 , w20705 , w20706 , w20707 , w20708 , w20709 , w20710 , w20711 , w20712 , w20713 , w20714 , w20715 , w20716 , w20717 , w20718 , w20719 , w20720 , w20721 , w20722 , w20723 , w20724 , w20725 , w20726 , w20727 , w20728 , w20729 , w20730 , w20731 , w20732 , w20733 , w20734 , w20735 , w20736 , w20737 , w20738 , w20739 , w20740 , w20741 , w20742 , w20743 , w20744 , w20745 , w20746 , w20747 , w20748 , w20749 , w20750 , w20751 , w20752 , w20753 , w20754 , w20755 , w20756 , w20757 , w20758 , w20759 , w20760 , w20761 , w20762 , w20763 , w20764 , w20765 , w20766 , w20767 , w20768 , w20769 , w20770 , w20771 , w20772 , w20773 , w20774 , w20775 , w20776 , w20777 , w20778 , w20779 , w20780 , w20781 , w20782 , w20783 , w20784 , w20785 , w20786 , w20787 , w20788 , w20789 , w20790 , w20791 , w20792 , w20793 , w20794 , w20795 , w20796 , w20797 , w20798 , w20799 , w20800 , w20801 , w20802 , w20803 , w20804 , w20805 , w20806 , w20807 , w20808 , w20809 , w20810 , w20811 , w20812 , w20813 , w20814 , w20815 , w20816 , w20817 , w20818 , w20819 , w20820 , w20821 , w20822 , w20823 , w20824 , w20825 , w20826 , w20827 , w20828 , w20829 , w20830 , w20831 , w20832 , w20833 , w20834 , w20835 , w20836 , w20837 , w20838 , w20839 , w20840 , w20841 , w20842 , w20843 , w20844 , w20845 , w20846 , w20847 , w20848 , w20849 , w20850 , w20851 , w20852 , w20853 , w20854 , w20855 , w20856 , w20857 , w20858 , w20859 , w20860 , w20861 , w20862 , w20863 , w20864 , w20865 , w20866 , w20867 , w20868 , w20869 , w20870 , w20871 , w20872 , w20873 , w20874 , w20875 , w20876 , w20877 , w20878 , w20879 , w20880 , w20881 , w20882 , w20883 , w20884 , w20885 , w20886 , w20887 , w20888 , w20889 , w20890 , w20891 , w20892 , w20893 , w20894 , w20895 , w20896 , w20897 , w20898 , w20899 , w20900 , w20901 , w20902 , w20903 , w20904 , w20905 , w20906 , w20907 , w20908 , w20909 , w20910 , w20911 , w20912 , w20913 , w20914 , w20915 , w20916 , w20917 , w20918 , w20919 , w20920 , w20921 , w20922 , w20923 , w20924 , w20925 , w20926 , w20927 , w20928 , w20929 , w20930 , w20931 , w20932 , w20933 , w20934 , w20935 , w20936 , w20937 , w20938 , w20939 , w20940 , w20941 , w20942 , w20943 , w20944 , w20945 , w20946 , w20947 , w20948 , w20949 , w20950 , w20951 , w20952 , w20953 , w20954 , w20955 , w20956 , w20957 , w20958 , w20959 , w20960 , w20961 , w20962 , w20963 , w20964 , w20965 , w20966 , w20967 , w20968 , w20969 , w20970 , w20971 , w20972 , w20973 , w20974 , w20975 , w20976 , w20977 , w20978 , w20979 , w20980 , w20981 , w20982 , w20983 , w20984 , w20985 , w20986 , w20987 , w20988 , w20989 , w20990 , w20991 , w20992 , w20993 , w20994 , w20995 , w20996 , w20997 , w20998 , w20999 , w21000 , w21001 , w21002 , w21003 , w21004 , w21005 , w21006 , w21007 , w21008 , w21009 , w21010 , w21011 , w21012 , w21013 , w21014 , w21015 , w21016 , w21017 , w21018 , w21019 , w21020 , w21021 , w21022 , w21023 , w21024 , w21025 , w21026 , w21027 , w21028 , w21029 , w21030 , w21031 , w21032 , w21033 , w21034 , w21035 , w21036 , w21037 , w21038 , w21039 , w21040 , w21041 , w21042 , w21043 , w21044 , w21045 , w21046 , w21047 , w21048 , w21049 , w21050 , w21051 , w21052 , w21053 , w21054 , w21055 , w21056 , w21057 , w21058 , w21059 , w21060 , w21061 , w21062 , w21063 , w21064 , w21065 , w21066 , w21067 , w21068 , w21069 , w21070 , w21071 , w21072 , w21073 , w21074 , w21075 , w21076 , w21077 , w21078 , w21079 , w21080 , w21081 , w21082 , w21083 , w21084 , w21085 , w21086 , w21087 , w21088 , w21089 , w21090 , w21091 , w21092 , w21093 , w21094 , w21095 , w21096 , w21097 , w21098 , w21099 , w21100 , w21101 , w21102 , w21103 , w21104 , w21105 , w21106 , w21107 , w21108 , w21109 , w21110 , w21111 , w21112 , w21113 , w21114 , w21115 , w21116 , w21117 , w21118 , w21119 , w21120 , w21121 , w21122 , w21123 , w21124 , w21125 , w21126 , w21127 , w21128 , w21129 , w21130 , w21131 , w21132 , w21133 , w21134 , w21135 , w21136 , w21137 , w21138 , w21139 , w21140 , w21141 , w21142 , w21143 , w21144 , w21145 , w21146 , w21147 , w21148 , w21149 , w21150 , w21151 , w21152 , w21153 , w21154 , w21155 , w21156 , w21157 , w21158 , w21159 , w21160 , w21161 , w21162 , w21163 , w21164 , w21165 , w21166 , w21167 , w21168 , w21169 , w21170 , w21171 , w21172 , w21173 , w21174 , w21175 , w21176 , w21177 , w21178 , w21179 , w21180 , w21181 , w21182 , w21183 , w21184 , w21185 , w21186 , w21187 , w21188 , w21189 , w21190 , w21191 , w21192 , w21193 , w21194 , w21195 , w21196 , w21197 , w21198 , w21199 , w21200 , w21201 , w21202 , w21203 , w21204 , w21205 , w21206 , w21207 , w21208 , w21209 , w21210 , w21211 , w21212 , w21213 , w21214 , w21215 , w21216 , w21217 , w21218 , w21219 , w21220 , w21221 , w21222 , w21223 , w21224 , w21225 , w21226 , w21227 , w21228 , w21229 , w21230 , w21231 , w21232 , w21233 , w21234 , w21235 , w21236 , w21237 , w21238 , w21239 , w21240 , w21241 , w21242 , w21243 , w21244 , w21245 , w21246 , w21247 , w21248 , w21249 , w21250 , w21251 , w21252 , w21253 , w21254 , w21255 , w21256 , w21257 , w21258 , w21259 , w21260 , w21261 , w21262 , w21263 , w21264 , w21265 , w21266 , w21267 , w21268 , w21269 , w21270 , w21271 , w21272 , w21273 , w21274 , w21275 , w21276 , w21277 , w21278 , w21279 , w21280 , w21281 , w21282 , w21283 , w21284 , w21285 , w21286 , w21287 , w21288 , w21289 , w21290 , w21291 , w21292 , w21293 , w21294 , w21295 , w21296 , w21297 , w21298 , w21299 , w21300 , w21301 , w21302 , w21303 , w21304 , w21305 , w21306 , w21307 , w21308 , w21309 , w21310 , w21311 , w21312 , w21313 , w21314 , w21315 , w21316 , w21317 , w21318 , w21319 , w21320 , w21321 , w21322 , w21323 , w21324 , w21325 , w21326 , w21327 , w21328 , w21329 , w21330 , w21331 , w21332 , w21333 , w21334 , w21335 , w21336 , w21337 , w21338 , w21339 , w21340 , w21341 , w21342 , w21343 , w21344 , w21345 , w21346 , w21347 , w21348 , w21349 , w21350 , w21351 , w21352 , w21353 , w21354 , w21355 , w21356 , w21357 , w21358 , w21359 , w21360 , w21361 , w21362 , w21363 , w21364 , w21365 , w21366 , w21367 , w21368 , w21369 , w21370 , w21371 , w21372 , w21373 , w21374 , w21375 , w21376 , w21377 , w21378 , w21379 , w21380 , w21381 , w21382 , w21383 , w21384 , w21385 , w21386 , w21387 , w21388 , w21389 , w21390 , w21391 , w21392 , w21393 , w21394 , w21395 , w21396 , w21397 , w21398 , w21399 , w21400 , w21401 , w21402 , w21403 , w21404 , w21405 , w21406 , w21407 , w21408 , w21409 , w21410 , w21411 , w21412 , w21413 , w21414 , w21415 , w21416 , w21417 , w21418 , w21419 , w21420 , w21421 , w21422 , w21423 , w21424 , w21425 , w21426 , w21427 , w21428 , w21429 , w21430 , w21431 , w21432 , w21433 , w21434 , w21435 , w21436 , w21437 , w21438 , w21439 , w21440 , w21441 , w21442 , w21443 , w21444 , w21445 , w21446 , w21447 , w21448 , w21449 , w21450 , w21451 , w21452 , w21453 , w21454 , w21455 , w21456 , w21457 , w21458 , w21459 , w21460 , w21461 , w21462 , w21463 , w21464 , w21465 , w21466 , w21467 , w21468 , w21469 , w21470 , w21471 , w21472 , w21473 , w21474 , w21475 , w21476 , w21477 , w21478 , w21479 , w21480 , w21481 , w21482 , w21483 , w21484 , w21485 , w21486 , w21487 , w21488 , w21489 , w21490 , w21491 , w21492 , w21493 , w21494 , w21495 , w21496 , w21497 , w21498 , w21499 , w21500 , w21501 , w21502 , w21503 , w21504 , w21505 , w21506 , w21507 , w21508 , w21509 , w21510 , w21511 , w21512 , w21513 , w21514 , w21515 , w21516 , w21517 , w21518 , w21519 , w21520 , w21521 , w21522 , w21523 , w21524 , w21525 , w21526 , w21527 , w21528 , w21529 , w21530 , w21531 , w21532 , w21533 , w21534 , w21535 , w21536 , w21537 , w21538 , w21539 , w21540 , w21541 , w21542 , w21543 , w21544 , w21545 , w21546 , w21547 , w21548 , w21549 , w21550 , w21551 , w21552 , w21553 , w21554 , w21555 , w21556 , w21557 , w21558 , w21559 , w21560 , w21561 , w21562 , w21563 , w21564 , w21565 , w21566 , w21567 , w21568 , w21569 , w21570 , w21571 , w21572 , w21573 , w21574 , w21575 , w21576 , w21577 , w21578 , w21579 , w21580 , w21581 , w21582 , w21583 , w21584 , w21585 , w21586 , w21587 , w21588 , w21589 , w21590 , w21591 , w21592 , w21593 , w21594 , w21595 , w21596 , w21597 , w21598 , w21599 , w21600 , w21601 , w21602 , w21603 , w21604 , w21605 , w21606 , w21607 , w21608 , w21609 , w21610 , w21611 , w21612 , w21613 , w21614 , w21615 , w21616 , w21617 , w21618 , w21619 , w21620 , w21621 , w21622 , w21623 , w21624 , w21625 , w21626 , w21627 , w21628 , w21629 , w21630 , w21631 , w21632 , w21633 , w21634 , w21635 , w21636 , w21637 , w21638 , w21639 , w21640 , w21641 , w21642 , w21643 , w21644 , w21645 , w21646 , w21647 , w21648 , w21649 , w21650 , w21651 , w21652 , w21653 , w21654 , w21655 , w21656 , w21657 , w21658 , w21659 , w21660 , w21661 , w21662 , w21663 , w21664 , w21665 , w21666 , w21667 , w21668 , w21669 , w21670 , w21671 , w21672 , w21673 , w21674 , w21675 , w21676 , w21677 , w21678 , w21679 , w21680 , w21681 , w21682 , w21683 , w21684 , w21685 , w21686 , w21687 , w21688 , w21689 , w21690 , w21691 , w21692 , w21693 , w21694 , w21695 , w21696 , w21697 , w21698 , w21699 , w21700 , w21701 , w21702 , w21703 , w21704 , w21705 , w21706 , w21707 , w21708 , w21709 , w21710 , w21711 , w21712 , w21713 , w21714 , w21715 , w21716 , w21717 , w21718 , w21719 , w21720 , w21721 , w21722 , w21723 , w21724 , w21725 , w21726 , w21727 , w21728 , w21729 , w21730 , w21731 , w21732 , w21733 , w21734 , w21735 , w21736 , w21737 , w21738 , w21739 , w21740 , w21741 , w21742 , w21743 , w21744 , w21745 , w21746 , w21747 , w21748 , w21749 , w21750 , w21751 , w21752 , w21753 , w21754 , w21755 , w21756 , w21757 , w21758 , w21759 , w21760 , w21761 , w21762 , w21763 , w21764 , w21765 , w21766 , w21767 , w21768 , w21769 , w21770 , w21771 , w21772 , w21773 , w21774 , w21775 , w21776 , w21777 , w21778 , w21779 , w21780 , w21781 , w21782 , w21783 , w21784 , w21785 , w21786 , w21787 , w21788 , w21789 , w21790 , w21791 , w21792 , w21793 , w21794 , w21795 , w21796 , w21797 , w21798 , w21799 , w21800 , w21801 , w21802 , w21803 , w21804 , w21805 , w21806 , w21807 , w21808 , w21809 , w21810 , w21811 , w21812 , w21813 , w21814 , w21815 , w21816 , w21817 , w21818 , w21819 , w21820 , w21821 , w21822 , w21823 , w21824 , w21825 , w21826 , w21827 , w21828 , w21829 , w21830 , w21831 , w21832 , w21833 , w21834 , w21835 , w21836 , w21837 , w21838 , w21839 , w21840 , w21841 , w21842 , w21843 , w21844 , w21845 , w21846 , w21847 , w21848 , w21849 , w21850 , w21851 , w21852 , w21853 , w21854 , w21855 , w21856 , w21857 , w21858 , w21859 , w21860 , w21861 , w21862 , w21863 , w21864 , w21865 , w21866 , w21867 , w21868 , w21869 , w21870 , w21871 , w21872 , w21873 , w21874 , w21875 , w21876 , w21877 , w21878 , w21879 , w21880 , w21881 , w21882 , w21883 , w21884 , w21885 , w21886 , w21887 , w21888 , w21889 , w21890 , w21891 , w21892 , w21893 , w21894 , w21895 , w21896 , w21897 , w21898 , w21899 , w21900 , w21901 , w21902 , w21903 , w21904 , w21905 , w21906 , w21907 , w21908 , w21909 , w21910 , w21911 , w21912 , w21913 , w21914 , w21915 , w21916 , w21917 , w21918 , w21919 , w21920 , w21921 , w21922 , w21923 , w21924 , w21925 , w21926 , w21927 , w21928 , w21929 , w21930 , w21931 , w21932 , w21933 , w21934 , w21935 , w21936 , w21937 , w21938 , w21939 , w21940 , w21941 , w21942 , w21943 , w21944 , w21945 , w21946 , w21947 , w21948 , w21949 , w21950 , w21951 , w21952 , w21953 , w21954 , w21955 , w21956 , w21957 , w21958 , w21959 , w21960 , w21961 , w21962 , w21963 , w21964 , w21965 , w21966 , w21967 , w21968 , w21969 , w21970 , w21971 , w21972 , w21973 , w21974 , w21975 , w21976 , w21977 , w21978 , w21979 , w21980 , w21981 , w21982 , w21983 , w21984 , w21985 , w21986 , w21987 , w21988 , w21989 , w21990 , w21991 , w21992 , w21993 , w21994 , w21995 , w21996 , w21997 , w21998 , w21999 , w22000 , w22001 , w22002 , w22003 , w22004 , w22005 , w22006 , w22007 , w22008 , w22009 , w22010 , w22011 , w22012 , w22013 , w22014 , w22015 , w22016 , w22017 , w22018 , w22019 , w22020 , w22021 , w22022 , w22023 , w22024 , w22025 , w22026 , w22027 , w22028 , w22029 , w22030 , w22031 , w22032 , w22033 , w22034 , w22035 , w22036 , w22037 , w22038 , w22039 , w22040 , w22041 , w22042 , w22043 , w22044 , w22045 , w22046 , w22047 , w22048 , w22049 , w22050 , w22051 , w22052 , w22053 , w22054 , w22055 , w22056 , w22057 , w22058 , w22059 , w22060 , w22061 , w22062 , w22063 , w22064 , w22065 , w22066 , w22067 , w22068 , w22069 , w22070 , w22071 , w22072 , w22073 , w22074 , w22075 , w22076 , w22077 , w22078 , w22079 , w22080 , w22081 , w22082 , w22083 , w22084 , w22085 , w22086 , w22087 , w22088 , w22089 , w22090 , w22091 , w22092 , w22093 , w22094 , w22095 , w22096 , w22097 , w22098 , w22099 , w22100 , w22101 , w22102 , w22103 , w22104 , w22105 , w22106 , w22107 , w22108 , w22109 , w22110 , w22111 , w22112 , w22113 , w22114 , w22115 , w22116 , w22117 , w22118 , w22119 , w22120 , w22121 , w22122 , w22123 , w22124 , w22125 , w22126 , w22127 , w22128 , w22129 , w22130 , w22131 , w22132 , w22133 , w22134 , w22135 , w22136 , w22137 , w22138 , w22139 , w22140 , w22141 , w22142 , w22143 , w22144 , w22145 , w22146 , w22147 , w22148 , w22149 , w22150 , w22151 , w22152 , w22153 , w22154 , w22155 , w22156 , w22157 , w22158 , w22159 , w22160 , w22161 , w22162 , w22163 , w22164 , w22165 , w22166 , w22167 , w22168 , w22169 , w22170 , w22171 , w22172 , w22173 , w22174 , w22175 , w22176 , w22177 , w22178 , w22179 , w22180 , w22181 , w22182 , w22183 , w22184 , w22185 , w22186 , w22187 , w22188 , w22189 , w22190 , w22191 , w22192 , w22193 , w22194 , w22195 , w22196 , w22197 , w22198 , w22199 , w22200 , w22201 , w22202 , w22203 , w22204 , w22205 , w22206 , w22207 , w22208 , w22209 , w22210 , w22211 , w22212 , w22213 , w22214 , w22215 , w22216 , w22217 , w22218 , w22219 , w22220 , w22221 , w22222 , w22223 , w22224 , w22225 , w22226 , w22227 , w22228 , w22229 , w22230 , w22231 , w22232 , w22233 , w22234 , w22235 , w22236 , w22237 , w22238 , w22239 , w22240 , w22241 , w22242 , w22243 , w22244 , w22245 , w22246 , w22247 , w22248 , w22249 , w22250 , w22251 , w22252 , w22253 , w22254 , w22255 , w22256 , w22257 , w22258 , w22259 , w22260 , w22261 , w22262 , w22263 , w22264 , w22265 , w22266 , w22267 , w22268 , w22269 , w22270 , w22271 , w22272 , w22273 , w22274 , w22275 , w22276 , w22277 , w22278 , w22279 , w22280 , w22281 , w22282 , w22283 , w22284 , w22285 , w22286 , w22287 , w22288 , w22289 , w22290 , w22291 , w22292 , w22293 , w22294 , w22295 , w22296 , w22297 , w22298 , w22299 , w22300 , w22301 , w22302 , w22303 , w22304 , w22305 , w22306 , w22307 , w22308 , w22309 , w22310 , w22311 , w22312 , w22313 , w22314 , w22315 , w22316 , w22317 , w22318 , w22319 , w22320 , w22321 , w22322 , w22323 , w22324 , w22325 , w22326 , w22327 , w22328 , w22329 , w22330 , w22331 , w22332 , w22333 , w22334 , w22335 , w22336 , w22337 , w22338 , w22339 , w22340 , w22341 , w22342 , w22343 , w22344 , w22345 , w22346 , w22347 , w22348 , w22349 , w22350 , w22351 , w22352 , w22353 , w22354 , w22355 , w22356 , w22357 , w22358 , w22359 , w22360 , w22361 , w22362 , w22363 , w22364 , w22365 , w22366 , w22367 , w22368 , w22369 , w22370 , w22371 , w22372 , w22373 , w22374 , w22375 , w22376 , w22377 , w22378 , w22379 , w22380 , w22381 , w22382 , w22383 , w22384 , w22385 , w22386 , w22387 , w22388 , w22389 , w22390 , w22391 , w22392 , w22393 , w22394 , w22395 , w22396 , w22397 , w22398 , w22399 , w22400 , w22401 , w22402 , w22403 , w22404 , w22405 , w22406 , w22407 , w22408 , w22409 , w22410 , w22411 , w22412 , w22413 , w22414 , w22415 , w22416 , w22417 , w22418 , w22419 , w22420 , w22421 , w22422 , w22423 , w22424 , w22425 , w22426 , w22427 , w22428 , w22429 , w22430 , w22431 , w22432 , w22433 , w22434 , w22435 , w22436 , w22437 , w22438 , w22439 , w22440 , w22441 , w22442 , w22443 , w22444 , w22445 , w22446 , w22447 , w22448 , w22449 , w22450 , w22451 , w22452 , w22453 , w22454 , w22455 , w22456 , w22457 , w22458 , w22459 , w22460 , w22461 , w22462 , w22463 , w22464 , w22465 , w22466 , w22467 , w22468 , w22469 , w22470 , w22471 , w22472 , w22473 , w22474 , w22475 , w22476 , w22477 , w22478 , w22479 , w22480 , w22481 , w22482 , w22483 , w22484 , w22485 , w22486 , w22487 , w22488 , w22489 , w22490 , w22491 , w22492 , w22493 , w22494 , w22495 , w22496 , w22497 , w22498 , w22499 , w22500 , w22501 , w22502 , w22503 , w22504 , w22505 , w22506 , w22507 , w22508 , w22509 , w22510 , w22511 , w22512 , w22513 , w22514 , w22515 , w22516 , w22517 , w22518 , w22519 , w22520 , w22521 , w22522 , w22523 , w22524 , w22525 , w22526 , w22527 , w22528 , w22529 , w22530 , w22531 , w22532 , w22533 , w22534 , w22535 , w22536 , w22537 , w22538 , w22539 , w22540 , w22541 , w22542 , w22543 , w22544 , w22545 , w22546 , w22547 , w22548 , w22549 , w22550 , w22551 , w22552 , w22553 , w22554 , w22555 , w22556 , w22557 , w22558 , w22559 , w22560 , w22561 , w22562 , w22563 , w22564 , w22565 , w22566 , w22567 , w22568 , w22569 , w22570 , w22571 , w22572 , w22573 , w22574 , w22575 , w22576 , w22577 , w22578 , w22579 , w22580 , w22581 , w22582 , w22583 , w22584 , w22585 , w22586 , w22587 , w22588 , w22589 , w22590 , w22591 , w22592 , w22593 , w22594 , w22595 , w22596 , w22597 , w22598 , w22599 , w22600 , w22601 , w22602 , w22603 , w22604 , w22605 , w22606 , w22607 , w22608 , w22609 , w22610 , w22611 , w22612 , w22613 , w22614 , w22615 , w22616 , w22617 , w22618 , w22619 , w22620 , w22621 , w22622 , w22623 , w22624 , w22625 , w22626 , w22627 , w22628 , w22629 , w22630 , w22631 , w22632 , w22633 , w22634 , w22635 , w22636 , w22637 , w22638 , w22639 , w22640 , w22641 , w22642 , w22643 , w22644 , w22645 , w22646 , w22647 , w22648 , w22649 , w22650 , w22651 , w22652 , w22653 , w22654 , w22655 , w22656 , w22657 , w22658 , w22659 , w22660 , w22661 , w22662 , w22663 , w22664 , w22665 , w22666 , w22667 , w22668 , w22669 , w22670 , w22671 , w22672 , w22673 , w22674 , w22675 , w22676 , w22677 , w22678 , w22679 , w22680 , w22681 , w22682 , w22683 , w22684 , w22685 , w22686 , w22687 , w22688 , w22689 , w22690 , w22691 , w22692 , w22693 , w22694 , w22695 , w22696 , w22697 , w22698 , w22699 , w22700 , w22701 , w22702 , w22703 , w22704 , w22705 , w22706 , w22707 , w22708 , w22709 , w22710 , w22711 , w22712 , w22713 , w22714 , w22715 , w22716 , w22717 , w22718 , w22719 , w22720 , w22721 , w22722 , w22723 , w22724 , w22725 , w22726 , w22727 , w22728 , w22729 , w22730 , w22731 , w22732 , w22733 , w22734 , w22735 , w22736 , w22737 , w22738 , w22739 , w22740 , w22741 , w22742 , w22743 , w22744 , w22745 , w22746 , w22747 , w22748 , w22749 , w22750 , w22751 , w22752 , w22753 , w22754 , w22755 , w22756 , w22757 , w22758 , w22759 , w22760 , w22761 , w22762 , w22763 , w22764 , w22765 , w22766 , w22767 , w22768 , w22769 , w22770 , w22771 , w22772 , w22773 , w22774 , w22775 , w22776 , w22777 , w22778 , w22779 , w22780 , w22781 , w22782 , w22783 , w22784 , w22785 , w22786 , w22787 , w22788 , w22789 , w22790 , w22791 , w22792 , w22793 , w22794 , w22795 , w22796 , w22797 , w22798 , w22799 , w22800 , w22801 , w22802 , w22803 , w22804 , w22805 , w22806 , w22807 , w22808 , w22809 , w22810 , w22811 , w22812 , w22813 , w22814 , w22815 , w22816 , w22817 , w22818 , w22819 , w22820 , w22821 , w22822 , w22823 , w22824 , w22825 , w22826 , w22827 , w22828 , w22829 , w22830 , w22831 , w22832 , w22833 , w22834 , w22835 , w22836 , w22837 , w22838 , w22839 , w22840 , w22841 , w22842 , w22843 , w22844 , w22845 , w22846 , w22847 , w22848 , w22849 , w22850 , w22851 , w22852 , w22853 , w22854 , w22855 , w22856 , w22857 , w22858 , w22859 , w22860 , w22861 , w22862 , w22863 , w22864 , w22865 , w22866 , w22867 , w22868 , w22869 , w22870 , w22871 , w22872 , w22873 , w22874 , w22875 , w22876 , w22877 , w22878 , w22879 , w22880 , w22881 , w22882 , w22883 , w22884 , w22885 , w22886 , w22887 , w22888 , w22889 , w22890 , w22891 , w22892 , w22893 , w22894 , w22895 , w22896 , w22897 , w22898 , w22899 , w22900 , w22901 , w22902 , w22903 , w22904 , w22905 , w22906 , w22907 , w22908 , w22909 , w22910 , w22911 , w22912 , w22913 , w22914 , w22915 , w22916 , w22917 , w22918 , w22919 , w22920 , w22921 , w22922 , w22923 , w22924 , w22925 , w22926 , w22927 , w22928 , w22929 , w22930 , w22931 , w22932 , w22933 , w22934 , w22935 , w22936 , w22937 , w22938 , w22939 , w22940 , w22941 , w22942 , w22943 , w22944 , w22945 , w22946 , w22947 , w22948 , w22949 , w22950 , w22951 , w22952 , w22953 , w22954 , w22955 , w22956 , w22957 , w22958 , w22959 , w22960 , w22961 , w22962 , w22963 , w22964 , w22965 , w22966 , w22967 , w22968 , w22969 , w22970 , w22971 , w22972 , w22973 , w22974 , w22975 , w22976 , w22977 , w22978 , w22979 , w22980 , w22981 , w22982 , w22983 , w22984 , w22985 , w22986 , w22987 , w22988 , w22989 , w22990 , w22991 , w22992 , w22993 , w22994 , w22995 , w22996 , w22997 , w22998 , w22999 , w23000 , w23001 , w23002 , w23003 , w23004 , w23005 , w23006 , w23007 , w23008 , w23009 , w23010 , w23011 , w23012 , w23013 , w23014 , w23015 , w23016 , w23017 , w23018 , w23019 , w23020 , w23021 , w23022 , w23023 , w23024 , w23025 , w23026 , w23027 , w23028 , w23029 , w23030 , w23031 , w23032 , w23033 , w23034 , w23035 , w23036 , w23037 , w23038 , w23039 , w23040 , w23041 , w23042 , w23043 , w23044 , w23045 , w23046 , w23047 , w23048 , w23049 , w23050 , w23051 , w23052 , w23053 , w23054 , w23055 , w23056 , w23057 , w23058 , w23059 , w23060 , w23061 , w23062 , w23063 , w23064 , w23065 , w23066 , w23067 , w23068 , w23069 , w23070 , w23071 , w23072 , w23073 , w23074 , w23075 , w23076 , w23077 , w23078 , w23079 , w23080 , w23081 , w23082 , w23083 , w23084 , w23085 , w23086 , w23087 , w23088 , w23089 , w23090 , w23091 , w23092 , w23093 , w23094 , w23095 , w23096 , w23097 , w23098 , w23099 , w23100 , w23101 , w23102 , w23103 , w23104 , w23105 , w23106 , w23107 , w23108 , w23109 , w23110 , w23111 , w23112 , w23113 , w23114 , w23115 , w23116 , w23117 , w23118 , w23119 , w23120 , w23121 , w23122 , w23123 , w23124 , w23125 , w23126 , w23127 , w23128 , w23129 , w23130 , w23131 , w23132 , w23133 , w23134 , w23135 , w23136 , w23137 , w23138 , w23139 , w23140 , w23141 , w23142 , w23143 , w23144 , w23145 , w23146 , w23147 , w23148 , w23149 , w23150 , w23151 , w23152 , w23153 , w23154 , w23155 , w23156 , w23157 , w23158 , w23159 , w23160 , w23161 , w23162 , w23163 , w23164 , w23165 , w23166 , w23167 , w23168 , w23169 , w23170 , w23171 , w23172 , w23173 , w23174 , w23175 , w23176 , w23177 , w23178 , w23179 , w23180 , w23181 , w23182 , w23183 , w23184 , w23185 , w23186 , w23187 , w23188 , w23189 , w23190 , w23191 , w23192 , w23193 , w23194 , w23195 , w23196 , w23197 , w23198 , w23199 , w23200 , w23201 , w23202 , w23203 , w23204 , w23205 , w23206 , w23207 , w23208 , w23209 , w23210 , w23211 , w23212 , w23213 , w23214 , w23215 , w23216 , w23217 , w23218 , w23219 , w23220 , w23221 , w23222 , w23223 , w23224 , w23225 , w23226 , w23227 , w23228 , w23229 , w23230 , w23231 , w23232 , w23233 , w23234 , w23235 , w23236 , w23237 , w23238 , w23239 , w23240 , w23241 , w23242 , w23243 , w23244 , w23245 , w23246 , w23247 , w23248 , w23249 , w23250 , w23251 , w23252 , w23253 , w23254 , w23255 , w23256 , w23257 , w23258 , w23259 , w23260 , w23261 , w23262 , w23263 , w23264 , w23265 , w23266 , w23267 , w23268 , w23269 , w23270 , w23271 , w23272 , w23273 , w23274 , w23275 , w23276 , w23277 , w23278 , w23279 , w23280 , w23281 , w23282 , w23283 , w23284 , w23285 , w23286 , w23287 , w23288 , w23289 , w23290 , w23291 , w23292 , w23293 , w23294 , w23295 , w23296 , w23297 , w23298 , w23299 , w23300 , w23301 , w23302 , w23303 , w23304 , w23305 , w23306 , w23307 , w23308 , w23309 , w23310 , w23311 , w23312 , w23313 , w23314 , w23315 , w23316 , w23317 , w23318 , w23319 , w23320 , w23321 , w23322 , w23323 , w23324 , w23325 , w23326 , w23327 , w23328 , w23329 , w23330 , w23331 , w23332 , w23333 , w23334 , w23335 , w23336 , w23337 , w23338 , w23339 , w23340 , w23341 , w23342 , w23343 , w23344 , w23345 , w23346 , w23347 , w23348 , w23349 , w23350 , w23351 , w23352 , w23353 , w23354 , w23355 , w23356 , w23357 , w23358 , w23359 , w23360 , w23361 , w23362 , w23363 , w23364 , w23365 , w23366 , w23367 , w23368 , w23369 , w23370 , w23371 , w23372 , w23373 , w23374 , w23375 , w23376 , w23377 , w23378 , w23379 , w23380 , w23381 , w23382 , w23383 , w23384 , w23385 , w23386 , w23387 , w23388 , w23389 , w23390 , w23391 , w23392 , w23393 , w23394 , w23395 , w23396 , w23397 , w23398 , w23399 , w23400 , w23401 , w23402 , w23403 , w23404 , w23405 , w23406 , w23407 , w23408 , w23409 , w23410 , w23411 , w23412 , w23413 , w23414 , w23415 , w23416 , w23417 , w23418 , w23419 , w23420 , w23421 , w23422 , w23423 , w23424 , w23425 , w23426 , w23427 , w23428 , w23429 , w23430 , w23431 , w23432 , w23433 , w23434 , w23435 , w23436 , w23437 , w23438 , w23439 , w23440 , w23441 , w23442 , w23443 , w23444 , w23445 , w23446 , w23447 , w23448 , w23449 , w23450 , w23451 , w23452 , w23453 , w23454 , w23455 , w23456 , w23457 , w23458 , w23459 , w23460 , w23461 , w23462 , w23463 , w23464 , w23465 , w23466 , w23467 , w23468 , w23469 , w23470 , w23471 , w23472 , w23473 , w23474 , w23475 , w23476 , w23477 , w23478 , w23479 , w23480 , w23481 , w23482 , w23483 , w23484 , w23485 , w23486 , w23487 , w23488 , w23489 , w23490 , w23491 , w23492 , w23493 , w23494 , w23495 , w23496 , w23497 , w23498 , w23499 , w23500 , w23501 , w23502 , w23503 , w23504 , w23505 , w23506 , w23507 , w23508 , w23509 , w23510 , w23511 , w23512 , w23513 , w23514 , w23515 , w23516 , w23517 , w23518 , w23519 , w23520 , w23521 , w23522 , w23523 , w23524 , w23525 , w23526 , w23527 , w23528 , w23529 , w23530 , w23531 , w23532 , w23533 , w23534 , w23535 , w23536 , w23537 , w23538 , w23539 , w23540 , w23541 , w23542 , w23543 , w23544 , w23545 , w23546 , w23547 , w23548 , w23549 , w23550 , w23551 , w23552 , w23553 , w23554 , w23555 , w23556 , w23557 , w23558 , w23559 , w23560 , w23561 , w23562 , w23563 , w23564 , w23565 , w23566 , w23567 , w23568 , w23569 , w23570 , w23571 , w23572 , w23573 , w23574 , w23575 , w23576 , w23577 , w23578 , w23579 , w23580 , w23581 , w23582 , w23583 , w23584 , w23585 , w23586 , w23587 , w23588 , w23589 , w23590 , w23591 , w23592 , w23593 , w23594 , w23595 , w23596 , w23597 , w23598 , w23599 , w23600 , w23601 , w23602 , w23603 , w23604 , w23605 , w23606 , w23607 , w23608 , w23609 , w23610 , w23611 , w23612 , w23613 , w23614 , w23615 , w23616 , w23617 , w23618 , w23619 , w23620 , w23621 , w23622 , w23623 , w23624 , w23625 , w23626 , w23627 , w23628 , w23629 , w23630 , w23631 , w23632 , w23633 , w23634 , w23635 , w23636 , w23637 , w23638 , w23639 , w23640 , w23641 , w23642 , w23643 , w23644 , w23645 , w23646 , w23647 , w23648 , w23649 , w23650 , w23651 , w23652 , w23653 , w23654 , w23655 , w23656 , w23657 , w23658 , w23659 , w23660 , w23661 , w23662 , w23663 , w23664 , w23665 , w23666 , w23667 , w23668 , w23669 , w23670 , w23671 , w23672 , w23673 , w23674 , w23675 , w23676 , w23677 , w23678 , w23679 , w23680 , w23681 , w23682 , w23683 , w23684 , w23685 , w23686 , w23687 , w23688 , w23689 , w23690 , w23691 , w23692 , w23693 , w23694 , w23695 , w23696 , w23697 , w23698 , w23699 , w23700 , w23701 , w23702 , w23703 , w23704 , w23705 , w23706 , w23707 , w23708 , w23709 , w23710 , w23711 , w23712 , w23713 , w23714 , w23715 , w23716 , w23717 , w23718 , w23719 , w23720 , w23721 , w23722 , w23723 , w23724 , w23725 , w23726 , w23727 , w23728 , w23729 , w23730 , w23731 , w23732 , w23733 , w23734 , w23735 , w23736 , w23737 , w23738 , w23739 , w23740 , w23741 , w23742 , w23743 , w23744 , w23745 , w23746 , w23747 , w23748 , w23749 , w23750 , w23751 , w23752 , w23753 , w23754 , w23755 , w23756 , w23757 , w23758 , w23759 , w23760 , w23761 , w23762 , w23763 , w23764 , w23765 , w23766 , w23767 , w23768 , w23769 , w23770 , w23771 , w23772 , w23773 , w23774 , w23775 , w23776 , w23777 , w23778 , w23779 , w23780 , w23781 , w23782 , w23783 , w23784 , w23785 , w23786 , w23787 , w23788 , w23789 , w23790 , w23791 , w23792 , w23793 , w23794 , w23795 , w23796 , w23797 , w23798 , w23799 , w23800 , w23801 , w23802 , w23803 , w23804 , w23805 , w23806 , w23807 , w23808 , w23809 , w23810 , w23811 , w23812 , w23813 , w23814 , w23815 , w23816 , w23817 , w23818 , w23819 , w23820 , w23821 , w23822 , w23823 , w23824 , w23825 , w23826 , w23827 , w23828 , w23829 , w23830 , w23831 , w23832 , w23833 , w23834 , w23835 , w23836 , w23837 , w23838 , w23839 , w23840 , w23841 , w23842 , w23843 , w23844 , w23845 , w23846 , w23847 , w23848 , w23849 , w23850 , w23851 , w23852 , w23853 , w23854 , w23855 , w23856 , w23857 , w23858 , w23859 , w23860 , w23861 , w23862 , w23863 , w23864 , w23865 , w23866 , w23867 , w23868 , w23869 , w23870 , w23871 , w23872 , w23873 , w23874 , w23875 , w23876 , w23877 , w23878 , w23879 , w23880 , w23881 , w23882 , w23883 , w23884 , w23885 , w23886 , w23887 , w23888 , w23889 , w23890 , w23891 , w23892 , w23893 , w23894 , w23895 , w23896 , w23897 , w23898 , w23899 , w23900 , w23901 , w23902 , w23903 , w23904 , w23905 , w23906 , w23907 , w23908 , w23909 , w23910 , w23911 , w23912 , w23913 , w23914 , w23915 , w23916 , w23917 , w23918 , w23919 , w23920 , w23921 , w23922 , w23923 , w23924 , w23925 , w23926 , w23927 , w23928 , w23929 , w23930 , w23931 , w23932 , w23933 , w23934 , w23935 , w23936 , w23937 , w23938 , w23939 , w23940 , w23941 , w23942 , w23943 , w23944 , w23945 , w23946 , w23947 , w23948 , w23949 , w23950 , w23951 , w23952 , w23953 , w23954 , w23955 , w23956 , w23957 , w23958 , w23959 , w23960 , w23961 , w23962 , w23963 , w23964 , w23965 , w23966 , w23967 , w23968 , w23969 , w23970 , w23971 , w23972 , w23973 , w23974 , w23975 , w23976 , w23977 , w23978 , w23979 , w23980 , w23981 , w23982 , w23983 , w23984 , w23985 , w23986 , w23987 , w23988 , w23989 , w23990 , w23991 , w23992 , w23993 , w23994 , w23995 , w23996 , w23997 , w23998 , w23999 , w24000 , w24001 , w24002 , w24003 , w24004 , w24005 , w24006 , w24007 , w24008 , w24009 , w24010 , w24011 , w24012 , w24013 , w24014 , w24015 , w24016 , w24017 , w24018 , w24019 , w24020 , w24021 , w24022 , w24023 , w24024 , w24025 , w24026 , w24027 , w24028 , w24029 , w24030 , w24031 , w24032 , w24033 , w24034 , w24035 , w24036 , w24037 , w24038 , w24039 , w24040 , w24041 , w24042 , w24043 , w24044 , w24045 , w24046 , w24047 , w24048 , w24049 , w24050 , w24051 , w24052 , w24053 , w24054 , w24055 , w24056 , w24057 , w24058 , w24059 , w24060 , w24061 , w24062 , w24063 , w24064 , w24065 , w24066 , w24067 , w24068 , w24069 , w24070 , w24071 , w24072 , w24073 , w24074 , w24075 , w24076 , w24077 , w24078 , w24079 , w24080 , w24081 , w24082 , w24083 , w24084 , w24085 , w24086 , w24087 , w24088 , w24089 , w24090 , w24091 , w24092 , w24093 , w24094 , w24095 , w24096 , w24097 , w24098 , w24099 , w24100 , w24101 , w24102 , w24103 , w24104 , w24105 , w24106 , w24107 , w24108 , w24109 , w24110 , w24111 , w24112 , w24113 , w24114 , w24115 , w24116 , w24117 , w24118 , w24119 , w24120 , w24121 , w24122 , w24123 , w24124 , w24125 , w24126 , w24127 , w24128 , w24129 , w24130 , w24131 , w24132 , w24133 , w24134 , w24135 , w24136 , w24137 , w24138 , w24139 , w24140 , w24141 , w24142 , w24143 , w24144 , w24145 , w24146 , w24147 , w24148 , w24149 , w24150 , w24151 , w24152 , w24153 , w24154 , w24155 , w24156 , w24157 , w24158 , w24159 , w24160 , w24161 , w24162 , w24163 , w24164 , w24165 , w24166 , w24167 , w24168 , w24169 , w24170 , w24171 , w24172 , w24173 , w24174 , w24175 , w24176 , w24177 , w24178 , w24179 , w24180 , w24181 , w24182 , w24183 , w24184 , w24185 , w24186 , w24187 , w24188 , w24189 , w24190 , w24191 , w24192 , w24193 , w24194 , w24195 , w24196 , w24197 , w24198 , w24199 , w24200 , w24201 , w24202 , w24203 , w24204 , w24205 , w24206 , w24207 , w24208 , w24209 , w24210 , w24211 , w24212 , w24213 , w24214 , w24215 , w24216 , w24217 , w24218 , w24219 , w24220 , w24221 , w24222 , w24223 , w24224 , w24225 , w24226 , w24227 , w24228 , w24229 , w24230 , w24231 , w24232 , w24233 , w24234 , w24235 , w24236 , w24237 , w24238 , w24239 , w24240 , w24241 , w24242 , w24243 , w24244 , w24245 , w24246 , w24247 , w24248 , w24249 , w24250 , w24251 , w24252 , w24253 , w24254 , w24255 , w24256 , w24257 , w24258 , w24259 , w24260 , w24261 , w24262 , w24263 , w24264 , w24265 , w24266 , w24267 , w24268 , w24269 , w24270 , w24271 , w24272 , w24273 , w24274 , w24275 , w24276 , w24277 , w24278 , w24279 , w24280 , w24281 , w24282 , w24283 , w24284 , w24285 , w24286 , w24287 , w24288 , w24289 , w24290 , w24291 , w24292 , w24293 , w24294 , w24295 , w24296 , w24297 , w24298 , w24299 , w24300 , w24301 , w24302 , w24303 , w24304 , w24305 , w24306 , w24307 , w24308 , w24309 , w24310 , w24311 , w24312 , w24313 , w24314 , w24315 , w24316 , w24317 , w24318 , w24319 , w24320 , w24321 , w24322 , w24323 , w24324 , w24325 , w24326 , w24327 , w24328 , w24329 , w24330 , w24331 , w24332 , w24333 , w24334 , w24335 , w24336 , w24337 , w24338 , w24339 , w24340 , w24341 , w24342 , w24343 , w24344 , w24345 , w24346 , w24347 , w24348 , w24349 , w24350 , w24351 , w24352 , w24353 , w24354 , w24355 , w24356 , w24357 , w24358 , w24359 , w24360 , w24361 , w24362 , w24363 , w24364 , w24365 , w24366 , w24367 , w24368 , w24369 , w24370 , w24371 , w24372 , w24373 , w24374 , w24375 , w24376 , w24377 , w24378 , w24379 , w24380 , w24381 , w24382 , w24383 , w24384 , w24385 , w24386 , w24387 , w24388 , w24389 , w24390 , w24391 , w24392 , w24393 , w24394 , w24395 , w24396 , w24397 , w24398 , w24399 , w24400 , w24401 , w24402 , w24403 , w24404 , w24405 , w24406 , w24407 , w24408 , w24409 , w24410 , w24411 , w24412 , w24413 , w24414 , w24415 , w24416 , w24417 , w24418 , w24419 , w24420 , w24421 , w24422 , w24423 , w24424 , w24425 , w24426 , w24427 , w24428 , w24429 , w24430 , w24431 , w24432 , w24433 , w24434 , w24435 , w24436 , w24437 , w24438 , w24439 , w24440 , w24441 , w24442 , w24443 , w24444 , w24445 , w24446 , w24447 , w24448 , w24449 , w24450 , w24451 , w24452 , w24453 , w24454 , w24455 , w24456 , w24457 , w24458 , w24459 , w24460 , w24461 , w24462 , w24463 , w24464 , w24465 , w24466 , w24467 , w24468 , w24469 , w24470 , w24471 , w24472 , w24473 , w24474 , w24475 , w24476 , w24477 , w24478 , w24479 , w24480 , w24481 , w24482 , w24483 , w24484 , w24485 , w24486 , w24487 , w24488 , w24489 , w24490 , w24491 , w24492 , w24493 , w24494 , w24495 , w24496 , w24497 , w24498 , w24499 , w24500 , w24501 , w24502 , w24503 , w24504 , w24505 , w24506 , w24507 , w24508 , w24509 , w24510 , w24511 , w24512 , w24513 , w24514 , w24515 , w24516 , w24517 , w24518 , w24519 , w24520 , w24521 , w24522 , w24523 , w24524 , w24525 , w24526 , w24527 , w24528 , w24529 , w24530 , w24531 , w24532 , w24533 , w24534 , w24535 , w24536 , w24537 , w24538 , w24539 , w24540 , w24541 , w24542 , w24543 , w24544 , w24545 , w24546 , w24547 , w24548 , w24549 , w24550 , w24551 , w24552 , w24553 , w24554 , w24555 , w24556 , w24557 , w24558 , w24559 , w24560 , w24561 , w24562 , w24563 , w24564 , w24565 , w24566 , w24567 , w24568 , w24569 , w24570 , w24571 , w24572 , w24573 , w24574 , w24575 , w24576 , w24577 , w24578 , w24579 , w24580 , w24581 , w24582 , w24583 , w24584 , w24585 , w24586 , w24587 , w24588 , w24589 , w24590 , w24591 , w24592 , w24593 , w24594 , w24595 , w24596 , w24597 , w24598 , w24599 , w24600 , w24601 , w24602 , w24603 , w24604 , w24605 , w24606 , w24607 , w24608 , w24609 , w24610 , w24611 , w24612 , w24613 , w24614 , w24615 , w24616 , w24617 , w24618 , w24619 , w24620 , w24621 , w24622 , w24623 , w24624 , w24625 , w24626 , w24627 , w24628 , w24629 , w24630 , w24631 , w24632 , w24633 , w24634 , w24635 , w24636 , w24637 , w24638 , w24639 , w24640 , w24641 , w24642 , w24643 , w24644 , w24645 , w24646 , w24647 , w24648 , w24649 , w24650 , w24651 , w24652 , w24653 , w24654 , w24655 , w24656 , w24657 , w24658 , w24659 , w24660 , w24661 , w24662 , w24663 , w24664 , w24665 , w24666 , w24667 , w24668 , w24669 , w24670 , w24671 , w24672 , w24673 , w24674 , w24675 , w24676 , w24677 , w24678 , w24679 , w24680 , w24681 , w24682 , w24683 , w24684 , w24685 , w24686 , w24687 , w24688 , w24689 , w24690 , w24691 , w24692 , w24693 , w24694 , w24695 , w24696 , w24697 , w24698 , w24699 , w24700 , w24701 , w24702 , w24703 , w24704 , w24705 , w24706 , w24707 , w24708 , w24709 , w24710 , w24711 , w24712 , w24713 , w24714 , w24715 , w24716 , w24717 , w24718 , w24719 , w24720 , w24721 , w24722 , w24723 , w24724 , w24725 , w24726 , w24727 , w24728 , w24729 , w24730 , w24731 , w24732 , w24733 , w24734 , w24735 , w24736 , w24737 , w24738 , w24739 , w24740 , w24741 , w24742 , w24743 , w24744 , w24745 , w24746 , w24747 , w24748 , w24749 , w24750 , w24751 , w24752 , w24753 , w24754 , w24755 , w24756 , w24757 , w24758 , w24759 , w24760 , w24761 , w24762 , w24763 , w24764 , w24765 , w24766 , w24767 , w24768 , w24769 , w24770 , w24771 , w24772 , w24773 , w24774 , w24775 , w24776 , w24777 , w24778 , w24779 , w24780 , w24781 , w24782 , w24783 , w24784 , w24785 , w24786 , w24787 , w24788 , w24789 , w24790 , w24791 , w24792 , w24793 , w24794 , w24795 , w24796 , w24797 , w24798 , w24799 , w24800 , w24801 , w24802 , w24803 , w24804 , w24805 , w24806 , w24807 , w24808 , w24809 , w24810 , w24811 , w24812 , w24813 , w24814 , w24815 , w24816 , w24817 , w24818 , w24819 , w24820 , w24821 , w24822 , w24823 , w24824 , w24825 , w24826 , w24827 , w24828 , w24829 , w24830 , w24831 , w24832 , w24833 , w24834 , w24835 , w24836 , w24837 , w24838 , w24839 , w24840 , w24841 , w24842 , w24843 , w24844 , w24845 , w24846 , w24847 , w24848 , w24849 , w24850 , w24851 , w24852 , w24853 , w24854 , w24855 , w24856 , w24857 , w24858 , w24859 , w24860 , w24861 , w24862 , w24863 , w24864 , w24865 , w24866 , w24867 , w24868 , w24869 , w24870 , w24871 , w24872 , w24873 , w24874 , w24875 , w24876 , w24877 , w24878 , w24879 , w24880 , w24881 , w24882 , w24883 , w24884 , w24885 , w24886 , w24887 , w24888 , w24889 , w24890 , w24891 , w24892 , w24893 , w24894 , w24895 , w24896 , w24897 , w24898 , w24899 , w24900 , w24901 , w24902 , w24903 , w24904 , w24905 , w24906 , w24907 , w24908 , w24909 , w24910 , w24911 , w24912 , w24913 , w24914 , w24915 , w24916 , w24917 , w24918 , w24919 , w24920 , w24921 , w24922 , w24923 , w24924 , w24925 , w24926 , w24927 , w24928 , w24929 , w24930 , w24931 , w24932 , w24933 , w24934 , w24935 , w24936 , w24937 , w24938 , w24939 , w24940 , w24941 , w24942 , w24943 , w24944 , w24945 , w24946 , w24947 , w24948 , w24949 , w24950 , w24951 , w24952 , w24953 , w24954 , w24955 , w24956 , w24957 , w24958 , w24959 , w24960 , w24961 , w24962 , w24963 , w24964 , w24965 , w24966 , w24967 , w24968 , w24969 , w24970 , w24971 , w24972 , w24973 , w24974 , w24975 , w24976 , w24977 , w24978 , w24979 , w24980 , w24981 , w24982 , w24983 , w24984 , w24985 , w24986 , w24987 , w24988 , w24989 , w24990 , w24991 , w24992 , w24993 , w24994 , w24995 , w24996 , w24997 , w24998 , w24999 , w25000 , w25001 , w25002 , w25003 , w25004 , w25005 , w25006 , w25007 , w25008 , w25009 , w25010 , w25011 , w25012 , w25013 , w25014 , w25015 , w25016 , w25017 , w25018 , w25019 , w25020 , w25021 , w25022 , w25023 , w25024 , w25025 , w25026 , w25027 , w25028 , w25029 , w25030 , w25031 , w25032 , w25033 , w25034 , w25035 , w25036 , w25037 , w25038 , w25039 , w25040 , w25041 , w25042 , w25043 , w25044 , w25045 , w25046 , w25047 , w25048 , w25049 , w25050 , w25051 , w25052 , w25053 , w25054 , w25055 , w25056 , w25057 , w25058 , w25059 , w25060 , w25061 , w25062 , w25063 , w25064 , w25065 , w25066 , w25067 , w25068 , w25069 , w25070 , w25071 , w25072 , w25073 , w25074 , w25075 , w25076 , w25077 , w25078 , w25079 , w25080 , w25081 , w25082 , w25083 , w25084 , w25085 , w25086 , w25087 , w25088 , w25089 , w25090 , w25091 , w25092 , w25093 , w25094 , w25095 , w25096 , w25097 , w25098 , w25099 , w25100 , w25101 , w25102 , w25103 , w25104 , w25105 , w25106 , w25107 , w25108 , w25109 , w25110 , w25111 , w25112 , w25113 , w25114 , w25115 , w25116 , w25117 , w25118 , w25119 , w25120 , w25121 , w25122 , w25123 , w25124 , w25125 , w25126 , w25127 , w25128 , w25129 , w25130 , w25131 , w25132 , w25133 , w25134 , w25135 , w25136 , w25137 , w25138 , w25139 , w25140 , w25141 , w25142 , w25143 , w25144 , w25145 , w25146 , w25147 , w25148 , w25149 , w25150 , w25151 , w25152 , w25153 , w25154 , w25155 , w25156 , w25157 , w25158 , w25159 , w25160 , w25161 , w25162 , w25163 , w25164 , w25165 , w25166 , w25167 , w25168 , w25169 , w25170 , w25171 , w25172 , w25173 , w25174 , w25175 , w25176 , w25177 , w25178 , w25179 , w25180 , w25181 , w25182 , w25183 , w25184 , w25185 , w25186 , w25187 , w25188 , w25189 , w25190 , w25191 , w25192 , w25193 , w25194 , w25195 , w25196 , w25197 , w25198 , w25199 , w25200 , w25201 , w25202 , w25203 , w25204 , w25205 , w25206 , w25207 , w25208 , w25209 , w25210 , w25211 , w25212 , w25213 , w25214 , w25215 , w25216 , w25217 , w25218 , w25219 , w25220 , w25221 , w25222 , w25223 , w25224 , w25225 , w25226 , w25227 , w25228 , w25229 , w25230 , w25231 , w25232 , w25233 , w25234 , w25235 , w25236 , w25237 , w25238 , w25239 , w25240 , w25241 , w25242 , w25243 , w25244 , w25245 , w25246 , w25247 , w25248 , w25249 , w25250 , w25251 , w25252 , w25253 , w25254 , w25255 , w25256 , w25257 , w25258 , w25259 , w25260 , w25261 , w25262 , w25263 , w25264 , w25265 , w25266 , w25267 , w25268 , w25269 , w25270 , w25271 , w25272 , w25273 , w25274 , w25275 , w25276 , w25277 , w25278 , w25279 , w25280 , w25281 , w25282 , w25283 , w25284 , w25285 , w25286 , w25287 , w25288 , w25289 , w25290 , w25291 , w25292 , w25293 , w25294 , w25295 , w25296 , w25297 , w25298 , w25299 , w25300 , w25301 , w25302 , w25303 , w25304 , w25305 , w25306 , w25307 , w25308 , w25309 , w25310 , w25311 , w25312 , w25313 , w25314 , w25315 , w25316 , w25317 , w25318 , w25319 , w25320 , w25321 , w25322 , w25323 , w25324 , w25325 , w25326 , w25327 , w25328 , w25329 , w25330 , w25331 , w25332 , w25333 , w25334 , w25335 , w25336 , w25337 , w25338 , w25339 , w25340 , w25341 , w25342 , w25343 , w25344 , w25345 , w25346 , w25347 , w25348 , w25349 , w25350 , w25351 , w25352 , w25353 , w25354 , w25355 , w25356 , w25357 , w25358 , w25359 , w25360 , w25361 , w25362 , w25363 , w25364 , w25365 , w25366 , w25367 , w25368 , w25369 , w25370 , w25371 , w25372 , w25373 , w25374 , w25375 , w25376 , w25377 , w25378 , w25379 , w25380 , w25381 , w25382 , w25383 , w25384 , w25385 , w25386 , w25387 , w25388 , w25389 , w25390 , w25391 , w25392 , w25393 , w25394 , w25395 , w25396 , w25397 , w25398 , w25399 , w25400 , w25401 , w25402 , w25403 , w25404 , w25405 , w25406 , w25407 , w25408 , w25409 , w25410 , w25411 , w25412 , w25413 , w25414 , w25415 , w25416 , w25417 , w25418 , w25419 , w25420 , w25421 , w25422 , w25423 , w25424 , w25425 , w25426 , w25427 , w25428 , w25429 , w25430 , w25431 , w25432 , w25433 , w25434 , w25435 , w25436 , w25437 , w25438 , w25439 , w25440 , w25441 , w25442 , w25443 , w25444 , w25445 , w25446 , w25447 , w25448 , w25449 , w25450 , w25451 , w25452 , w25453 , w25454 , w25455 , w25456 , w25457 , w25458 , w25459 , w25460 , w25461 , w25462 , w25463 , w25464 , w25465 , w25466 , w25467 , w25468 , w25469 , w25470 , w25471 , w25472 , w25473 , w25474 , w25475 , w25476 , w25477 , w25478 , w25479 , w25480 , w25481 , w25482 , w25483 , w25484 , w25485 , w25486 , w25487 , w25488 , w25489 , w25490 , w25491 , w25492 , w25493 , w25494 , w25495 , w25496 , w25497 , w25498 , w25499 , w25500 , w25501 , w25502 , w25503 , w25504 , w25505 , w25506 , w25507 , w25508 , w25509 , w25510 , w25511 , w25512 , w25513 , w25514 , w25515 , w25516 , w25517 , w25518 , w25519 , w25520 , w25521 , w25522 , w25523 , w25524 , w25525 , w25526 , w25527 , w25528 , w25529 , w25530 , w25531 , w25532 , w25533 , w25534 , w25535 , w25536 , w25537 , w25538 , w25539 , w25540 , w25541 , w25542 , w25543 , w25544 , w25545 , w25546 , w25547 , w25548 , w25549 , w25550 , w25551 , w25552 , w25553 , w25554 , w25555 , w25556 , w25557 , w25558 , w25559 , w25560 , w25561 , w25562 , w25563 , w25564 , w25565 , w25566 , w25567 , w25568 , w25569 , w25570 , w25571 , w25572 , w25573 , w25574 , w25575 , w25576 , w25577 , w25578 , w25579 , w25580 , w25581 , w25582 , w25583 , w25584 , w25585 , w25586 , w25587 , w25588 , w25589 , w25590 , w25591 , w25592 , w25593 , w25594 , w25595 , w25596 , w25597 , w25598 , w25599 , w25600 , w25601 , w25602 , w25603 , w25604 , w25605 , w25606 , w25607 , w25608 , w25609 , w25610 , w25611 , w25612 , w25613 , w25614 , w25615 , w25616 , w25617 , w25618 , w25619 , w25620 , w25621 , w25622 , w25623 , w25624 , w25625 , w25626 , w25627 , w25628 , w25629 , w25630 , w25631 , w25632 , w25633 , w25634 , w25635 , w25636 , w25637 , w25638 , w25639 , w25640 , w25641 , w25642 , w25643 , w25644 , w25645 , w25646 , w25647 , w25648 , w25649 , w25650 , w25651 , w25652 , w25653 , w25654 , w25655 , w25656 , w25657 , w25658 , w25659 , w25660 , w25661 , w25662 , w25663 , w25664 , w25665 , w25666 , w25667 , w25668 , w25669 , w25670 , w25671 , w25672 , w25673 , w25674 , w25675 , w25676 , w25677 , w25678 , w25679 , w25680 , w25681 , w25682 , w25683 , w25684 , w25685 , w25686 , w25687 , w25688 , w25689 , w25690 , w25691 , w25692 , w25693 , w25694 , w25695 , w25696 , w25697 , w25698 , w25699 , w25700 , w25701 , w25702 , w25703 , w25704 , w25705 , w25706 , w25707 , w25708 , w25709 , w25710 , w25711 , w25712 , w25713 , w25714 , w25715 , w25716 , w25717 , w25718 , w25719 , w25720 , w25721 , w25722 , w25723 , w25724 , w25725 , w25726 , w25727 , w25728 , w25729 , w25730 , w25731 , w25732 , w25733 , w25734 , w25735 , w25736 , w25737 , w25738 , w25739 , w25740 , w25741 , w25742 , w25743 , w25744 , w25745 , w25746 , w25747 , w25748 , w25749 , w25750 , w25751 , w25752 , w25753 , w25754 , w25755 , w25756 , w25757 , w25758 , w25759 , w25760 , w25761 , w25762 , w25763 , w25764 , w25765 , w25766 , w25767 , w25768 , w25769 , w25770 , w25771 , w25772 , w25773 , w25774 , w25775 , w25776 , w25777 , w25778 , w25779 , w25780 , w25781 , w25782 , w25783 , w25784 , w25785 , w25786 , w25787 , w25788 , w25789 , w25790 , w25791 , w25792 , w25793 , w25794 , w25795 , w25796 , w25797 , w25798 , w25799 , w25800 , w25801 , w25802 , w25803 , w25804 , w25805 , w25806 , w25807 , w25808 , w25809 , w25810 , w25811 , w25812 , w25813 , w25814 , w25815 , w25816 , w25817 , w25818 , w25819 , w25820 , w25821 , w25822 , w25823 , w25824 , w25825 , w25826 , w25827 , w25828 , w25829 , w25830 , w25831 , w25832 , w25833 , w25834 , w25835 , w25836 , w25837 , w25838 , w25839 , w25840 , w25841 , w25842 , w25843 , w25844 , w25845 , w25846 , w25847 , w25848 , w25849 , w25850 , w25851 , w25852 , w25853 , w25854 , w25855 , w25856 , w25857 , w25858 , w25859 , w25860 , w25861 , w25862 , w25863 , w25864 , w25865 , w25866 , w25867 , w25868 , w25869 , w25870 , w25871 , w25872 , w25873 , w25874 , w25875 , w25876 , w25877 , w25878 , w25879 , w25880 , w25881 , w25882 , w25883 , w25884 , w25885 , w25886 , w25887 , w25888 , w25889 , w25890 , w25891 , w25892 , w25893 , w25894 , w25895 , w25896 , w25897 , w25898 , w25899 , w25900 , w25901 , w25902 , w25903 , w25904 , w25905 , w25906 , w25907 , w25908 , w25909 , w25910 , w25911 , w25912 , w25913 , w25914 , w25915 , w25916 , w25917 , w25918 , w25919 , w25920 , w25921 , w25922 , w25923 , w25924 , w25925 , w25926 , w25927 , w25928 , w25929 , w25930 , w25931 , w25932 , w25933 , w25934 , w25935 , w25936 , w25937 , w25938 , w25939 , w25940 , w25941 , w25942 , w25943 , w25944 , w25945 , w25946 , w25947 , w25948 , w25949 , w25950 , w25951 , w25952 , w25953 , w25954 , w25955 , w25956 , w25957 , w25958 , w25959 , w25960 , w25961 , w25962 , w25963 , w25964 , w25965 , w25966 , w25967 , w25968 , w25969 , w25970 , w25971 , w25972 , w25973 , w25974 , w25975 , w25976 , w25977 , w25978 , w25979 , w25980 , w25981 , w25982 , w25983 , w25984 , w25985 , w25986 , w25987 , w25988 , w25989 , w25990 , w25991 , w25992 , w25993 , w25994 , w25995 , w25996 , w25997 , w25998 , w25999 , w26000 , w26001 , w26002 , w26003 , w26004 , w26005 , w26006 , w26007 , w26008 , w26009 , w26010 , w26011 , w26012 , w26013 , w26014 , w26015 , w26016 , w26017 , w26018 , w26019 , w26020 , w26021 , w26022 , w26023 , w26024 , w26025 , w26026 , w26027 , w26028 , w26029 , w26030 , w26031 , w26032 , w26033 , w26034 , w26035 , w26036 , w26037 , w26038 , w26039 , w26040 , w26041 , w26042 , w26043 , w26044 , w26045 , w26046 , w26047 , w26048 , w26049 , w26050 , w26051 , w26052 , w26053 , w26054 , w26055 , w26056 , w26057 , w26058 , w26059 , w26060 , w26061 , w26062 , w26063 , w26064 , w26065 , w26066 , w26067 , w26068 , w26069 , w26070 , w26071 , w26072 , w26073 , w26074 , w26075 , w26076 , w26077 , w26078 , w26079 , w26080 , w26081 , w26082 , w26083 , w26084 , w26085 , w26086 , w26087 , w26088 , w26089 , w26090 , w26091 , w26092 , w26093 , w26094 , w26095 , w26096 , w26097 , w26098 , w26099 , w26100 , w26101 , w26102 , w26103 , w26104 , w26105 , w26106 , w26107 , w26108 , w26109 , w26110 , w26111 , w26112 , w26113 , w26114 , w26115 , w26116 , w26117 , w26118 , w26119 , w26120 , w26121 , w26122 , w26123 , w26124 , w26125 , w26126 , w26127 , w26128 , w26129 , w26130 , w26131 , w26132 , w26133 , w26134 , w26135 , w26136 , w26137 , w26138 , w26139 , w26140 , w26141 , w26142 , w26143 , w26144 , w26145 , w26146 , w26147 , w26148 , w26149 , w26150 , w26151 , w26152 , w26153 , w26154 , w26155 , w26156 , w26157 , w26158 , w26159 , w26160 , w26161 , w26162 , w26163 , w26164 , w26165 , w26166 , w26167 , w26168 , w26169 , w26170 , w26171 , w26172 , w26173 , w26174 , w26175 , w26176 , w26177 , w26178 , w26179 , w26180 , w26181 , w26182 , w26183 , w26184 , w26185 , w26186 , w26187 , w26188 , w26189 , w26190 , w26191 , w26192 , w26193 , w26194 , w26195 , w26196 , w26197 , w26198 , w26199 , w26200 , w26201 , w26202 , w26203 , w26204 , w26205 , w26206 , w26207 , w26208 , w26209 , w26210 , w26211 , w26212 , w26213 , w26214 , w26215 , w26216 , w26217 , w26218 , w26219 , w26220 , w26221 , w26222 , w26223 , w26224 , w26225 , w26226 , w26227 , w26228 , w26229 , w26230 , w26231 , w26232 , w26233 , w26234 , w26235 , w26236 , w26237 , w26238 , w26239 , w26240 , w26241 , w26242 , w26243 , w26244 , w26245 , w26246 , w26247 , w26248 , w26249 , w26250 , w26251 , w26252 , w26253 , w26254 , w26255 , w26256 , w26257 , w26258 , w26259 , w26260 , w26261 , w26262 , w26263 , w26264 , w26265 , w26266 , w26267 , w26268 , w26269 , w26270 , w26271 , w26272 , w26273 , w26274 , w26275 , w26276 , w26277 , w26278 , w26279 , w26280 , w26281 , w26282 , w26283 , w26284 , w26285 , w26286 , w26287 , w26288 , w26289 , w26290 , w26291 , w26292 , w26293 , w26294 , w26295 , w26296 , w26297 , w26298 , w26299 , w26300 , w26301 , w26302 , w26303 , w26304 , w26305 , w26306 , w26307 , w26308 , w26309 , w26310 , w26311 , w26312 , w26313 , w26314 , w26315 , w26316 , w26317 , w26318 , w26319 , w26320 , w26321 , w26322 , w26323 , w26324 , w26325 , w26326 , w26327 , w26328 , w26329 , w26330 , w26331 , w26332 , w26333 , w26334 , w26335 , w26336 , w26337 , w26338 , w26339 , w26340 , w26341 , w26342 , w26343 , w26344 , w26345 , w26346 , w26347 , w26348 , w26349 , w26350 , w26351 , w26352 , w26353 , w26354 , w26355 , w26356 , w26357 , w26358 , w26359 , w26360 , w26361 , w26362 , w26363 , w26364 , w26365 , w26366 , w26367 , w26368 , w26369 , w26370 , w26371 , w26372 , w26373 , w26374 , w26375 , w26376 , w26377 , w26378 , w26379 , w26380 , w26381 , w26382 , w26383 , w26384 , w26385 , w26386 , w26387 , w26388 , w26389 , w26390 , w26391 , w26392 , w26393 , w26394 , w26395 , w26396 , w26397 , w26398 , w26399 , w26400 , w26401 , w26402 , w26403 , w26404 , w26405 , w26406 , w26407 , w26408 , w26409 , w26410 , w26411 , w26412 , w26413 , w26414 , w26415 , w26416 , w26417 , w26418 , w26419 , w26420 , w26421 , w26422 , w26423 , w26424 , w26425 , w26426 , w26427 , w26428 , w26429 , w26430 , w26431 , w26432 , w26433 , w26434 , w26435 , w26436 , w26437 , w26438 , w26439 , w26440 , w26441 , w26442 , w26443 , w26444 , w26445 , w26446 , w26447 , w26448 , w26449 , w26450 , w26451 , w26452 , w26453 , w26454 , w26455 , w26456 , w26457 , w26458 , w26459 , w26460 , w26461 , w26462 , w26463 , w26464 , w26465 , w26466 , w26467 , w26468 , w26469 , w26470 , w26471 , w26472 , w26473 , w26474 , w26475 , w26476 , w26477 , w26478 , w26479 , w26480 , w26481 , w26482 , w26483 , w26484 , w26485 , w26486 , w26487 , w26488 , w26489 , w26490 , w26491 , w26492 , w26493 , w26494 , w26495 , w26496 , w26497 , w26498 , w26499 , w26500 , w26501 , w26502 , w26503 , w26504 , w26505 , w26506 , w26507 , w26508 , w26509 , w26510 , w26511 , w26512 , w26513 , w26514 , w26515 , w26516 , w26517 , w26518 , w26519 , w26520 , w26521 , w26522 , w26523 , w26524 , w26525 , w26526 , w26527 , w26528 , w26529 , w26530 , w26531 , w26532 , w26533 , w26534 , w26535 , w26536 , w26537 , w26538 , w26539 , w26540 , w26541 , w26542 , w26543 , w26544 , w26545 , w26546 , w26547 , w26548 , w26549 , w26550 , w26551 , w26552 , w26553 , w26554 , w26555 , w26556 , w26557 , w26558 , w26559 , w26560 , w26561 , w26562 , w26563 , w26564 , w26565 , w26566 , w26567 , w26568 , w26569 , w26570 , w26571 , w26572 , w26573 , w26574 , w26575 , w26576 , w26577 , w26578 , w26579 , w26580 , w26581 , w26582 , w26583 , w26584 , w26585 , w26586 , w26587 , w26588 , w26589 , w26590 , w26591 , w26592 , w26593 , w26594 , w26595 , w26596 , w26597 , w26598 , w26599 , w26600 , w26601 , w26602 , w26603 , w26604 , w26605 , w26606 , w26607 , w26608 , w26609 , w26610 , w26611 , w26612 , w26613 , w26614 , w26615 , w26616 , w26617 , w26618 , w26619 , w26620 , w26621 , w26622 , w26623 , w26624 , w26625 , w26626 , w26627 , w26628 , w26629 , w26630 , w26631 , w26632 , w26633 , w26634 , w26635 , w26636 , w26637 , w26638 , w26639 , w26640 , w26641 , w26642 , w26643 , w26644 , w26645 , w26646 , w26647 , w26648 , w26649 , w26650 , w26651 , w26652 , w26653 , w26654 , w26655 , w26656 , w26657 , w26658 , w26659 , w26660 , w26661 , w26662 , w26663 , w26664 , w26665 , w26666 , w26667 , w26668 , w26669 , w26670 , w26671 , w26672 , w26673 , w26674 , w26675 , w26676 , w26677 , w26678 , w26679 , w26680 , w26681 , w26682 , w26683 , w26684 , w26685 , w26686 , w26687 , w26688 , w26689 , w26690 , w26691 , w26692 , w26693 , w26694 , w26695 , w26696 , w26697 , w26698 , w26699 , w26700 , w26701 , w26702 , w26703 , w26704 , w26705 , w26706 , w26707 , w26708 , w26709 , w26710 , w26711 , w26712 , w26713 , w26714 , w26715 , w26716 , w26717 , w26718 , w26719 , w26720 , w26721 , w26722 , w26723 , w26724 , w26725 , w26726 , w26727 , w26728 , w26729 , w26730 , w26731 , w26732 , w26733 , w26734 , w26735 , w26736 , w26737 , w26738 , w26739 , w26740 , w26741 , w26742 , w26743 , w26744 , w26745 , w26746 , w26747 , w26748 , w26749 , w26750 , w26751 , w26752 , w26753 , w26754 , w26755 , w26756 , w26757 , w26758 , w26759 , w26760 , w26761 , w26762 , w26763 , w26764 , w26765 , w26766 , w26767 , w26768 , w26769 , w26770 , w26771 , w26772 , w26773 , w26774 , w26775 , w26776 , w26777 , w26778 , w26779 , w26780 , w26781 , w26782 , w26783 , w26784 , w26785 , w26786 , w26787 , w26788 , w26789 , w26790 , w26791 , w26792 , w26793 , w26794 , w26795 , w26796 , w26797 , w26798 , w26799 , w26800 , w26801 , w26802 , w26803 , w26804 , w26805 , w26806 , w26807 , w26808 , w26809 , w26810 , w26811 , w26812 , w26813 , w26814 , w26815 , w26816 , w26817 , w26818 , w26819 , w26820 , w26821 , w26822 , w26823 , w26824 , w26825 , w26826 , w26827 , w26828 , w26829 , w26830 , w26831 , w26832 , w26833 , w26834 , w26835 , w26836 , w26837 , w26838 , w26839 , w26840 , w26841 , w26842 , w26843 , w26844 , w26845 , w26846 , w26847 , w26848 , w26849 , w26850 , w26851 , w26852 , w26853 , w26854 , w26855 , w26856 , w26857 , w26858 , w26859 , w26860 , w26861 , w26862 , w26863 , w26864 , w26865 , w26866 , w26867 , w26868 , w26869 , w26870 , w26871 , w26872 , w26873 , w26874 , w26875 , w26876 , w26877 , w26878 , w26879 , w26880 , w26881 , w26882 , w26883 , w26884 , w26885 , w26886 , w26887 , w26888 , w26889 , w26890 , w26891 , w26892 , w26893 , w26894 , w26895 , w26896 , w26897 , w26898 , w26899 , w26900 , w26901 , w26902 , w26903 , w26904 , w26905 , w26906 , w26907 , w26908 , w26909 , w26910 , w26911 , w26912 , w26913 , w26914 , w26915 , w26916 , w26917 , w26918 , w26919 , w26920 , w26921 , w26922 , w26923 , w26924 , w26925 , w26926 , w26927 , w26928 , w26929 , w26930 , w26931 , w26932 , w26933 , w26934 , w26935 , w26936 , w26937 , w26938 , w26939 , w26940 , w26941 , w26942 , w26943 , w26944 , w26945 , w26946 , w26947 , w26948 , w26949 , w26950 , w26951 , w26952 , w26953 , w26954 , w26955 , w26956 , w26957 , w26958 , w26959 , w26960 , w26961 , w26962 , w26963 , w26964 , w26965 , w26966 , w26967 , w26968 , w26969 , w26970 , w26971 , w26972 , w26973 , w26974 , w26975 , w26976 , w26977 , w26978 , w26979 , w26980 , w26981 , w26982 , w26983 , w26984 , w26985 , w26986 , w26987 , w26988 , w26989 , w26990 , w26991 , w26992 , w26993 , w26994 , w26995 , w26996 , w26997 , w26998 , w26999 , w27000 , w27001 , w27002 , w27003 , w27004 , w27005 , w27006 , w27007 , w27008 , w27009 , w27010 , w27011 , w27012 , w27013 , w27014 , w27015 , w27016 , w27017 , w27018 , w27019 , w27020 , w27021 , w27022 , w27023 , w27024 , w27025 , w27026 , w27027 , w27028 , w27029 , w27030 , w27031 , w27032 , w27033 , w27034 , w27035 , w27036 , w27037 , w27038 , w27039 , w27040 , w27041 , w27042 , w27043 , w27044 , w27045 , w27046 , w27047 , w27048 , w27049 , w27050 , w27051 , w27052 , w27053 , w27054 , w27055 , w27056 , w27057 , w27058 , w27059 , w27060 , w27061 , w27062 , w27063 , w27064 , w27065 , w27066 , w27067 , w27068 , w27069 , w27070 , w27071 , w27072 , w27073 , w27074 , w27075 , w27076 , w27077 , w27078 , w27079 , w27080 , w27081 , w27082 , w27083 , w27084 , w27085 , w27086 , w27087 , w27088 , w27089 , w27090 , w27091 , w27092 , w27093 , w27094 , w27095 , w27096 , w27097 , w27098 , w27099 , w27100 , w27101 , w27102 , w27103 , w27104 , w27105 , w27106 , w27107 , w27108 , w27109 , w27110 , w27111 , w27112 , w27113 , w27114 , w27115 , w27116 , w27117 , w27118 , w27119 , w27120 , w27121 , w27122 , w27123 , w27124 , w27125 , w27126 , w27127 , w27128 , w27129 , w27130 , w27131 , w27132 , w27133 , w27134 , w27135 , w27136 , w27137 , w27138 , w27139 , w27140 , w27141 , w27142 , w27143 , w27144 , w27145 , w27146 , w27147 , w27148 , w27149 , w27150 , w27151 , w27152 , w27153 , w27154 , w27155 , w27156 , w27157 , w27158 , w27159 , w27160 , w27161 , w27162 , w27163 , w27164 , w27165 , w27166 , w27167 , w27168 , w27169 , w27170 , w27171 , w27172 , w27173 , w27174 , w27175 , w27176 , w27177 , w27178 , w27179 , w27180 , w27181 , w27182 , w27183 , w27184 , w27185 , w27186 , w27187 , w27188 , w27189 , w27190 , w27191 , w27192 , w27193 , w27194 , w27195 , w27196 , w27197 , w27198 , w27199 , w27200 , w27201 , w27202 , w27203 , w27204 , w27205 , w27206 , w27207 , w27208 , w27209 , w27210 , w27211 , w27212 , w27213 , w27214 , w27215 , w27216 , w27217 , w27218 , w27219 , w27220 , w27221 , w27222 , w27223 , w27224 , w27225 , w27226 , w27227 , w27228 , w27229 , w27230 , w27231 , w27232 , w27233 , w27234 , w27235 , w27236 , w27237 , w27238 , w27239 , w27240 , w27241 , w27242 , w27243 , w27244 , w27245 , w27246 , w27247 , w27248 , w27249 , w27250 , w27251 , w27252 , w27253 , w27254 , w27255 , w27256 , w27257 , w27258 , w27259 , w27260 , w27261 , w27262 , w27263 , w27264 , w27265 , w27266 , w27267 , w27268 , w27269 , w27270 , w27271 , w27272 , w27273 , w27274 , w27275 , w27276 , w27277 , w27278 , w27279 , w27280 , w27281 , w27282 , w27283 , w27284 , w27285 , w27286 , w27287 , w27288 , w27289 , w27290 , w27291 , w27292 , w27293 , w27294 , w27295 , w27296 , w27297 , w27298 , w27299 , w27300 , w27301 , w27302 , w27303 , w27304 , w27305 , w27306 , w27307 , w27308 , w27309 , w27310 , w27311 , w27312 , w27313 , w27314 , w27315 , w27316 , w27317 , w27318 , w27319 , w27320 , w27321 , w27322 , w27323 , w27324 , w27325 , w27326 , w27327 , w27328 , w27329 , w27330 , w27331 , w27332 , w27333 , w27334 , w27335 , w27336 , w27337 , w27338 , w27339 , w27340 , w27341 , w27342 , w27343 , w27344 , w27345 , w27346 , w27347 , w27348 , w27349 , w27350 , w27351 , w27352 , w27353 , w27354 , w27355 , w27356 , w27357 , w27358 , w27359 , w27360 , w27361 , w27362 , w27363 , w27364 , w27365 , w27366 , w27367 , w27368 , w27369 , w27370 , w27371 , w27372 , w27373 , w27374 , w27375 , w27376 , w27377 , w27378 , w27379 , w27380 , w27381 , w27382 , w27383 , w27384 , w27385 , w27386 , w27387 , w27388 , w27389 , w27390 , w27391 , w27392 , w27393 , w27394 , w27395 , w27396 , w27397 , w27398 , w27399 , w27400 , w27401 , w27402 , w27403 , w27404 , w27405 , w27406 , w27407 , w27408 , w27409 , w27410 , w27411 , w27412 , w27413 , w27414 , w27415 , w27416 , w27417 , w27418 , w27419 , w27420 , w27421 , w27422 , w27423 , w27424 , w27425 , w27426 , w27427 , w27428 , w27429 , w27430 , w27431 , w27432 , w27433 , w27434 , w27435 , w27436 , w27437 , w27438 , w27439 , w27440 , w27441 , w27442 , w27443 , w27444 , w27445 , w27446 , w27447 , w27448 , w27449 , w27450 , w27451 , w27452 , w27453 , w27454 , w27455 , w27456 , w27457 , w27458 , w27459 , w27460 , w27461 , w27462 , w27463 , w27464 , w27465 , w27466 , w27467 , w27468 , w27469 , w27470 , w27471 , w27472 , w27473 , w27474 , w27475 , w27476 , w27477 , w27478 , w27479 , w27480 , w27481 , w27482 , w27483 , w27484 , w27485 , w27486 , w27487 , w27488 , w27489 , w27490 , w27491 , w27492 , w27493 , w27494 , w27495 , w27496 , w27497 , w27498 , w27499 , w27500 , w27501 , w27502 , w27503 , w27504 , w27505 , w27506 , w27507 , w27508 , w27509 , w27510 , w27511 , w27512 , w27513 , w27514 , w27515 , w27516 , w27517 , w27518 , w27519 , w27520 , w27521 , w27522 , w27523 , w27524 , w27525 , w27526 , w27527 , w27528 , w27529 , w27530 , w27531 , w27532 , w27533 , w27534 , w27535 , w27536 , w27537 , w27538 , w27539 , w27540 , w27541 , w27542 , w27543 , w27544 , w27545 , w27546 , w27547 , w27548 , w27549 , w27550 , w27551 , w27552 , w27553 , w27554 , w27555 , w27556 , w27557 , w27558 , w27559 , w27560 , w27561 , w27562 , w27563 , w27564 , w27565 , w27566 , w27567 , w27568 , w27569 , w27570 , w27571 , w27572 , w27573 , w27574 , w27575 , w27576 , w27577 , w27578 , w27579 , w27580 , w27581 , w27582 , w27583 , w27584 , w27585 , w27586 , w27587 , w27588 , w27589 , w27590 , w27591 , w27592 , w27593 , w27594 , w27595 , w27596 , w27597 , w27598 , w27599 , w27600 , w27601 , w27602 , w27603 , w27604 , w27605 , w27606 , w27607 , w27608 , w27609 , w27610 , w27611 , w27612 , w27613 , w27614 , w27615 , w27616 , w27617 , w27618 , w27619 , w27620 , w27621 , w27622 , w27623 , w27624 , w27625 , w27626 , w27627 , w27628 , w27629 , w27630 , w27631 , w27632 , w27633 , w27634 , w27635 , w27636 , w27637 , w27638 , w27639 , w27640 , w27641 , w27642 , w27643 , w27644 , w27645 , w27646 , w27647 , w27648 , w27649 , w27650 , w27651 , w27652 , w27653 , w27654 , w27655 , w27656 , w27657 , w27658 , w27659 , w27660 , w27661 , w27662 , w27663 , w27664 , w27665 , w27666 , w27667 , w27668 , w27669 , w27670 , w27671 , w27672 , w27673 , w27674 , w27675 , w27676 , w27677 , w27678 , w27679 , w27680 , w27681 , w27682 , w27683 , w27684 , w27685 , w27686 , w27687 , w27688 , w27689 , w27690 , w27691 , w27692 , w27693 , w27694 , w27695 , w27696 , w27697 , w27698 , w27699 , w27700 , w27701 , w27702 , w27703 , w27704 , w27705 , w27706 , w27707 , w27708 , w27709 , w27710 , w27711 , w27712 , w27713 , w27714 , w27715 , w27716 , w27717 , w27718 , w27719 , w27720 , w27721 , w27722 , w27723 , w27724 , w27725 , w27726 , w27727 , w27728 , w27729 , w27730 , w27731 , w27732 , w27733 , w27734 , w27735 , w27736 , w27737 , w27738 , w27739 , w27740 , w27741 , w27742 , w27743 , w27744 , w27745 , w27746 , w27747 , w27748 , w27749 , w27750 , w27751 , w27752 , w27753 , w27754 , w27755 , w27756 , w27757 , w27758 , w27759 , w27760 , w27761 , w27762 , w27763 , w27764 , w27765 , w27766 , w27767 , w27768 , w27769 , w27770 , w27771 , w27772 , w27773 , w27774 , w27775 , w27776 , w27777 , w27778 , w27779 , w27780 , w27781 , w27782 , w27783 , w27784 , w27785 , w27786 , w27787 , w27788 , w27789 , w27790 , w27791 , w27792 , w27793 , w27794 , w27795 , w27796 , w27797 , w27798 , w27799 , w27800 , w27801 , w27802 , w27803 , w27804 , w27805 , w27806 , w27807 , w27808 , w27809 , w27810 , w27811 , w27812 , w27813 , w27814 , w27815 , w27816 , w27817 , w27818 , w27819 , w27820 , w27821 , w27822 , w27823 , w27824 , w27825 , w27826 , w27827 , w27828 , w27829 , w27830 , w27831 , w27832 , w27833 , w27834 , w27835 , w27836 , w27837 , w27838 , w27839 , w27840 , w27841 , w27842 , w27843 , w27844 , w27845 , w27846 , w27847 , w27848 , w27849 , w27850 , w27851 , w27852 , w27853 , w27854 , w27855 , w27856 , w27857 , w27858 , w27859 , w27860 , w27861 , w27862 , w27863 , w27864 , w27865 , w27866 , w27867 , w27868 , w27869 , w27870 , w27871 , w27872 , w27873 , w27874 , w27875 , w27876 , w27877 , w27878 , w27879 , w27880 , w27881 , w27882 , w27883 , w27884 , w27885 , w27886 , w27887 , w27888 , w27889 , w27890 , w27891 , w27892 , w27893 , w27894 , w27895 , w27896 , w27897 , w27898 , w27899 , w27900 , w27901 , w27902 , w27903 , w27904 , w27905 , w27906 , w27907 , w27908 , w27909 , w27910 , w27911 , w27912 , w27913 , w27914 , w27915 , w27916 , w27917 , w27918 , w27919 , w27920 , w27921 , w27922 , w27923 , w27924 , w27925 , w27926 , w27927 , w27928 , w27929 , w27930 , w27931 , w27932 , w27933 , w27934 , w27935 , w27936 , w27937 , w27938 , w27939 , w27940 , w27941 , w27942 , w27943 , w27944 , w27945 , w27946 , w27947 , w27948 , w27949 , w27950 , w27951 , w27952 , w27953 , w27954 , w27955 , w27956 , w27957 , w27958 , w27959 , w27960 , w27961 , w27962 , w27963 , w27964 , w27965 , w27966 , w27967 , w27968 , w27969 , w27970 , w27971 , w27972 , w27973 , w27974 , w27975 , w27976 , w27977 , w27978 , w27979 , w27980 , w27981 , w27982 , w27983 , w27984 , w27985 , w27986 , w27987 , w27988 , w27989 , w27990 , w27991 , w27992 , w27993 , w27994 , w27995 , w27996 , w27997 , w27998 , w27999 , w28000 , w28001 , w28002 , w28003 , w28004 , w28005 , w28006 , w28007 , w28008 , w28009 , w28010 , w28011 , w28012 , w28013 , w28014 , w28015 , w28016 , w28017 , w28018 , w28019 , w28020 , w28021 , w28022 , w28023 , w28024 , w28025 , w28026 , w28027 , w28028 , w28029 , w28030 , w28031 , w28032 , w28033 , w28034 , w28035 , w28036 , w28037 , w28038 , w28039 , w28040 , w28041 , w28042 , w28043 , w28044 , w28045 , w28046 , w28047 , w28048 , w28049 , w28050 , w28051 , w28052 , w28053 , w28054 , w28055 , w28056 , w28057 , w28058 , w28059 , w28060 , w28061 , w28062 , w28063 , w28064 , w28065 , w28066 , w28067 , w28068 , w28069 , w28070 , w28071 , w28072 , w28073 , w28074 , w28075 , w28076 , w28077 , w28078 , w28079 , w28080 , w28081 , w28082 , w28083 , w28084 , w28085 , w28086 , w28087 , w28088 , w28089 , w28090 , w28091 , w28092 , w28093 , w28094 , w28095 , w28096 , w28097 , w28098 , w28099 , w28100 , w28101 , w28102 , w28103 , w28104 , w28105 , w28106 , w28107 , w28108 , w28109 , w28110 , w28111 , w28112 , w28113 , w28114 , w28115 , w28116 , w28117 , w28118 , w28119 , w28120 , w28121 , w28122 , w28123 , w28124 , w28125 , w28126 , w28127 , w28128 , w28129 , w28130 , w28131 , w28132 , w28133 , w28134 , w28135 , w28136 , w28137 , w28138 , w28139 , w28140 , w28141 , w28142 , w28143 , w28144 , w28145 , w28146 , w28147 , w28148 , w28149 , w28150 , w28151 , w28152 , w28153 , w28154 , w28155 , w28156 , w28157 , w28158 , w28159 , w28160 , w28161 , w28162 , w28163 , w28164 , w28165 , w28166 , w28167 , w28168 , w28169 , w28170 , w28171 , w28172 , w28173 , w28174 , w28175 , w28176 , w28177 , w28178 , w28179 , w28180 , w28181 , w28182 , w28183 , w28184 , w28185 , w28186 , w28187 , w28188 , w28189 , w28190 , w28191 , w28192 , w28193 , w28194 , w28195 , w28196 , w28197 , w28198 , w28199 , w28200 , w28201 , w28202 , w28203 , w28204 , w28205 , w28206 , w28207 , w28208 , w28209 , w28210 , w28211 , w28212 , w28213 , w28214 , w28215 , w28216 , w28217 , w28218 , w28219 , w28220 , w28221 , w28222 , w28223 , w28224 , w28225 , w28226 , w28227 , w28228 , w28229 , w28230 , w28231 , w28232 , w28233 , w28234 , w28235 , w28236 , w28237 , w28238 , w28239 , w28240 , w28241 , w28242 , w28243 , w28244 , w28245 , w28246 , w28247 , w28248 , w28249 , w28250 , w28251 , w28252 , w28253 , w28254 , w28255 , w28256 , w28257 , w28258 , w28259 , w28260 , w28261 , w28262 , w28263 , w28264 , w28265 , w28266 , w28267 , w28268 , w28269 , w28270 , w28271 , w28272 , w28273 , w28274 , w28275 , w28276 , w28277 , w28278 , w28279 , w28280 , w28281 , w28282 , w28283 , w28284 , w28285 , w28286 , w28287 , w28288 , w28289 , w28290 , w28291 , w28292 , w28293 , w28294 , w28295 , w28296 , w28297 , w28298 , w28299 , w28300 , w28301 , w28302 , w28303 , w28304 , w28305 , w28306 , w28307 , w28308 , w28309 , w28310 , w28311 , w28312 , w28313 , w28314 , w28315 , w28316 , w28317 , w28318 , w28319 , w28320 , w28321 , w28322 , w28323 , w28324 , w28325 , w28326 , w28327 , w28328 , w28329 , w28330 , w28331 , w28332 , w28333 , w28334 , w28335 , w28336 , w28337 , w28338 , w28339 , w28340 , w28341 , w28342 , w28343 , w28344 , w28345 , w28346 , w28347 , w28348 , w28349 , w28350 , w28351 , w28352 , w28353 , w28354 , w28355 , w28356 , w28357 , w28358 , w28359 , w28360 , w28361 , w28362 , w28363 , w28364 , w28365 , w28366 , w28367 , w28368 , w28369 , w28370 , w28371 , w28372 , w28373 , w28374 , w28375 , w28376 , w28377 , w28378 , w28379 , w28380 , w28381 , w28382 , w28383 , w28384 , w28385 , w28386 , w28387 , w28388 , w28389 , w28390 , w28391 , w28392 , w28393 , w28394 , w28395 , w28396 , w28397 , w28398 , w28399 , w28400 , w28401 , w28402 , w28403 , w28404 , w28405 , w28406 , w28407 , w28408 , w28409 , w28410 , w28411 , w28412 , w28413 , w28414 , w28415 , w28416 , w28417 , w28418 , w28419 , w28420 , w28421 , w28422 , w28423 , w28424 , w28425 , w28426 , w28427 , w28428 , w28429 , w28430 , w28431 , w28432 , w28433 , w28434 , w28435 , w28436 , w28437 , w28438 , w28439 , w28440 , w28441 , w28442 , w28443 , w28444 , w28445 , w28446 , w28447 , w28448 , w28449 , w28450 , w28451 , w28452 , w28453 , w28454 , w28455 , w28456 , w28457 , w28458 , w28459 , w28460 , w28461 , w28462 , w28463 , w28464 , w28465 , w28466 , w28467 , w28468 , w28469 , w28470 , w28471 , w28472 , w28473 , w28474 , w28475 , w28476 , w28477 , w28478 , w28479 , w28480 , w28481 , w28482 , w28483 , w28484 , w28485 , w28486 , w28487 , w28488 , w28489 , w28490 , w28491 , w28492 , w28493 , w28494 , w28495 , w28496 , w28497 , w28498 , w28499 , w28500 , w28501 , w28502 , w28503 , w28504 , w28505 , w28506 , w28507 , w28508 , w28509 , w28510 , w28511 , w28512 , w28513 , w28514 , w28515 , w28516 , w28517 , w28518 , w28519 , w28520 , w28521 , w28522 , w28523 , w28524 , w28525 , w28526 , w28527 , w28528 , w28529 , w28530 , w28531 , w28532 , w28533 , w28534 , w28535 , w28536 , w28537 , w28538 , w28539 , w28540 , w28541 , w28542 , w28543 , w28544 , w28545 , w28546 , w28547 , w28548 , w28549 , w28550 , w28551 , w28552 , w28553 , w28554 , w28555 , w28556 , w28557 , w28558 , w28559 , w28560 , w28561 , w28562 , w28563 , w28564 , w28565 , w28566 , w28567 , w28568 , w28569 , w28570 , w28571 , w28572 , w28573 , w28574 , w28575 , w28576 , w28577 , w28578 , w28579 , w28580 , w28581 , w28582 , w28583 , w28584 , w28585 , w28586 , w28587 , w28588 , w28589 , w28590 , w28591 , w28592 , w28593 , w28594 , w28595 , w28596 , w28597 , w28598 , w28599 , w28600 , w28601 , w28602 , w28603 , w28604 , w28605 , w28606 , w28607 , w28608 , w28609 , w28610 , w28611 , w28612 , w28613 , w28614 , w28615 , w28616 , w28617 , w28618 , w28619 , w28620 , w28621 , w28622 , w28623 , w28624 , w28625 , w28626 , w28627 , w28628 , w28629 , w28630 , w28631 , w28632 , w28633 , w28634 , w28635 , w28636 , w28637 , w28638 , w28639 , w28640 , w28641 , w28642 , w28643 , w28644 , w28645 , w28646 , w28647 , w28648 , w28649 , w28650 , w28651 , w28652 , w28653 , w28654 , w28655 , w28656 , w28657 , w28658 , w28659 , w28660 , w28661 , w28662 , w28663 , w28664 , w28665 , w28666 , w28667 , w28668 , w28669 , w28670 , w28671 , w28672 , w28673 , w28674 , w28675 , w28676 , w28677 , w28678 , w28679 , w28680 , w28681 , w28682 , w28683 , w28684 , w28685 , w28686 , w28687 , w28688 , w28689 , w28690 , w28691 , w28692 , w28693 , w28694 , w28695 , w28696 , w28697 , w28698 , w28699 , w28700 , w28701 , w28702 , w28703 , w28704 , w28705 , w28706 , w28707 , w28708 , w28709 , w28710 , w28711 , w28712 , w28713 , w28714 , w28715 , w28716 , w28717 , w28718 , w28719 , w28720 , w28721 , w28722 , w28723 , w28724 , w28725 , w28726 , w28727 , w28728 , w28729 , w28730 , w28731 , w28732 , w28733 , w28734 , w28735 , w28736 , w28737 , w28738 , w28739 , w28740 , w28741 , w28742 , w28743 , w28744 , w28745 , w28746 , w28747 , w28748 , w28749 , w28750 , w28751 , w28752 , w28753 , w28754 , w28755 , w28756 , w28757 , w28758 , w28759 , w28760 , w28761 , w28762 , w28763 , w28764 , w28765 , w28766 , w28767 , w28768 , w28769 , w28770 , w28771 , w28772 , w28773 , w28774 , w28775 , w28776 , w28777 , w28778 , w28779 , w28780 , w28781 , w28782 , w28783 , w28784 , w28785 , w28786 , w28787 , w28788 , w28789 , w28790 , w28791 , w28792 , w28793 , w28794 , w28795 , w28796 , w28797 , w28798 , w28799 , w28800 , w28801 , w28802 , w28803 , w28804 , w28805 , w28806 , w28807 , w28808 , w28809 , w28810 , w28811 , w28812 , w28813 , w28814 , w28815 , w28816 , w28817 , w28818 , w28819 , w28820 , w28821 , w28822 , w28823 , w28824 , w28825 , w28826 , w28827 , w28828 , w28829 , w28830 , w28831 , w28832 , w28833 , w28834 , w28835 , w28836 , w28837 , w28838 , w28839 , w28840 , w28841 , w28842 , w28843 , w28844 , w28845 , w28846 , w28847 , w28848 , w28849 , w28850 , w28851 , w28852 , w28853 , w28854 , w28855 , w28856 , w28857 , w28858 , w28859 , w28860 , w28861 , w28862 , w28863 , w28864 , w28865 , w28866 , w28867 , w28868 , w28869 , w28870 , w28871 , w28872 , w28873 , w28874 , w28875 , w28876 , w28877 , w28878 , w28879 , w28880 , w28881 , w28882 , w28883 , w28884 , w28885 , w28886 , w28887 , w28888 , w28889 , w28890 , w28891 , w28892 , w28893 , w28894 , w28895 , w28896 , w28897 , w28898 , w28899 , w28900 , w28901 , w28902 , w28903 , w28904 , w28905 , w28906 , w28907 , w28908 , w28909 , w28910 , w28911 , w28912 , w28913 , w28914 , w28915 , w28916 , w28917 , w28918 , w28919 , w28920 , w28921 , w28922 , w28923 , w28924 , w28925 , w28926 , w28927 , w28928 , w28929 , w28930 , w28931 , w28932 , w28933 , w28934 , w28935 , w28936 , w28937 , w28938 , w28939 , w28940 , w28941 , w28942 , w28943 , w28944 , w28945 , w28946 , w28947 , w28948 , w28949 , w28950 , w28951 , w28952 , w28953 , w28954 , w28955 , w28956 , w28957 , w28958 , w28959 , w28960 , w28961 , w28962 , w28963 , w28964 , w28965 , w28966 , w28967 , w28968 , w28969 , w28970 , w28971 , w28972 , w28973 , w28974 , w28975 , w28976 , w28977 , w28978 , w28979 , w28980 , w28981 , w28982 , w28983 , w28984 , w28985 , w28986 , w28987 , w28988 , w28989 , w28990 , w28991 , w28992 , w28993 , w28994 , w28995 , w28996 , w28997 , w28998 , w28999 , w29000 , w29001 , w29002 , w29003 , w29004 , w29005 , w29006 , w29007 , w29008 , w29009 , w29010 , w29011 , w29012 , w29013 , w29014 , w29015 , w29016 , w29017 , w29018 , w29019 , w29020 , w29021 , w29022 , w29023 , w29024 , w29025 , w29026 , w29027 , w29028 , w29029 , w29030 , w29031 , w29032 , w29033 , w29034 , w29035 , w29036 , w29037 , w29038 , w29039 , w29040 , w29041 , w29042 , w29043 , w29044 , w29045 , w29046 , w29047 , w29048 , w29049 , w29050 , w29051 , w29052 , w29053 , w29054 , w29055 , w29056 , w29057 , w29058 , w29059 , w29060 , w29061 , w29062 , w29063 , w29064 , w29065 , w29066 , w29067 , w29068 , w29069 , w29070 , w29071 , w29072 , w29073 , w29074 , w29075 , w29076 , w29077 , w29078 , w29079 , w29080 , w29081 , w29082 , w29083 , w29084 , w29085 , w29086 , w29087 , w29088 , w29089 , w29090 , w29091 , w29092 , w29093 , w29094 , w29095 , w29096 , w29097 , w29098 , w29099 , w29100 , w29101 , w29102 , w29103 , w29104 , w29105 , w29106 , w29107 , w29108 , w29109 , w29110 , w29111 , w29112 , w29113 , w29114 , w29115 , w29116 , w29117 , w29118 , w29119 , w29120 , w29121 , w29122 , w29123 , w29124 , w29125 , w29126 , w29127 , w29128 , w29129 , w29130 , w29131 , w29132 , w29133 , w29134 , w29135 , w29136 , w29137 , w29138 , w29139 , w29140 , w29141 , w29142 , w29143 , w29144 , w29145 , w29146 , w29147 , w29148 , w29149 , w29150 , w29151 , w29152 , w29153 , w29154 , w29155 , w29156 , w29157 , w29158 , w29159 , w29160 , w29161 , w29162 , w29163 , w29164 , w29165 , w29166 , w29167 , w29168 , w29169 , w29170 , w29171 , w29172 , w29173 , w29174 , w29175 , w29176 , w29177 , w29178 , w29179 , w29180 , w29181 , w29182 , w29183 , w29184 , w29185 , w29186 , w29187 , w29188 , w29189 , w29190 , w29191 , w29192 , w29193 , w29194 , w29195 , w29196 , w29197 , w29198 , w29199 , w29200 , w29201 , w29202 , w29203 , w29204 , w29205 , w29206 , w29207 , w29208 , w29209 , w29210 , w29211 , w29212 , w29213 , w29214 , w29215 , w29216 , w29217 , w29218 , w29219 , w29220 , w29221 , w29222 , w29223 , w29224 , w29225 , w29226 , w29227 , w29228 , w29229 , w29230 , w29231 , w29232 , w29233 , w29234 , w29235 , w29236 , w29237 , w29238 , w29239 , w29240 , w29241 , w29242 , w29243 , w29244 , w29245 , w29246 , w29247 , w29248 , w29249 , w29250 , w29251 , w29252 , w29253 , w29254 , w29255 , w29256 , w29257 , w29258 , w29259 , w29260 , w29261 , w29262 , w29263 , w29264 , w29265 , w29266 , w29267 , w29268 , w29269 , w29270 , w29271 , w29272 , w29273 , w29274 , w29275 , w29276 , w29277 , w29278 , w29279 , w29280 , w29281 , w29282 , w29283 , w29284 , w29285 , w29286 , w29287 , w29288 , w29289 , w29290 , w29291 , w29292 , w29293 , w29294 , w29295 , w29296 , w29297 , w29298 , w29299 , w29300 , w29301 , w29302 , w29303 , w29304 , w29305 , w29306 , w29307 , w29308 , w29309 , w29310 , w29311 , w29312 , w29313 , w29314 , w29315 , w29316 , w29317 , w29318 , w29319 , w29320 , w29321 , w29322 , w29323 , w29324 , w29325 , w29326 , w29327 , w29328 , w29329 , w29330 , w29331 , w29332 , w29333 , w29334 , w29335 , w29336 , w29337 , w29338 , w29339 , w29340 , w29341 , w29342 , w29343 , w29344 , w29345 , w29346 , w29347 , w29348 , w29349 , w29350 , w29351 , w29352 , w29353 , w29354 , w29355 , w29356 , w29357 , w29358 , w29359 , w29360 , w29361 , w29362 , w29363 , w29364 , w29365 , w29366 , w29367 , w29368 , w29369 , w29370 , w29371 , w29372 , w29373 , w29374 , w29375 , w29376 , w29377 , w29378 , w29379 , w29380 , w29381 , w29382 , w29383 , w29384 , w29385 , w29386 , w29387 , w29388 , w29389 , w29390 , w29391 , w29392 , w29393 , w29394 , w29395 , w29396 , w29397 , w29398 , w29399 , w29400 , w29401 , w29402 , w29403 , w29404 , w29405 , w29406 , w29407 , w29408 , w29409 , w29410 , w29411 , w29412 , w29413 , w29414 , w29415 , w29416 , w29417 , w29418 , w29419 , w29420 , w29421 , w29422 , w29423 , w29424 , w29425 , w29426 , w29427 , w29428 , w29429 , w29430 , w29431 , w29432 , w29433 , w29434 , w29435 , w29436 , w29437 , w29438 , w29439 , w29440 , w29441 , w29442 , w29443 , w29444 , w29445 , w29446 , w29447 , w29448 , w29449 , w29450 , w29451 , w29452 , w29453 , w29454 , w29455 , w29456 , w29457 , w29458 , w29459 , w29460 , w29461 , w29462 , w29463 , w29464 , w29465 , w29466 , w29467 , w29468 , w29469 , w29470 , w29471 , w29472 , w29473 , w29474 , w29475 , w29476 , w29477 , w29478 , w29479 , w29480 , w29481 , w29482 , w29483 , w29484 , w29485 , w29486 , w29487 , w29488 , w29489 , w29490 , w29491 , w29492 , w29493 , w29494 , w29495 , w29496 , w29497 , w29498 , w29499 , w29500 , w29501 , w29502 , w29503 , w29504 , w29505 , w29506 , w29507 , w29508 , w29509 , w29510 , w29511 , w29512 , w29513 , w29514 , w29515 , w29516 , w29517 , w29518 , w29519 , w29520 , w29521 , w29522 , w29523 , w29524 , w29525 , w29526 , w29527 , w29528 , w29529 , w29530 , w29531 , w29532 , w29533 , w29534 , w29535 , w29536 , w29537 , w29538 , w29539 , w29540 , w29541 , w29542 , w29543 , w29544 , w29545 , w29546 , w29547 , w29548 , w29549 , w29550 , w29551 , w29552 , w29553 , w29554 , w29555 , w29556 , w29557 , w29558 , w29559 , w29560 , w29561 , w29562 , w29563 , w29564 , w29565 , w29566 , w29567 , w29568 , w29569 , w29570 , w29571 , w29572 , w29573 , w29574 , w29575 , w29576 , w29577 , w29578 , w29579 , w29580 , w29581 , w29582 , w29583 , w29584 , w29585 , w29586 , w29587 , w29588 , w29589 , w29590 , w29591 , w29592 , w29593 , w29594 , w29595 , w29596 , w29597 , w29598 , w29599 , w29600 , w29601 , w29602 , w29603 , w29604 , w29605 , w29606 , w29607 , w29608 , w29609 , w29610 , w29611 , w29612 , w29613 , w29614 , w29615 , w29616 , w29617 , w29618 , w29619 , w29620 , w29621 , w29622 , w29623 , w29624 , w29625 , w29626 , w29627 , w29628 , w29629 , w29630 , w29631 , w29632 , w29633 , w29634 , w29635 , w29636 , w29637 , w29638 , w29639 , w29640 , w29641 , w29642 , w29643 , w29644 , w29645 , w29646 , w29647 , w29648 , w29649 , w29650 , w29651 , w29652 , w29653 , w29654 , w29655 , w29656 , w29657 , w29658 , w29659 , w29660 , w29661 , w29662 , w29663 , w29664 , w29665 , w29666 , w29667 , w29668 , w29669 , w29670 , w29671 , w29672 , w29673 , w29674 , w29675 , w29676 , w29677 , w29678 , w29679 , w29680 , w29681 , w29682 , w29683 , w29684 , w29685 , w29686 , w29687 , w29688 , w29689 , w29690 , w29691 , w29692 , w29693 , w29694 , w29695 , w29696 , w29697 , w29698 , w29699 , w29700 , w29701 , w29702 , w29703 , w29704 , w29705 , w29706 , w29707 , w29708 , w29709 , w29710 , w29711 , w29712 , w29713 , w29714 , w29715 , w29716 , w29717 , w29718 , w29719 , w29720 , w29721 , w29722 , w29723 , w29724 , w29725 , w29726 , w29727 , w29728 , w29729 , w29730 , w29731 , w29732 , w29733 , w29734 , w29735 , w29736 , w29737 , w29738 , w29739 , w29740 , w29741 , w29742 , w29743 , w29744 , w29745 , w29746 , w29747 , w29748 , w29749 , w29750 , w29751 , w29752 , w29753 , w29754 , w29755 , w29756 , w29757 , w29758 , w29759 , w29760 , w29761 , w29762 , w29763 , w29764 , w29765 , w29766 , w29767 , w29768 , w29769 , w29770 , w29771 , w29772 , w29773 , w29774 , w29775 , w29776 , w29777 , w29778 , w29779 , w29780 , w29781 , w29782 , w29783 , w29784 , w29785 , w29786 , w29787 , w29788 , w29789 , w29790 , w29791 , w29792 , w29793 , w29794 , w29795 , w29796 , w29797 , w29798 , w29799 , w29800 , w29801 , w29802 , w29803 , w29804 , w29805 , w29806 , w29807 , w29808 , w29809 , w29810 , w29811 , w29812 , w29813 , w29814 , w29815 , w29816 , w29817 , w29818 , w29819 , w29820 , w29821 , w29822 , w29823 , w29824 , w29825 , w29826 , w29827 , w29828 , w29829 , w29830 , w29831 , w29832 , w29833 , w29834 , w29835 , w29836 , w29837 , w29838 , w29839 , w29840 , w29841 , w29842 , w29843 , w29844 , w29845 , w29846 , w29847 , w29848 , w29849 , w29850 , w29851 , w29852 , w29853 , w29854 , w29855 , w29856 , w29857 , w29858 , w29859 , w29860 , w29861 , w29862 , w29863 , w29864 , w29865 , w29866 , w29867 , w29868 , w29869 , w29870 , w29871 , w29872 , w29873 , w29874 , w29875 , w29876 , w29877 , w29878 , w29879 , w29880 , w29881 , w29882 , w29883 , w29884 , w29885 , w29886 , w29887 , w29888 , w29889 , w29890 , w29891 , w29892 , w29893 , w29894 , w29895 , w29896 , w29897 , w29898 , w29899 , w29900 , w29901 , w29902 , w29903 , w29904 , w29905 , w29906 , w29907 , w29908 , w29909 , w29910 , w29911 , w29912 , w29913 , w29914 , w29915 , w29916 , w29917 , w29918 , w29919 , w29920 , w29921 , w29922 , w29923 , w29924 , w29925 , w29926 , w29927 , w29928 , w29929 , w29930 , w29931 , w29932 , w29933 , w29934 , w29935 , w29936 , w29937 , w29938 , w29939 , w29940 , w29941 , w29942 , w29943 , w29944 , w29945 , w29946 , w29947 , w29948 , w29949 , w29950 , w29951 , w29952 , w29953 , w29954 , w29955 , w29956 , w29957 , w29958 , w29959 , w29960 , w29961 , w29962 , w29963 , w29964 , w29965 , w29966 , w29967 , w29968 , w29969 , w29970 , w29971 , w29972 , w29973 , w29974 , w29975 , w29976 , w29977 , w29978 , w29979 , w29980 , w29981 , w29982 , w29983 , w29984 , w29985 , w29986 , w29987 , w29988 , w29989 , w29990 , w29991 , w29992 , w29993 , w29994 , w29995 , w29996 , w29997 , w29998 , w29999 , w30000 , w30001 , w30002 , w30003 , w30004 , w30005 , w30006 , w30007 , w30008 , w30009 , w30010 , w30011 , w30012 , w30013 , w30014 , w30015 , w30016 , w30017 , w30018 , w30019 , w30020 , w30021 , w30022 , w30023 , w30024 , w30025 , w30026 , w30027 , w30028 , w30029 , w30030 , w30031 , w30032 , w30033 , w30034 , w30035 , w30036 , w30037 , w30038 , w30039 , w30040 , w30041 , w30042 , w30043 , w30044 , w30045 , w30046 , w30047 , w30048 , w30049 , w30050 , w30051 , w30052 , w30053 , w30054 , w30055 , w30056 , w30057 , w30058 , w30059 , w30060 , w30061 , w30062 , w30063 , w30064 , w30065 , w30066 , w30067 , w30068 , w30069 , w30070 , w30071 , w30072 , w30073 , w30074 , w30075 , w30076 , w30077 , w30078 , w30079 , w30080 , w30081 , w30082 , w30083 , w30084 , w30085 , w30086 , w30087 , w30088 , w30089 , w30090 , w30091 , w30092 , w30093 , w30094 , w30095 , w30096 , w30097 , w30098 , w30099 , w30100 , w30101 , w30102 , w30103 , w30104 , w30105 , w30106 , w30107 , w30108 , w30109 , w30110 , w30111 , w30112 , w30113 , w30114 , w30115 , w30116 , w30117 , w30118 , w30119 , w30120 , w30121 , w30122 , w30123 , w30124 , w30125 , w30126 , w30127 , w30128 , w30129 , w30130 , w30131 , w30132 , w30133 , w30134 , w30135 , w30136 , w30137 , w30138 , w30139 , w30140 , w30141 , w30142 , w30143 , w30144 , w30145 , w30146 , w30147 , w30148 , w30149 , w30150 , w30151 , w30152 , w30153 , w30154 , w30155 , w30156 , w30157 , w30158 , w30159 , w30160 , w30161 , w30162 , w30163 , w30164 , w30165 , w30166 , w30167 , w30168 , w30169 , w30170 , w30171 , w30172 , w30173 , w30174 , w30175 , w30176 , w30177 , w30178 , w30179 , w30180 , w30181 , w30182 , w30183 , w30184 , w30185 , w30186 , w30187 , w30188 , w30189 , w30190 , w30191 , w30192 , w30193 , w30194 , w30195 , w30196 , w30197 , w30198 , w30199 , w30200 , w30201 , w30202 , w30203 , w30204 , w30205 , w30206 , w30207 , w30208 , w30209 , w30210 , w30211 , w30212 , w30213 , w30214 , w30215 , w30216 , w30217 , w30218 , w30219 , w30220 , w30221 , w30222 , w30223 , w30224 , w30225 , w30226 , w30227 , w30228 , w30229 , w30230 , w30231 , w30232 , w30233 , w30234 , w30235 , w30236 , w30237 , w30238 , w30239 , w30240 , w30241 , w30242 , w30243 , w30244 , w30245 , w30246 , w30247 , w30248 , w30249 , w30250 , w30251 , w30252 , w30253 , w30254 , w30255 , w30256 , w30257 , w30258 , w30259 , w30260 , w30261 , w30262 , w30263 , w30264 , w30265 , w30266 , w30267 , w30268 , w30269 , w30270 , w30271 , w30272 , w30273 , w30274 , w30275 , w30276 , w30277 , w30278 , w30279 , w30280 , w30281 , w30282 , w30283 , w30284 , w30285 , w30286 , w30287 , w30288 , w30289 , w30290 , w30291 , w30292 , w30293 , w30294 , w30295 , w30296 , w30297 , w30298 , w30299 , w30300 , w30301 , w30302 , w30303 , w30304 , w30305 , w30306 , w30307 , w30308 , w30309 , w30310 , w30311 , w30312 , w30313 , w30314 , w30315 , w30316 , w30317 , w30318 , w30319 , w30320 , w30321 , w30322 , w30323 , w30324 , w30325 , w30326 , w30327 , w30328 , w30329 , w30330 , w30331 , w30332 , w30333 , w30334 , w30335 , w30336 , w30337 , w30338 , w30339 , w30340 , w30341 , w30342 , w30343 , w30344 , w30345 , w30346 , w30347 , w30348 , w30349 , w30350 , w30351 , w30352 , w30353 , w30354 , w30355 , w30356 , w30357 , w30358 , w30359 , w30360 , w30361 , w30362 , w30363 , w30364 , w30365 , w30366 , w30367 , w30368 , w30369 , w30370 , w30371 , w30372 , w30373 , w30374 , w30375 , w30376 , w30377 , w30378 , w30379 , w30380 , w30381 , w30382 , w30383 , w30384 , w30385 , w30386 , w30387 , w30388 , w30389 , w30390 , w30391 , w30392 , w30393 , w30394 , w30395 , w30396 , w30397 , w30398 , w30399 , w30400 , w30401 , w30402 , w30403 , w30404 , w30405 , w30406 , w30407 , w30408 , w30409 , w30410 , w30411 , w30412 , w30413 , w30414 , w30415 , w30416 , w30417 , w30418 , w30419 , w30420 , w30421 , w30422 , w30423 , w30424 , w30425 , w30426 , w30427 , w30428 , w30429 , w30430 , w30431 , w30432 , w30433 , w30434 , w30435 , w30436 , w30437 , w30438 , w30439 , w30440 , w30441 , w30442 , w30443 , w30444 , w30445 , w30446 , w30447 , w30448 , w30449 , w30450 , w30451 , w30452 , w30453 , w30454 , w30455 , w30456 , w30457 , w30458 , w30459 , w30460 , w30461 , w30462 , w30463 , w30464 , w30465 , w30466 , w30467 , w30468 , w30469 , w30470 , w30471 , w30472 , w30473 , w30474 , w30475 , w30476 , w30477 , w30478 , w30479 , w30480 , w30481 , w30482 , w30483 , w30484 , w30485 , w30486 , w30487 , w30488 , w30489 , w30490 , w30491 , w30492 , w30493 , w30494 , w30495 , w30496 , w30497 , w30498 , w30499 , w30500 , w30501 , w30502 , w30503 , w30504 , w30505 , w30506 , w30507 , w30508 , w30509 , w30510 , w30511 , w30512 , w30513 , w30514 , w30515 , w30516 , w30517 , w30518 , w30519 , w30520 , w30521 , w30522 , w30523 , w30524 , w30525 , w30526 , w30527 , w30528 , w30529 , w30530 , w30531 , w30532 , w30533 , w30534 , w30535 , w30536 , w30537 , w30538 , w30539 , w30540 , w30541 , w30542 , w30543 , w30544 , w30545 , w30546 , w30547 , w30548 , w30549 , w30550 , w30551 , w30552 , w30553 , w30554 , w30555 , w30556 , w30557 , w30558 , w30559 , w30560 , w30561 , w30562 , w30563 , w30564 , w30565 , w30566 , w30567 , w30568 , w30569 , w30570 , w30571 , w30572 , w30573 , w30574 , w30575 , w30576 , w30577 , w30578 , w30579 , w30580 , w30581 , w30582 , w30583 , w30584 , w30585 , w30586 , w30587 , w30588 , w30589 , w30590 , w30591 , w30592 , w30593 , w30594 , w30595 , w30596 , w30597 , w30598 , w30599 , w30600 , w30601 , w30602 , w30603 , w30604 , w30605 , w30606 , w30607 , w30608 , w30609 , w30610 , w30611 , w30612 , w30613 , w30614 , w30615 , w30616 , w30617 , w30618 , w30619 , w30620 , w30621 , w30622 , w30623 , w30624 , w30625 , w30626 , w30627 , w30628 , w30629 , w30630 , w30631 , w30632 , w30633 , w30634 , w30635 , w30636 , w30637 , w30638 , w30639 , w30640 , w30641 , w30642 , w30643 , w30644 , w30645 , w30646 , w30647 , w30648 , w30649 , w30650 , w30651 , w30652 , w30653 , w30654 , w30655 , w30656 , w30657 , w30658 , w30659 , w30660 , w30661 , w30662 , w30663 , w30664 , w30665 , w30666 , w30667 , w30668 , w30669 , w30670 , w30671 , w30672 , w30673 , w30674 , w30675 , w30676 , w30677 , w30678 , w30679 , w30680 , w30681 , w30682 , w30683 , w30684 , w30685 , w30686 , w30687 , w30688 , w30689 , w30690 , w30691 , w30692 , w30693 , w30694 , w30695 , w30696 , w30697 , w30698 , w30699 , w30700 , w30701 , w30702 , w30703 , w30704 , w30705 , w30706 , w30707 , w30708 , w30709 , w30710 , w30711 , w30712 , w30713 , w30714 , w30715 , w30716 , w30717 , w30718 , w30719 , w30720 , w30721 , w30722 , w30723 , w30724 , w30725 , w30726 , w30727 , w30728 , w30729 , w30730 , w30731 , w30732 , w30733 , w30734 , w30735 , w30736 , w30737 , w30738 , w30739 , w30740 , w30741 , w30742 , w30743 , w30744 , w30745 , w30746 , w30747 , w30748 , w30749 , w30750 , w30751 , w30752 , w30753 , w30754 , w30755 , w30756 , w30757 , w30758 , w30759 , w30760 , w30761 , w30762 , w30763 , w30764 , w30765 , w30766 , w30767 , w30768 , w30769 , w30770 , w30771 , w30772 , w30773 , w30774 , w30775 , w30776 , w30777 , w30778 , w30779 , w30780 , w30781 , w30782 , w30783 , w30784 , w30785 , w30786 , w30787 , w30788 , w30789 , w30790 , w30791 , w30792 , w30793 , w30794 , w30795 , w30796 , w30797 , w30798 , w30799 , w30800 , w30801 , w30802 , w30803 , w30804 , w30805 , w30806 , w30807 , w30808 , w30809 , w30810 , w30811 , w30812 , w30813 , w30814 , w30815 , w30816 , w30817 , w30818 , w30819 , w30820 , w30821 , w30822 , w30823 , w30824 , w30825 , w30826 , w30827 , w30828 , w30829 , w30830 , w30831 , w30832 , w30833 , w30834 , w30835 , w30836 , w30837 , w30838 , w30839 , w30840 , w30841 , w30842 , w30843 , w30844 , w30845 , w30846 , w30847 , w30848 , w30849 , w30850 , w30851 , w30852 , w30853 , w30854 , w30855 , w30856 , w30857 , w30858 , w30859 , w30860 , w30861 , w30862 , w30863 , w30864 , w30865 , w30866 , w30867 , w30868 , w30869 , w30870 , w30871 , w30872 , w30873 , w30874 , w30875 , w30876 , w30877 , w30878 , w30879 , w30880 , w30881 , w30882 , w30883 , w30884 , w30885 , w30886 , w30887 , w30888 , w30889 , w30890 , w30891 , w30892 , w30893 , w30894 , w30895 , w30896 , w30897 , w30898 , w30899 , w30900 , w30901 , w30902 , w30903 , w30904 , w30905 , w30906 , w30907 , w30908 , w30909 , w30910 , w30911 , w30912 , w30913 , w30914 , w30915 , w30916 , w30917 , w30918 , w30919 , w30920 , w30921 , w30922 , w30923 , w30924 , w30925 , w30926 , w30927 , w30928 , w30929 , w30930 , w30931 , w30932 , w30933 , w30934 , w30935 , w30936 , w30937 , w30938 , w30939 , w30940 , w30941 , w30942 , w30943 , w30944 , w30945 , w30946 , w30947 , w30948 , w30949 , w30950 , w30951 , w30952 , w30953 , w30954 , w30955 , w30956 , w30957 , w30958 , w30959 , w30960 , w30961 , w30962 , w30963 , w30964 , w30965 , w30966 , w30967 , w30968 , w30969 , w30970 , w30971 , w30972 , w30973 , w30974 , w30975 , w30976 , w30977 , w30978 , w30979 , w30980 , w30981 , w30982 , w30983 , w30984 , w30985 , w30986 , w30987 , w30988 , w30989 , w30990 , w30991 , w30992 , w30993 , w30994 , w30995 , w30996 , w30997 , w30998 , w30999 , w31000 , w31001 , w31002 , w31003 , w31004 , w31005 , w31006 , w31007 , w31008 , w31009 , w31010 , w31011 , w31012 , w31013 , w31014 , w31015 , w31016 , w31017 , w31018 , w31019 , w31020 , w31021 , w31022 , w31023 , w31024 , w31025 , w31026 , w31027 , w31028 , w31029 , w31030 , w31031 , w31032 , w31033 , w31034 , w31035 , w31036 , w31037 , w31038 , w31039 , w31040 , w31041 , w31042 , w31043 , w31044 , w31045 , w31046 , w31047 , w31048 , w31049 , w31050 , w31051 , w31052 , w31053 , w31054 , w31055 , w31056 , w31057 , w31058 , w31059 , w31060 , w31061 , w31062 , w31063 , w31064 , w31065 , w31066 , w31067 , w31068 , w31069 , w31070 , w31071 , w31072 , w31073 , w31074 , w31075 , w31076 , w31077 , w31078 , w31079 , w31080 , w31081 , w31082 , w31083 , w31084 , w31085 , w31086 , w31087 , w31088 , w31089 , w31090 , w31091 , w31092 , w31093 , w31094 , w31095 , w31096 , w31097 , w31098 , w31099 , w31100 , w31101 , w31102 , w31103 , w31104 , w31105 , w31106 , w31107 , w31108 , w31109 , w31110 , w31111 , w31112 , w31113 , w31114 , w31115 , w31116 , w31117 , w31118 , w31119 , w31120 , w31121 , w31122 , w31123 , w31124 , w31125 , w31126 , w31127 , w31128 , w31129 , w31130 , w31131 , w31132 , w31133 , w31134 , w31135 , w31136 , w31137 , w31138 , w31139 , w31140 , w31141 , w31142 , w31143 , w31144 , w31145 , w31146 , w31147 , w31148 , w31149 , w31150 , w31151 , w31152 , w31153 , w31154 , w31155 , w31156 , w31157 , w31158 , w31159 , w31160 , w31161 , w31162 , w31163 , w31164 , w31165 , w31166 , w31167 , w31168 , w31169 , w31170 , w31171 , w31172 , w31173 , w31174 , w31175 , w31176 , w31177 , w31178 , w31179 , w31180 , w31181 , w31182 , w31183 , w31184 , w31185 , w31186 , w31187 , w31188 , w31189 , w31190 , w31191 , w31192 , w31193 , w31194 , w31195 , w31196 , w31197 , w31198 , w31199 , w31200 , w31201 , w31202 , w31203 , w31204 , w31205 , w31206 , w31207 , w31208 , w31209 , w31210 , w31211 , w31212 , w31213 , w31214 , w31215 , w31216 , w31217 , w31218 , w31219 , w31220 , w31221 , w31222 , w31223 , w31224 , w31225 , w31226 , w31227 , w31228 , w31229 , w31230 , w31231 , w31232 , w31233 , w31234 , w31235 , w31236 , w31237 , w31238 , w31239 , w31240 , w31241 , w31242 , w31243 , w31244 , w31245 , w31246 , w31247 , w31248 , w31249 , w31250 , w31251 , w31252 , w31253 , w31254 , w31255 , w31256 , w31257 , w31258 , w31259 , w31260 , w31261 , w31262 , w31263 , w31264 , w31265 , w31266 , w31267 , w31268 , w31269 , w31270 , w31271 , w31272 , w31273 , w31274 , w31275 , w31276 , w31277 , w31278 , w31279 , w31280 , w31281 , w31282 , w31283 , w31284 , w31285 , w31286 , w31287 , w31288 , w31289 , w31290 , w31291 , w31292 , w31293 , w31294 , w31295 , w31296 , w31297 , w31298 , w31299 , w31300 , w31301 , w31302 , w31303 , w31304 , w31305 , w31306 , w31307 , w31308 , w31309 , w31310 , w31311 , w31312 , w31313 , w31314 , w31315 , w31316 , w31317 , w31318 , w31319 , w31320 , w31321 , w31322 , w31323 , w31324 , w31325 , w31326 , w31327 , w31328 , w31329 , w31330 , w31331 , w31332 , w31333 , w31334 , w31335 , w31336 , w31337 , w31338 , w31339 , w31340 , w31341 , w31342 , w31343 , w31344 , w31345 , w31346 , w31347 , w31348 , w31349 , w31350 , w31351 , w31352 , w31353 , w31354 , w31355 , w31356 , w31357 , w31358 , w31359 , w31360 , w31361 , w31362 , w31363 , w31364 , w31365 , w31366 , w31367 , w31368 , w31369 , w31370 , w31371 , w31372 , w31373 , w31374 , w31375 , w31376 , w31377 , w31378 , w31379 , w31380 , w31381 , w31382 , w31383 , w31384 , w31385 , w31386 , w31387 , w31388 , w31389 , w31390 , w31391 , w31392 , w31393 , w31394 , w31395 , w31396 , w31397 , w31398 , w31399 , w31400 , w31401 , w31402 , w31403 , w31404 , w31405 , w31406 , w31407 , w31408 , w31409 , w31410 , w31411 , w31412 , w31413 , w31414 , w31415 , w31416 , w31417 , w31418 , w31419 , w31420 , w31421 , w31422 , w31423 , w31424 , w31425 , w31426 , w31427 , w31428 , w31429 , w31430 , w31431 , w31432 , w31433 , w31434 , w31435 , w31436 , w31437 , w31438 , w31439 , w31440 , w31441 , w31442 , w31443 , w31444 , w31445 , w31446 , w31447 , w31448 , w31449 , w31450 , w31451 , w31452 , w31453 , w31454 , w31455 , w31456 , w31457 , w31458 , w31459 , w31460 , w31461 , w31462 , w31463 , w31464 , w31465 , w31466 , w31467 , w31468 , w31469 , w31470 , w31471 , w31472 , w31473 , w31474 , w31475 , w31476 , w31477 , w31478 , w31479 , w31480 , w31481 , w31482 , w31483 , w31484 , w31485 , w31486 , w31487 , w31488 , w31489 , w31490 , w31491 , w31492 , w31493 , w31494 , w31495 , w31496 , w31497 , w31498 , w31499 , w31500 , w31501 , w31502 , w31503 , w31504 , w31505 , w31506 , w31507 , w31508 , w31509 , w31510 , w31511 , w31512 , w31513 , w31514 , w31515 , w31516 , w31517 , w31518 , w31519 , w31520 , w31521 , w31522 , w31523 , w31524 , w31525 , w31526 , w31527 , w31528 , w31529 , w31530 , w31531 , w31532 , w31533 , w31534 , w31535 , w31536 , w31537 , w31538 , w31539 , w31540 , w31541 , w31542 , w31543 , w31544 , w31545 , w31546 , w31547 , w31548 , w31549 , w31550 , w31551 , w31552 , w31553 , w31554 , w31555 , w31556 , w31557 , w31558 , w31559 , w31560 , w31561 , w31562 , w31563 , w31564 , w31565 , w31566 , w31567 , w31568 , w31569 , w31570 , w31571 , w31572 , w31573 , w31574 , w31575 , w31576 , w31577 , w31578 , w31579 , w31580 , w31581 , w31582 , w31583 , w31584 , w31585 , w31586 , w31587 , w31588 , w31589 , w31590 , w31591 , w31592 , w31593 , w31594 , w31595 , w31596 , w31597 , w31598 , w31599 , w31600 , w31601 , w31602 , w31603 , w31604 , w31605 , w31606 , w31607 , w31608 , w31609 , w31610 , w31611 , w31612 , w31613 , w31614 , w31615 , w31616 , w31617 , w31618 , w31619 , w31620 , w31621 , w31622 , w31623 , w31624 , w31625 , w31626 , w31627 , w31628 , w31629 , w31630 , w31631 , w31632 , w31633 , w31634 , w31635 , w31636 , w31637 , w31638 , w31639 , w31640 , w31641 , w31642 , w31643 , w31644 , w31645 , w31646 , w31647 , w31648 , w31649 , w31650 , w31651 , w31652 , w31653 , w31654 , w31655 , w31656 , w31657 , w31658 , w31659 , w31660 , w31661 , w31662 , w31663 , w31664 , w31665 , w31666 , w31667 , w31668 , w31669 , w31670 , w31671 , w31672 , w31673 , w31674 , w31675 , w31676 , w31677 , w31678 , w31679 , w31680 , w31681 , w31682 , w31683 , w31684 , w31685 , w31686 , w31687 , w31688 , w31689 , w31690 , w31691 , w31692 , w31693 , w31694 , w31695 , w31696 , w31697 , w31698 , w31699 , w31700 , w31701 , w31702 , w31703 , w31704 , w31705 , w31706 , w31707 , w31708 , w31709 , w31710 , w31711 , w31712 , w31713 , w31714 , w31715 , w31716 , w31717 , w31718 , w31719 , w31720 , w31721 , w31722 , w31723 , w31724 , w31725 , w31726 , w31727 , w31728 , w31729 , w31730 , w31731 , w31732 , w31733 , w31734 , w31735 , w31736 , w31737 , w31738 , w31739 , w31740 , w31741 , w31742 , w31743 , w31744 , w31745 , w31746 , w31747 , w31748 , w31749 , w31750 , w31751 , w31752 , w31753 , w31754 , w31755 , w31756 , w31757 , w31758 , w31759 , w31760 , w31761 , w31762 , w31763 , w31764 , w31765 , w31766 , w31767 , w31768 , w31769 , w31770 , w31771 , w31772 , w31773 , w31774 , w31775 , w31776 , w31777 , w31778 , w31779 , w31780 , w31781 , w31782 , w31783 , w31784 , w31785 , w31786 , w31787 , w31788 , w31789 , w31790 , w31791 , w31792 , w31793 , w31794 , w31795 , w31796 , w31797 , w31798 , w31799 , w31800 , w31801 , w31802 , w31803 , w31804 , w31805 , w31806 , w31807 , w31808 , w31809 , w31810 , w31811 , w31812 , w31813 , w31814 , w31815 , w31816 , w31817 , w31818 , w31819 , w31820 , w31821 , w31822 , w31823 , w31824 , w31825 , w31826 , w31827 , w31828 , w31829 , w31830 , w31831 , w31832 , w31833 , w31834 , w31835 , w31836 , w31837 , w31838 , w31839 , w31840 , w31841 , w31842 , w31843 , w31844 , w31845 , w31846 , w31847 , w31848 , w31849 , w31850 , w31851 , w31852 , w31853 , w31854 , w31855 , w31856 , w31857 , w31858 , w31859 , w31860 , w31861 , w31862 , w31863 , w31864 , w31865 , w31866 , w31867 , w31868 , w31869 , w31870 , w31871 , w31872 , w31873 , w31874 , w31875 , w31876 , w31877 , w31878 , w31879 , w31880 , w31881 , w31882 , w31883 , w31884 , w31885 , w31886 , w31887 , w31888 , w31889 , w31890 , w31891 , w31892 , w31893 , w31894 , w31895 , w31896 , w31897 , w31898 , w31899 , w31900 , w31901 , w31902 , w31903 , w31904 , w31905 , w31906 , w31907 , w31908 , w31909 , w31910 , w31911 , w31912 , w31913 , w31914 , w31915 , w31916 , w31917 , w31918 , w31919 , w31920 , w31921 , w31922 , w31923 , w31924 , w31925 , w31926 , w31927 , w31928 , w31929 , w31930 , w31931 , w31932 , w31933 , w31934 , w31935 , w31936 , w31937 , w31938 , w31939 , w31940 , w31941 , w31942 , w31943 , w31944 , w31945 , w31946 , w31947 , w31948 , w31949 , w31950 , w31951 , w31952 , w31953 , w31954 , w31955 , w31956 , w31957 , w31958 , w31959 , w31960 , w31961 , w31962 , w31963 , w31964 , w31965 , w31966 , w31967 , w31968 , w31969 , w31970 , w31971 , w31972 , w31973 , w31974 , w31975 , w31976 , w31977 , w31978 , w31979 , w31980 , w31981 , w31982 , w31983 , w31984 , w31985 , w31986 , w31987 , w31988 , w31989 , w31990 , w31991 , w31992 , w31993 , w31994 , w31995 , w31996 , w31997 , w31998 , w31999 , w32000 , w32001 , w32002 , w32003 , w32004 , w32005 , w32006 , w32007 , w32008 , w32009 , w32010 , w32011 , w32012 , w32013 , w32014 , w32015 , w32016 , w32017 , w32018 , w32019 , w32020 , w32021 , w32022 , w32023 , w32024 , w32025 , w32026 , w32027 , w32028 , w32029 , w32030 , w32031 , w32032 , w32033 , w32034 , w32035 , w32036 , w32037 , w32038 , w32039 , w32040 , w32041 , w32042 , w32043 , w32044 , w32045 , w32046 , w32047 , w32048 , w32049 , w32050 , w32051 , w32052 , w32053 , w32054 , w32055 , w32056 , w32057 , w32058 , w32059 , w32060 , w32061 , w32062 , w32063 , w32064 , w32065 , w32066 , w32067 , w32068 , w32069 , w32070 , w32071 , w32072 , w32073 , w32074 , w32075 , w32076 , w32077 , w32078 , w32079 , w32080 , w32081 , w32082 , w32083 , w32084 , w32085 , w32086 , w32087 , w32088 , w32089 , w32090 , w32091 , w32092 , w32093 , w32094 , w32095 , w32096 , w32097 , w32098 , w32099 , w32100 , w32101 , w32102 , w32103 , w32104 , w32105 , w32106 , w32107 , w32108 , w32109 , w32110 , w32111 , w32112 , w32113 , w32114 , w32115 , w32116 , w32117 , w32118 , w32119 , w32120 , w32121 , w32122 , w32123 , w32124 , w32125 , w32126 , w32127 , w32128 , w32129 , w32130 , w32131 , w32132 , w32133 , w32134 , w32135 , w32136 , w32137 , w32138 , w32139 , w32140 , w32141 , w32142 , w32143 , w32144 , w32145 , w32146 , w32147 , w32148 , w32149 , w32150 , w32151 , w32152 , w32153 , w32154 , w32155 , w32156 , w32157 , w32158 , w32159 , w32160 , w32161 , w32162 , w32163 , w32164 , w32165 , w32166 , w32167 , w32168 , w32169 , w32170 , w32171 , w32172 , w32173 , w32174 , w32175 , w32176 , w32177 , w32178 , w32179 , w32180 , w32181 , w32182 , w32183 , w32184 , w32185 , w32186 , w32187 , w32188 , w32189 , w32190 , w32191 , w32192 , w32193 , w32194 , w32195 , w32196 , w32197 , w32198 , w32199 , w32200 , w32201 , w32202 , w32203 , w32204 , w32205 , w32206 , w32207 , w32208 , w32209 , w32210 , w32211 , w32212 , w32213 , w32214 , w32215 , w32216 , w32217 , w32218 , w32219 , w32220 , w32221 , w32222 , w32223 , w32224 , w32225 , w32226 , w32227 , w32228 , w32229 , w32230 , w32231 , w32232 , w32233 , w32234 , w32235 , w32236 , w32237 , w32238 , w32239 , w32240 , w32241 , w32242 , w32243 , w32244 , w32245 , w32246 , w32247 , w32248 , w32249 , w32250 , w32251 , w32252 , w32253 , w32254 , w32255 , w32256 , w32257 , w32258 , w32259 , w32260 , w32261 , w32262 , w32263 , w32264 , w32265 , w32266 , w32267 , w32268 , w32269 , w32270 , w32271 , w32272 , w32273 , w32274 , w32275 , w32276 , w32277 , w32278 , w32279 , w32280 , w32281 , w32282 , w32283 , w32284 , w32285 , w32286 , w32287 , w32288 , w32289 , w32290 , w32291 , w32292 , w32293 , w32294 , w32295 , w32296 , w32297 , w32298 , w32299 , w32300 , w32301 , w32302 , w32303 , w32304 , w32305 , w32306 , w32307 , w32308 , w32309 , w32310 , w32311 , w32312 , w32313 , w32314 , w32315 , w32316 , w32317 , w32318 , w32319 , w32320 , w32321 , w32322 , w32323 , w32324 , w32325 , w32326 , w32327 , w32328 , w32329 , w32330 , w32331 , w32332 , w32333 , w32334 , w32335 , w32336 , w32337 , w32338 , w32339 , w32340 , w32341 , w32342 , w32343 , w32344 , w32345 , w32346 , w32347 , w32348 , w32349 , w32350 , w32351 , w32352 , w32353 , w32354 , w32355 , w32356 , w32357 , w32358 , w32359 , w32360 , w32361 , w32362 , w32363 , w32364 , w32365 , w32366 , w32367 , w32368 , w32369 , w32370 , w32371 , w32372 , w32373 , w32374 , w32375 , w32376 , w32377 , w32378 , w32379 , w32380 , w32381 , w32382 , w32383 , w32384 , w32385 , w32386 , w32387 , w32388 , w32389 , w32390 , w32391 , w32392 , w32393 , w32394 , w32395 , w32396 , w32397 , w32398 , w32399 , w32400 , w32401 , w32402 , w32403 , w32404 , w32405 , w32406 , w32407 , w32408 , w32409 , w32410 , w32411 , w32412 , w32413 , w32414 , w32415 , w32416 , w32417 , w32418 , w32419 , w32420 , w32421 , w32422 , w32423 , w32424 , w32425 , w32426 , w32427 , w32428 , w32429 , w32430 , w32431 , w32432 , w32433 , w32434 , w32435 , w32436 , w32437 , w32438 , w32439 , w32440 , w32441 , w32442 , w32443 , w32444 , w32445 , w32446 , w32447 , w32448 , w32449 , w32450 , w32451 , w32452 , w32453 , w32454 , w32455 , w32456 , w32457 , w32458 , w32459 , w32460 , w32461 , w32462 , w32463 , w32464 , w32465 , w32466 , w32467 , w32468 , w32469 , w32470 , w32471 , w32472 , w32473 , w32474 , w32475 , w32476 , w32477 , w32478 , w32479 , w32480 , w32481 , w32482 , w32483 , w32484 , w32485 , w32486 , w32487 , w32488 , w32489 , w32490 , w32491 , w32492 , w32493 , w32494 , w32495 , w32496 , w32497 , w32498 , w32499 , w32500 , w32501 , w32502 , w32503 , w32504 , w32505 , w32506 , w32507 , w32508 , w32509 , w32510 , w32511 , w32512 , w32513 , w32514 , w32515 , w32516 , w32517 , w32518 , w32519 , w32520 , w32521 , w32522 , w32523 , w32524 , w32525 , w32526 , w32527 , w32528 , w32529 , w32530 , w32531 , w32532 , w32533 , w32534 , w32535 , w32536 , w32537 , w32538 , w32539 , w32540 , w32541 , w32542 , w32543 , w32544 , w32545 , w32546 , w32547 , w32548 , w32549 , w32550 , w32551 , w32552 , w32553 , w32554 , w32555 , w32556 , w32557 , w32558 , w32559 , w32560 , w32561 , w32562 , w32563 , w32564 , w32565 , w32566 , w32567 , w32568 , w32569 , w32570 , w32571 , w32572 , w32573 , w32574 , w32575 , w32576 , w32577 , w32578 , w32579 , w32580 , w32581 , w32582 , w32583 , w32584 , w32585 , w32586 , w32587 , w32588 , w32589 , w32590 , w32591 , w32592 , w32593 , w32594 , w32595 , w32596 , w32597 , w32598 , w32599 , w32600 , w32601 , w32602 , w32603 , w32604 , w32605 , w32606 , w32607 , w32608 , w32609 , w32610 , w32611 , w32612 , w32613 , w32614 , w32615 , w32616 , w32617 , w32618 , w32619 , w32620 , w32621 , w32622 , w32623 , w32624 , w32625 , w32626 , w32627 , w32628 , w32629 , w32630 , w32631 , w32632 , w32633 , w32634 , w32635 , w32636 , w32637 , w32638 , w32639 , w32640 , w32641 , w32642 , w32643 , w32644 , w32645 , w32646 , w32647 , w32648 , w32649 , w32650 , w32651 , w32652 , w32653 , w32654 , w32655 , w32656 , w32657 , w32658 , w32659 , w32660 , w32661 , w32662 , w32663 , w32664 , w32665 , w32666 , w32667 , w32668 , w32669 , w32670 , w32671 , w32672 , w32673 , w32674 , w32675 , w32676 , w32677 , w32678 , w32679 , w32680 , w32681 , w32682 , w32683 , w32684 , w32685 , w32686 , w32687 , w32688 , w32689 , w32690 , w32691 , w32692 , w32693 , w32694 , w32695 , w32696 , w32697 , w32698 , w32699 , w32700 , w32701 , w32702 , w32703 , w32704 , w32705 , w32706 , w32707 , w32708 , w32709 , w32710 , w32711 , w32712 , w32713 , w32714 , w32715 , w32716 , w32717 , w32718 , w32719 , w32720 , w32721 , w32722 , w32723 , w32724 , w32725 , w32726 , w32727 , w32728 , w32729 , w32730 , w32731 , w32732 , w32733 , w32734 , w32735 , w32736 , w32737 , w32738 , w32739 , w32740 , w32741 , w32742 , w32743 , w32744 , w32745 , w32746 , w32747 , w32748 , w32749 , w32750 , w32751 , w32752 , w32753 , w32754 , w32755 , w32756 , w32757 , w32758 , w32759 , w32760 , w32761 , w32762 , w32763 , w32764 , w32765 , w32766 , w32767 , w32768 , w32769 , w32770 , w32771 , w32772 , w32773 , w32774 , w32775 , w32776 , w32777 , w32778 , w32779 , w32780 , w32781 , w32782 , w32783 , w32784 , w32785 , w32786 , w32787 , w32788 , w32789 , w32790 , w32791 , w32792 , w32793 , w32794 , w32795 , w32796 , w32797 , w32798 , w32799 , w32800 , w32801 , w32802 , w32803 , w32804 , w32805 , w32806 , w32807 , w32808 , w32809 , w32810 , w32811 , w32812 , w32813 , w32814 , w32815 , w32816 , w32817 , w32818 , w32819 , w32820 , w32821 , w32822 , w32823 , w32824 , w32825 , w32826 , w32827 , w32828 , w32829 , w32830 , w32831 , w32832 , w32833 , w32834 , w32835 , w32836 , w32837 , w32838 , w32839 , w32840 , w32841 , w32842 , w32843 , w32844 , w32845 , w32846 , w32847 , w32848 , w32849 , w32850 , w32851 , w32852 , w32853 , w32854 , w32855 , w32856 , w32857 , w32858 , w32859 , w32860 , w32861 , w32862 , w32863 , w32864 , w32865 , w32866 , w32867 , w32868 , w32869 , w32870 , w32871 , w32872 , w32873 , w32874 , w32875 , w32876 , w32877 , w32878 , w32879 , w32880 , w32881 , w32882 , w32883 , w32884 , w32885 , w32886 , w32887 , w32888 , w32889 , w32890 , w32891 , w32892 , w32893 , w32894 , w32895 , w32896 , w32897 , w32898 , w32899 , w32900 , w32901 , w32902 , w32903 , w32904 , w32905 , w32906 , w32907 , w32908 , w32909 , w32910 , w32911 , w32912 , w32913 , w32914 , w32915 , w32916 , w32917 , w32918 , w32919 , w32920 , w32921 , w32922 , w32923 , w32924 , w32925 , w32926 , w32927 , w32928 , w32929 , w32930 , w32931 , w32932 , w32933 , w32934 , w32935 , w32936 , w32937 , w32938 , w32939 , w32940 , w32941 , w32942 , w32943 , w32944 , w32945 , w32946 , w32947 , w32948 , w32949 , w32950 , w32951 , w32952 , w32953 , w32954 , w32955 , w32956 , w32957 , w32958 , w32959 , w32960 , w32961 , w32962 , w32963 , w32964 , w32965 , w32966 , w32967 , w32968 , w32969 , w32970 , w32971 , w32972 , w32973 , w32974 , w32975 , w32976 , w32977 , w32978 , w32979 , w32980 , w32981 , w32982 , w32983 , w32984 , w32985 , w32986 , w32987 , w32988 , w32989 , w32990 , w32991 , w32992 , w32993 , w32994 , w32995 , w32996 , w32997 , w32998 , w32999 , w33000 , w33001 , w33002 , w33003 , w33004 , w33005 , w33006 , w33007 , w33008 , w33009 , w33010 , w33011 , w33012 , w33013 , w33014 , w33015 , w33016 , w33017 , w33018 , w33019 , w33020 , w33021 , w33022 , w33023 , w33024 , w33025 , w33026 , w33027 , w33028 , w33029 , w33030 , w33031 , w33032 , w33033 , w33034 , w33035 , w33036 , w33037 , w33038 , w33039 , w33040 , w33041 , w33042 , w33043 , w33044 , w33045 , w33046 , w33047 , w33048 , w33049 , w33050 , w33051 , w33052 , w33053 , w33054 , w33055 , w33056 , w33057 , w33058 , w33059 , w33060 , w33061 , w33062 , w33063 , w33064 , w33065 , w33066 , w33067 , w33068 , w33069 , w33070 , w33071 , w33072 , w33073 , w33074 , w33075 , w33076 , w33077 , w33078 , w33079 , w33080 , w33081 , w33082 , w33083 , w33084 , w33085 , w33086 , w33087 , w33088 , w33089 , w33090 , w33091 , w33092 , w33093 , w33094 , w33095 , w33096 , w33097 , w33098 , w33099 , w33100 , w33101 , w33102 , w33103 , w33104 , w33105 , w33106 , w33107 , w33108 , w33109 , w33110 , w33111 , w33112 , w33113 , w33114 , w33115 , w33116 , w33117 , w33118 , w33119 , w33120 , w33121 , w33122 , w33123 , w33124 , w33125 , w33126 , w33127 , w33128 , w33129 , w33130 , w33131 , w33132 , w33133 , w33134 , w33135 , w33136 , w33137 , w33138 , w33139 , w33140 , w33141 , w33142 , w33143 , w33144 , w33145 , w33146 , w33147 , w33148 , w33149 , w33150 , w33151 , w33152 , w33153 , w33154 , w33155 , w33156 , w33157 , w33158 , w33159 , w33160 , w33161 , w33162 , w33163 , w33164 , w33165 , w33166 , w33167 , w33168 , w33169 , w33170 , w33171 , w33172 , w33173 , w33174 , w33175 , w33176 , w33177 , w33178 , w33179 , w33180 , w33181 , w33182 , w33183 , w33184 , w33185 , w33186 , w33187 , w33188 , w33189 , w33190 , w33191 , w33192 , w33193 , w33194 , w33195 , w33196 , w33197 , w33198 , w33199 , w33200 , w33201 , w33202 , w33203 , w33204 , w33205 , w33206 , w33207 , w33208 , w33209 , w33210 , w33211 , w33212 , w33213 , w33214 , w33215 , w33216 , w33217 , w33218 , w33219 , w33220 , w33221 , w33222 , w33223 , w33224 , w33225 , w33226 , w33227 , w33228 , w33229 , w33230 , w33231 , w33232 , w33233 , w33234 , w33235 , w33236 , w33237 , w33238 , w33239 , w33240 , w33241 , w33242 , w33243 , w33244 , w33245 , w33246 , w33247 , w33248 , w33249 , w33250 , w33251 , w33252 , w33253 , w33254 , w33255 , w33256 , w33257 , w33258 , w33259 , w33260 , w33261 , w33262 , w33263 , w33264 , w33265 , w33266 , w33267 , w33268 , w33269 , w33270 , w33271 , w33272 , w33273 , w33274 , w33275 , w33276 , w33277 , w33278 , w33279 , w33280 , w33281 , w33282 , w33283 , w33284 , w33285 , w33286 , w33287 , w33288 , w33289 , w33290 , w33291 , w33292 , w33293 , w33294 , w33295 , w33296 , w33297 , w33298 , w33299 , w33300 , w33301 , w33302 , w33303 , w33304 , w33305 , w33306 , w33307 , w33308 , w33309 , w33310 , w33311 , w33312 , w33313 , w33314 , w33315 , w33316 , w33317 , w33318 , w33319 , w33320 , w33321 , w33322 , w33323 , w33324 , w33325 , w33326 , w33327 , w33328 , w33329 , w33330 , w33331 , w33332 , w33333 , w33334 , w33335 , w33336 , w33337 , w33338 , w33339 , w33340 , w33341 , w33342 , w33343 , w33344 , w33345 , w33346 , w33347 , w33348 , w33349 , w33350 , w33351 , w33352 , w33353 , w33354 , w33355 , w33356 , w33357 , w33358 , w33359 , w33360 , w33361 , w33362 , w33363 , w33364 , w33365 , w33366 , w33367 , w33368 , w33369 , w33370 , w33371 , w33372 , w33373 , w33374 , w33375 , w33376 , w33377 , w33378 , w33379 , w33380 , w33381 , w33382 , w33383 , w33384 , w33385 , w33386 , w33387 , w33388 , w33389 , w33390 , w33391 , w33392 , w33393 , w33394 , w33395 , w33396 , w33397 , w33398 , w33399 , w33400 , w33401 , w33402 , w33403 , w33404 , w33405 , w33406 , w33407 , w33408 , w33409 , w33410 , w33411 , w33412 , w33413 , w33414 , w33415 , w33416 , w33417 , w33418 , w33419 , w33420 , w33421 , w33422 , w33423 , w33424 , w33425 , w33426 , w33427 , w33428 , w33429 , w33430 , w33431 , w33432 , w33433 , w33434 , w33435 , w33436 , w33437 , w33438 , w33439 , w33440 , w33441 , w33442 , w33443 , w33444 , w33445 , w33446 , w33447 , w33448 , w33449 , w33450 , w33451 , w33452 , w33453 , w33454 , w33455 , w33456 , w33457 , w33458 , w33459 , w33460 , w33461 , w33462 , w33463 , w33464 , w33465 , w33466 , w33467 , w33468 , w33469 , w33470 , w33471 , w33472 , w33473 , w33474 , w33475 , w33476 , w33477 , w33478 , w33479 , w33480 , w33481 , w33482 , w33483 , w33484 , w33485 , w33486 , w33487 , w33488 , w33489 , w33490 , w33491 , w33492 , w33493 , w33494 , w33495 , w33496 , w33497 , w33498 , w33499 , w33500 , w33501 , w33502 , w33503 , w33504 , w33505 , w33506 , w33507 , w33508 , w33509 , w33510 , w33511 , w33512 , w33513 , w33514 , w33515 , w33516 , w33517 , w33518 , w33519 , w33520 , w33521 , w33522 , w33523 , w33524 , w33525 , w33526 , w33527 , w33528 , w33529 , w33530 , w33531 , w33532 , w33533 , w33534 , w33535 , w33536 , w33537 , w33538 , w33539 , w33540 , w33541 , w33542 , w33543 , w33544 , w33545 , w33546 , w33547 , w33548 , w33549 , w33550 , w33551 , w33552 , w33553 , w33554 , w33555 , w33556 , w33557 , w33558 , w33559 , w33560 , w33561 , w33562 , w33563 , w33564 , w33565 , w33566 , w33567 , w33568 , w33569 , w33570 , w33571 , w33572 , w33573 , w33574 , w33575 , w33576 , w33577 , w33578 , w33579 , w33580 , w33581 , w33582 , w33583 , w33584 , w33585 , w33586 , w33587 , w33588 , w33589 , w33590 , w33591 , w33592 , w33593 , w33594 , w33595 , w33596 , w33597 , w33598 , w33599 , w33600 , w33601 , w33602 , w33603 , w33604 , w33605 , w33606 , w33607 , w33608 , w33609 , w33610 , w33611 , w33612 , w33613 , w33614 , w33615 , w33616 , w33617 , w33618 , w33619 , w33620 , w33621 , w33622 , w33623 , w33624 , w33625 , w33626 , w33627 , w33628 , w33629 , w33630 , w33631 , w33632 , w33633 , w33634 , w33635 , w33636 , w33637 , w33638 , w33639 , w33640 , w33641 , w33642 , w33643 , w33644 , w33645 , w33646 , w33647 , w33648 , w33649 , w33650 , w33651 , w33652 , w33653 , w33654 , w33655 , w33656 , w33657 , w33658 , w33659 , w33660 , w33661 , w33662 , w33663 , w33664 , w33665 , w33666 , w33667 , w33668 , w33669 , w33670 , w33671 , w33672 , w33673 , w33674 , w33675 , w33676 , w33677 , w33678 , w33679 , w33680 , w33681 , w33682 , w33683 , w33684 , w33685 , w33686 , w33687 , w33688 , w33689 , w33690 , w33691 , w33692 , w33693 , w33694 , w33695 , w33696 , w33697 , w33698 , w33699 , w33700 , w33701 , w33702 , w33703 , w33704 , w33705 , w33706 , w33707 , w33708 , w33709 , w33710 , w33711 , w33712 , w33713 , w33714 , w33715 , w33716 , w33717 , w33718 , w33719 , w33720 , w33721 , w33722 , w33723 , w33724 , w33725 , w33726 , w33727 , w33728 , w33729 , w33730 , w33731 , w33732 , w33733 , w33734 , w33735 , w33736 , w33737 , w33738 , w33739 , w33740 , w33741 , w33742 , w33743 , w33744 , w33745 , w33746 , w33747 , w33748 , w33749 , w33750 , w33751 , w33752 , w33753 , w33754 , w33755 , w33756 , w33757 , w33758 , w33759 , w33760 , w33761 , w33762 , w33763 , w33764 , w33765 , w33766 , w33767 , w33768 , w33769 , w33770 , w33771 , w33772 , w33773 , w33774 , w33775 , w33776 , w33777 , w33778 , w33779 , w33780 , w33781 , w33782 , w33783 , w33784 , w33785 , w33786 , w33787 , w33788 , w33789 , w33790 , w33791 , w33792 , w33793 , w33794 , w33795 , w33796 , w33797 , w33798 , w33799 , w33800 , w33801 , w33802 , w33803 , w33804 , w33805 , w33806 , w33807 , w33808 , w33809 , w33810 , w33811 , w33812 , w33813 , w33814 , w33815 , w33816 , w33817 , w33818 , w33819 , w33820 , w33821 , w33822 , w33823 , w33824 , w33825 , w33826 , w33827 , w33828 , w33829 , w33830 , w33831 , w33832 , w33833 , w33834 , w33835 , w33836 , w33837 , w33838 , w33839 , w33840 , w33841 , w33842 , w33843 , w33844 , w33845 , w33846 , w33847 , w33848 , w33849 , w33850 , w33851 , w33852 , w33853 , w33854 , w33855 , w33856 , w33857 , w33858 , w33859 , w33860 , w33861 , w33862 , w33863 , w33864 , w33865 , w33866 , w33867 , w33868 , w33869 , w33870 , w33871 , w33872 , w33873 , w33874 , w33875 , w33876 , w33877 , w33878 , w33879 , w33880 , w33881 , w33882 , w33883 , w33884 , w33885 , w33886 , w33887 , w33888 , w33889 , w33890 , w33891 , w33892 , w33893 , w33894 , w33895 , w33896 , w33897 , w33898 , w33899 , w33900 , w33901 , w33902 , w33903 , w33904 , w33905 , w33906 , w33907 , w33908 , w33909 , w33910 , w33911 , w33912 , w33913 , w33914 , w33915 , w33916 , w33917 , w33918 , w33919 , w33920 , w33921 , w33922 , w33923 , w33924 , w33925 , w33926 , w33927 , w33928 , w33929 , w33930 , w33931 , w33932 , w33933 , w33934 , w33935 , w33936 , w33937 , w33938 , w33939 , w33940 , w33941 , w33942 , w33943 , w33944 , w33945 , w33946 , w33947 , w33948 , w33949 , w33950 , w33951 , w33952 , w33953 , w33954 , w33955 , w33956 , w33957 , w33958 , w33959 , w33960 , w33961 , w33962 , w33963 , w33964 , w33965 , w33966 , w33967 , w33968 , w33969 , w33970 , w33971 , w33972 , w33973 , w33974 , w33975 , w33976 , w33977 , w33978 , w33979 , w33980 , w33981 , w33982 , w33983 , w33984 , w33985 , w33986 , w33987 , w33988 , w33989 , w33990 , w33991 , w33992 , w33993 , w33994 , w33995 , w33996 , w33997 , w33998 , w33999 , w34000 , w34001 , w34002 , w34003 , w34004 , w34005 , w34006 , w34007 , w34008 , w34009 , w34010 , w34011 , w34012 , w34013 , w34014 , w34015 , w34016 , w34017 , w34018 , w34019 , w34020 , w34021 , w34022 , w34023 , w34024 , w34025 , w34026 , w34027 , w34028 , w34029 , w34030 , w34031 , w34032 , w34033 , w34034 , w34035 , w34036 , w34037 , w34038 , w34039 , w34040 , w34041 , w34042 , w34043 , w34044 , w34045 , w34046 , w34047 , w34048 , w34049 , w34050 , w34051 , w34052 , w34053 , w34054 , w34055 , w34056 , w34057 , w34058 , w34059 , w34060 , w34061 , w34062 , w34063 , w34064 , w34065 , w34066 , w34067 , w34068 , w34069 , w34070 , w34071 , w34072 , w34073 , w34074 , w34075 , w34076 , w34077 , w34078 , w34079 , w34080 , w34081 , w34082 , w34083 , w34084 , w34085 , w34086 , w34087 , w34088 , w34089 , w34090 , w34091 , w34092 , w34093 , w34094 , w34095 , w34096 , w34097 , w34098 , w34099 , w34100 , w34101 , w34102 , w34103 , w34104 , w34105 , w34106 , w34107 , w34108 , w34109 , w34110 , w34111 , w34112 , w34113 , w34114 , w34115 , w34116 , w34117 , w34118 , w34119 , w34120 , w34121 , w34122 , w34123 , w34124 , w34125 , w34126 , w34127 , w34128 , w34129 , w34130 , w34131 , w34132 , w34133 , w34134 , w34135 , w34136 , w34137 , w34138 , w34139 , w34140 , w34141 , w34142 , w34143 , w34144 , w34145 , w34146 , w34147 , w34148 , w34149 , w34150 , w34151 , w34152 , w34153 , w34154 , w34155 , w34156 , w34157 , w34158 , w34159 , w34160 , w34161 , w34162 , w34163 , w34164 , w34165 , w34166 , w34167 , w34168 , w34169 , w34170 , w34171 , w34172 , w34173 , w34174 , w34175 , w34176 , w34177 , w34178 , w34179 , w34180 , w34181 , w34182 , w34183 , w34184 , w34185 , w34186 , w34187 , w34188 , w34189 , w34190 , w34191 , w34192 , w34193 , w34194 , w34195 , w34196 , w34197 , w34198 , w34199 , w34200 , w34201 , w34202 , w34203 , w34204 , w34205 , w34206 , w34207 , w34208 , w34209 , w34210 , w34211 , w34212 , w34213 , w34214 , w34215 , w34216 , w34217 , w34218 , w34219 , w34220 , w34221 , w34222 , w34223 , w34224 , w34225 , w34226 , w34227 , w34228 , w34229 , w34230 , w34231 , w34232 , w34233 , w34234 , w34235 , w34236 , w34237 , w34238 , w34239 , w34240 , w34241 , w34242 , w34243 , w34244 , w34245 , w34246 , w34247 , w34248 , w34249 , w34250 , w34251 , w34252 , w34253 , w34254 , w34255 , w34256 , w34257 , w34258 , w34259 , w34260 , w34261 , w34262 , w34263 , w34264 , w34265 , w34266 , w34267 , w34268 , w34269 , w34270 , w34271 , w34272 , w34273 , w34274 , w34275 , w34276 , w34277 , w34278 , w34279 , w34280 , w34281 , w34282 , w34283 , w34284 , w34285 , w34286 , w34287 , w34288 , w34289 , w34290 , w34291 , w34292 , w34293 , w34294 , w34295 , w34296 , w34297 , w34298 , w34299 , w34300 , w34301 , w34302 , w34303 , w34304 , w34305 , w34306 , w34307 , w34308 , w34309 , w34310 , w34311 , w34312 , w34313 , w34314 , w34315 , w34316 , w34317 , w34318 , w34319 , w34320 , w34321 , w34322 , w34323 , w34324 , w34325 , w34326 , w34327 , w34328 , w34329 , w34330 , w34331 , w34332 , w34333 , w34334 , w34335 , w34336 , w34337 , w34338 , w34339 , w34340 , w34341 , w34342 , w34343 , w34344 , w34345 , w34346 , w34347 , w34348 , w34349 , w34350 , w34351 , w34352 , w34353 , w34354 , w34355 , w34356 , w34357 , w34358 , w34359 , w34360 , w34361 , w34362 , w34363 , w34364 , w34365 , w34366 , w34367 , w34368 , w34369 , w34370 , w34371 , w34372 , w34373 , w34374 , w34375 , w34376 , w34377 , w34378 , w34379 , w34380 , w34381 , w34382 , w34383 , w34384 , w34385 , w34386 , w34387 , w34388 , w34389 , w34390 , w34391 , w34392 , w34393 , w34394 , w34395 , w34396 , w34397 , w34398 , w34399 , w34400 , w34401 , w34402 , w34403 , w34404 , w34405 , w34406 , w34407 , w34408 , w34409 , w34410 , w34411 , w34412 , w34413 , w34414 , w34415 , w34416 , w34417 , w34418 , w34419 , w34420 , w34421 , w34422 , w34423 , w34424 , w34425 , w34426 , w34427 , w34428 , w34429 , w34430 , w34431 , w34432 , w34433 , w34434 , w34435 , w34436 , w34437 , w34438 , w34439 , w34440 , w34441 , w34442 , w34443 , w34444 , w34445 , w34446 , w34447 , w34448 , w34449 , w34450 , w34451 , w34452 , w34453 , w34454 , w34455 , w34456 , w34457 , w34458 , w34459 , w34460 , w34461 , w34462 , w34463 , w34464 , w34465 , w34466 , w34467 , w34468 , w34469 , w34470 , w34471 , w34472 , w34473 , w34474 , w34475 , w34476 , w34477 , w34478 , w34479 , w34480 , w34481 , w34482 , w34483 , w34484 , w34485 , w34486 , w34487 , w34488 , w34489 , w34490 , w34491 , w34492 , w34493 , w34494 , w34495 , w34496 , w34497 , w34498 , w34499 , w34500 , w34501 , w34502 , w34503 , w34504 , w34505 , w34506 , w34507 , w34508 , w34509 , w34510 , w34511 , w34512 , w34513 , w34514 , w34515 , w34516 , w34517 , w34518 , w34519 , w34520 , w34521 , w34522 , w34523 , w34524 , w34525 , w34526 , w34527 , w34528 , w34529 , w34530 , w34531 , w34532 , w34533 , w34534 , w34535 , w34536 , w34537 , w34538 , w34539 , w34540 , w34541 , w34542 , w34543 , w34544 , w34545 , w34546 , w34547 , w34548 , w34549 , w34550 , w34551 , w34552 , w34553 , w34554 , w34555 , w34556 , w34557 , w34558 , w34559 , w34560 , w34561 , w34562 , w34563 , w34564 , w34565 , w34566 , w34567 , w34568 , w34569 , w34570 , w34571 , w34572 , w34573 , w34574 , w34575 , w34576 , w34577 , w34578 , w34579 , w34580 , w34581 , w34582 , w34583 , w34584 , w34585 , w34586 , w34587 , w34588 , w34589 , w34590 , w34591 , w34592 , w34593 , w34594 , w34595 , w34596 , w34597 , w34598 , w34599 , w34600 , w34601 , w34602 , w34603 , w34604 , w34605 , w34606 , w34607 , w34608 , w34609 , w34610 , w34611 , w34612 , w34613 , w34614 , w34615 , w34616 , w34617 , w34618 , w34619 , w34620 , w34621 , w34622 , w34623 , w34624 , w34625 , w34626 , w34627 , w34628 , w34629 , w34630 , w34631 , w34632 , w34633 , w34634 , w34635 , w34636 , w34637 , w34638 , w34639 , w34640 , w34641 , w34642 , w34643 , w34644 , w34645 , w34646 , w34647 , w34648 , w34649 , w34650 , w34651 , w34652 , w34653 , w34654 , w34655 , w34656 , w34657 , w34658 , w34659 , w34660 , w34661 , w34662 , w34663 , w34664 , w34665 , w34666 , w34667 , w34668 , w34669 , w34670 , w34671 , w34672 , w34673 , w34674 , w34675 , w34676 , w34677 , w34678 , w34679 , w34680 , w34681 , w34682 , w34683 , w34684 , w34685 , w34686 , w34687 , w34688 , w34689 , w34690 , w34691 , w34692 , w34693 , w34694 , w34695 , w34696 , w34697 , w34698 , w34699 , w34700 , w34701 , w34702 , w34703 , w34704 , w34705 , w34706 , w34707 , w34708 , w34709 , w34710 , w34711 , w34712 , w34713 , w34714 , w34715 , w34716 , w34717 , w34718 , w34719 , w34720 , w34721 , w34722 , w34723 , w34724 , w34725 , w34726 , w34727 , w34728 , w34729 , w34730 , w34731 , w34732 , w34733 , w34734 , w34735 , w34736 , w34737 , w34738 , w34739 , w34740 , w34741 , w34742 , w34743 , w34744 , w34745 , w34746 , w34747 , w34748 , w34749 , w34750 , w34751 , w34752 , w34753 , w34754 , w34755 , w34756 , w34757 , w34758 , w34759 , w34760 , w34761 , w34762 , w34763 , w34764 , w34765 , w34766 , w34767 , w34768 , w34769 , w34770 , w34771 , w34772 , w34773 , w34774 , w34775 , w34776 , w34777 , w34778 , w34779 , w34780 , w34781 , w34782 , w34783 , w34784 , w34785 , w34786 , w34787 , w34788 , w34789 , w34790 , w34791 , w34792 , w34793 , w34794 , w34795 , w34796 , w34797 , w34798 , w34799 , w34800 , w34801 , w34802 , w34803 , w34804 , w34805 , w34806 , w34807 , w34808 , w34809 , w34810 , w34811 , w34812 , w34813 , w34814 , w34815 , w34816 , w34817 , w34818 , w34819 , w34820 , w34821 , w34822 , w34823 , w34824 , w34825 , w34826 , w34827 , w34828 , w34829 , w34830 , w34831 , w34832 , w34833 , w34834 , w34835 , w34836 , w34837 , w34838 , w34839 , w34840 , w34841 , w34842 , w34843 , w34844 , w34845 , w34846 , w34847 , w34848 , w34849 , w34850 , w34851 , w34852 , w34853 , w34854 , w34855 , w34856 , w34857 , w34858 , w34859 , w34860 , w34861 , w34862 , w34863 , w34864 , w34865 , w34866 , w34867 , w34868 , w34869 , w34870 , w34871 , w34872 , w34873 , w34874 , w34875 , w34876 , w34877 , w34878 , w34879 , w34880 , w34881 , w34882 , w34883 , w34884 , w34885 , w34886 , w34887 , w34888 , w34889 , w34890 , w34891 , w34892 , w34893 , w34894 , w34895 , w34896 , w34897 , w34898 , w34899 , w34900 , w34901 , w34902 , w34903 , w34904 , w34905 , w34906 , w34907 , w34908 , w34909 , w34910 , w34911 , w34912 , w34913 , w34914 , w34915 , w34916 , w34917 , w34918 , w34919 , w34920 , w34921 , w34922 , w34923 , w34924 , w34925 , w34926 , w34927 , w34928 , w34929 , w34930 , w34931 , w34932 , w34933 , w34934 , w34935 , w34936 , w34937 , w34938 , w34939 , w34940 , w34941 , w34942 , w34943 , w34944 , w34945 , w34946 , w34947 , w34948 , w34949 , w34950 , w34951 , w34952 , w34953 , w34954 , w34955 , w34956 , w34957 , w34958 , w34959 , w34960 , w34961 , w34962 , w34963 , w34964 , w34965 , w34966 , w34967 , w34968 , w34969 , w34970 , w34971 , w34972 , w34973 , w34974 , w34975 , w34976 , w34977 , w34978 , w34979 , w34980 , w34981 , w34982 , w34983 , w34984 , w34985 , w34986 , w34987 , w34988 , w34989 , w34990 , w34991 , w34992 , w34993 , w34994 , w34995 , w34996 , w34997 , w34998 , w34999 , w35000 , w35001 , w35002 , w35003 , w35004 , w35005 , w35006 , w35007 , w35008 , w35009 , w35010 , w35011 , w35012 , w35013 , w35014 , w35015 , w35016 , w35017 , w35018 , w35019 , w35020 , w35021 , w35022 , w35023 , w35024 , w35025 , w35026 , w35027 , w35028 , w35029 , w35030 , w35031 , w35032 , w35033 , w35034 , w35035 , w35036 , w35037 , w35038 , w35039 , w35040 , w35041 , w35042 , w35043 , w35044 , w35045 , w35046 , w35047 , w35048 , w35049 , w35050 , w35051 , w35052 , w35053 , w35054 , w35055 , w35056 , w35057 , w35058 , w35059 , w35060 , w35061 , w35062 , w35063 , w35064 , w35065 , w35066 , w35067 , w35068 , w35069 , w35070 , w35071 , w35072 , w35073 , w35074 , w35075 , w35076 , w35077 , w35078 , w35079 , w35080 , w35081 , w35082 , w35083 , w35084 , w35085 , w35086 , w35087 , w35088 , w35089 , w35090 , w35091 , w35092 , w35093 , w35094 , w35095 , w35096 , w35097 , w35098 , w35099 , w35100 , w35101 , w35102 , w35103 , w35104 , w35105 , w35106 , w35107 , w35108 , w35109 , w35110 , w35111 , w35112 , w35113 , w35114 , w35115 , w35116 , w35117 , w35118 , w35119 , w35120 , w35121 , w35122 , w35123 , w35124 , w35125 , w35126 , w35127 , w35128 , w35129 , w35130 , w35131 , w35132 , w35133 , w35134 , w35135 , w35136 , w35137 , w35138 , w35139 , w35140 , w35141 , w35142 , w35143 , w35144 , w35145 , w35146 , w35147 , w35148 , w35149 , w35150 , w35151 , w35152 , w35153 , w35154 , w35155 , w35156 , w35157 , w35158 , w35159 , w35160 , w35161 , w35162 , w35163 , w35164 , w35165 , w35166 , w35167 , w35168 , w35169 , w35170 , w35171 , w35172 , w35173 , w35174 , w35175 , w35176 , w35177 , w35178 , w35179 , w35180 , w35181 , w35182 , w35183 , w35184 , w35185 , w35186 , w35187 , w35188 , w35189 , w35190 , w35191 , w35192 , w35193 , w35194 , w35195 , w35196 , w35197 , w35198 , w35199 , w35200 , w35201 , w35202 , w35203 , w35204 , w35205 , w35206 , w35207 , w35208 , w35209 , w35210 , w35211 , w35212 , w35213 , w35214 , w35215 , w35216 , w35217 , w35218 , w35219 , w35220 , w35221 , w35222 , w35223 , w35224 , w35225 , w35226 , w35227 , w35228 , w35229 , w35230 , w35231 , w35232 , w35233 , w35234 , w35235 , w35236 , w35237 , w35238 , w35239 , w35240 , w35241 , w35242 , w35243 , w35244 , w35245 , w35246 , w35247 , w35248 , w35249 , w35250 , w35251 , w35252 , w35253 , w35254 , w35255 , w35256 , w35257 , w35258 , w35259 , w35260 , w35261 , w35262 , w35263 , w35264 , w35265 , w35266 , w35267 , w35268 , w35269 , w35270 , w35271 , w35272 , w35273 , w35274 , w35275 , w35276 , w35277 , w35278 , w35279 , w35280 , w35281 , w35282 , w35283 , w35284 , w35285 , w35286 , w35287 , w35288 , w35289 , w35290 , w35291 , w35292 , w35293 , w35294 , w35295 , w35296 , w35297 , w35298 , w35299 , w35300 , w35301 , w35302 , w35303 , w35304 , w35305 , w35306 , w35307 , w35308 , w35309 , w35310 , w35311 , w35312 , w35313 , w35314 , w35315 , w35316 , w35317 , w35318 , w35319 , w35320 , w35321 , w35322 , w35323 , w35324 , w35325 , w35326 , w35327 , w35328 , w35329 , w35330 , w35331 , w35332 , w35333 , w35334 , w35335 , w35336 , w35337 , w35338 , w35339 , w35340 , w35341 , w35342 , w35343 , w35344 , w35345 , w35346 , w35347 , w35348 , w35349 , w35350 , w35351 , w35352 , w35353 , w35354 , w35355 , w35356 , w35357 , w35358 , w35359 , w35360 , w35361 , w35362 , w35363 , w35364 , w35365 , w35366 , w35367 , w35368 , w35369 , w35370 , w35371 , w35372 , w35373 , w35374 , w35375 , w35376 , w35377 , w35378 , w35379 , w35380 , w35381 , w35382 , w35383 , w35384 , w35385 , w35386 , w35387 , w35388 , w35389 , w35390 , w35391 , w35392 , w35393 , w35394 , w35395 , w35396 , w35397 , w35398 , w35399 , w35400 , w35401 , w35402 , w35403 , w35404 , w35405 , w35406 , w35407 , w35408 , w35409 , w35410 , w35411 , w35412 , w35413 , w35414 , w35415 , w35416 , w35417 , w35418 , w35419 , w35420 , w35421 , w35422 , w35423 , w35424 , w35425 , w35426 , w35427 , w35428 , w35429 , w35430 , w35431 , w35432 , w35433 , w35434 , w35435 , w35436 , w35437 , w35438 , w35439 , w35440 , w35441 , w35442 , w35443 , w35444 , w35445 , w35446 , w35447 , w35448 , w35449 , w35450 , w35451 , w35452 , w35453 , w35454 , w35455 , w35456 , w35457 , w35458 , w35459 , w35460 , w35461 , w35462 , w35463 , w35464 , w35465 , w35466 , w35467 , w35468 , w35469 , w35470 , w35471 , w35472 , w35473 , w35474 , w35475 , w35476 , w35477 , w35478 , w35479 , w35480 , w35481 , w35482 , w35483 , w35484 , w35485 , w35486 , w35487 , w35488 , w35489 , w35490 , w35491 , w35492 , w35493 , w35494 , w35495 , w35496 , w35497 , w35498 , w35499 , w35500 , w35501 , w35502 , w35503 , w35504 , w35505 , w35506 , w35507 , w35508 , w35509 , w35510 , w35511 , w35512 , w35513 , w35514 , w35515 , w35516 , w35517 , w35518 , w35519 , w35520 , w35521 , w35522 , w35523 , w35524 , w35525 , w35526 , w35527 , w35528 , w35529 , w35530 , w35531 , w35532 , w35533 , w35534 , w35535 , w35536 , w35537 , w35538 , w35539 , w35540 , w35541 , w35542 , w35543 , w35544 , w35545 , w35546 , w35547 , w35548 , w35549 , w35550 , w35551 , w35552 , w35553 , w35554 , w35555 , w35556 , w35557 , w35558 , w35559 , w35560 , w35561 , w35562 , w35563 , w35564 , w35565 , w35566 , w35567 , w35568 , w35569 , w35570 , w35571 , w35572 , w35573 , w35574 , w35575 , w35576 , w35577 , w35578 , w35579 , w35580 , w35581 , w35582 , w35583 , w35584 , w35585 , w35586 , w35587 , w35588 , w35589 , w35590 , w35591 , w35592 , w35593 , w35594 , w35595 , w35596 , w35597 , w35598 , w35599 , w35600 , w35601 , w35602 , w35603 , w35604 , w35605 , w35606 , w35607 , w35608 , w35609 , w35610 , w35611 , w35612 , w35613 , w35614 , w35615 , w35616 , w35617 , w35618 , w35619 , w35620 , w35621 , w35622 , w35623 , w35624 , w35625 , w35626 , w35627 , w35628 , w35629 , w35630 , w35631 , w35632 , w35633 , w35634 , w35635 , w35636 , w35637 , w35638 , w35639 , w35640 , w35641 , w35642 , w35643 , w35644 , w35645 , w35646 , w35647 , w35648 , w35649 , w35650 , w35651 , w35652 , w35653 , w35654 , w35655 , w35656 , w35657 , w35658 , w35659 , w35660 , w35661 , w35662 , w35663 , w35664 , w35665 , w35666 , w35667 , w35668 , w35669 , w35670 , w35671 , w35672 , w35673 , w35674 , w35675 , w35676 , w35677 , w35678 , w35679 , w35680 , w35681 , w35682 , w35683 , w35684 , w35685 , w35686 , w35687 , w35688 , w35689 , w35690 , w35691 , w35692 , w35693 , w35694 , w35695 , w35696 , w35697 , w35698 , w35699 , w35700 , w35701 , w35702 , w35703 , w35704 , w35705 , w35706 , w35707 , w35708 , w35709 , w35710 , w35711 , w35712 , w35713 , w35714 , w35715 , w35716 , w35717 , w35718 , w35719 , w35720 , w35721 , w35722 , w35723 , w35724 , w35725 , w35726 , w35727 , w35728 , w35729 , w35730 , w35731 , w35732 , w35733 , w35734 , w35735 , w35736 , w35737 , w35738 , w35739 , w35740 , w35741 , w35742 , w35743 , w35744 , w35745 , w35746 , w35747 , w35748 , w35749 , w35750 , w35751 , w35752 , w35753 , w35754 , w35755 , w35756 , w35757 , w35758 , w35759 , w35760 , w35761 , w35762 , w35763 , w35764 , w35765 , w35766 , w35767 , w35768 , w35769 , w35770 , w35771 , w35772 , w35773 , w35774 , w35775 , w35776 , w35777 , w35778 , w35779 , w35780 , w35781 , w35782 , w35783 , w35784 , w35785 , w35786 , w35787 , w35788 , w35789 , w35790 , w35791 , w35792 , w35793 , w35794 , w35795 , w35796 , w35797 , w35798 , w35799 , w35800 , w35801 , w35802 , w35803 , w35804 , w35805 , w35806 , w35807 , w35808 , w35809 , w35810 , w35811 , w35812 , w35813 , w35814 , w35815 , w35816 , w35817 , w35818 , w35819 , w35820 , w35821 , w35822 , w35823 , w35824 , w35825 , w35826 , w35827 , w35828 , w35829 , w35830 , w35831 , w35832 , w35833 , w35834 , w35835 , w35836 , w35837 , w35838 , w35839 , w35840 , w35841 , w35842 , w35843 , w35844 , w35845 , w35846 , w35847 , w35848 , w35849 , w35850 , w35851 , w35852 , w35853 , w35854 , w35855 , w35856 , w35857 , w35858 , w35859 , w35860 , w35861 , w35862 , w35863 , w35864 , w35865 , w35866 , w35867 , w35868 , w35869 , w35870 , w35871 , w35872 , w35873 , w35874 , w35875 , w35876 , w35877 , w35878 , w35879 , w35880 , w35881 , w35882 , w35883 , w35884 , w35885 , w35886 , w35887 , w35888 , w35889 , w35890 , w35891 , w35892 , w35893 , w35894 , w35895 , w35896 , w35897 , w35898 , w35899 , w35900 , w35901 , w35902 , w35903 , w35904 , w35905 , w35906 , w35907 , w35908 , w35909 , w35910 , w35911 , w35912 , w35913 , w35914 , w35915 , w35916 , w35917 , w35918 , w35919 , w35920 , w35921 , w35922 , w35923 , w35924 , w35925 , w35926 , w35927 , w35928 , w35929 , w35930 , w35931 , w35932 , w35933 , w35934 , w35935 , w35936 , w35937 , w35938 , w35939 , w35940 , w35941 , w35942 , w35943 , w35944 , w35945 , w35946 , w35947 , w35948 , w35949 , w35950 , w35951 , w35952 , w35953 , w35954 , w35955 , w35956 , w35957 , w35958 , w35959 , w35960 , w35961 , w35962 , w35963 , w35964 , w35965 , w35966 , w35967 , w35968 , w35969 , w35970 , w35971 , w35972 , w35973 , w35974 , w35975 , w35976 , w35977 , w35978 , w35979 , w35980 , w35981 , w35982 , w35983 , w35984 , w35985 , w35986 , w35987 , w35988 , w35989 , w35990 , w35991 , w35992 , w35993 , w35994 , w35995 , w35996 , w35997 , w35998 , w35999 , w36000 , w36001 , w36002 , w36003 , w36004 , w36005 , w36006 , w36007 , w36008 , w36009 , w36010 , w36011 , w36012 , w36013 , w36014 , w36015 , w36016 , w36017 , w36018 , w36019 , w36020 , w36021 , w36022 , w36023 , w36024 , w36025 , w36026 , w36027 , w36028 , w36029 , w36030 , w36031 , w36032 , w36033 , w36034 , w36035 , w36036 , w36037 , w36038 , w36039 , w36040 , w36041 , w36042 , w36043 , w36044 , w36045 , w36046 , w36047 , w36048 , w36049 , w36050 , w36051 , w36052 , w36053 , w36054 , w36055 , w36056 , w36057 , w36058 , w36059 , w36060 , w36061 , w36062 , w36063 , w36064 , w36065 , w36066 , w36067 , w36068 , w36069 , w36070 , w36071 , w36072 , w36073 , w36074 , w36075 , w36076 , w36077 , w36078 , w36079 , w36080 , w36081 , w36082 , w36083 , w36084 , w36085 , w36086 , w36087 , w36088 , w36089 , w36090 , w36091 , w36092 , w36093 , w36094 , w36095 , w36096 , w36097 , w36098 , w36099 , w36100 , w36101 , w36102 , w36103 , w36104 , w36105 , w36106 , w36107 , w36108 , w36109 , w36110 , w36111 , w36112 , w36113 , w36114 , w36115 , w36116 , w36117 , w36118 , w36119 , w36120 , w36121 , w36122 , w36123 , w36124 , w36125 , w36126 , w36127 , w36128 , w36129 , w36130 , w36131 , w36132 , w36133 , w36134 , w36135 , w36136 , w36137 , w36138 , w36139 , w36140 , w36141 , w36142 , w36143 , w36144 , w36145 , w36146 , w36147 , w36148 , w36149 , w36150 , w36151 , w36152 , w36153 , w36154 , w36155 , w36156 , w36157 , w36158 , w36159 , w36160 , w36161 , w36162 , w36163 , w36164 , w36165 , w36166 , w36167 , w36168 , w36169 , w36170 , w36171 , w36172 , w36173 , w36174 , w36175 , w36176 , w36177 , w36178 , w36179 , w36180 , w36181 , w36182 , w36183 , w36184 , w36185 , w36186 , w36187 , w36188 , w36189 , w36190 , w36191 , w36192 , w36193 , w36194 , w36195 , w36196 , w36197 , w36198 , w36199 , w36200 , w36201 , w36202 , w36203 , w36204 , w36205 , w36206 , w36207 , w36208 , w36209 , w36210 , w36211 , w36212 , w36213 , w36214 , w36215 , w36216 , w36217 , w36218 , w36219 , w36220 , w36221 , w36222 , w36223 , w36224 , w36225 , w36226 , w36227 , w36228 , w36229 , w36230 , w36231 , w36232 , w36233 , w36234 , w36235 , w36236 , w36237 , w36238 , w36239 , w36240 , w36241 , w36242 , w36243 , w36244 , w36245 , w36246 , w36247 , w36248 , w36249 , w36250 , w36251 , w36252 , w36253 , w36254 , w36255 , w36256 , w36257 , w36258 , w36259 , w36260 , w36261 , w36262 , w36263 , w36264 , w36265 , w36266 , w36267 , w36268 , w36269 , w36270 , w36271 , w36272 , w36273 , w36274 , w36275 , w36276 , w36277 , w36278 , w36279 , w36280 , w36281 , w36282 , w36283 , w36284 , w36285 , w36286 , w36287 , w36288 , w36289 , w36290 , w36291 , w36292 , w36293 , w36294 , w36295 , w36296 , w36297 , w36298 , w36299 , w36300 , w36301 , w36302 , w36303 , w36304 , w36305 , w36306 , w36307 , w36308 , w36309 , w36310 , w36311 , w36312 , w36313 , w36314 , w36315 , w36316 , w36317 , w36318 , w36319 , w36320 , w36321 , w36322 , w36323 , w36324 , w36325 , w36326 , w36327 , w36328 , w36329 , w36330 , w36331 , w36332 , w36333 , w36334 , w36335 , w36336 , w36337 , w36338 , w36339 , w36340 , w36341 , w36342 , w36343 , w36344 , w36345 , w36346 , w36347 , w36348 , w36349 , w36350 , w36351 , w36352 , w36353 , w36354 , w36355 , w36356 , w36357 , w36358 , w36359 , w36360 , w36361 , w36362 , w36363 , w36364 , w36365 , w36366 , w36367 , w36368 , w36369 , w36370 , w36371 , w36372 , w36373 , w36374 , w36375 , w36376 , w36377 , w36378 , w36379 , w36380 , w36381 , w36382 , w36383 , w36384 , w36385 , w36386 , w36387 , w36388 , w36389 , w36390 , w36391 , w36392 , w36393 , w36394 , w36395 , w36396 , w36397 , w36398 , w36399 , w36400 , w36401 , w36402 , w36403 , w36404 , w36405 , w36406 , w36407 , w36408 , w36409 , w36410 , w36411 , w36412 , w36413 , w36414 , w36415 , w36416 , w36417 , w36418 , w36419 , w36420 , w36421 , w36422 , w36423 , w36424 , w36425 , w36426 , w36427 , w36428 , w36429 , w36430 , w36431 , w36432 , w36433 , w36434 , w36435 , w36436 , w36437 , w36438 , w36439 , w36440 , w36441 , w36442 , w36443 , w36444 , w36445 , w36446 , w36447 , w36448 , w36449 , w36450 , w36451 , w36452 , w36453 , w36454 , w36455 , w36456 , w36457 , w36458 , w36459 , w36460 , w36461 , w36462 , w36463 , w36464 , w36465 , w36466 , w36467 , w36468 , w36469 , w36470 , w36471 , w36472 , w36473 , w36474 , w36475 , w36476 , w36477 , w36478 , w36479 , w36480 , w36481 , w36482 , w36483 , w36484 , w36485 , w36486 , w36487 , w36488 , w36489 , w36490 , w36491 , w36492 , w36493 , w36494 , w36495 , w36496 , w36497 , w36498 , w36499 , w36500 , w36501 , w36502 , w36503 , w36504 , w36505 , w36506 , w36507 , w36508 , w36509 , w36510 , w36511 , w36512 , w36513 , w36514 , w36515 , w36516 , w36517 , w36518 , w36519 , w36520 , w36521 , w36522 , w36523 , w36524 , w36525 , w36526 , w36527 , w36528 , w36529 , w36530 , w36531 , w36532 , w36533 , w36534 , w36535 , w36536 , w36537 , w36538 , w36539 , w36540 , w36541 , w36542 , w36543 , w36544 , w36545 , w36546 , w36547 , w36548 , w36549 , w36550 , w36551 , w36552 , w36553 , w36554 , w36555 , w36556 , w36557 , w36558 , w36559 , w36560 , w36561 , w36562 , w36563 , w36564 , w36565 , w36566 , w36567 , w36568 , w36569 , w36570 , w36571 , w36572 , w36573 , w36574 , w36575 , w36576 , w36577 , w36578 , w36579 , w36580 , w36581 , w36582 , w36583 , w36584 , w36585 , w36586 , w36587 , w36588 , w36589 , w36590 , w36591 , w36592 , w36593 , w36594 , w36595 , w36596 , w36597 , w36598 , w36599 , w36600 , w36601 , w36602 , w36603 , w36604 , w36605 , w36606 , w36607 , w36608 , w36609 , w36610 , w36611 , w36612 , w36613 , w36614 , w36615 , w36616 , w36617 , w36618 , w36619 , w36620 , w36621 , w36622 , w36623 , w36624 , w36625 , w36626 , w36627 , w36628 , w36629 , w36630 , w36631 , w36632 , w36633 , w36634 , w36635 , w36636 , w36637 , w36638 , w36639 , w36640 , w36641 , w36642 , w36643 , w36644 , w36645 , w36646 , w36647 , w36648 , w36649 , w36650 , w36651 , w36652 , w36653 , w36654 , w36655 , w36656 , w36657 , w36658 , w36659 , w36660 , w36661 , w36662 , w36663 , w36664 , w36665 , w36666 , w36667 , w36668 , w36669 , w36670 , w36671 , w36672 , w36673 , w36674 , w36675 , w36676 , w36677 , w36678 , w36679 , w36680 , w36681 , w36682 , w36683 , w36684 , w36685 , w36686 , w36687 , w36688 , w36689 , w36690 , w36691 , w36692 , w36693 , w36694 , w36695 , w36696 , w36697 , w36698 , w36699 , w36700 , w36701 , w36702 , w36703 , w36704 , w36705 , w36706 , w36707 , w36708 , w36709 , w36710 , w36711 , w36712 , w36713 , w36714 , w36715 , w36716 , w36717 , w36718 , w36719 , w36720 , w36721 , w36722 , w36723 , w36724 , w36725 , w36726 , w36727 , w36728 , w36729 , w36730 , w36731 , w36732 , w36733 , w36734 , w36735 , w36736 , w36737 , w36738 , w36739 , w36740 , w36741 , w36742 , w36743 , w36744 , w36745 , w36746 , w36747 , w36748 , w36749 , w36750 , w36751 , w36752 , w36753 , w36754 , w36755 , w36756 , w36757 , w36758 , w36759 , w36760 , w36761 , w36762 , w36763 , w36764 , w36765 , w36766 , w36767 , w36768 , w36769 , w36770 , w36771 , w36772 , w36773 , w36774 , w36775 , w36776 , w36777 , w36778 , w36779 , w36780 , w36781 , w36782 , w36783 , w36784 , w36785 , w36786 , w36787 , w36788 , w36789 , w36790 , w36791 , w36792 , w36793 , w36794 , w36795 , w36796 , w36797 , w36798 , w36799 , w36800 , w36801 , w36802 , w36803 , w36804 , w36805 , w36806 , w36807 , w36808 , w36809 , w36810 , w36811 , w36812 , w36813 , w36814 , w36815 , w36816 , w36817 , w36818 , w36819 , w36820 , w36821 , w36822 , w36823 , w36824 , w36825 , w36826 , w36827 , w36828 , w36829 , w36830 , w36831 , w36832 , w36833 , w36834 , w36835 , w36836 , w36837 , w36838 , w36839 , w36840 , w36841 , w36842 , w36843 , w36844 , w36845 , w36846 , w36847 , w36848 , w36849 , w36850 , w36851 , w36852 , w36853 , w36854 , w36855 , w36856 , w36857 , w36858 , w36859 , w36860 , w36861 , w36862 , w36863 , w36864 , w36865 , w36866 , w36867 , w36868 , w36869 , w36870 , w36871 , w36872 , w36873 , w36874 , w36875 , w36876 , w36877 , w36878 , w36879 , w36880 , w36881 , w36882 , w36883 , w36884 , w36885 , w36886 , w36887 , w36888 , w36889 , w36890 , w36891 , w36892 , w36893 , w36894 , w36895 , w36896 , w36897 , w36898 , w36899 , w36900 , w36901 , w36902 , w36903 , w36904 , w36905 , w36906 , w36907 , w36908 , w36909 , w36910 , w36911 , w36912 , w36913 , w36914 , w36915 , w36916 , w36917 , w36918 , w36919 , w36920 , w36921 , w36922 , w36923 , w36924 , w36925 , w36926 , w36927 , w36928 , w36929 , w36930 , w36931 , w36932 , w36933 , w36934 , w36935 , w36936 , w36937 , w36938 , w36939 , w36940 , w36941 , w36942 , w36943 , w36944 , w36945 , w36946 , w36947 , w36948 , w36949 , w36950 , w36951 , w36952 , w36953 , w36954 , w36955 , w36956 , w36957 , w36958 , w36959 , w36960 , w36961 , w36962 , w36963 , w36964 , w36965 , w36966 , w36967 , w36968 , w36969 , w36970 , w36971 , w36972 , w36973 , w36974 , w36975 , w36976 , w36977 , w36978 , w36979 , w36980 , w36981 , w36982 , w36983 , w36984 , w36985 , w36986 , w36987 , w36988 , w36989 , w36990 , w36991 , w36992 , w36993 , w36994 , w36995 , w36996 , w36997 , w36998 , w36999 , w37000 , w37001 , w37002 , w37003 , w37004 , w37005 , w37006 , w37007 , w37008 , w37009 , w37010 , w37011 , w37012 , w37013 , w37014 , w37015 , w37016 , w37017 , w37018 , w37019 , w37020 , w37021 , w37022 , w37023 , w37024 , w37025 , w37026 , w37027 , w37028 , w37029 , w37030 , w37031 , w37032 , w37033 , w37034 , w37035 , w37036 , w37037 , w37038 , w37039 , w37040 , w37041 , w37042 , w37043 , w37044 , w37045 , w37046 , w37047 , w37048 , w37049 , w37050 , w37051 , w37052 , w37053 , w37054 , w37055 , w37056 , w37057 , w37058 , w37059 , w37060 , w37061 , w37062 , w37063 , w37064 , w37065 , w37066 , w37067 , w37068 , w37069 , w37070 , w37071 , w37072 , w37073 , w37074 , w37075 , w37076 , w37077 , w37078 , w37079 , w37080 , w37081 , w37082 , w37083 , w37084 , w37085 , w37086 , w37087 , w37088 , w37089 , w37090 , w37091 , w37092 , w37093 , w37094 , w37095 , w37096 , w37097 , w37098 , w37099 , w37100 , w37101 , w37102 , w37103 , w37104 , w37105 , w37106 , w37107 , w37108 , w37109 , w37110 , w37111 , w37112 , w37113 , w37114 , w37115 , w37116 , w37117 , w37118 , w37119 , w37120 , w37121 , w37122 , w37123 , w37124 , w37125 , w37126 , w37127 , w37128 , w37129 , w37130 , w37131 , w37132 , w37133 , w37134 , w37135 , w37136 , w37137 , w37138 , w37139 , w37140 , w37141 , w37142 , w37143 , w37144 , w37145 , w37146 , w37147 , w37148 , w37149 , w37150 , w37151 , w37152 , w37153 , w37154 , w37155 , w37156 , w37157 , w37158 , w37159 , w37160 , w37161 , w37162 , w37163 , w37164 , w37165 , w37166 , w37167 , w37168 , w37169 , w37170 , w37171 , w37172 , w37173 , w37174 , w37175 , w37176 , w37177 , w37178 , w37179 , w37180 , w37181 , w37182 , w37183 , w37184 , w37185 , w37186 , w37187 , w37188 , w37189 , w37190 , w37191 , w37192 , w37193 , w37194 , w37195 , w37196 , w37197 , w37198 , w37199 , w37200 , w37201 , w37202 , w37203 , w37204 , w37205 , w37206 , w37207 , w37208 , w37209 , w37210 , w37211 , w37212 , w37213 , w37214 , w37215 , w37216 , w37217 , w37218 , w37219 , w37220 , w37221 , w37222 , w37223 , w37224 , w37225 , w37226 , w37227 , w37228 , w37229 , w37230 , w37231 , w37232 , w37233 , w37234 , w37235 , w37236 , w37237 , w37238 , w37239 , w37240 , w37241 , w37242 , w37243 , w37244 , w37245 , w37246 , w37247 , w37248 , w37249 , w37250 , w37251 , w37252 , w37253 , w37254 , w37255 , w37256 , w37257 , w37258 , w37259 , w37260 , w37261 , w37262 , w37263 , w37264 , w37265 , w37266 , w37267 , w37268 , w37269 , w37270 , w37271 , w37272 , w37273 , w37274 , w37275 , w37276 , w37277 , w37278 , w37279 , w37280 , w37281 , w37282 , w37283 , w37284 , w37285 , w37286 , w37287 , w37288 , w37289 , w37290 , w37291 , w37292 , w37293 , w37294 , w37295 , w37296 , w37297 , w37298 , w37299 , w37300 , w37301 , w37302 , w37303 , w37304 , w37305 , w37306 , w37307 , w37308 , w37309 , w37310 , w37311 , w37312 , w37313 , w37314 , w37315 , w37316 , w37317 , w37318 , w37319 , w37320 , w37321 , w37322 , w37323 , w37324 , w37325 , w37326 , w37327 , w37328 , w37329 , w37330 , w37331 , w37332 , w37333 , w37334 , w37335 , w37336 , w37337 , w37338 , w37339 , w37340 , w37341 , w37342 , w37343 , w37344 , w37345 , w37346 , w37347 , w37348 , w37349 , w37350 , w37351 , w37352 , w37353 , w37354 , w37355 , w37356 , w37357 , w37358 , w37359 , w37360 , w37361 , w37362 , w37363 , w37364 , w37365 , w37366 , w37367 , w37368 , w37369 , w37370 , w37371 , w37372 , w37373 , w37374 , w37375 , w37376 , w37377 , w37378 , w37379 , w37380 , w37381 , w37382 , w37383 , w37384 , w37385 , w37386 , w37387 , w37388 , w37389 , w37390 , w37391 , w37392 , w37393 , w37394 , w37395 , w37396 , w37397 , w37398 , w37399 , w37400 , w37401 , w37402 , w37403 , w37404 , w37405 , w37406 , w37407 , w37408 , w37409 , w37410 , w37411 , w37412 , w37413 , w37414 , w37415 , w37416 , w37417 , w37418 , w37419 , w37420 , w37421 , w37422 , w37423 , w37424 , w37425 , w37426 , w37427 , w37428 , w37429 , w37430 , w37431 , w37432 , w37433 , w37434 , w37435 , w37436 , w37437 , w37438 , w37439 , w37440 , w37441 , w37442 , w37443 , w37444 , w37445 , w37446 , w37447 , w37448 , w37449 , w37450 , w37451 , w37452 , w37453 , w37454 , w37455 , w37456 , w37457 , w37458 , w37459 , w37460 , w37461 , w37462 , w37463 , w37464 , w37465 , w37466 , w37467 , w37468 , w37469 , w37470 , w37471 , w37472 , w37473 , w37474 , w37475 , w37476 , w37477 , w37478 , w37479 , w37480 , w37481 , w37482 , w37483 , w37484 , w37485 , w37486 , w37487 , w37488 , w37489 , w37490 , w37491 , w37492 , w37493 , w37494 , w37495 , w37496 , w37497 , w37498 , w37499 , w37500 , w37501 , w37502 , w37503 , w37504 , w37505 , w37506 , w37507 , w37508 , w37509 , w37510 , w37511 , w37512 , w37513 , w37514 , w37515 , w37516 , w37517 , w37518 , w37519 , w37520 , w37521 , w37522 , w37523 , w37524 , w37525 , w37526 , w37527 , w37528 , w37529 , w37530 , w37531 , w37532 , w37533 , w37534 , w37535 , w37536 , w37537 , w37538 , w37539 , w37540 , w37541 , w37542 , w37543 , w37544 , w37545 , w37546 , w37547 , w37548 , w37549 , w37550 , w37551 , w37552 , w37553 , w37554 , w37555 , w37556 , w37557 , w37558 , w37559 , w37560 , w37561 , w37562 , w37563 , w37564 , w37565 , w37566 , w37567 , w37568 , w37569 , w37570 , w37571 , w37572 , w37573 , w37574 , w37575 , w37576 , w37577 , w37578 , w37579 , w37580 , w37581 , w37582 , w37583 , w37584 , w37585 , w37586 , w37587 , w37588 , w37589 , w37590 , w37591 , w37592 , w37593 , w37594 , w37595 , w37596 , w37597 , w37598 , w37599 , w37600 , w37601 , w37602 , w37603 , w37604 , w37605 , w37606 , w37607 , w37608 , w37609 , w37610 , w37611 , w37612 , w37613 , w37614 , w37615 , w37616 , w37617 , w37618 , w37619 , w37620 , w37621 , w37622 , w37623 , w37624 , w37625 , w37626 , w37627 , w37628 , w37629 , w37630 , w37631 , w37632 , w37633 , w37634 , w37635 , w37636 , w37637 , w37638 , w37639 , w37640 , w37641 , w37642 , w37643 , w37644 , w37645 , w37646 , w37647 , w37648 , w37649 , w37650 , w37651 , w37652 , w37653 , w37654 , w37655 , w37656 , w37657 , w37658 , w37659 , w37660 , w37661 , w37662 , w37663 , w37664 , w37665 , w37666 , w37667 , w37668 , w37669 , w37670 , w37671 , w37672 , w37673 , w37674 , w37675 , w37676 , w37677 , w37678 , w37679 , w37680 , w37681 , w37682 , w37683 , w37684 , w37685 , w37686 , w37687 , w37688 , w37689 , w37690 , w37691 , w37692 , w37693 , w37694 , w37695 , w37696 , w37697 , w37698 , w37699 , w37700 , w37701 , w37702 , w37703 , w37704 , w37705 , w37706 , w37707 , w37708 , w37709 , w37710 , w37711 , w37712 , w37713 , w37714 , w37715 , w37716 , w37717 , w37718 , w37719 , w37720 , w37721 , w37722 , w37723 , w37724 , w37725 , w37726 , w37727 , w37728 , w37729 , w37730 , w37731 , w37732 , w37733 , w37734 , w37735 , w37736 , w37737 , w37738 , w37739 , w37740 , w37741 , w37742 , w37743 , w37744 , w37745 , w37746 , w37747 , w37748 , w37749 , w37750 , w37751 , w37752 , w37753 , w37754 , w37755 , w37756 , w37757 , w37758 , w37759 , w37760 , w37761 , w37762 , w37763 , w37764 , w37765 , w37766 , w37767 , w37768 , w37769 , w37770 , w37771 , w37772 , w37773 , w37774 , w37775 , w37776 , w37777 , w37778 , w37779 , w37780 , w37781 , w37782 , w37783 , w37784 , w37785 , w37786 , w37787 , w37788 , w37789 , w37790 , w37791 , w37792 , w37793 , w37794 , w37795 , w37796 , w37797 , w37798 , w37799 , w37800 , w37801 , w37802 , w37803 , w37804 , w37805 , w37806 , w37807 , w37808 , w37809 , w37810 , w37811 , w37812 , w37813 , w37814 , w37815 , w37816 , w37817 , w37818 , w37819 , w37820 , w37821 , w37822 , w37823 , w37824 , w37825 , w37826 , w37827 , w37828 , w37829 , w37830 , w37831 , w37832 , w37833 , w37834 , w37835 , w37836 , w37837 , w37838 , w37839 , w37840 , w37841 , w37842 , w37843 , w37844 , w37845 , w37846 , w37847 , w37848 , w37849 , w37850 , w37851 , w37852 , w37853 , w37854 , w37855 , w37856 , w37857 , w37858 , w37859 , w37860 , w37861 , w37862 , w37863 , w37864 , w37865 , w37866 , w37867 , w37868 , w37869 , w37870 , w37871 , w37872 , w37873 , w37874 , w37875 , w37876 , w37877 , w37878 , w37879 , w37880 , w37881 , w37882 , w37883 , w37884 , w37885 , w37886 , w37887 , w37888 , w37889 , w37890 , w37891 , w37892 , w37893 , w37894 , w37895 , w37896 , w37897 , w37898 , w37899 , w37900 , w37901 , w37902 , w37903 , w37904 , w37905 , w37906 , w37907 , w37908 , w37909 , w37910 , w37911 , w37912 , w37913 , w37914 , w37915 , w37916 , w37917 , w37918 , w37919 , w37920 , w37921 , w37922 , w37923 , w37924 , w37925 , w37926 , w37927 , w37928 , w37929 , w37930 , w37931 , w37932 , w37933 , w37934 , w37935 , w37936 , w37937 , w37938 , w37939 , w37940 , w37941 , w37942 , w37943 , w37944 , w37945 , w37946 , w37947 , w37948 , w37949 , w37950 , w37951 , w37952 , w37953 , w37954 , w37955 , w37956 , w37957 , w37958 , w37959 , w37960 , w37961 , w37962 , w37963 , w37964 , w37965 , w37966 , w37967 , w37968 , w37969 , w37970 , w37971 , w37972 , w37973 , w37974 , w37975 , w37976 , w37977 , w37978 , w37979 , w37980 , w37981 , w37982 , w37983 , w37984 , w37985 , w37986 , w37987 , w37988 , w37989 , w37990 , w37991 , w37992 , w37993 , w37994 , w37995 , w37996 , w37997 , w37998 , w37999 , w38000 , w38001 , w38002 , w38003 , w38004 , w38005 , w38006 , w38007 , w38008 , w38009 , w38010 , w38011 , w38012 , w38013 , w38014 , w38015 , w38016 , w38017 , w38018 , w38019 , w38020 , w38021 , w38022 , w38023 , w38024 , w38025 , w38026 , w38027 , w38028 , w38029 , w38030 , w38031 , w38032 , w38033 , w38034 , w38035 , w38036 , w38037 , w38038 , w38039 , w38040 , w38041 , w38042 , w38043 , w38044 , w38045 , w38046 , w38047 , w38048 , w38049 , w38050 , w38051 , w38052 , w38053 , w38054 , w38055 , w38056 , w38057 , w38058 , w38059 , w38060 , w38061 , w38062 , w38063 , w38064 , w38065 , w38066 , w38067 , w38068 , w38069 , w38070 , w38071 , w38072 , w38073 , w38074 , w38075 , w38076 , w38077 , w38078 , w38079 , w38080 , w38081 , w38082 , w38083 , w38084 , w38085 , w38086 , w38087 , w38088 , w38089 , w38090 , w38091 , w38092 , w38093 , w38094 , w38095 , w38096 , w38097 , w38098 , w38099 , w38100 , w38101 , w38102 , w38103 , w38104 , w38105 , w38106 , w38107 , w38108 , w38109 , w38110 , w38111 , w38112 , w38113 , w38114 , w38115 , w38116 , w38117 , w38118 , w38119 , w38120 , w38121 , w38122 , w38123 , w38124 , w38125 , w38126 , w38127 , w38128 , w38129 , w38130 , w38131 , w38132 , w38133 , w38134 , w38135 , w38136 , w38137 , w38138 , w38139 , w38140 , w38141 , w38142 , w38143 , w38144 , w38145 , w38146 , w38147 , w38148 , w38149 , w38150 , w38151 , w38152 , w38153 , w38154 , w38155 , w38156 , w38157 , w38158 , w38159 , w38160 , w38161 , w38162 , w38163 , w38164 , w38165 , w38166 , w38167 , w38168 , w38169 , w38170 , w38171 , w38172 , w38173 , w38174 , w38175 , w38176 , w38177 , w38178 , w38179 , w38180 , w38181 , w38182 , w38183 , w38184 , w38185 , w38186 , w38187 , w38188 , w38189 , w38190 , w38191 , w38192 , w38193 , w38194 , w38195 , w38196 , w38197 , w38198 , w38199 , w38200 , w38201 , w38202 , w38203 , w38204 , w38205 , w38206 , w38207 , w38208 , w38209 , w38210 , w38211 , w38212 , w38213 , w38214 , w38215 , w38216 , w38217 , w38218 , w38219 , w38220 , w38221 , w38222 , w38223 , w38224 , w38225 , w38226 , w38227 , w38228 , w38229 , w38230 , w38231 , w38232 , w38233 , w38234 , w38235 , w38236 , w38237 , w38238 , w38239 , w38240 , w38241 , w38242 , w38243 , w38244 , w38245 , w38246 , w38247 , w38248 , w38249 , w38250 , w38251 , w38252 , w38253 , w38254 , w38255 , w38256 , w38257 , w38258 , w38259 , w38260 , w38261 , w38262 , w38263 , w38264 , w38265 , w38266 , w38267 , w38268 , w38269 , w38270 , w38271 , w38272 , w38273 , w38274 , w38275 , w38276 , w38277 , w38278 , w38279 , w38280 , w38281 , w38282 , w38283 , w38284 , w38285 , w38286 , w38287 , w38288 , w38289 , w38290 , w38291 , w38292 , w38293 , w38294 , w38295 , w38296 , w38297 , w38298 , w38299 , w38300 , w38301 , w38302 , w38303 , w38304 , w38305 , w38306 , w38307 , w38308 , w38309 , w38310 , w38311 , w38312 , w38313 , w38314 , w38315 , w38316 , w38317 , w38318 , w38319 , w38320 , w38321 , w38322 , w38323 , w38324 , w38325 , w38326 , w38327 , w38328 , w38329 , w38330 , w38331 , w38332 , w38333 , w38334 , w38335 , w38336 , w38337 , w38338 , w38339 , w38340 , w38341 , w38342 , w38343 , w38344 , w38345 , w38346 , w38347 , w38348 , w38349 , w38350 , w38351 , w38352 , w38353 , w38354 , w38355 , w38356 , w38357 , w38358 , w38359 , w38360 , w38361 , w38362 , w38363 , w38364 , w38365 , w38366 , w38367 , w38368 , w38369 , w38370 , w38371 , w38372 , w38373 , w38374 , w38375 , w38376 , w38377 , w38378 , w38379 , w38380 , w38381 , w38382 , w38383 , w38384 , w38385 , w38386 , w38387 , w38388 , w38389 , w38390 , w38391 , w38392 , w38393 , w38394 , w38395 , w38396 , w38397 , w38398 , w38399 , w38400 , w38401 , w38402 , w38403 , w38404 , w38405 , w38406 , w38407 , w38408 , w38409 , w38410 , w38411 , w38412 , w38413 , w38414 , w38415 , w38416 , w38417 , w38418 , w38419 , w38420 , w38421 , w38422 , w38423 , w38424 , w38425 , w38426 , w38427 , w38428 , w38429 , w38430 , w38431 , w38432 , w38433 , w38434 , w38435 , w38436 , w38437 , w38438 , w38439 , w38440 , w38441 , w38442 , w38443 , w38444 , w38445 , w38446 , w38447 , w38448 , w38449 , w38450 , w38451 , w38452 , w38453 , w38454 , w38455 , w38456 , w38457 , w38458 , w38459 , w38460 , w38461 , w38462 , w38463 , w38464 , w38465 , w38466 , w38467 , w38468 , w38469 , w38470 , w38471 , w38472 , w38473 , w38474 , w38475 , w38476 , w38477 , w38478 , w38479 , w38480 , w38481 , w38482 , w38483 , w38484 , w38485 , w38486 , w38487 , w38488 , w38489 , w38490 , w38491 , w38492 , w38493 , w38494 , w38495 , w38496 , w38497 , w38498 , w38499 , w38500 , w38501 , w38502 , w38503 , w38504 , w38505 , w38506 , w38507 , w38508 , w38509 , w38510 , w38511 , w38512 , w38513 , w38514 , w38515 , w38516 , w38517 , w38518 , w38519 , w38520 , w38521 , w38522 , w38523 , w38524 , w38525 , w38526 , w38527 , w38528 , w38529 , w38530 , w38531 , w38532 , w38533 , w38534 , w38535 , w38536 , w38537 , w38538 , w38539 , w38540 , w38541 , w38542 , w38543 , w38544 , w38545 , w38546 , w38547 , w38548 , w38549 , w38550 , w38551 , w38552 , w38553 , w38554 , w38555 , w38556 , w38557 , w38558 , w38559 , w38560 , w38561 , w38562 , w38563 , w38564 , w38565 , w38566 , w38567 , w38568 , w38569 , w38570 , w38571 , w38572 , w38573 , w38574 , w38575 , w38576 , w38577 , w38578 , w38579 , w38580 , w38581 , w38582 , w38583 , w38584 , w38585 , w38586 , w38587 , w38588 , w38589 , w38590 , w38591 , w38592 , w38593 , w38594 , w38595 , w38596 , w38597 , w38598 , w38599 , w38600 , w38601 , w38602 , w38603 , w38604 , w38605 , w38606 , w38607 , w38608 , w38609 , w38610 , w38611 , w38612 , w38613 , w38614 , w38615 , w38616 , w38617 , w38618 , w38619 , w38620 , w38621 , w38622 , w38623 , w38624 , w38625 , w38626 , w38627 , w38628 , w38629 , w38630 , w38631 , w38632 , w38633 , w38634 , w38635 , w38636 , w38637 , w38638 , w38639 , w38640 , w38641 , w38642 , w38643 , w38644 , w38645 , w38646 , w38647 , w38648 , w38649 , w38650 , w38651 , w38652 , w38653 , w38654 , w38655 , w38656 , w38657 , w38658 , w38659 , w38660 , w38661 , w38662 , w38663 , w38664 , w38665 , w38666 , w38667 , w38668 , w38669 , w38670 , w38671 , w38672 , w38673 , w38674 , w38675 , w38676 , w38677 , w38678 , w38679 , w38680 , w38681 , w38682 , w38683 , w38684 , w38685 , w38686 , w38687 , w38688 , w38689 , w38690 , w38691 , w38692 , w38693 , w38694 , w38695 , w38696 , w38697 , w38698 , w38699 , w38700 , w38701 , w38702 , w38703 , w38704 , w38705 , w38706 , w38707 , w38708 , w38709 , w38710 , w38711 , w38712 , w38713 , w38714 , w38715 , w38716 , w38717 , w38718 , w38719 , w38720 , w38721 , w38722 , w38723 , w38724 , w38725 , w38726 , w38727 , w38728 , w38729 , w38730 , w38731 , w38732 , w38733 , w38734 , w38735 , w38736 , w38737 , w38738 , w38739 , w38740 , w38741 , w38742 , w38743 , w38744 , w38745 , w38746 , w38747 , w38748 , w38749 , w38750 , w38751 , w38752 , w38753 , w38754 , w38755 , w38756 , w38757 , w38758 , w38759 , w38760 , w38761 , w38762 , w38763 , w38764 , w38765 , w38766 , w38767 , w38768 , w38769 , w38770 , w38771 , w38772 , w38773 , w38774 , w38775 , w38776 , w38777 , w38778 , w38779 , w38780 , w38781 , w38782 , w38783 , w38784 , w38785 , w38786 , w38787 , w38788 , w38789 , w38790 , w38791 , w38792 , w38793 , w38794 , w38795 , w38796 , w38797 , w38798 , w38799 , w38800 , w38801 , w38802 , w38803 , w38804 , w38805 , w38806 , w38807 , w38808 , w38809 , w38810 , w38811 , w38812 , w38813 , w38814 , w38815 , w38816 , w38817 , w38818 , w38819 , w38820 , w38821 , w38822 , w38823 , w38824 , w38825 , w38826 , w38827 , w38828 , w38829 , w38830 , w38831 , w38832 , w38833 , w38834 , w38835 , w38836 , w38837 , w38838 , w38839 , w38840 , w38841 , w38842 , w38843 , w38844 , w38845 , w38846 , w38847 , w38848 , w38849 , w38850 , w38851 , w38852 , w38853 , w38854 , w38855 , w38856 , w38857 , w38858 , w38859 , w38860 , w38861 , w38862 , w38863 , w38864 , w38865 , w38866 , w38867 , w38868 , w38869 , w38870 , w38871 , w38872 , w38873 , w38874 , w38875 , w38876 , w38877 , w38878 , w38879 , w38880 , w38881 , w38882 , w38883 , w38884 , w38885 , w38886 , w38887 , w38888 , w38889 , w38890 , w38891 , w38892 , w38893 , w38894 , w38895 , w38896 , w38897 , w38898 , w38899 , w38900 , w38901 , w38902 , w38903 , w38904 , w38905 , w38906 , w38907 , w38908 , w38909 , w38910 , w38911 , w38912 , w38913 , w38914 , w38915 , w38916 , w38917 , w38918 , w38919 , w38920 , w38921 , w38922 , w38923 , w38924 , w38925 , w38926 , w38927 , w38928 , w38929 , w38930 , w38931 , w38932 , w38933 , w38934 , w38935 , w38936 , w38937 , w38938 , w38939 , w38940 , w38941 , w38942 , w38943 , w38944 , w38945 , w38946 , w38947 , w38948 , w38949 , w38950 , w38951 , w38952 , w38953 , w38954 , w38955 , w38956 , w38957 , w38958 , w38959 , w38960 , w38961 , w38962 , w38963 , w38964 , w38965 , w38966 , w38967 , w38968 , w38969 , w38970 , w38971 , w38972 , w38973 , w38974 , w38975 , w38976 , w38977 , w38978 , w38979 , w38980 , w38981 , w38982 , w38983 , w38984 , w38985 , w38986 , w38987 , w38988 , w38989 , w38990 , w38991 , w38992 , w38993 , w38994 , w38995 , w38996 , w38997 , w38998 , w38999 , w39000 , w39001 , w39002 , w39003 , w39004 , w39005 , w39006 , w39007 , w39008 , w39009 , w39010 , w39011 , w39012 , w39013 , w39014 , w39015 , w39016 , w39017 , w39018 , w39019 , w39020 , w39021 , w39022 , w39023 , w39024 , w39025 , w39026 , w39027 , w39028 , w39029 , w39030 , w39031 , w39032 , w39033 , w39034 , w39035 , w39036 , w39037 , w39038 , w39039 , w39040 , w39041 , w39042 , w39043 , w39044 , w39045 , w39046 , w39047 , w39048 , w39049 , w39050 , w39051 , w39052 , w39053 , w39054 , w39055 , w39056 , w39057 , w39058 , w39059 , w39060 , w39061 , w39062 , w39063 , w39064 , w39065 , w39066 , w39067 , w39068 , w39069 , w39070 , w39071 , w39072 , w39073 , w39074 , w39075 , w39076 , w39077 , w39078 , w39079 , w39080 , w39081 , w39082 , w39083 , w39084 , w39085 , w39086 , w39087 , w39088 , w39089 , w39090 , w39091 , w39092 , w39093 , w39094 , w39095 , w39096 , w39097 , w39098 , w39099 , w39100 , w39101 , w39102 , w39103 , w39104 , w39105 , w39106 , w39107 , w39108 , w39109 , w39110 , w39111 , w39112 , w39113 , w39114 , w39115 , w39116 , w39117 , w39118 , w39119 , w39120 , w39121 , w39122 , w39123 , w39124 , w39125 , w39126 , w39127 , w39128 , w39129 , w39130 , w39131 , w39132 , w39133 , w39134 , w39135 , w39136 , w39137 , w39138 , w39139 , w39140 , w39141 , w39142 , w39143 , w39144 , w39145 , w39146 , w39147 , w39148 , w39149 , w39150 , w39151 , w39152 , w39153 , w39154 , w39155 , w39156 , w39157 , w39158 , w39159 , w39160 , w39161 , w39162 , w39163 , w39164 , w39165 , w39166 , w39167 , w39168 , w39169 , w39170 , w39171 , w39172 , w39173 , w39174 , w39175 , w39176 , w39177 , w39178 , w39179 , w39180 , w39181 , w39182 , w39183 , w39184 , w39185 , w39186 , w39187 , w39188 , w39189 , w39190 , w39191 , w39192 , w39193 , w39194 , w39195 , w39196 , w39197 , w39198 , w39199 , w39200 , w39201 , w39202 , w39203 , w39204 , w39205 , w39206 , w39207 , w39208 , w39209 , w39210 , w39211 , w39212 , w39213 , w39214 , w39215 , w39216 , w39217 , w39218 , w39219 , w39220 , w39221 , w39222 , w39223 , w39224 , w39225 , w39226 , w39227 , w39228 , w39229 , w39230 , w39231 , w39232 , w39233 , w39234 , w39235 , w39236 , w39237 , w39238 , w39239 , w39240 , w39241 , w39242 , w39243 , w39244 , w39245 , w39246 , w39247 , w39248 , w39249 , w39250 , w39251 , w39252 , w39253 , w39254 , w39255 , w39256 , w39257 , w39258 , w39259 , w39260 , w39261 , w39262 , w39263 , w39264 , w39265 , w39266 , w39267 , w39268 , w39269 , w39270 , w39271 , w39272 , w39273 , w39274 , w39275 , w39276 , w39277 , w39278 , w39279 , w39280 , w39281 , w39282 , w39283 , w39284 , w39285 , w39286 , w39287 , w39288 , w39289 , w39290 , w39291 , w39292 , w39293 , w39294 , w39295 , w39296 , w39297 , w39298 , w39299 , w39300 , w39301 , w39302 , w39303 , w39304 , w39305 , w39306 , w39307 , w39308 , w39309 , w39310 , w39311 , w39312 , w39313 , w39314 , w39315 , w39316 , w39317 , w39318 , w39319 , w39320 , w39321 , w39322 , w39323 , w39324 , w39325 , w39326 , w39327 , w39328 , w39329 , w39330 , w39331 , w39332 , w39333 , w39334 , w39335 , w39336 , w39337 , w39338 , w39339 , w39340 , w39341 , w39342 , w39343 , w39344 , w39345 , w39346 , w39347 , w39348 , w39349 , w39350 , w39351 , w39352 , w39353 , w39354 , w39355 , w39356 , w39357 , w39358 , w39359 , w39360 , w39361 , w39362 , w39363 , w39364 , w39365 , w39366 , w39367 , w39368 , w39369 , w39370 , w39371 , w39372 , w39373 , w39374 , w39375 , w39376 , w39377 , w39378 , w39379 , w39380 , w39381 , w39382 , w39383 , w39384 , w39385 , w39386 , w39387 , w39388 , w39389 , w39390 , w39391 , w39392 , w39393 , w39394 , w39395 , w39396 , w39397 , w39398 , w39399 , w39400 , w39401 , w39402 , w39403 , w39404 , w39405 , w39406 , w39407 , w39408 , w39409 , w39410 , w39411 , w39412 , w39413 , w39414 , w39415 , w39416 , w39417 , w39418 , w39419 , w39420 , w39421 , w39422 , w39423 , w39424 , w39425 , w39426 , w39427 , w39428 , w39429 , w39430 , w39431 , w39432 , w39433 , w39434 , w39435 , w39436 , w39437 , w39438 , w39439 , w39440 , w39441 , w39442 , w39443 , w39444 , w39445 , w39446 , w39447 , w39448 , w39449 , w39450 , w39451 , w39452 , w39453 , w39454 , w39455 , w39456 , w39457 , w39458 , w39459 , w39460 , w39461 , w39462 , w39463 , w39464 , w39465 , w39466 , w39467 , w39468 , w39469 , w39470 , w39471 , w39472 , w39473 , w39474 , w39475 , w39476 , w39477 , w39478 , w39479 , w39480 , w39481 , w39482 , w39483 , w39484 , w39485 , w39486 , w39487 , w39488 , w39489 , w39490 , w39491 , w39492 , w39493 , w39494 , w39495 , w39496 , w39497 , w39498 , w39499 , w39500 , w39501 , w39502 , w39503 , w39504 , w39505 , w39506 , w39507 , w39508 , w39509 , w39510 , w39511 , w39512 , w39513 , w39514 , w39515 , w39516 , w39517 , w39518 , w39519 , w39520 , w39521 , w39522 , w39523 , w39524 , w39525 , w39526 , w39527 , w39528 , w39529 , w39530 , w39531 , w39532 , w39533 , w39534 , w39535 , w39536 , w39537 , w39538 , w39539 , w39540 , w39541 , w39542 , w39543 , w39544 , w39545 , w39546 , w39547 , w39548 , w39549 , w39550 , w39551 , w39552 , w39553 , w39554 , w39555 , w39556 , w39557 , w39558 , w39559 , w39560 , w39561 , w39562 , w39563 , w39564 , w39565 , w39566 , w39567 , w39568 , w39569 , w39570 , w39571 , w39572 , w39573 , w39574 , w39575 , w39576 , w39577 , w39578 , w39579 , w39580 , w39581 , w39582 , w39583 , w39584 , w39585 , w39586 , w39587 , w39588 , w39589 , w39590 , w39591 , w39592 , w39593 , w39594 , w39595 , w39596 , w39597 , w39598 , w39599 , w39600 , w39601 , w39602 , w39603 , w39604 , w39605 , w39606 , w39607 , w39608 , w39609 , w39610 , w39611 , w39612 , w39613 , w39614 , w39615 , w39616 , w39617 , w39618 , w39619 , w39620 , w39621 , w39622 , w39623 , w39624 , w39625 , w39626 , w39627 , w39628 , w39629 , w39630 , w39631 , w39632 , w39633 , w39634 , w39635 , w39636 , w39637 , w39638 , w39639 , w39640 , w39641 , w39642 , w39643 , w39644 , w39645 , w39646 , w39647 , w39648 , w39649 , w39650 , w39651 , w39652 , w39653 , w39654 , w39655 , w39656 , w39657 , w39658 , w39659 , w39660 , w39661 , w39662 , w39663 , w39664 , w39665 , w39666 , w39667 , w39668 , w39669 , w39670 , w39671 , w39672 , w39673 , w39674 , w39675 , w39676 , w39677 , w39678 , w39679 , w39680 , w39681 , w39682 , w39683 , w39684 , w39685 , w39686 , w39687 , w39688 , w39689 , w39690 , w39691 , w39692 , w39693 , w39694 , w39695 , w39696 , w39697 , w39698 , w39699 , w39700 , w39701 , w39702 , w39703 , w39704 , w39705 , w39706 , w39707 , w39708 , w39709 , w39710 , w39711 , w39712 , w39713 , w39714 , w39715 , w39716 , w39717 , w39718 , w39719 , w39720 , w39721 , w39722 , w39723 , w39724 , w39725 , w39726 , w39727 , w39728 , w39729 , w39730 , w39731 , w39732 , w39733 , w39734 , w39735 , w39736 , w39737 , w39738 , w39739 , w39740 , w39741 , w39742 , w39743 , w39744 , w39745 , w39746 , w39747 , w39748 , w39749 , w39750 , w39751 , w39752 , w39753 , w39754 , w39755 , w39756 , w39757 , w39758 , w39759 , w39760 , w39761 , w39762 , w39763 , w39764 , w39765 , w39766 , w39767 , w39768 , w39769 , w39770 , w39771 , w39772 , w39773 , w39774 , w39775 , w39776 , w39777 , w39778 , w39779 , w39780 , w39781 , w39782 , w39783 , w39784 , w39785 , w39786 , w39787 , w39788 , w39789 , w39790 , w39791 , w39792 , w39793 , w39794 , w39795 , w39796 , w39797 , w39798 , w39799 , w39800 , w39801 , w39802 , w39803 , w39804 , w39805 , w39806 , w39807 , w39808 , w39809 , w39810 , w39811 , w39812 , w39813 , w39814 , w39815 , w39816 , w39817 , w39818 , w39819 , w39820 , w39821 , w39822 , w39823 , w39824 , w39825 , w39826 , w39827 , w39828 , w39829 , w39830 , w39831 , w39832 , w39833 , w39834 , w39835 , w39836 , w39837 , w39838 , w39839 , w39840 , w39841 , w39842 , w39843 , w39844 , w39845 , w39846 , w39847 , w39848 , w39849 , w39850 , w39851 , w39852 , w39853 , w39854 , w39855 , w39856 , w39857 , w39858 , w39859 , w39860 , w39861 , w39862 , w39863 , w39864 , w39865 , w39866 , w39867 , w39868 , w39869 , w39870 , w39871 , w39872 , w39873 , w39874 , w39875 , w39876 , w39877 , w39878 , w39879 , w39880 , w39881 , w39882 , w39883 , w39884 , w39885 , w39886 , w39887 , w39888 , w39889 , w39890 , w39891 , w39892 , w39893 , w39894 , w39895 , w39896 ;
  assign zero = 0;
  assign w129 = \pi066 | \pi067 ;
  assign w130 = \pi073 | \pi075 ;
  assign w131 = ( \pi072 & ~\pi073 ) | ( \pi072 & \pi074 ) | ( ~\pi073 & \pi074 ) ;
  assign w132 = w130 | w131 ;
  assign w133 = \pi069 | \pi071 ;
  assign w134 = ( \pi068 & ~\pi069 ) | ( \pi068 & \pi070 ) | ( ~\pi069 & \pi070 ) ;
  assign w135 = w133 | w134 ;
  assign w136 = \pi081 | \pi083 ;
  assign w137 = ( \pi080 & ~\pi081 ) | ( \pi080 & \pi082 ) | ( ~\pi081 & \pi082 ) ;
  assign w138 = w136 | w137 ;
  assign w139 = \pi077 | \pi079 ;
  assign w140 = ( \pi076 & ~\pi077 ) | ( \pi076 & \pi078 ) | ( ~\pi077 & \pi078 ) ;
  assign w141 = w139 | w140 ;
  assign w142 = w138 | w141 ;
  assign w143 = ( ~w132 & w135 ) | ( ~w132 & w142 ) | ( w135 & w142 ) ;
  assign w144 = w132 | w143 ;
  assign w145 = \pi125 | \pi127 ;
  assign w146 = ( \pi124 & ~\pi125 ) | ( \pi124 & \pi126 ) | ( ~\pi125 & \pi126 ) ;
  assign w147 = w145 | w146 ;
  assign w148 = \pi121 | \pi123 ;
  assign w149 = ( \pi120 & ~\pi121 ) | ( \pi120 & \pi122 ) | ( ~\pi121 & \pi122 ) ;
  assign w150 = w148 | w149 ;
  assign w151 = \pi117 | \pi119 ;
  assign w152 = ( \pi116 & ~\pi117 ) | ( \pi116 & \pi118 ) | ( ~\pi117 & \pi118 ) ;
  assign w153 = w151 | w152 ;
  assign w154 = ( w147 & ~w150 ) | ( w147 & w153 ) | ( ~w150 & w153 ) ;
  assign w155 = w150 | w154 ;
  assign w156 = \pi105 | \pi107 ;
  assign w157 = ( \pi104 & ~\pi105 ) | ( \pi104 & \pi106 ) | ( ~\pi105 & \pi106 ) ;
  assign w158 = w156 | w157 ;
  assign w159 = \pi101 | \pi103 ;
  assign w160 = ( \pi100 & ~\pi101 ) | ( \pi100 & \pi102 ) | ( ~\pi101 & \pi102 ) ;
  assign w161 = w159 | w160 ;
  assign w162 = \pi113 | \pi115 ;
  assign w163 = ( \pi112 & ~\pi113 ) | ( \pi112 & \pi114 ) | ( ~\pi113 & \pi114 ) ;
  assign w164 = w162 | w163 ;
  assign w165 = \pi109 | \pi111 ;
  assign w166 = ( \pi108 & ~\pi109 ) | ( \pi108 & \pi110 ) | ( ~\pi109 & \pi110 ) ;
  assign w167 = w165 | w166 ;
  assign w168 = w164 | w167 ;
  assign w169 = ( ~w158 & w161 ) | ( ~w158 & w168 ) | ( w161 & w168 ) ;
  assign w170 = w158 | w169 ;
  assign w171 = \pi089 | \pi091 ;
  assign w172 = ( \pi088 & ~\pi089 ) | ( \pi088 & \pi090 ) | ( ~\pi089 & \pi090 ) ;
  assign w173 = w171 | w172 ;
  assign w174 = \pi085 | \pi087 ;
  assign w175 = ( \pi084 & ~\pi085 ) | ( \pi084 & \pi086 ) | ( ~\pi085 & \pi086 ) ;
  assign w176 = w174 | w175 ;
  assign w177 = \pi097 | \pi099 ;
  assign w178 = ( \pi096 & ~\pi097 ) | ( \pi096 & \pi098 ) | ( ~\pi097 & \pi098 ) ;
  assign w179 = w177 | w178 ;
  assign w180 = \pi093 | \pi095 ;
  assign w181 = ( \pi092 & ~\pi093 ) | ( \pi092 & \pi094 ) | ( ~\pi093 & \pi094 ) ;
  assign w182 = w180 | w181 ;
  assign w183 = w179 | w182 ;
  assign w184 = ( ~w173 & w176 ) | ( ~w173 & w183 ) | ( w176 & w183 ) ;
  assign w185 = w173 | w184 ;
  assign w186 = ( w155 & w170 ) | ( w155 & ~w185 ) | ( w170 & ~w185 ) ;
  assign w187 = w185 | w186 ;
  assign w188 = ( ~\pi063 & \pi064 ) | ( ~\pi063 & w129 ) | ( \pi064 & w129 ) ;
  assign w189 = w144 | w187 ;
  assign w190 = ( \pi064 & ~\pi065 ) | ( \pi064 & w144 ) | ( ~\pi065 & w144 ) ;
  assign w191 = ~w189 & w190 ;
  assign w192 = ~w188 & w191 ;
  assign w193 = \pi063 & ~w192 ;
  assign w194 = ~\pi062 & \pi064 ;
  assign w195 = ( \pi065 & ~w193 ) | ( \pi065 & w194 ) | ( ~w193 & w194 ) ;
  assign w196 = w132 | w141 ;
  assign w197 = ( ~w129 & w135 ) | ( ~w129 & w196 ) | ( w135 & w196 ) ;
  assign w198 = w129 | w197 ;
  assign w199 = w147 | w150 ;
  assign w200 = ( ~w153 & w164 ) | ( ~w153 & w199 ) | ( w164 & w199 ) ;
  assign w201 = w153 | w200 ;
  assign w202 = w158 | w167 ;
  assign w203 = ( ~w161 & w179 ) | ( ~w161 & w202 ) | ( w179 & w202 ) ;
  assign w204 = w161 | w203 ;
  assign w205 = w173 | w182 ;
  assign w206 = ( ~w138 & w176 ) | ( ~w138 & w205 ) | ( w176 & w205 ) ;
  assign w207 = w138 | w206 ;
  assign w208 = ( w201 & ~w204 ) | ( w201 & w207 ) | ( ~w204 & w207 ) ;
  assign w209 = w204 | w208 ;
  assign w210 = w198 | w209 ;
  assign w211 = \pi065 ^ w194 ;
  assign w212 = ~w210 & w211 ;
  assign w213 = ~w195 & w212 ;
  assign w214 = ( \pi063 & ~w192 ) | ( \pi063 & w195 ) | ( ~w192 & w195 ) ;
  assign w215 = w213 & ~w214 ;
  assign w216 = w138 | w176 ;
  assign w217 = w129 | w216 ;
  assign w218 = w197 | w217 ;
  assign w219 = ( w153 & w161 ) | ( w153 & ~w164 ) | ( w161 & ~w164 ) ;
  assign w220 = w202 | w205 ;
  assign w221 = ( w164 & w179 ) | ( w164 & ~w205 ) | ( w179 & ~w205 ) ;
  assign w222 = w220 | w221 ;
  assign w223 = w219 | w222 ;
  assign w224 = ( ~\pi062 & \pi064 ) | ( ~\pi062 & w218 ) | ( \pi064 & w218 ) ;
  assign w225 = \pi065 ^ w224 ;
  assign w226 = ( w199 & ~w223 ) | ( w199 & w225 ) | ( ~w223 & w225 ) ;
  assign w227 = ( ~w199 & w218 ) | ( ~w199 & w226 ) | ( w218 & w226 ) ;
  assign w228 = ~w218 & w227 ;
  assign w229 = ( w192 & ~w195 ) | ( w192 & w228 ) | ( ~w195 & w228 ) ;
  assign w230 = w193 & ~w229 ;
  assign w231 = ~\pi061 & \pi064 ;
  assign w232 = \pi086 | \pi088 ;
  assign w233 = ( \pi085 & ~\pi086 ) | ( \pi085 & \pi087 ) | ( ~\pi086 & \pi087 ) ;
  assign w234 = w232 | w233 ;
  assign w235 = \pi082 | \pi084 ;
  assign w236 = ( \pi081 & ~\pi082 ) | ( \pi081 & \pi083 ) | ( ~\pi082 & \pi083 ) ;
  assign w237 = w235 | w236 ;
  assign w238 = \pi094 | \pi096 ;
  assign w239 = ( \pi093 & ~\pi094 ) | ( \pi093 & \pi095 ) | ( ~\pi094 & \pi095 ) ;
  assign w240 = w238 | w239 ;
  assign w241 = \pi090 | \pi092 ;
  assign w242 = ( \pi089 & ~\pi090 ) | ( \pi089 & \pi091 ) | ( ~\pi090 & \pi091 ) ;
  assign w243 = w241 | w242 ;
  assign w244 = w240 | w243 ;
  assign w245 = ( ~w234 & w237 ) | ( ~w234 & w244 ) | ( w237 & w244 ) ;
  assign w246 = w234 | w245 ;
  assign w247 = \pi070 | \pi072 ;
  assign w248 = ( \pi069 & ~\pi070 ) | ( \pi069 & \pi071 ) | ( ~\pi070 & \pi071 ) ;
  assign w249 = w247 | w248 ;
  assign w250 = \pi067 | \pi068 ;
  assign w251 = \pi078 | \pi080 ;
  assign w252 = ( \pi077 & ~\pi078 ) | ( \pi077 & \pi079 ) | ( ~\pi078 & \pi079 ) ;
  assign w253 = w251 | w252 ;
  assign w254 = \pi074 | \pi076 ;
  assign w255 = ( \pi073 & ~\pi074 ) | ( \pi073 & \pi075 ) | ( ~\pi074 & \pi075 ) ;
  assign w256 = w254 | w255 ;
  assign w257 = w253 | w256 ;
  assign w258 = \pi064 & ~\pi066 ;
  assign w259 = ~w249 & w258 ;
  assign w260 = ( ~w249 & w250 ) | ( ~w249 & w257 ) | ( w250 & w257 ) ;
  assign w261 = w259 & ~w260 ;
  assign w262 = \pi118 | \pi120 ;
  assign w263 = ( \pi117 & ~\pi118 ) | ( \pi117 & \pi119 ) | ( ~\pi118 & \pi119 ) ;
  assign w264 = w262 | w263 ;
  assign w265 = \pi114 | \pi116 ;
  assign w266 = ( \pi113 & ~\pi114 ) | ( \pi113 & \pi115 ) | ( ~\pi114 & \pi115 ) ;
  assign w267 = w265 | w266 ;
  assign w268 = ( \pi125 & ~\pi126 ) | ( \pi125 & \pi127 ) | ( ~\pi126 & \pi127 ) ;
  assign w269 = \pi126 | w268 ;
  assign w270 = \pi123 | \pi124 ;
  assign w271 = ( ~\pi121 & \pi122 ) | ( ~\pi121 & w270 ) | ( \pi122 & w270 ) ;
  assign w272 = \pi121 | w271 ;
  assign w273 = w269 | w272 ;
  assign w274 = ( ~w264 & w267 ) | ( ~w264 & w273 ) | ( w267 & w273 ) ;
  assign w275 = w264 | w274 ;
  assign w276 = \pi102 | \pi104 ;
  assign w277 = ( \pi101 & ~\pi102 ) | ( \pi101 & \pi103 ) | ( ~\pi102 & \pi103 ) ;
  assign w278 = w276 | w277 ;
  assign w279 = \pi098 | \pi100 ;
  assign w280 = ( \pi097 & ~\pi098 ) | ( \pi097 & \pi099 ) | ( ~\pi098 & \pi099 ) ;
  assign w281 = w279 | w280 ;
  assign w282 = \pi110 | \pi112 ;
  assign w283 = ( \pi109 & ~\pi110 ) | ( \pi109 & \pi111 ) | ( ~\pi110 & \pi111 ) ;
  assign w284 = w282 | w283 ;
  assign w285 = \pi106 | \pi108 ;
  assign w286 = ( \pi105 & ~\pi106 ) | ( \pi105 & \pi107 ) | ( ~\pi106 & \pi107 ) ;
  assign w287 = w285 | w286 ;
  assign w288 = w284 | w287 ;
  assign w289 = ( ~w278 & w281 ) | ( ~w278 & w288 ) | ( w281 & w288 ) ;
  assign w290 = w278 | w289 ;
  assign w291 = w275 | w290 ;
  assign w292 = ( w246 & w261 ) | ( w246 & ~w291 ) | ( w261 & ~w291 ) ;
  assign w293 = ~w246 & w292 ;
  assign w294 = ( \pi062 & w195 ) | ( \pi062 & ~w293 ) | ( w195 & ~w293 ) ;
  assign w295 = \pi062 & w294 ;
  assign w296 = ~w129 & w194 ;
  assign w297 = ~w197 & w296 ;
  assign w298 = w201 | w204 ;
  assign w299 = ( w207 & w297 ) | ( w207 & ~w298 ) | ( w297 & ~w298 ) ;
  assign w300 = ~w207 & w299 ;
  assign w301 = ~w195 & w300 ;
  assign w302 = w295 | w301 ;
  assign w303 = ( \pi065 & w231 ) | ( \pi065 & ~w302 ) | ( w231 & ~w302 ) ;
  assign w304 = w215 | w230 ;
  assign w305 = ( \pi066 & w303 ) | ( \pi066 & ~w304 ) | ( w303 & ~w304 ) ;
  assign w306 = w249 | w250 ;
  assign w307 = w246 | w306 ;
  assign w308 = ( ~w246 & w257 ) | ( ~w246 & w291 ) | ( w257 & w291 ) ;
  assign w309 = w307 | w308 ;
  assign w310 = w305 | w309 ;
  assign w311 = ( \pi067 & w215 ) | ( \pi067 & w230 ) | ( w215 & w230 ) ;
  assign w312 = \pi067 & ~w311 ;
  assign w313 = \pi066 ^ w303 ;
  assign w314 = ( ~\pi067 & w309 ) | ( ~\pi067 & w313 ) | ( w309 & w313 ) ;
  assign w315 = ( w312 & w313 ) | ( w312 & ~w314 ) | ( w313 & ~w314 ) ;
  assign w316 = w234 | w306 ;
  assign w317 = ( ~w234 & w237 ) | ( ~w234 & w257 ) | ( w237 & w257 ) ;
  assign w318 = w316 | w317 ;
  assign w319 = ( w264 & w267 ) | ( w264 & ~w278 ) | ( w267 & ~w278 ) ;
  assign w320 = w244 | w288 ;
  assign w321 = ( w278 & w281 ) | ( w278 & ~w288 ) | ( w281 & ~w288 ) ;
  assign w322 = w320 | w321 ;
  assign w323 = w319 | w322 ;
  assign w324 = ( \pi065 & w231 ) | ( \pi065 & ~w318 ) | ( w231 & ~w318 ) ;
  assign w325 = w273 | w323 ;
  assign w326 = ( \pi065 & w231 ) | ( \pi065 & w325 ) | ( w231 & w325 ) ;
  assign w327 = w324 & ~w326 ;
  assign w328 = ( w302 & w305 ) | ( w302 & ~w327 ) | ( w305 & ~w327 ) ;
  assign w329 = w302 & w328 ;
  assign w330 = ( ~w246 & w275 ) | ( ~w246 & w290 ) | ( w275 & w290 ) ;
  assign w331 = w246 | w330 ;
  assign w332 = \pi065 ^ w231 ;
  assign w333 = ( ~w257 & w331 ) | ( ~w257 & w332 ) | ( w331 & w332 ) ;
  assign w334 = ( w249 & ~w250 ) | ( w249 & w331 ) | ( ~w250 & w331 ) ;
  assign w335 = ( w250 & w333 ) | ( w250 & w334 ) | ( w333 & w334 ) ;
  assign w336 = w333 & ~w335 ;
  assign w337 = ~w295 & w336 ;
  assign w338 = ( ~w295 & w301 ) | ( ~w295 & w305 ) | ( w301 & w305 ) ;
  assign w339 = w337 & ~w338 ;
  assign w340 = w329 | w339 ;
  assign w341 = ~\pi066 & w340 ;
  assign w342 = ( \pi066 & ~w329 ) | ( \pi066 & w339 ) | ( ~w329 & w339 ) ;
  assign w343 = ~w339 & w342 ;
  assign w344 = ( \pi064 & w135 ) | ( \pi064 & w196 ) | ( w135 & w196 ) ;
  assign w345 = w207 | w298 ;
  assign w346 = ( \pi064 & ~\pi067 ) | ( \pi064 & w207 ) | ( ~\pi067 & w207 ) ;
  assign w347 = ~w345 & w346 ;
  assign w348 = ~w344 & w347 ;
  assign w349 = ( w231 & w249 ) | ( w231 & ~w257 ) | ( w249 & ~w257 ) ;
  assign w350 = w246 | w291 ;
  assign w351 = ( ~w246 & w249 ) | ( ~w246 & w250 ) | ( w249 & w250 ) ;
  assign w352 = w350 | w351 ;
  assign w353 = w349 & ~w352 ;
  assign w354 = ( \pi061 & w305 ) | ( \pi061 & ~w348 ) | ( w305 & ~w348 ) ;
  assign w355 = \pi061 & w354 ;
  assign w356 = w305 | w353 ;
  assign w357 = ( ~w305 & w355 ) | ( ~w305 & w356 ) | ( w355 & w356 ) ;
  assign w358 = ~\pi060 & \pi064 ;
  assign w359 = ( \pi065 & ~w357 ) | ( \pi065 & w358 ) | ( ~w357 & w358 ) ;
  assign w360 = w343 | w359 ;
  assign w361 = ~w341 & w360 ;
  assign w362 = ( \pi066 & w303 ) | ( \pi066 & ~w309 ) | ( w303 & ~w309 ) ;
  assign w363 = \pi066 & w303 ;
  assign w364 = ( w304 & ~w362 ) | ( w304 & w363 ) | ( ~w362 & w363 ) ;
  assign w365 = ~\pi067 & w364 ;
  assign w366 = ( w315 & w361 ) | ( w315 & ~w365 ) | ( w361 & ~w365 ) ;
  assign w367 = ~w365 & w366 ;
  assign w368 = w155 | w170 ;
  assign w369 = ( ~w144 & w185 ) | ( ~w144 & w368 ) | ( w185 & w368 ) ;
  assign w370 = w144 | w369 ;
  assign w371 = ~w361 & w365 ;
  assign w372 = ~w370 & w371 ;
  assign w373 = w367 | w370 ;
  assign w374 = w364 & w373 ;
  assign w375 = ( \pi068 & w372 ) | ( \pi068 & ~w374 ) | ( w372 & ~w374 ) ;
  assign w376 = ~w372 & w375 ;
  assign w377 = ( w341 & w343 ) | ( w341 & w359 ) | ( w343 & w359 ) ;
  assign w378 = w359 & w377 ;
  assign w379 = w370 | w378 ;
  assign w380 = ( w360 & ~w367 ) | ( w360 & w378 ) | ( ~w367 & w378 ) ;
  assign w381 = ~w379 & w380 ;
  assign w382 = ( \pi066 & ~w370 ) | ( \pi066 & w378 ) | ( ~w370 & w378 ) ;
  assign w383 = w370 & w382 ;
  assign w384 = ( w367 & w382 ) | ( w367 & w383 ) | ( w382 & w383 ) ;
  assign w385 = ( w340 & ~w382 ) | ( w340 & w384 ) | ( ~w382 & w384 ) ;
  assign w386 = w381 | w385 ;
  assign w387 = ~\pi067 & w386 ;
  assign w388 = ( \pi067 & ~w381 ) | ( \pi067 & w385 ) | ( ~w381 & w385 ) ;
  assign w389 = ~w385 & w388 ;
  assign w390 = w173 | w176 ;
  assign w391 = w132 | w390 ;
  assign w392 = w143 | w391 ;
  assign w393 = ( w150 & w153 ) | ( w150 & ~w158 ) | ( w153 & ~w158 ) ;
  assign w394 = w168 | w183 ;
  assign w395 = ( w158 & w161 ) | ( w158 & ~w183 ) | ( w161 & ~w183 ) ;
  assign w396 = w394 | w395 ;
  assign w397 = w393 | w396 ;
  assign w398 = ( ~\pi060 & \pi064 ) | ( ~\pi060 & w392 ) | ( \pi064 & w392 ) ;
  assign w399 = \pi065 ^ w398 ;
  assign w400 = ( w147 & ~w397 ) | ( w147 & w399 ) | ( ~w397 & w399 ) ;
  assign w401 = ( ~w147 & w392 ) | ( ~w147 & w400 ) | ( w392 & w400 ) ;
  assign w402 = ~w392 & w401 ;
  assign w403 = ( w357 & w367 ) | ( w357 & ~w402 ) | ( w367 & ~w402 ) ;
  assign w404 = w357 & w403 ;
  assign w405 = \pi065 ^ w358 ;
  assign w406 = ~w189 & w405 ;
  assign w407 = ( w305 & w367 ) | ( w305 & w406 ) | ( w367 & w406 ) ;
  assign w408 = w348 & ~w407 ;
  assign w409 = ( \pi061 & w367 ) | ( \pi061 & ~w408 ) | ( w367 & ~w408 ) ;
  assign w410 = ( ~w353 & w406 ) | ( ~w353 & w407 ) | ( w406 & w407 ) ;
  assign w411 = ~w409 & w410 ;
  assign w412 = w404 | w411 ;
  assign w413 = ~\pi066 & w412 ;
  assign w414 = ( \pi066 & ~w404 ) | ( \pi066 & w411 ) | ( ~w404 & w411 ) ;
  assign w415 = ~w411 & w414 ;
  assign w416 = ~\pi059 & \pi064 ;
  assign w417 = ( \pi064 & w249 ) | ( \pi064 & w257 ) | ( w249 & w257 ) ;
  assign w418 = ( \pi064 & ~\pi068 ) | ( \pi064 & w246 ) | ( ~\pi068 & w246 ) ;
  assign w419 = ~w350 & w418 ;
  assign w420 = ~w417 & w419 ;
  assign w421 = ( ~\pi060 & w135 ) | ( ~\pi060 & w196 ) | ( w135 & w196 ) ;
  assign w422 = ( ~\pi060 & \pi064 ) | ( ~\pi060 & w207 ) | ( \pi064 & w207 ) ;
  assign w423 = ~w345 & w422 ;
  assign w424 = ~w421 & w423 ;
  assign w425 = ( \pi060 & w367 ) | ( \pi060 & ~w420 ) | ( w367 & ~w420 ) ;
  assign w426 = \pi060 & w425 ;
  assign w427 = w367 | w424 ;
  assign w428 = ( ~w367 & w426 ) | ( ~w367 & w427 ) | ( w426 & w427 ) ;
  assign w429 = ( \pi065 & w416 ) | ( \pi065 & ~w428 ) | ( w416 & ~w428 ) ;
  assign w430 = w415 | w429 ;
  assign w431 = ( w389 & ~w413 ) | ( w389 & w430 ) | ( ~w413 & w430 ) ;
  assign w432 = w389 | w431 ;
  assign w433 = ( ~\pi068 & w372 ) | ( ~\pi068 & w374 ) | ( w372 & w374 ) ;
  assign w434 = ~\pi068 & w433 ;
  assign w435 = ~w387 & w432 ;
  assign w436 = w376 & ~w435 ;
  assign w437 = ( ~w434 & w435 ) | ( ~w434 & w436 ) | ( w435 & w436 ) ;
  assign w438 = ~w413 & w430 ;
  assign w439 = ( w387 & w389 ) | ( w387 & w430 ) | ( w389 & w430 ) ;
  assign w440 = w438 & w439 ;
  assign w441 = w240 | w281 ;
  assign w442 = ( ~w234 & w243 ) | ( ~w234 & w441 ) | ( w243 & w441 ) ;
  assign w443 = w234 | w442 ;
  assign w444 = w237 | w253 ;
  assign w445 = ( ~w249 & w256 ) | ( ~w249 & w444 ) | ( w256 & w444 ) ;
  assign w446 = w249 | w445 ;
  assign w447 = ( ~w264 & w269 ) | ( ~w264 & w272 ) | ( w269 & w272 ) ;
  assign w448 = w264 | w447 ;
  assign w449 = w267 | w284 ;
  assign w450 = ( ~w278 & w287 ) | ( ~w278 & w449 ) | ( w287 & w449 ) ;
  assign w451 = w278 | w450 ;
  assign w452 = w448 | w451 ;
  assign w453 = ( ~w443 & w446 ) | ( ~w443 & w452 ) | ( w446 & w452 ) ;
  assign w454 = w443 | w453 ;
  assign w455 = w432 & ~w454 ;
  assign w456 = ( w432 & w437 ) | ( w432 & w440 ) | ( w437 & w440 ) ;
  assign w457 = w455 & ~w456 ;
  assign w458 = ( \pi067 & w440 ) | ( \pi067 & ~w454 ) | ( w440 & ~w454 ) ;
  assign w459 = w454 & w458 ;
  assign w460 = ( w437 & w458 ) | ( w437 & w459 ) | ( w458 & w459 ) ;
  assign w461 = ( w386 & ~w458 ) | ( w386 & w460 ) | ( ~w458 & w460 ) ;
  assign w462 = w457 | w461 ;
  assign w463 = \pi068 ^ w462 ;
  assign w464 = ( w413 & w415 ) | ( w413 & w429 ) | ( w415 & w429 ) ;
  assign w465 = w429 & w464 ;
  assign w466 = w454 | w465 ;
  assign w467 = ( w430 & ~w437 ) | ( w430 & w465 ) | ( ~w437 & w465 ) ;
  assign w468 = ~w466 & w467 ;
  assign w469 = ( \pi066 & ~w454 ) | ( \pi066 & w465 ) | ( ~w454 & w465 ) ;
  assign w470 = w454 & w469 ;
  assign w471 = ( w437 & w469 ) | ( w437 & w470 ) | ( w469 & w470 ) ;
  assign w472 = ( w412 & ~w469 ) | ( w412 & w471 ) | ( ~w469 & w471 ) ;
  assign w473 = w468 | w472 ;
  assign w474 = \pi067 ^ w473 ;
  assign w475 = w249 | w256 ;
  assign w476 = w234 | w475 ;
  assign w477 = ( ~w234 & w243 ) | ( ~w234 & w444 ) | ( w243 & w444 ) ;
  assign w478 = w476 | w477 ;
  assign w479 = ( w264 & ~w278 ) | ( w264 & w449 ) | ( ~w278 & w449 ) ;
  assign w480 = w272 | w441 ;
  assign w481 = ( w278 & w287 ) | ( w278 & ~w441 ) | ( w287 & ~w441 ) ;
  assign w482 = w480 | w481 ;
  assign w483 = w479 | w482 ;
  assign w484 = ( \pi065 & w416 ) | ( \pi065 & ~w483 ) | ( w416 & ~w483 ) ;
  assign w485 = w269 | w478 ;
  assign w486 = ( \pi065 & w416 ) | ( \pi065 & w485 ) | ( w416 & w485 ) ;
  assign w487 = w484 & ~w486 ;
  assign w488 = ( w428 & w437 ) | ( w428 & ~w487 ) | ( w437 & ~w487 ) ;
  assign w489 = w428 & w488 ;
  assign w490 = ( w443 & ~w448 ) | ( w443 & w451 ) | ( ~w448 & w451 ) ;
  assign w491 = w448 | w490 ;
  assign w492 = \pi065 ^ w416 ;
  assign w493 = ( w446 & ~w491 ) | ( w446 & w492 ) | ( ~w491 & w492 ) ;
  assign w494 = ~w446 & w493 ;
  assign w495 = ( w367 & w437 ) | ( w367 & w494 ) | ( w437 & w494 ) ;
  assign w496 = w420 & ~w495 ;
  assign w497 = ( \pi060 & w437 ) | ( \pi060 & ~w496 ) | ( w437 & ~w496 ) ;
  assign w498 = ( ~w424 & w494 ) | ( ~w424 & w495 ) | ( w494 & w495 ) ;
  assign w499 = ~w497 & w498 ;
  assign w500 = w489 | w499 ;
  assign w501 = ~\pi066 & w500 ;
  assign w502 = ( \pi064 & ~\pi069 ) | ( \pi064 & \pi070 ) | ( ~\pi069 & \pi070 ) ;
  assign w503 = w132 | w142 ;
  assign w504 = ( \pi070 & \pi071 ) | ( \pi070 & ~w132 ) | ( \pi071 & ~w132 ) ;
  assign w505 = w503 | w504 ;
  assign w506 = w502 & ~w505 ;
  assign w507 = ( w185 & ~w368 ) | ( w185 & w506 ) | ( ~w368 & w506 ) ;
  assign w508 = ~w185 & w507 ;
  assign w509 = ( \pi059 & w437 ) | ( \pi059 & ~w508 ) | ( w437 & ~w508 ) ;
  assign w510 = \pi059 & w509 ;
  assign w511 = ( w246 & ~w249 ) | ( w246 & w257 ) | ( ~w249 & w257 ) ;
  assign w512 = w291 | w437 ;
  assign w513 = ( ~w249 & w291 ) | ( ~w249 & w416 ) | ( w291 & w416 ) ;
  assign w514 = ~w512 & w513 ;
  assign w515 = ~w511 & w514 ;
  assign w516 = w510 | w515 ;
  assign w517 = ~\pi058 & \pi064 ;
  assign w518 = ( w510 & w515 ) | ( w510 & ~w517 ) | ( w515 & ~w517 ) ;
  assign w519 = \pi065 ^ w518 ;
  assign w520 = w517 | w519 ;
  assign w521 = ~\pi065 & w516 ;
  assign w522 = \pi066 ^ w500 ;
  assign w523 = ( w520 & ~w521 ) | ( w520 & w522 ) | ( ~w521 & w522 ) ;
  assign w524 = w522 | w523 ;
  assign w525 = ( w474 & ~w501 ) | ( w474 & w524 ) | ( ~w501 & w524 ) ;
  assign w526 = w474 | w525 ;
  assign w527 = ~\pi067 & w473 ;
  assign w528 = ( w463 & w526 ) | ( w463 & ~w527 ) | ( w526 & ~w527 ) ;
  assign w529 = w463 | w528 ;
  assign w530 = ~\pi068 & w462 ;
  assign w531 = w376 & w434 ;
  assign w532 = ( w387 & ~w432 ) | ( w387 & w531 ) | ( ~w432 & w531 ) ;
  assign w533 = ( w454 & w531 ) | ( w454 & ~w532 ) | ( w531 & ~w532 ) ;
  assign w534 = w531 & ~w533 ;
  assign w535 = w372 | w374 ;
  assign w536 = ( ~w387 & w432 ) | ( ~w387 & w454 ) | ( w432 & w454 ) ;
  assign w537 = \pi068 ^ w536 ;
  assign w538 = ( w454 & w535 ) | ( w454 & ~w537 ) | ( w535 & ~w537 ) ;
  assign w539 = w535 & w538 ;
  assign w540 = w534 | w539 ;
  assign w541 = \pi069 ^ w540 ;
  assign w542 = ( ~\pi070 & w132 ) | ( ~\pi070 & w142 ) | ( w132 & w142 ) ;
  assign w543 = w185 | w368 ;
  assign w544 = ( \pi070 & \pi071 ) | ( \pi070 & ~w185 ) | ( \pi071 & ~w185 ) ;
  assign w545 = w543 | w544 ;
  assign w546 = w542 | w545 ;
  assign w547 = w541 | w546 ;
  assign w548 = ( w529 & ~w530 ) | ( w529 & w546 ) | ( ~w530 & w546 ) ;
  assign w549 = w547 | w548 ;
  assign w550 = ~w454 & w540 ;
  assign w551 = w549 & ~w550 ;
  assign w552 = w526 & ~w527 ;
  assign w553 = w463 ^ w552 ;
  assign w554 = ~w551 & w553 ;
  assign w555 = ( w462 & ~w549 ) | ( w462 & w550 ) | ( ~w549 & w550 ) ;
  assign w556 = w462 & ~w555 ;
  assign w557 = w554 | w556 ;
  assign w558 = w529 & ~w530 ;
  assign w559 = w541 ^ w558 ;
  assign w560 = ~w551 & w559 ;
  assign w561 = ( w454 & ~w540 ) | ( w454 & w549 ) | ( ~w540 & w549 ) ;
  assign w562 = w540 & w561 ;
  assign w563 = w560 | w562 ;
  assign w564 = ~\pi069 & w557 ;
  assign w565 = ~w501 & w524 ;
  assign w566 = w474 ^ w565 ;
  assign w567 = ~w551 & w566 ;
  assign w568 = ( w473 & ~w549 ) | ( w473 & w550 ) | ( ~w549 & w550 ) ;
  assign w569 = w473 & ~w568 ;
  assign w570 = w567 | w569 ;
  assign w571 = ~\pi068 & w570 ;
  assign w572 = w520 & ~w521 ;
  assign w573 = w522 ^ w572 ;
  assign w574 = ~w551 & w573 ;
  assign w575 = ( w500 & ~w549 ) | ( w500 & w550 ) | ( ~w549 & w550 ) ;
  assign w576 = w500 & ~w575 ;
  assign w577 = w574 | w576 ;
  assign w578 = ~\pi067 & w577 ;
  assign w579 = ( w510 & w515 ) | ( w510 & ~w551 ) | ( w515 & ~w551 ) ;
  assign w580 = ( ~\pi058 & \pi064 ) | ( ~\pi058 & w551 ) | ( \pi064 & w551 ) ;
  assign w581 = w579 ^ w580 ;
  assign w582 = \pi065 ^ w581 ;
  assign w583 = ~w551 & w582 ;
  assign w584 = ( w516 & ~w549 ) | ( w516 & w550 ) | ( ~w549 & w550 ) ;
  assign w585 = w516 & ~w584 ;
  assign w586 = w583 | w585 ;
  assign w587 = ~\pi066 & w586 ;
  assign w588 = \pi066 ^ w586 ;
  assign w589 = \pi064 & ~w551 ;
  assign w590 = \pi058 ^ w589 ;
  assign w591 = ( ~\pi057 & \pi064 ) | ( ~\pi057 & w588 ) | ( \pi064 & w588 ) ;
  assign w592 = ( \pi065 & ~w590 ) | ( \pi065 & w591 ) | ( ~w590 & w591 ) ;
  assign w593 = w588 | w592 ;
  assign w594 = \pi067 ^ w577 ;
  assign w595 = ( ~w587 & w593 ) | ( ~w587 & w594 ) | ( w593 & w594 ) ;
  assign w596 = w594 | w595 ;
  assign w597 = \pi068 ^ w570 ;
  assign w598 = ( ~w578 & w596 ) | ( ~w578 & w597 ) | ( w596 & w597 ) ;
  assign w599 = w597 | w598 ;
  assign w600 = \pi069 ^ w557 ;
  assign w601 = ( ~w571 & w599 ) | ( ~w571 & w600 ) | ( w599 & w600 ) ;
  assign w602 = w600 | w601 ;
  assign w603 = \pi070 ^ w563 ;
  assign w604 = w564 & ~w603 ;
  assign w605 = ( w602 & w603 ) | ( w602 & ~w604 ) | ( w603 & ~w604 ) ;
  assign w606 = ~\pi070 & w563 ;
  assign w607 = w605 & ~w606 ;
  assign w608 = ( ~\pi071 & w256 ) | ( ~\pi071 & w444 ) | ( w256 & w444 ) ;
  assign w609 = w443 | w452 ;
  assign w610 = ( \pi071 & \pi072 ) | ( \pi071 & ~w443 ) | ( \pi072 & ~w443 ) ;
  assign w611 = w609 | w610 ;
  assign w612 = w608 | w611 ;
  assign w613 = w607 | w612 ;
  assign w614 = w557 & w613 ;
  assign w615 = ~w571 & w599 ;
  assign w616 = w600 ^ w615 ;
  assign w617 = ~w613 & w616 ;
  assign w618 = w614 | w617 ;
  assign w619 = w563 & w613 ;
  assign w620 = ~w564 & w602 ;
  assign w621 = w603 ^ w620 ;
  assign w622 = ~w613 & w621 ;
  assign w623 = w619 | w622 ;
  assign w624 = ~\pi070 & w618 ;
  assign w625 = w570 & w613 ;
  assign w626 = ~w578 & w596 ;
  assign w627 = w597 ^ w626 ;
  assign w628 = ~w613 & w627 ;
  assign w629 = w625 | w628 ;
  assign w630 = ~\pi069 & w629 ;
  assign w631 = w577 & w613 ;
  assign w632 = ~w587 & w593 ;
  assign w633 = w594 ^ w632 ;
  assign w634 = ~w613 & w633 ;
  assign w635 = w631 | w634 ;
  assign w636 = ~\pi068 & w635 ;
  assign w637 = w586 & w613 ;
  assign w638 = ~\pi057 & \pi064 ;
  assign w639 = ( \pi065 & ~w590 ) | ( \pi065 & w638 ) | ( ~w590 & w638 ) ;
  assign w640 = w588 ^ w639 ;
  assign w641 = ( w607 & w612 ) | ( w607 & w640 ) | ( w612 & w640 ) ;
  assign w642 = w640 & ~w641 ;
  assign w643 = w637 | w642 ;
  assign w644 = ~\pi067 & w643 ;
  assign w645 = \pi058 ^ \pi065 ;
  assign w646 = \pi057 ^ w551 ;
  assign w647 = ( \pi064 & w612 ) | ( \pi064 & w646 ) | ( w612 & w646 ) ;
  assign w648 = w645 ^ w647 ;
  assign w649 = ~w612 & w648 ;
  assign w650 = ~w607 & w649 ;
  assign w651 = ( ~\pi064 & w551 ) | ( ~\pi064 & w613 ) | ( w551 & w613 ) ;
  assign w652 = \pi058 ^ w651 ;
  assign w653 = w613 & ~w652 ;
  assign w654 = w650 | w653 ;
  assign w655 = ~\pi066 & w654 ;
  assign w656 = ( \pi064 & w132 ) | ( \pi064 & w142 ) | ( w132 & w142 ) ;
  assign w657 = ( \pi064 & ~\pi071 ) | ( \pi064 & w185 ) | ( ~\pi071 & w185 ) ;
  assign w658 = ~w543 & w657 ;
  assign w659 = ~w656 & w658 ;
  assign w660 = ( ~\pi057 & \pi064 ) | ( ~\pi057 & \pi071 ) | ( \pi064 & \pi071 ) ;
  assign w661 = w256 | w444 ;
  assign w662 = ( \pi071 & \pi072 ) | ( \pi071 & ~w256 ) | ( \pi072 & ~w256 ) ;
  assign w663 = w661 | w662 ;
  assign w664 = w660 & ~w663 ;
  assign w665 = ( w443 & ~w452 ) | ( w443 & w664 ) | ( ~w452 & w664 ) ;
  assign w666 = ~w443 & w665 ;
  assign w667 = ( \pi057 & w607 ) | ( \pi057 & ~w659 ) | ( w607 & ~w659 ) ;
  assign w668 = \pi057 & w667 ;
  assign w669 = w607 | w666 ;
  assign w670 = ( ~w607 & w668 ) | ( ~w607 & w669 ) | ( w668 & w669 ) ;
  assign w671 = \pi065 & w670 ;
  assign w672 = ( \pi065 & ~w607 ) | ( \pi065 & w666 ) | ( ~w607 & w666 ) ;
  assign w673 = ~w607 & w659 ;
  assign w674 = ( \pi057 & \pi065 ) | ( \pi057 & ~w673 ) | ( \pi065 & ~w673 ) ;
  assign w675 = w672 | w674 ;
  assign w676 = \pi056 & \pi064 ;
  assign w677 = ~w671 & w675 ;
  assign w678 = ( \pi064 & ~w676 ) | ( \pi064 & w677 ) | ( ~w676 & w677 ) ;
  assign w679 = ~\pi065 & w670 ;
  assign w680 = w613 | w650 ;
  assign w681 = ( w590 & w650 ) | ( w590 & w680 ) | ( w650 & w680 ) ;
  assign w682 = \pi066 ^ w681 ;
  assign w683 = ( w678 & ~w679 ) | ( w678 & w682 ) | ( ~w679 & w682 ) ;
  assign w684 = w682 | w683 ;
  assign w685 = \pi067 ^ w643 ;
  assign w686 = ( ~w655 & w684 ) | ( ~w655 & w685 ) | ( w684 & w685 ) ;
  assign w687 = w685 | w686 ;
  assign w688 = \pi068 ^ w635 ;
  assign w689 = ( ~w644 & w687 ) | ( ~w644 & w688 ) | ( w687 & w688 ) ;
  assign w690 = w688 | w689 ;
  assign w691 = \pi069 ^ w629 ;
  assign w692 = ( ~w636 & w690 ) | ( ~w636 & w691 ) | ( w690 & w691 ) ;
  assign w693 = w691 | w692 ;
  assign w694 = \pi070 ^ w618 ;
  assign w695 = ( ~w630 & w693 ) | ( ~w630 & w694 ) | ( w693 & w694 ) ;
  assign w696 = w694 | w695 ;
  assign w697 = \pi071 ^ w623 ;
  assign w698 = w624 & ~w697 ;
  assign w699 = ( w696 & w697 ) | ( w696 & ~w698 ) | ( w697 & ~w698 ) ;
  assign w700 = ~\pi071 & w623 ;
  assign w701 = w699 & ~w700 ;
  assign w702 = ( w196 & ~w207 ) | ( w196 & w298 ) | ( ~w207 & w298 ) ;
  assign w703 = w207 | w702 ;
  assign w704 = w701 | w703 ;
  assign w705 = w618 & w704 ;
  assign w706 = ~w630 & w693 ;
  assign w707 = w694 ^ w706 ;
  assign w708 = ~w704 & w707 ;
  assign w709 = w705 | w708 ;
  assign w710 = ~\pi071 & w709 ;
  assign w711 = w629 & w704 ;
  assign w712 = ~w636 & w690 ;
  assign w713 = w691 ^ w712 ;
  assign w714 = ~w704 & w713 ;
  assign w715 = w711 | w714 ;
  assign w716 = ~\pi070 & w715 ;
  assign w717 = w635 & w704 ;
  assign w718 = ~w644 & w687 ;
  assign w719 = w688 ^ w718 ;
  assign w720 = ~w704 & w719 ;
  assign w721 = w717 | w720 ;
  assign w722 = ~\pi069 & w721 ;
  assign w723 = w643 & w704 ;
  assign w724 = ~w655 & w684 ;
  assign w725 = w685 ^ w724 ;
  assign w726 = ~w704 & w725 ;
  assign w727 = w723 | w726 ;
  assign w728 = ~\pi068 & w727 ;
  assign w729 = w654 & w704 ;
  assign w730 = w678 & ~w679 ;
  assign w731 = w682 ^ w730 ;
  assign w732 = ~w704 & w731 ;
  assign w733 = w729 | w732 ;
  assign w734 = ~\pi067 & w733 ;
  assign w735 = w670 & w704 ;
  assign w736 = ( ~\pi056 & \pi064 ) | ( ~\pi056 & w701 ) | ( \pi064 & w701 ) ;
  assign w737 = ( ~w671 & w675 ) | ( ~w671 & w703 ) | ( w675 & w703 ) ;
  assign w738 = w736 ^ w737 ;
  assign w739 = ( ~w701 & w703 ) | ( ~w701 & w738 ) | ( w703 & w738 ) ;
  assign w740 = ~w703 & w739 ;
  assign w741 = w735 | w740 ;
  assign w742 = ~\pi066 & w741 ;
  assign w743 = ( \pi064 & w256 ) | ( \pi064 & w444 ) | ( w256 & w444 ) ;
  assign w744 = ( \pi064 & ~\pi072 ) | ( \pi064 & w443 ) | ( ~\pi072 & w443 ) ;
  assign w745 = ~w609 & w744 ;
  assign w746 = ~w743 & w745 ;
  assign w747 = ( ~\pi056 & w132 ) | ( ~\pi056 & w142 ) | ( w132 & w142 ) ;
  assign w748 = ( ~\pi056 & \pi064 ) | ( ~\pi056 & w185 ) | ( \pi064 & w185 ) ;
  assign w749 = ~w543 & w748 ;
  assign w750 = ~w747 & w749 ;
  assign w751 = ( \pi056 & w701 ) | ( \pi056 & ~w746 ) | ( w701 & ~w746 ) ;
  assign w752 = \pi056 & w751 ;
  assign w753 = w701 | w750 ;
  assign w754 = ( ~w701 & w752 ) | ( ~w701 & w753 ) | ( w752 & w753 ) ;
  assign w755 = ~\pi055 & \pi064 ;
  assign w756 = w746 & ~w753 ;
  assign w757 = \pi056 & ~w756 ;
  assign w758 = ( ~w701 & w753 ) | ( ~w701 & w757 ) | ( w753 & w757 ) ;
  assign w759 = \pi065 ^ w758 ;
  assign w760 = w755 | w759 ;
  assign w761 = ~\pi065 & w754 ;
  assign w762 = \pi066 ^ w741 ;
  assign w763 = ( w760 & ~w761 ) | ( w760 & w762 ) | ( ~w761 & w762 ) ;
  assign w764 = w762 | w763 ;
  assign w765 = \pi067 ^ w733 ;
  assign w766 = ( ~w742 & w764 ) | ( ~w742 & w765 ) | ( w764 & w765 ) ;
  assign w767 = w765 | w766 ;
  assign w768 = \pi068 ^ w727 ;
  assign w769 = ( ~w734 & w767 ) | ( ~w734 & w768 ) | ( w767 & w768 ) ;
  assign w770 = w768 | w769 ;
  assign w771 = \pi069 ^ w721 ;
  assign w772 = ( ~w728 & w770 ) | ( ~w728 & w771 ) | ( w770 & w771 ) ;
  assign w773 = w771 | w772 ;
  assign w774 = \pi070 ^ w715 ;
  assign w775 = ( ~w722 & w773 ) | ( ~w722 & w774 ) | ( w773 & w774 ) ;
  assign w776 = w774 | w775 ;
  assign w777 = \pi071 ^ w709 ;
  assign w778 = ( ~w716 & w776 ) | ( ~w716 & w777 ) | ( w776 & w777 ) ;
  assign w779 = w777 | w778 ;
  assign w780 = w623 & w704 ;
  assign w781 = ~w624 & w696 ;
  assign w782 = w697 ^ w781 ;
  assign w783 = ~w704 & w782 ;
  assign w784 = w780 | w783 ;
  assign w785 = ~\pi072 & w784 ;
  assign w786 = ( \pi072 & ~w780 ) | ( \pi072 & w783 ) | ( ~w780 & w783 ) ;
  assign w787 = ~w783 & w786 ;
  assign w788 = w246 | w257 ;
  assign w789 = w787 | w788 ;
  assign w790 = ( w291 & w785 ) | ( w291 & ~w787 ) | ( w785 & ~w787 ) ;
  assign w791 = w789 | w790 ;
  assign w792 = ( ~w710 & w779 ) | ( ~w710 & w791 ) | ( w779 & w791 ) ;
  assign w793 = w791 | w792 ;
  assign w794 = ~w703 & w784 ;
  assign w795 = w793 & ~w794 ;
  assign w796 = ~w716 & w776 ;
  assign w797 = w777 ^ w796 ;
  assign w798 = ~w795 & w797 ;
  assign w799 = ( w709 & w793 ) | ( w709 & w794 ) | ( w793 & w794 ) ;
  assign w800 = ~w794 & w799 ;
  assign w801 = w798 | w800 ;
  assign w802 = w785 | w787 ;
  assign w803 = ( ~w710 & w779 ) | ( ~w710 & w795 ) | ( w779 & w795 ) ;
  assign w804 = w802 ^ w803 ;
  assign w805 = ~w795 & w804 ;
  assign w806 = ( w703 & ~w784 ) | ( w703 & w793 ) | ( ~w784 & w793 ) ;
  assign w807 = w784 & w806 ;
  assign w808 = w805 | w807 ;
  assign w809 = ~\pi072 & w801 ;
  assign w810 = ~w722 & w773 ;
  assign w811 = w774 ^ w810 ;
  assign w812 = ~w795 & w811 ;
  assign w813 = ( w715 & w793 ) | ( w715 & w794 ) | ( w793 & w794 ) ;
  assign w814 = ~w794 & w813 ;
  assign w815 = w812 | w814 ;
  assign w816 = ~\pi071 & w815 ;
  assign w817 = ~w728 & w770 ;
  assign w818 = w771 ^ w817 ;
  assign w819 = ~w795 & w818 ;
  assign w820 = ( w721 & w793 ) | ( w721 & w794 ) | ( w793 & w794 ) ;
  assign w821 = ~w794 & w820 ;
  assign w822 = w819 | w821 ;
  assign w823 = ~\pi070 & w822 ;
  assign w824 = ~w734 & w767 ;
  assign w825 = w768 ^ w824 ;
  assign w826 = ~w795 & w825 ;
  assign w827 = ( w727 & w793 ) | ( w727 & w794 ) | ( w793 & w794 ) ;
  assign w828 = ~w794 & w827 ;
  assign w829 = w826 | w828 ;
  assign w830 = ~\pi069 & w829 ;
  assign w831 = ~w742 & w764 ;
  assign w832 = w765 ^ w831 ;
  assign w833 = ~w795 & w832 ;
  assign w834 = ( w733 & w793 ) | ( w733 & w794 ) | ( w793 & w794 ) ;
  assign w835 = ~w794 & w834 ;
  assign w836 = w833 | w835 ;
  assign w837 = ~\pi068 & w836 ;
  assign w838 = w760 & ~w761 ;
  assign w839 = w762 ^ w838 ;
  assign w840 = ~w795 & w839 ;
  assign w841 = ( w741 & w793 ) | ( w741 & w794 ) | ( w793 & w794 ) ;
  assign w842 = ~w794 & w841 ;
  assign w843 = w840 | w842 ;
  assign w844 = ~\pi067 & w843 ;
  assign w845 = w746 & ~w750 ;
  assign w846 = w701 ^ w750 ;
  assign w847 = ( \pi056 & ~w845 ) | ( \pi056 & w846 ) | ( ~w845 & w846 ) ;
  assign w848 = ( \pi056 & w750 ) | ( \pi056 & w847 ) | ( w750 & w847 ) ;
  assign w849 = w755 ^ w848 ;
  assign w850 = \pi065 ^ w849 ;
  assign w851 = ~w795 & w850 ;
  assign w852 = ( w754 & w793 ) | ( w754 & w794 ) | ( w793 & w794 ) ;
  assign w853 = ~w794 & w852 ;
  assign w854 = w851 | w853 ;
  assign w855 = ~\pi066 & w854 ;
  assign w856 = ~\pi054 & \pi064 ;
  assign w857 = \pi066 ^ w854 ;
  assign w858 = \pi064 & ~w795 ;
  assign w859 = \pi055 ^ w858 ;
  assign w860 = ( ~\pi054 & \pi064 ) | ( ~\pi054 & w857 ) | ( \pi064 & w857 ) ;
  assign w861 = ( \pi065 & ~w859 ) | ( \pi065 & w860 ) | ( ~w859 & w860 ) ;
  assign w862 = w857 | w861 ;
  assign w863 = \pi067 ^ w843 ;
  assign w864 = ( ~w855 & w862 ) | ( ~w855 & w863 ) | ( w862 & w863 ) ;
  assign w865 = w863 | w864 ;
  assign w866 = \pi068 ^ w836 ;
  assign w867 = ( ~w844 & w865 ) | ( ~w844 & w866 ) | ( w865 & w866 ) ;
  assign w868 = w866 | w867 ;
  assign w869 = \pi069 ^ w829 ;
  assign w870 = ( ~w837 & w868 ) | ( ~w837 & w869 ) | ( w868 & w869 ) ;
  assign w871 = w869 | w870 ;
  assign w872 = \pi070 ^ w822 ;
  assign w873 = ( ~w830 & w871 ) | ( ~w830 & w872 ) | ( w871 & w872 ) ;
  assign w874 = w872 | w873 ;
  assign w875 = \pi071 ^ w815 ;
  assign w876 = ( ~w823 & w874 ) | ( ~w823 & w875 ) | ( w874 & w875 ) ;
  assign w877 = w875 | w876 ;
  assign w878 = \pi072 ^ w801 ;
  assign w879 = ( ~w816 & w877 ) | ( ~w816 & w878 ) | ( w877 & w878 ) ;
  assign w880 = w878 | w879 ;
  assign w881 = \pi073 ^ w808 ;
  assign w882 = w809 & ~w881 ;
  assign w883 = ( w880 & w881 ) | ( w880 & ~w882 ) | ( w881 & ~w882 ) ;
  assign w884 = ~\pi073 & w808 ;
  assign w885 = w883 & ~w884 ;
  assign w886 = \pi074 | \pi075 ;
  assign w887 = w207 | w886 ;
  assign w888 = ( w141 & ~w207 ) | ( w141 & w298 ) | ( ~w207 & w298 ) ;
  assign w889 = w887 | w888 ;
  assign w890 = w885 | w889 ;
  assign w891 = w801 & w890 ;
  assign w892 = ~w816 & w877 ;
  assign w893 = w878 ^ w892 ;
  assign w894 = ~w890 & w893 ;
  assign w895 = w891 | w894 ;
  assign w896 = w808 & w890 ;
  assign w897 = ~w809 & w880 ;
  assign w898 = w881 ^ w897 ;
  assign w899 = ~w890 & w898 ;
  assign w900 = w896 | w899 ;
  assign w901 = ~\pi073 & w895 ;
  assign w902 = w815 & w890 ;
  assign w903 = ~w823 & w874 ;
  assign w904 = w875 ^ w903 ;
  assign w905 = ~w890 & w904 ;
  assign w906 = w902 | w905 ;
  assign w907 = ~\pi072 & w906 ;
  assign w908 = w822 & w890 ;
  assign w909 = ~w830 & w871 ;
  assign w910 = w872 ^ w909 ;
  assign w911 = ~w890 & w910 ;
  assign w912 = w908 | w911 ;
  assign w913 = ~\pi071 & w912 ;
  assign w914 = w829 & w890 ;
  assign w915 = ~w837 & w868 ;
  assign w916 = w869 ^ w915 ;
  assign w917 = ~w890 & w916 ;
  assign w918 = w914 | w917 ;
  assign w919 = ~\pi070 & w918 ;
  assign w920 = w836 & w890 ;
  assign w921 = ~w844 & w865 ;
  assign w922 = w866 ^ w921 ;
  assign w923 = ~w890 & w922 ;
  assign w924 = w920 | w923 ;
  assign w925 = ~\pi069 & w924 ;
  assign w926 = w843 & w890 ;
  assign w927 = ~w855 & w862 ;
  assign w928 = w863 ^ w927 ;
  assign w929 = ~w890 & w928 ;
  assign w930 = w926 | w929 ;
  assign w931 = ~\pi068 & w930 ;
  assign w932 = w854 & w890 ;
  assign w933 = ( \pi065 & w856 ) | ( \pi065 & ~w859 ) | ( w856 & ~w859 ) ;
  assign w934 = w857 ^ w933 ;
  assign w935 = ( w885 & w889 ) | ( w885 & w934 ) | ( w889 & w934 ) ;
  assign w936 = w934 & ~w935 ;
  assign w937 = w932 | w936 ;
  assign w938 = ~\pi067 & w937 ;
  assign w939 = \pi055 ^ \pi065 ;
  assign w940 = \pi054 ^ w795 ;
  assign w941 = ( \pi064 & w889 ) | ( \pi064 & w940 ) | ( w889 & w940 ) ;
  assign w942 = w939 ^ w941 ;
  assign w943 = ~w889 & w942 ;
  assign w944 = ~w885 & w943 ;
  assign w945 = ( ~\pi064 & w795 ) | ( ~\pi064 & w890 ) | ( w795 & w890 ) ;
  assign w946 = \pi055 ^ w945 ;
  assign w947 = w890 & ~w946 ;
  assign w948 = w944 | w947 ;
  assign w949 = ~\pi066 & w948 ;
  assign w950 = ( \pi064 & ~\pi074 ) | ( \pi064 & \pi075 ) | ( ~\pi074 & \pi075 ) ;
  assign w951 = w246 | w253 ;
  assign w952 = ( \pi075 & \pi076 ) | ( \pi075 & ~w253 ) | ( \pi076 & ~w253 ) ;
  assign w953 = w951 | w952 ;
  assign w954 = w950 & ~w953 ;
  assign w955 = ~w291 & w954 ;
  assign w956 = ( \pi074 & ~w141 ) | ( \pi074 & w856 ) | ( ~w141 & w856 ) ;
  assign w957 = ( \pi074 & \pi075 ) | ( \pi074 & ~w207 ) | ( \pi075 & ~w207 ) ;
  assign w958 = w345 | w957 ;
  assign w959 = w956 & ~w958 ;
  assign w960 = ( \pi054 & w885 ) | ( \pi054 & ~w955 ) | ( w885 & ~w955 ) ;
  assign w961 = \pi054 & w960 ;
  assign w962 = w885 | w959 ;
  assign w963 = ( ~w885 & w961 ) | ( ~w885 & w962 ) | ( w961 & w962 ) ;
  assign w964 = ( \pi065 & ~w885 ) | ( \pi065 & w959 ) | ( ~w885 & w959 ) ;
  assign w965 = ~w885 & w955 ;
  assign w966 = ( \pi054 & \pi065 ) | ( \pi054 & ~w965 ) | ( \pi065 & ~w965 ) ;
  assign w967 = w964 | w966 ;
  assign w968 = ~\pi053 & \pi064 ;
  assign w969 = \pi065 & w963 ;
  assign w970 = w967 | w969 ;
  assign w971 = ( w968 & ~w969 ) | ( w968 & w970 ) | ( ~w969 & w970 ) ;
  assign w972 = ~\pi065 & w963 ;
  assign w973 = w890 | w944 ;
  assign w974 = ( w859 & w944 ) | ( w859 & w973 ) | ( w944 & w973 ) ;
  assign w975 = \pi066 ^ w974 ;
  assign w976 = ( w971 & ~w972 ) | ( w971 & w975 ) | ( ~w972 & w975 ) ;
  assign w977 = w975 | w976 ;
  assign w978 = \pi067 ^ w937 ;
  assign w979 = ( ~w949 & w977 ) | ( ~w949 & w978 ) | ( w977 & w978 ) ;
  assign w980 = w978 | w979 ;
  assign w981 = \pi068 ^ w930 ;
  assign w982 = ( ~w938 & w980 ) | ( ~w938 & w981 ) | ( w980 & w981 ) ;
  assign w983 = w981 | w982 ;
  assign w984 = \pi069 ^ w924 ;
  assign w985 = ( ~w931 & w983 ) | ( ~w931 & w984 ) | ( w983 & w984 ) ;
  assign w986 = w984 | w985 ;
  assign w987 = \pi070 ^ w918 ;
  assign w988 = ( ~w925 & w986 ) | ( ~w925 & w987 ) | ( w986 & w987 ) ;
  assign w989 = w987 | w988 ;
  assign w990 = \pi071 ^ w912 ;
  assign w991 = ( ~w919 & w989 ) | ( ~w919 & w990 ) | ( w989 & w990 ) ;
  assign w992 = w990 | w991 ;
  assign w993 = \pi072 ^ w906 ;
  assign w994 = ( ~w913 & w992 ) | ( ~w913 & w993 ) | ( w992 & w993 ) ;
  assign w995 = w993 | w994 ;
  assign w996 = \pi073 ^ w895 ;
  assign w997 = ( ~w907 & w995 ) | ( ~w907 & w996 ) | ( w995 & w996 ) ;
  assign w998 = w996 | w997 ;
  assign w999 = \pi074 ^ w900 ;
  assign w1000 = w901 & ~w999 ;
  assign w1001 = ( w998 & w999 ) | ( w998 & ~w1000 ) | ( w999 & ~w1000 ) ;
  assign w1002 = ~\pi074 & w900 ;
  assign w1003 = w1001 & ~w1002 ;
  assign w1004 = \pi075 | \pi076 ;
  assign w1005 = w246 | w1004 ;
  assign w1006 = ( ~w246 & w253 ) | ( ~w246 & w291 ) | ( w253 & w291 ) ;
  assign w1007 = w1005 | w1006 ;
  assign w1008 = w1003 | w1007 ;
  assign w1009 = w895 & w1008 ;
  assign w1010 = ~w907 & w995 ;
  assign w1011 = w996 ^ w1010 ;
  assign w1012 = ~w1008 & w1011 ;
  assign w1013 = w1009 | w1012 ;
  assign w1014 = ~\pi074 & w1013 ;
  assign w1015 = w906 & w1008 ;
  assign w1016 = ~w913 & w992 ;
  assign w1017 = w993 ^ w1016 ;
  assign w1018 = ~w1008 & w1017 ;
  assign w1019 = w1015 | w1018 ;
  assign w1020 = ~\pi073 & w1019 ;
  assign w1021 = w912 & w1008 ;
  assign w1022 = ~w919 & w989 ;
  assign w1023 = w990 ^ w1022 ;
  assign w1024 = ~w1008 & w1023 ;
  assign w1025 = w1021 | w1024 ;
  assign w1026 = ~\pi072 & w1025 ;
  assign w1027 = w918 & w1008 ;
  assign w1028 = ~w925 & w986 ;
  assign w1029 = w987 ^ w1028 ;
  assign w1030 = ~w1008 & w1029 ;
  assign w1031 = w1027 | w1030 ;
  assign w1032 = ~\pi071 & w1031 ;
  assign w1033 = w924 & w1008 ;
  assign w1034 = ~w931 & w983 ;
  assign w1035 = w984 ^ w1034 ;
  assign w1036 = ~w1008 & w1035 ;
  assign w1037 = w1033 | w1036 ;
  assign w1038 = ~\pi070 & w1037 ;
  assign w1039 = w930 & w1008 ;
  assign w1040 = ~w938 & w980 ;
  assign w1041 = w981 ^ w1040 ;
  assign w1042 = ~w1008 & w1041 ;
  assign w1043 = w1039 | w1042 ;
  assign w1044 = ~\pi069 & w1043 ;
  assign w1045 = w937 & w1008 ;
  assign w1046 = ~w949 & w977 ;
  assign w1047 = w978 ^ w1046 ;
  assign w1048 = ~w1008 & w1047 ;
  assign w1049 = w1045 | w1048 ;
  assign w1050 = ~\pi068 & w1049 ;
  assign w1051 = w948 & w1008 ;
  assign w1052 = w971 & ~w972 ;
  assign w1053 = w975 ^ w1052 ;
  assign w1054 = ~w1008 & w1053 ;
  assign w1055 = w1051 | w1054 ;
  assign w1056 = ~\pi067 & w1055 ;
  assign w1057 = w963 & w1008 ;
  assign w1058 = ~w963 & w967 ;
  assign w1059 = ( ~\pi065 & w967 ) | ( ~\pi065 & w1058 ) | ( w967 & w1058 ) ;
  assign w1060 = w968 ^ w1059 ;
  assign w1061 = ~w1008 & w1060 ;
  assign w1062 = w1057 | w1061 ;
  assign w1063 = ~\pi066 & w1062 ;
  assign w1064 = \pi064 & ~\pi075 ;
  assign w1065 = ~w207 & w1064 ;
  assign w1066 = ~w888 & w1065 ;
  assign w1067 = ( \pi075 & ~w253 ) | ( \pi075 & w968 ) | ( ~w253 & w968 ) ;
  assign w1068 = ( \pi075 & \pi076 ) | ( \pi075 & ~w246 ) | ( \pi076 & ~w246 ) ;
  assign w1069 = w350 | w1068 ;
  assign w1070 = w1067 & ~w1069 ;
  assign w1071 = ( \pi053 & w1003 ) | ( \pi053 & ~w1066 ) | ( w1003 & ~w1066 ) ;
  assign w1072 = \pi053 & w1071 ;
  assign w1073 = w1003 | w1070 ;
  assign w1074 = ( ~w1003 & w1072 ) | ( ~w1003 & w1073 ) | ( w1072 & w1073 ) ;
  assign w1075 = ~\pi052 & \pi064 ;
  assign w1076 = w1066 & ~w1073 ;
  assign w1077 = \pi053 & ~w1076 ;
  assign w1078 = ( ~w1003 & w1073 ) | ( ~w1003 & w1077 ) | ( w1073 & w1077 ) ;
  assign w1079 = \pi065 ^ w1078 ;
  assign w1080 = w1075 | w1079 ;
  assign w1081 = ~\pi065 & w1074 ;
  assign w1082 = \pi066 ^ w1062 ;
  assign w1083 = ( w1080 & ~w1081 ) | ( w1080 & w1082 ) | ( ~w1081 & w1082 ) ;
  assign w1084 = w1082 | w1083 ;
  assign w1085 = \pi067 ^ w1055 ;
  assign w1086 = ( ~w1063 & w1084 ) | ( ~w1063 & w1085 ) | ( w1084 & w1085 ) ;
  assign w1087 = w1085 | w1086 ;
  assign w1088 = \pi068 ^ w1049 ;
  assign w1089 = ( ~w1056 & w1087 ) | ( ~w1056 & w1088 ) | ( w1087 & w1088 ) ;
  assign w1090 = w1088 | w1089 ;
  assign w1091 = \pi069 ^ w1043 ;
  assign w1092 = ( ~w1050 & w1090 ) | ( ~w1050 & w1091 ) | ( w1090 & w1091 ) ;
  assign w1093 = w1091 | w1092 ;
  assign w1094 = \pi070 ^ w1037 ;
  assign w1095 = ( ~w1044 & w1093 ) | ( ~w1044 & w1094 ) | ( w1093 & w1094 ) ;
  assign w1096 = w1094 | w1095 ;
  assign w1097 = \pi071 ^ w1031 ;
  assign w1098 = ( ~w1038 & w1096 ) | ( ~w1038 & w1097 ) | ( w1096 & w1097 ) ;
  assign w1099 = w1097 | w1098 ;
  assign w1100 = \pi072 ^ w1025 ;
  assign w1101 = ( ~w1032 & w1099 ) | ( ~w1032 & w1100 ) | ( w1099 & w1100 ) ;
  assign w1102 = w1100 | w1101 ;
  assign w1103 = \pi073 ^ w1019 ;
  assign w1104 = ( ~w1026 & w1102 ) | ( ~w1026 & w1103 ) | ( w1102 & w1103 ) ;
  assign w1105 = w1103 | w1104 ;
  assign w1106 = \pi074 ^ w1013 ;
  assign w1107 = ( ~w1020 & w1105 ) | ( ~w1020 & w1106 ) | ( w1105 & w1106 ) ;
  assign w1108 = w1106 | w1107 ;
  assign w1109 = w900 & w1008 ;
  assign w1110 = ~w901 & w998 ;
  assign w1111 = w999 ^ w1110 ;
  assign w1112 = ~w1008 & w1111 ;
  assign w1113 = w1109 | w1112 ;
  assign w1114 = ~\pi075 & w1113 ;
  assign w1115 = ( \pi075 & ~w1109 ) | ( \pi075 & w1112 ) | ( ~w1109 & w1112 ) ;
  assign w1116 = ~w1112 & w1115 ;
  assign w1117 = w142 | w185 ;
  assign w1118 = w1116 | w1117 ;
  assign w1119 = ( w368 & w1114 ) | ( w368 & ~w1116 ) | ( w1114 & ~w1116 ) ;
  assign w1120 = w1118 | w1119 ;
  assign w1121 = ( ~w1014 & w1108 ) | ( ~w1014 & w1120 ) | ( w1108 & w1120 ) ;
  assign w1122 = w1120 | w1121 ;
  assign w1123 = ~w1007 & w1113 ;
  assign w1124 = w1122 & ~w1123 ;
  assign w1125 = ~w1020 & w1105 ;
  assign w1126 = w1106 ^ w1125 ;
  assign w1127 = ~w1124 & w1126 ;
  assign w1128 = ( w1013 & w1122 ) | ( w1013 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1129 = ~w1123 & w1128 ;
  assign w1130 = w1127 | w1129 ;
  assign w1131 = w1114 | w1116 ;
  assign w1132 = ( ~w1014 & w1108 ) | ( ~w1014 & w1124 ) | ( w1108 & w1124 ) ;
  assign w1133 = w1131 ^ w1132 ;
  assign w1134 = ~w1124 & w1133 ;
  assign w1135 = ( w1007 & ~w1113 ) | ( w1007 & w1122 ) | ( ~w1113 & w1122 ) ;
  assign w1136 = w1113 & w1135 ;
  assign w1137 = w1134 | w1136 ;
  assign w1138 = ~\pi075 & w1130 ;
  assign w1139 = ~w1026 & w1102 ;
  assign w1140 = w1103 ^ w1139 ;
  assign w1141 = ~w1124 & w1140 ;
  assign w1142 = ( w1019 & w1122 ) | ( w1019 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1143 = ~w1123 & w1142 ;
  assign w1144 = w1141 | w1143 ;
  assign w1145 = ~\pi074 & w1144 ;
  assign w1146 = ~w1032 & w1099 ;
  assign w1147 = w1100 ^ w1146 ;
  assign w1148 = ~w1124 & w1147 ;
  assign w1149 = ( w1025 & w1122 ) | ( w1025 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1150 = ~w1123 & w1149 ;
  assign w1151 = w1148 | w1150 ;
  assign w1152 = ~\pi073 & w1151 ;
  assign w1153 = ~w1038 & w1096 ;
  assign w1154 = w1097 ^ w1153 ;
  assign w1155 = ~w1124 & w1154 ;
  assign w1156 = ( w1031 & w1122 ) | ( w1031 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1157 = ~w1123 & w1156 ;
  assign w1158 = w1155 | w1157 ;
  assign w1159 = ~\pi072 & w1158 ;
  assign w1160 = ~w1044 & w1093 ;
  assign w1161 = w1094 ^ w1160 ;
  assign w1162 = ~w1124 & w1161 ;
  assign w1163 = ( w1037 & w1122 ) | ( w1037 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1164 = ~w1123 & w1163 ;
  assign w1165 = w1162 | w1164 ;
  assign w1166 = ~\pi071 & w1165 ;
  assign w1167 = ~w1050 & w1090 ;
  assign w1168 = w1091 ^ w1167 ;
  assign w1169 = ~w1124 & w1168 ;
  assign w1170 = ( w1043 & w1122 ) | ( w1043 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1171 = ~w1123 & w1170 ;
  assign w1172 = w1169 | w1171 ;
  assign w1173 = ~\pi070 & w1172 ;
  assign w1174 = ~w1056 & w1087 ;
  assign w1175 = w1088 ^ w1174 ;
  assign w1176 = ~w1124 & w1175 ;
  assign w1177 = ( w1049 & w1122 ) | ( w1049 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1178 = ~w1123 & w1177 ;
  assign w1179 = w1176 | w1178 ;
  assign w1180 = ~\pi069 & w1179 ;
  assign w1181 = ~w1063 & w1084 ;
  assign w1182 = w1085 ^ w1181 ;
  assign w1183 = ~w1124 & w1182 ;
  assign w1184 = ( w1055 & w1122 ) | ( w1055 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1185 = ~w1123 & w1184 ;
  assign w1186 = w1183 | w1185 ;
  assign w1187 = ~\pi068 & w1186 ;
  assign w1188 = w1080 & ~w1081 ;
  assign w1189 = w1082 ^ w1188 ;
  assign w1190 = ~w1124 & w1189 ;
  assign w1191 = ( w1062 & w1122 ) | ( w1062 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1192 = ~w1123 & w1191 ;
  assign w1193 = w1190 | w1192 ;
  assign w1194 = ~\pi067 & w1193 ;
  assign w1195 = w1066 & ~w1070 ;
  assign w1196 = w1003 ^ w1070 ;
  assign w1197 = ( \pi053 & ~w1195 ) | ( \pi053 & w1196 ) | ( ~w1195 & w1196 ) ;
  assign w1198 = ( \pi053 & w1070 ) | ( \pi053 & w1197 ) | ( w1070 & w1197 ) ;
  assign w1199 = w1075 ^ w1198 ;
  assign w1200 = \pi065 ^ w1199 ;
  assign w1201 = ~w1124 & w1200 ;
  assign w1202 = ( w1074 & w1122 ) | ( w1074 & w1123 ) | ( w1122 & w1123 ) ;
  assign w1203 = ~w1123 & w1202 ;
  assign w1204 = w1201 | w1203 ;
  assign w1205 = ~\pi066 & w1204 ;
  assign w1206 = \pi066 ^ w1204 ;
  assign w1207 = \pi064 & ~w1124 ;
  assign w1208 = \pi052 ^ w1207 ;
  assign w1209 = ( ~\pi051 & \pi064 ) | ( ~\pi051 & w1206 ) | ( \pi064 & w1206 ) ;
  assign w1210 = ( \pi065 & ~w1208 ) | ( \pi065 & w1209 ) | ( ~w1208 & w1209 ) ;
  assign w1211 = w1206 | w1210 ;
  assign w1212 = \pi067 ^ w1193 ;
  assign w1213 = ( ~w1205 & w1211 ) | ( ~w1205 & w1212 ) | ( w1211 & w1212 ) ;
  assign w1214 = w1212 | w1213 ;
  assign w1215 = \pi068 ^ w1186 ;
  assign w1216 = ( ~w1194 & w1214 ) | ( ~w1194 & w1215 ) | ( w1214 & w1215 ) ;
  assign w1217 = w1215 | w1216 ;
  assign w1218 = \pi069 ^ w1179 ;
  assign w1219 = ( ~w1187 & w1217 ) | ( ~w1187 & w1218 ) | ( w1217 & w1218 ) ;
  assign w1220 = w1218 | w1219 ;
  assign w1221 = \pi070 ^ w1172 ;
  assign w1222 = ( ~w1180 & w1220 ) | ( ~w1180 & w1221 ) | ( w1220 & w1221 ) ;
  assign w1223 = w1221 | w1222 ;
  assign w1224 = \pi071 ^ w1165 ;
  assign w1225 = ( ~w1173 & w1223 ) | ( ~w1173 & w1224 ) | ( w1223 & w1224 ) ;
  assign w1226 = w1224 | w1225 ;
  assign w1227 = \pi072 ^ w1158 ;
  assign w1228 = ( ~w1166 & w1226 ) | ( ~w1166 & w1227 ) | ( w1226 & w1227 ) ;
  assign w1229 = w1227 | w1228 ;
  assign w1230 = \pi073 ^ w1151 ;
  assign w1231 = ( ~w1159 & w1229 ) | ( ~w1159 & w1230 ) | ( w1229 & w1230 ) ;
  assign w1232 = w1230 | w1231 ;
  assign w1233 = \pi074 ^ w1144 ;
  assign w1234 = ( ~w1152 & w1232 ) | ( ~w1152 & w1233 ) | ( w1232 & w1233 ) ;
  assign w1235 = w1233 | w1234 ;
  assign w1236 = \pi075 ^ w1130 ;
  assign w1237 = ( ~w1145 & w1235 ) | ( ~w1145 & w1236 ) | ( w1235 & w1236 ) ;
  assign w1238 = w1236 | w1237 ;
  assign w1239 = \pi076 ^ w1137 ;
  assign w1240 = w1138 & ~w1239 ;
  assign w1241 = ( w1238 & w1239 ) | ( w1238 & ~w1240 ) | ( w1239 & ~w1240 ) ;
  assign w1242 = ~\pi076 & w1137 ;
  assign w1243 = w1241 & ~w1242 ;
  assign w1244 = ( ~w443 & w444 ) | ( ~w443 & w452 ) | ( w444 & w452 ) ;
  assign w1245 = w443 | w1244 ;
  assign w1246 = w1243 | w1245 ;
  assign w1247 = w1130 & w1246 ;
  assign w1248 = ~w1145 & w1235 ;
  assign w1249 = w1236 ^ w1248 ;
  assign w1250 = ~w1246 & w1249 ;
  assign w1251 = w1247 | w1250 ;
  assign w1252 = w1137 & w1246 ;
  assign w1253 = ~w1138 & w1238 ;
  assign w1254 = w1239 ^ w1253 ;
  assign w1255 = ~w1246 & w1254 ;
  assign w1256 = w1252 | w1255 ;
  assign w1257 = ~\pi076 & w1251 ;
  assign w1258 = w1144 & w1246 ;
  assign w1259 = ~w1152 & w1232 ;
  assign w1260 = w1233 ^ w1259 ;
  assign w1261 = ~w1246 & w1260 ;
  assign w1262 = w1258 | w1261 ;
  assign w1263 = ~\pi075 & w1262 ;
  assign w1264 = w1151 & w1246 ;
  assign w1265 = ~w1159 & w1229 ;
  assign w1266 = w1230 ^ w1265 ;
  assign w1267 = ~w1246 & w1266 ;
  assign w1268 = w1264 | w1267 ;
  assign w1269 = ~\pi074 & w1268 ;
  assign w1270 = w1158 & w1246 ;
  assign w1271 = ~w1166 & w1226 ;
  assign w1272 = w1227 ^ w1271 ;
  assign w1273 = ~w1246 & w1272 ;
  assign w1274 = w1270 | w1273 ;
  assign w1275 = ~\pi073 & w1274 ;
  assign w1276 = w1165 & w1246 ;
  assign w1277 = ~w1173 & w1223 ;
  assign w1278 = w1224 ^ w1277 ;
  assign w1279 = ~w1246 & w1278 ;
  assign w1280 = w1276 | w1279 ;
  assign w1281 = ~\pi072 & w1280 ;
  assign w1282 = w1172 & w1246 ;
  assign w1283 = ~w1180 & w1220 ;
  assign w1284 = w1221 ^ w1283 ;
  assign w1285 = ~w1246 & w1284 ;
  assign w1286 = w1282 | w1285 ;
  assign w1287 = ~\pi071 & w1286 ;
  assign w1288 = w1179 & w1246 ;
  assign w1289 = ~w1187 & w1217 ;
  assign w1290 = w1218 ^ w1289 ;
  assign w1291 = ~w1246 & w1290 ;
  assign w1292 = w1288 | w1291 ;
  assign w1293 = ~\pi070 & w1292 ;
  assign w1294 = w1186 & w1246 ;
  assign w1295 = ~w1194 & w1214 ;
  assign w1296 = w1215 ^ w1295 ;
  assign w1297 = ~w1246 & w1296 ;
  assign w1298 = w1294 | w1297 ;
  assign w1299 = ~\pi069 & w1298 ;
  assign w1300 = w1193 & w1246 ;
  assign w1301 = ~w1205 & w1211 ;
  assign w1302 = w1212 ^ w1301 ;
  assign w1303 = ~w1246 & w1302 ;
  assign w1304 = w1300 | w1303 ;
  assign w1305 = ~\pi068 & w1304 ;
  assign w1306 = w1204 & w1246 ;
  assign w1307 = ~\pi051 & \pi064 ;
  assign w1308 = ( \pi065 & ~w1208 ) | ( \pi065 & w1307 ) | ( ~w1208 & w1307 ) ;
  assign w1309 = w1206 ^ w1308 ;
  assign w1310 = ( w1243 & w1245 ) | ( w1243 & w1309 ) | ( w1245 & w1309 ) ;
  assign w1311 = w1309 & ~w1310 ;
  assign w1312 = w1306 | w1311 ;
  assign w1313 = ~\pi067 & w1312 ;
  assign w1314 = \pi052 ^ \pi065 ;
  assign w1315 = \pi051 ^ w1124 ;
  assign w1316 = ( \pi064 & w1245 ) | ( \pi064 & w1315 ) | ( w1245 & w1315 ) ;
  assign w1317 = w1314 ^ w1316 ;
  assign w1318 = ~w1245 & w1317 ;
  assign w1319 = ~w1243 & w1318 ;
  assign w1320 = ( ~\pi064 & w1124 ) | ( ~\pi064 & w1246 ) | ( w1124 & w1246 ) ;
  assign w1321 = \pi052 ^ w1320 ;
  assign w1322 = w1246 & ~w1321 ;
  assign w1323 = w1319 | w1322 ;
  assign w1324 = ~\pi066 & w1323 ;
  assign w1325 = ( \pi064 & ~\pi077 ) | ( \pi064 & \pi078 ) | ( ~\pi077 & \pi078 ) ;
  assign w1326 = w138 | w185 ;
  assign w1327 = ( \pi078 & \pi079 ) | ( \pi078 & ~w138 ) | ( \pi079 & ~w138 ) ;
  assign w1328 = w1326 | w1327 ;
  assign w1329 = w1325 & ~w1328 ;
  assign w1330 = ~w368 & w1329 ;
  assign w1331 = ( \pi051 & w1243 ) | ( \pi051 & ~w1330 ) | ( w1243 & ~w1330 ) ;
  assign w1332 = \pi051 & w1331 ;
  assign w1333 = ~w246 & w1307 ;
  assign w1334 = ~w1006 & w1333 ;
  assign w1335 = ~w1243 & w1334 ;
  assign w1336 = w1332 | w1335 ;
  assign w1337 = ~\pi050 & \pi064 ;
  assign w1338 = \pi065 ^ w1336 ;
  assign w1339 = w1337 | w1338 ;
  assign w1340 = ~\pi065 & w1336 ;
  assign w1341 = w1246 | w1319 ;
  assign w1342 = ( w1208 & w1319 ) | ( w1208 & w1341 ) | ( w1319 & w1341 ) ;
  assign w1343 = \pi066 ^ w1342 ;
  assign w1344 = ( w1339 & ~w1340 ) | ( w1339 & w1343 ) | ( ~w1340 & w1343 ) ;
  assign w1345 = w1343 | w1344 ;
  assign w1346 = \pi067 ^ w1312 ;
  assign w1347 = ( ~w1324 & w1345 ) | ( ~w1324 & w1346 ) | ( w1345 & w1346 ) ;
  assign w1348 = w1346 | w1347 ;
  assign w1349 = \pi068 ^ w1304 ;
  assign w1350 = ( ~w1313 & w1348 ) | ( ~w1313 & w1349 ) | ( w1348 & w1349 ) ;
  assign w1351 = w1349 | w1350 ;
  assign w1352 = \pi069 ^ w1298 ;
  assign w1353 = ( ~w1305 & w1351 ) | ( ~w1305 & w1352 ) | ( w1351 & w1352 ) ;
  assign w1354 = w1352 | w1353 ;
  assign w1355 = \pi070 ^ w1292 ;
  assign w1356 = ( ~w1299 & w1354 ) | ( ~w1299 & w1355 ) | ( w1354 & w1355 ) ;
  assign w1357 = w1355 | w1356 ;
  assign w1358 = \pi071 ^ w1286 ;
  assign w1359 = ( ~w1293 & w1357 ) | ( ~w1293 & w1358 ) | ( w1357 & w1358 ) ;
  assign w1360 = w1358 | w1359 ;
  assign w1361 = \pi072 ^ w1280 ;
  assign w1362 = ( ~w1287 & w1360 ) | ( ~w1287 & w1361 ) | ( w1360 & w1361 ) ;
  assign w1363 = w1361 | w1362 ;
  assign w1364 = \pi073 ^ w1274 ;
  assign w1365 = ( ~w1281 & w1363 ) | ( ~w1281 & w1364 ) | ( w1363 & w1364 ) ;
  assign w1366 = w1364 | w1365 ;
  assign w1367 = \pi074 ^ w1268 ;
  assign w1368 = ( ~w1275 & w1366 ) | ( ~w1275 & w1367 ) | ( w1366 & w1367 ) ;
  assign w1369 = w1367 | w1368 ;
  assign w1370 = \pi075 ^ w1262 ;
  assign w1371 = ( ~w1269 & w1369 ) | ( ~w1269 & w1370 ) | ( w1369 & w1370 ) ;
  assign w1372 = w1370 | w1371 ;
  assign w1373 = \pi076 ^ w1251 ;
  assign w1374 = ( ~w1263 & w1372 ) | ( ~w1263 & w1373 ) | ( w1372 & w1373 ) ;
  assign w1375 = w1373 | w1374 ;
  assign w1376 = \pi077 ^ w1256 ;
  assign w1377 = w1257 & ~w1376 ;
  assign w1378 = ( w1375 & w1376 ) | ( w1375 & ~w1377 ) | ( w1376 & ~w1377 ) ;
  assign w1379 = ~\pi077 & w1256 ;
  assign w1380 = w1378 & ~w1379 ;
  assign w1381 = \pi078 | \pi079 ;
  assign w1382 = w185 | w1381 ;
  assign w1383 = ( w138 & ~w185 ) | ( w138 & w368 ) | ( ~w185 & w368 ) ;
  assign w1384 = w1382 | w1383 ;
  assign w1385 = w1380 | w1384 ;
  assign w1386 = w1251 & w1385 ;
  assign w1387 = ~w1263 & w1372 ;
  assign w1388 = w1373 ^ w1387 ;
  assign w1389 = ~w1385 & w1388 ;
  assign w1390 = w1386 | w1389 ;
  assign w1391 = ~\pi077 & w1390 ;
  assign w1392 = w1262 & w1385 ;
  assign w1393 = ~w1269 & w1369 ;
  assign w1394 = w1370 ^ w1393 ;
  assign w1395 = ~w1385 & w1394 ;
  assign w1396 = w1392 | w1395 ;
  assign w1397 = ~\pi076 & w1396 ;
  assign w1398 = w1268 & w1385 ;
  assign w1399 = ~w1275 & w1366 ;
  assign w1400 = w1367 ^ w1399 ;
  assign w1401 = ~w1385 & w1400 ;
  assign w1402 = w1398 | w1401 ;
  assign w1403 = ~\pi075 & w1402 ;
  assign w1404 = w1274 & w1385 ;
  assign w1405 = ~w1281 & w1363 ;
  assign w1406 = w1364 ^ w1405 ;
  assign w1407 = ~w1385 & w1406 ;
  assign w1408 = w1404 | w1407 ;
  assign w1409 = ~\pi074 & w1408 ;
  assign w1410 = w1280 & w1385 ;
  assign w1411 = ~w1287 & w1360 ;
  assign w1412 = w1361 ^ w1411 ;
  assign w1413 = ~w1385 & w1412 ;
  assign w1414 = w1410 | w1413 ;
  assign w1415 = ~\pi073 & w1414 ;
  assign w1416 = w1286 & w1385 ;
  assign w1417 = ~w1293 & w1357 ;
  assign w1418 = w1358 ^ w1417 ;
  assign w1419 = ~w1385 & w1418 ;
  assign w1420 = w1416 | w1419 ;
  assign w1421 = ~\pi072 & w1420 ;
  assign w1422 = w1292 & w1385 ;
  assign w1423 = ~w1299 & w1354 ;
  assign w1424 = w1355 ^ w1423 ;
  assign w1425 = ~w1385 & w1424 ;
  assign w1426 = w1422 | w1425 ;
  assign w1427 = ~\pi071 & w1426 ;
  assign w1428 = w1298 & w1385 ;
  assign w1429 = ~w1305 & w1351 ;
  assign w1430 = w1352 ^ w1429 ;
  assign w1431 = ~w1385 & w1430 ;
  assign w1432 = w1428 | w1431 ;
  assign w1433 = ~\pi070 & w1432 ;
  assign w1434 = w1304 & w1385 ;
  assign w1435 = ~w1313 & w1348 ;
  assign w1436 = w1349 ^ w1435 ;
  assign w1437 = ~w1385 & w1436 ;
  assign w1438 = w1434 | w1437 ;
  assign w1439 = ~\pi069 & w1438 ;
  assign w1440 = w1312 & w1385 ;
  assign w1441 = ~w1324 & w1345 ;
  assign w1442 = w1346 ^ w1441 ;
  assign w1443 = ~w1385 & w1442 ;
  assign w1444 = w1440 | w1443 ;
  assign w1445 = ~\pi068 & w1444 ;
  assign w1446 = w1323 & w1385 ;
  assign w1447 = w1339 & ~w1340 ;
  assign w1448 = w1343 ^ w1447 ;
  assign w1449 = ~w1385 & w1448 ;
  assign w1450 = w1446 | w1449 ;
  assign w1451 = ~\pi067 & w1450 ;
  assign w1452 = w1336 & w1385 ;
  assign w1453 = ( w1332 & w1335 ) | ( w1332 & ~w1384 ) | ( w1335 & ~w1384 ) ;
  assign w1454 = \pi065 ^ w1453 ;
  assign w1455 = ( w1337 & ~w1384 ) | ( w1337 & w1454 ) | ( ~w1384 & w1454 ) ;
  assign w1456 = ( w1337 & w1380 ) | ( w1337 & w1454 ) | ( w1380 & w1454 ) ;
  assign w1457 = w1455 & ~w1456 ;
  assign w1458 = w1452 | w1457 ;
  assign w1459 = ~\pi066 & w1458 ;
  assign w1460 = ( \pi064 & ~\pi078 ) | ( \pi064 & \pi079 ) | ( ~\pi078 & \pi079 ) ;
  assign w1461 = w237 | w443 ;
  assign w1462 = ( \pi079 & \pi080 ) | ( \pi079 & ~w237 ) | ( \pi080 & ~w237 ) ;
  assign w1463 = w1461 | w1462 ;
  assign w1464 = w1460 & ~w1463 ;
  assign w1465 = ~w452 & w1464 ;
  assign w1466 = ( \pi078 & ~w138 ) | ( \pi078 & w1337 ) | ( ~w138 & w1337 ) ;
  assign w1467 = ( \pi078 & \pi079 ) | ( \pi078 & ~w185 ) | ( \pi079 & ~w185 ) ;
  assign w1468 = w543 | w1467 ;
  assign w1469 = w1466 & ~w1468 ;
  assign w1470 = ( \pi050 & w1380 ) | ( \pi050 & ~w1465 ) | ( w1380 & ~w1465 ) ;
  assign w1471 = \pi050 & w1470 ;
  assign w1472 = w1380 | w1469 ;
  assign w1473 = ( ~w1380 & w1471 ) | ( ~w1380 & w1472 ) | ( w1471 & w1472 ) ;
  assign w1474 = ~\pi049 & \pi064 ;
  assign w1475 = w1465 & ~w1472 ;
  assign w1476 = \pi050 & ~w1475 ;
  assign w1477 = ( ~w1380 & w1472 ) | ( ~w1380 & w1476 ) | ( w1472 & w1476 ) ;
  assign w1478 = \pi065 ^ w1477 ;
  assign w1479 = w1474 | w1478 ;
  assign w1480 = ~\pi065 & w1473 ;
  assign w1481 = \pi066 ^ w1458 ;
  assign w1482 = ( w1479 & ~w1480 ) | ( w1479 & w1481 ) | ( ~w1480 & w1481 ) ;
  assign w1483 = w1481 | w1482 ;
  assign w1484 = \pi067 ^ w1450 ;
  assign w1485 = ( ~w1459 & w1483 ) | ( ~w1459 & w1484 ) | ( w1483 & w1484 ) ;
  assign w1486 = w1484 | w1485 ;
  assign w1487 = \pi068 ^ w1444 ;
  assign w1488 = ( ~w1451 & w1486 ) | ( ~w1451 & w1487 ) | ( w1486 & w1487 ) ;
  assign w1489 = w1487 | w1488 ;
  assign w1490 = \pi069 ^ w1438 ;
  assign w1491 = ( ~w1445 & w1489 ) | ( ~w1445 & w1490 ) | ( w1489 & w1490 ) ;
  assign w1492 = w1490 | w1491 ;
  assign w1493 = \pi070 ^ w1432 ;
  assign w1494 = ( ~w1439 & w1492 ) | ( ~w1439 & w1493 ) | ( w1492 & w1493 ) ;
  assign w1495 = w1493 | w1494 ;
  assign w1496 = \pi071 ^ w1426 ;
  assign w1497 = ( ~w1433 & w1495 ) | ( ~w1433 & w1496 ) | ( w1495 & w1496 ) ;
  assign w1498 = w1496 | w1497 ;
  assign w1499 = \pi072 ^ w1420 ;
  assign w1500 = ( ~w1427 & w1498 ) | ( ~w1427 & w1499 ) | ( w1498 & w1499 ) ;
  assign w1501 = w1499 | w1500 ;
  assign w1502 = \pi073 ^ w1414 ;
  assign w1503 = ( ~w1421 & w1501 ) | ( ~w1421 & w1502 ) | ( w1501 & w1502 ) ;
  assign w1504 = w1502 | w1503 ;
  assign w1505 = \pi074 ^ w1408 ;
  assign w1506 = ( ~w1415 & w1504 ) | ( ~w1415 & w1505 ) | ( w1504 & w1505 ) ;
  assign w1507 = w1505 | w1506 ;
  assign w1508 = \pi075 ^ w1402 ;
  assign w1509 = ( ~w1409 & w1507 ) | ( ~w1409 & w1508 ) | ( w1507 & w1508 ) ;
  assign w1510 = w1508 | w1509 ;
  assign w1511 = \pi076 ^ w1396 ;
  assign w1512 = ( ~w1403 & w1510 ) | ( ~w1403 & w1511 ) | ( w1510 & w1511 ) ;
  assign w1513 = w1511 | w1512 ;
  assign w1514 = \pi077 ^ w1390 ;
  assign w1515 = ( ~w1397 & w1513 ) | ( ~w1397 & w1514 ) | ( w1513 & w1514 ) ;
  assign w1516 = w1514 | w1515 ;
  assign w1517 = w1256 & w1385 ;
  assign w1518 = ~w1257 & w1375 ;
  assign w1519 = w1376 ^ w1518 ;
  assign w1520 = ~w1385 & w1519 ;
  assign w1521 = w1517 | w1520 ;
  assign w1522 = ~\pi078 & w1521 ;
  assign w1523 = ( \pi078 & ~w1517 ) | ( \pi078 & w1520 ) | ( ~w1517 & w1520 ) ;
  assign w1524 = ~w1520 & w1523 ;
  assign w1525 = \pi079 | \pi080 ;
  assign w1526 = w443 | w1525 ;
  assign w1527 = ( w237 & ~w443 ) | ( w237 & w452 ) | ( ~w443 & w452 ) ;
  assign w1528 = w1526 | w1527 ;
  assign w1529 = w1522 | w1524 ;
  assign w1530 = ( ~w1391 & w1516 ) | ( ~w1391 & w1529 ) | ( w1516 & w1529 ) ;
  assign w1531 = ( w1528 & ~w1529 ) | ( w1528 & w1530 ) | ( ~w1529 & w1530 ) ;
  assign w1532 = w1529 | w1531 ;
  assign w1533 = ~w1384 & w1521 ;
  assign w1534 = w1532 & ~w1533 ;
  assign w1535 = ~w1397 & w1513 ;
  assign w1536 = w1514 ^ w1535 ;
  assign w1537 = ~w1534 & w1536 ;
  assign w1538 = ( w1390 & w1532 ) | ( w1390 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1539 = ~w1533 & w1538 ;
  assign w1540 = w1537 | w1539 ;
  assign w1541 = ( ~w1391 & w1516 ) | ( ~w1391 & w1534 ) | ( w1516 & w1534 ) ;
  assign w1542 = w1529 ^ w1541 ;
  assign w1543 = ~w1534 & w1542 ;
  assign w1544 = ( w1384 & ~w1521 ) | ( w1384 & w1532 ) | ( ~w1521 & w1532 ) ;
  assign w1545 = w1521 & w1544 ;
  assign w1546 = w1543 | w1545 ;
  assign w1547 = ~\pi078 & w1540 ;
  assign w1548 = ~w1403 & w1510 ;
  assign w1549 = w1511 ^ w1548 ;
  assign w1550 = ~w1534 & w1549 ;
  assign w1551 = ( w1396 & w1532 ) | ( w1396 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1552 = ~w1533 & w1551 ;
  assign w1553 = w1550 | w1552 ;
  assign w1554 = ~\pi077 & w1553 ;
  assign w1555 = ~w1409 & w1507 ;
  assign w1556 = w1508 ^ w1555 ;
  assign w1557 = ~w1534 & w1556 ;
  assign w1558 = ( w1402 & w1532 ) | ( w1402 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1559 = ~w1533 & w1558 ;
  assign w1560 = w1557 | w1559 ;
  assign w1561 = ~\pi076 & w1560 ;
  assign w1562 = ~w1415 & w1504 ;
  assign w1563 = w1505 ^ w1562 ;
  assign w1564 = ~w1534 & w1563 ;
  assign w1565 = ( w1408 & w1532 ) | ( w1408 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1566 = ~w1533 & w1565 ;
  assign w1567 = w1564 | w1566 ;
  assign w1568 = ~\pi075 & w1567 ;
  assign w1569 = ~w1421 & w1501 ;
  assign w1570 = w1502 ^ w1569 ;
  assign w1571 = ~w1534 & w1570 ;
  assign w1572 = ( w1414 & w1532 ) | ( w1414 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1573 = ~w1533 & w1572 ;
  assign w1574 = w1571 | w1573 ;
  assign w1575 = ~\pi074 & w1574 ;
  assign w1576 = ~w1427 & w1498 ;
  assign w1577 = w1499 ^ w1576 ;
  assign w1578 = ~w1534 & w1577 ;
  assign w1579 = ( w1420 & w1532 ) | ( w1420 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1580 = ~w1533 & w1579 ;
  assign w1581 = w1578 | w1580 ;
  assign w1582 = ~\pi073 & w1581 ;
  assign w1583 = ~w1433 & w1495 ;
  assign w1584 = w1496 ^ w1583 ;
  assign w1585 = ~w1534 & w1584 ;
  assign w1586 = ( w1426 & w1532 ) | ( w1426 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1587 = ~w1533 & w1586 ;
  assign w1588 = w1585 | w1587 ;
  assign w1589 = ~\pi072 & w1588 ;
  assign w1590 = ~w1439 & w1492 ;
  assign w1591 = w1493 ^ w1590 ;
  assign w1592 = ~w1534 & w1591 ;
  assign w1593 = ( w1432 & w1532 ) | ( w1432 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1594 = ~w1533 & w1593 ;
  assign w1595 = w1592 | w1594 ;
  assign w1596 = ~\pi071 & w1595 ;
  assign w1597 = ~w1445 & w1489 ;
  assign w1598 = w1490 ^ w1597 ;
  assign w1599 = ~w1534 & w1598 ;
  assign w1600 = ( w1438 & w1532 ) | ( w1438 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1601 = ~w1533 & w1600 ;
  assign w1602 = w1599 | w1601 ;
  assign w1603 = ~\pi070 & w1602 ;
  assign w1604 = ~w1451 & w1486 ;
  assign w1605 = w1487 ^ w1604 ;
  assign w1606 = ~w1534 & w1605 ;
  assign w1607 = ( w1444 & w1532 ) | ( w1444 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1608 = ~w1533 & w1607 ;
  assign w1609 = w1606 | w1608 ;
  assign w1610 = ~\pi069 & w1609 ;
  assign w1611 = ~w1459 & w1483 ;
  assign w1612 = w1484 ^ w1611 ;
  assign w1613 = ~w1534 & w1612 ;
  assign w1614 = ( w1450 & w1532 ) | ( w1450 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1615 = ~w1533 & w1614 ;
  assign w1616 = w1613 | w1615 ;
  assign w1617 = ~\pi068 & w1616 ;
  assign w1618 = w1479 & ~w1480 ;
  assign w1619 = w1481 ^ w1618 ;
  assign w1620 = ~w1534 & w1619 ;
  assign w1621 = ( w1458 & w1532 ) | ( w1458 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1622 = ~w1533 & w1621 ;
  assign w1623 = w1620 | w1622 ;
  assign w1624 = ~\pi067 & w1623 ;
  assign w1625 = w1465 & ~w1469 ;
  assign w1626 = w1380 ^ w1469 ;
  assign w1627 = ( \pi050 & ~w1625 ) | ( \pi050 & w1626 ) | ( ~w1625 & w1626 ) ;
  assign w1628 = ( \pi050 & w1469 ) | ( \pi050 & w1627 ) | ( w1469 & w1627 ) ;
  assign w1629 = w1474 ^ w1628 ;
  assign w1630 = \pi065 ^ w1629 ;
  assign w1631 = ~w1534 & w1630 ;
  assign w1632 = ( w1473 & w1532 ) | ( w1473 & w1533 ) | ( w1532 & w1533 ) ;
  assign w1633 = ~w1533 & w1632 ;
  assign w1634 = w1631 | w1633 ;
  assign w1635 = ~\pi066 & w1634 ;
  assign w1636 = \pi066 ^ w1634 ;
  assign w1637 = \pi064 & ~w1534 ;
  assign w1638 = \pi049 ^ w1637 ;
  assign w1639 = ( ~\pi048 & \pi064 ) | ( ~\pi048 & w1636 ) | ( \pi064 & w1636 ) ;
  assign w1640 = ( \pi065 & ~w1638 ) | ( \pi065 & w1639 ) | ( ~w1638 & w1639 ) ;
  assign w1641 = w1636 | w1640 ;
  assign w1642 = \pi067 ^ w1623 ;
  assign w1643 = ( ~w1635 & w1641 ) | ( ~w1635 & w1642 ) | ( w1641 & w1642 ) ;
  assign w1644 = w1642 | w1643 ;
  assign w1645 = \pi068 ^ w1616 ;
  assign w1646 = ( ~w1624 & w1644 ) | ( ~w1624 & w1645 ) | ( w1644 & w1645 ) ;
  assign w1647 = w1645 | w1646 ;
  assign w1648 = \pi069 ^ w1609 ;
  assign w1649 = ( ~w1617 & w1647 ) | ( ~w1617 & w1648 ) | ( w1647 & w1648 ) ;
  assign w1650 = w1648 | w1649 ;
  assign w1651 = \pi070 ^ w1602 ;
  assign w1652 = ( ~w1610 & w1650 ) | ( ~w1610 & w1651 ) | ( w1650 & w1651 ) ;
  assign w1653 = w1651 | w1652 ;
  assign w1654 = \pi071 ^ w1595 ;
  assign w1655 = ( ~w1603 & w1653 ) | ( ~w1603 & w1654 ) | ( w1653 & w1654 ) ;
  assign w1656 = w1654 | w1655 ;
  assign w1657 = \pi072 ^ w1588 ;
  assign w1658 = ( ~w1596 & w1656 ) | ( ~w1596 & w1657 ) | ( w1656 & w1657 ) ;
  assign w1659 = w1657 | w1658 ;
  assign w1660 = \pi073 ^ w1581 ;
  assign w1661 = ( ~w1589 & w1659 ) | ( ~w1589 & w1660 ) | ( w1659 & w1660 ) ;
  assign w1662 = w1660 | w1661 ;
  assign w1663 = \pi074 ^ w1574 ;
  assign w1664 = ( ~w1582 & w1662 ) | ( ~w1582 & w1663 ) | ( w1662 & w1663 ) ;
  assign w1665 = w1663 | w1664 ;
  assign w1666 = \pi075 ^ w1567 ;
  assign w1667 = ( ~w1575 & w1665 ) | ( ~w1575 & w1666 ) | ( w1665 & w1666 ) ;
  assign w1668 = w1666 | w1667 ;
  assign w1669 = \pi076 ^ w1560 ;
  assign w1670 = ( ~w1568 & w1668 ) | ( ~w1568 & w1669 ) | ( w1668 & w1669 ) ;
  assign w1671 = w1669 | w1670 ;
  assign w1672 = \pi077 ^ w1553 ;
  assign w1673 = ( ~w1561 & w1671 ) | ( ~w1561 & w1672 ) | ( w1671 & w1672 ) ;
  assign w1674 = w1672 | w1673 ;
  assign w1675 = \pi078 ^ w1540 ;
  assign w1676 = ( ~w1554 & w1674 ) | ( ~w1554 & w1675 ) | ( w1674 & w1675 ) ;
  assign w1677 = w1675 | w1676 ;
  assign w1678 = \pi079 ^ w1546 ;
  assign w1679 = w1547 & ~w1678 ;
  assign w1680 = ( w1677 & w1678 ) | ( w1677 & ~w1679 ) | ( w1678 & ~w1679 ) ;
  assign w1681 = ~\pi079 & w1546 ;
  assign w1682 = w1680 & ~w1681 ;
  assign w1683 = w209 | w1682 ;
  assign w1684 = w1540 & w1683 ;
  assign w1685 = ~w1554 & w1674 ;
  assign w1686 = w1675 ^ w1685 ;
  assign w1687 = ~w1683 & w1686 ;
  assign w1688 = w1684 | w1687 ;
  assign w1689 = w1546 & w1683 ;
  assign w1690 = ~w1547 & w1677 ;
  assign w1691 = w1678 ^ w1690 ;
  assign w1692 = ~w1683 & w1691 ;
  assign w1693 = w1689 | w1692 ;
  assign w1694 = ~\pi079 & w1688 ;
  assign w1695 = w1553 & w1683 ;
  assign w1696 = ~w1561 & w1671 ;
  assign w1697 = w1672 ^ w1696 ;
  assign w1698 = ~w1683 & w1697 ;
  assign w1699 = w1695 | w1698 ;
  assign w1700 = ~\pi078 & w1699 ;
  assign w1701 = w1560 & w1683 ;
  assign w1702 = ~w1568 & w1668 ;
  assign w1703 = w1669 ^ w1702 ;
  assign w1704 = ~w1683 & w1703 ;
  assign w1705 = w1701 | w1704 ;
  assign w1706 = ~\pi077 & w1705 ;
  assign w1707 = w1567 & w1683 ;
  assign w1708 = ~w1575 & w1665 ;
  assign w1709 = w1666 ^ w1708 ;
  assign w1710 = ~w1683 & w1709 ;
  assign w1711 = w1707 | w1710 ;
  assign w1712 = ~\pi076 & w1711 ;
  assign w1713 = w1574 & w1683 ;
  assign w1714 = ~w1582 & w1662 ;
  assign w1715 = w1663 ^ w1714 ;
  assign w1716 = ~w1683 & w1715 ;
  assign w1717 = w1713 | w1716 ;
  assign w1718 = ~\pi075 & w1717 ;
  assign w1719 = w1581 & w1683 ;
  assign w1720 = ~w1589 & w1659 ;
  assign w1721 = w1660 ^ w1720 ;
  assign w1722 = ~w1683 & w1721 ;
  assign w1723 = w1719 | w1722 ;
  assign w1724 = ~\pi074 & w1723 ;
  assign w1725 = w1588 & w1683 ;
  assign w1726 = ~w1596 & w1656 ;
  assign w1727 = w1657 ^ w1726 ;
  assign w1728 = ~w1683 & w1727 ;
  assign w1729 = w1725 | w1728 ;
  assign w1730 = ~\pi073 & w1729 ;
  assign w1731 = w1595 & w1683 ;
  assign w1732 = ~w1603 & w1653 ;
  assign w1733 = w1654 ^ w1732 ;
  assign w1734 = ~w1683 & w1733 ;
  assign w1735 = w1731 | w1734 ;
  assign w1736 = ~\pi072 & w1735 ;
  assign w1737 = w1602 & w1683 ;
  assign w1738 = ~w1610 & w1650 ;
  assign w1739 = w1651 ^ w1738 ;
  assign w1740 = ~w1683 & w1739 ;
  assign w1741 = w1737 | w1740 ;
  assign w1742 = ~\pi071 & w1741 ;
  assign w1743 = w1609 & w1683 ;
  assign w1744 = ~w1617 & w1647 ;
  assign w1745 = w1648 ^ w1744 ;
  assign w1746 = ~w1683 & w1745 ;
  assign w1747 = w1743 | w1746 ;
  assign w1748 = ~\pi070 & w1747 ;
  assign w1749 = w1616 & w1683 ;
  assign w1750 = ~w1624 & w1644 ;
  assign w1751 = w1645 ^ w1750 ;
  assign w1752 = ~w1683 & w1751 ;
  assign w1753 = w1749 | w1752 ;
  assign w1754 = ~\pi069 & w1753 ;
  assign w1755 = w1623 & w1683 ;
  assign w1756 = ~w1635 & w1641 ;
  assign w1757 = w1642 ^ w1756 ;
  assign w1758 = ~w1683 & w1757 ;
  assign w1759 = w1755 | w1758 ;
  assign w1760 = ~\pi068 & w1759 ;
  assign w1761 = w1634 & w1683 ;
  assign w1762 = ~\pi048 & \pi064 ;
  assign w1763 = ( \pi065 & ~w1638 ) | ( \pi065 & w1762 ) | ( ~w1638 & w1762 ) ;
  assign w1764 = w1636 ^ w1763 ;
  assign w1765 = ( w209 & w1682 ) | ( w209 & w1764 ) | ( w1682 & w1764 ) ;
  assign w1766 = w1764 & ~w1765 ;
  assign w1767 = w1761 | w1766 ;
  assign w1768 = ~\pi067 & w1767 ;
  assign w1769 = \pi049 ^ \pi065 ;
  assign w1770 = \pi048 ^ w1534 ;
  assign w1771 = ( \pi064 & w209 ) | ( \pi064 & w1770 ) | ( w209 & w1770 ) ;
  assign w1772 = w1769 ^ w1771 ;
  assign w1773 = ~w209 & w1772 ;
  assign w1774 = ~w1682 & w1773 ;
  assign w1775 = ( ~\pi064 & w1534 ) | ( ~\pi064 & w1683 ) | ( w1534 & w1683 ) ;
  assign w1776 = \pi049 ^ w1775 ;
  assign w1777 = w1683 & ~w1776 ;
  assign w1778 = w1774 | w1777 ;
  assign w1779 = ~\pi066 & w1778 ;
  assign w1780 = \pi064 & ~\pi080 ;
  assign w1781 = ~w443 & w1780 ;
  assign w1782 = ~w1527 & w1781 ;
  assign w1783 = ( \pi048 & w1682 ) | ( \pi048 & ~w1782 ) | ( w1682 & ~w1782 ) ;
  assign w1784 = \pi048 & w1783 ;
  assign w1785 = ~w185 & w1762 ;
  assign w1786 = ~w1383 & w1785 ;
  assign w1787 = ~w1682 & w1786 ;
  assign w1788 = w1784 | w1787 ;
  assign w1789 = ~\pi047 & \pi064 ;
  assign w1790 = \pi065 ^ w1788 ;
  assign w1791 = w1789 | w1790 ;
  assign w1792 = w1683 | w1774 ;
  assign w1793 = ( w1638 & w1774 ) | ( w1638 & w1792 ) | ( w1774 & w1792 ) ;
  assign w1794 = \pi066 ^ w1793 ;
  assign w1795 = ~\pi065 & w1788 ;
  assign w1796 = w1791 | w1795 ;
  assign w1797 = ( w1794 & ~w1795 ) | ( w1794 & w1796 ) | ( ~w1795 & w1796 ) ;
  assign w1798 = \pi067 ^ w1767 ;
  assign w1799 = ( ~w1779 & w1797 ) | ( ~w1779 & w1798 ) | ( w1797 & w1798 ) ;
  assign w1800 = w1798 | w1799 ;
  assign w1801 = \pi068 ^ w1759 ;
  assign w1802 = ( ~w1768 & w1800 ) | ( ~w1768 & w1801 ) | ( w1800 & w1801 ) ;
  assign w1803 = w1801 | w1802 ;
  assign w1804 = \pi069 ^ w1753 ;
  assign w1805 = ( ~w1760 & w1803 ) | ( ~w1760 & w1804 ) | ( w1803 & w1804 ) ;
  assign w1806 = w1804 | w1805 ;
  assign w1807 = \pi070 ^ w1747 ;
  assign w1808 = ( ~w1754 & w1806 ) | ( ~w1754 & w1807 ) | ( w1806 & w1807 ) ;
  assign w1809 = w1807 | w1808 ;
  assign w1810 = \pi071 ^ w1741 ;
  assign w1811 = ( ~w1748 & w1809 ) | ( ~w1748 & w1810 ) | ( w1809 & w1810 ) ;
  assign w1812 = w1810 | w1811 ;
  assign w1813 = \pi072 ^ w1735 ;
  assign w1814 = ( ~w1742 & w1812 ) | ( ~w1742 & w1813 ) | ( w1812 & w1813 ) ;
  assign w1815 = w1813 | w1814 ;
  assign w1816 = \pi073 ^ w1729 ;
  assign w1817 = ( ~w1736 & w1815 ) | ( ~w1736 & w1816 ) | ( w1815 & w1816 ) ;
  assign w1818 = w1816 | w1817 ;
  assign w1819 = \pi074 ^ w1723 ;
  assign w1820 = ( ~w1730 & w1818 ) | ( ~w1730 & w1819 ) | ( w1818 & w1819 ) ;
  assign w1821 = w1819 | w1820 ;
  assign w1822 = \pi075 ^ w1717 ;
  assign w1823 = ( ~w1724 & w1821 ) | ( ~w1724 & w1822 ) | ( w1821 & w1822 ) ;
  assign w1824 = w1822 | w1823 ;
  assign w1825 = \pi076 ^ w1711 ;
  assign w1826 = ( ~w1718 & w1824 ) | ( ~w1718 & w1825 ) | ( w1824 & w1825 ) ;
  assign w1827 = w1825 | w1826 ;
  assign w1828 = \pi077 ^ w1705 ;
  assign w1829 = ( ~w1712 & w1827 ) | ( ~w1712 & w1828 ) | ( w1827 & w1828 ) ;
  assign w1830 = w1828 | w1829 ;
  assign w1831 = \pi078 ^ w1699 ;
  assign w1832 = ( ~w1706 & w1830 ) | ( ~w1706 & w1831 ) | ( w1830 & w1831 ) ;
  assign w1833 = w1831 | w1832 ;
  assign w1834 = \pi079 ^ w1688 ;
  assign w1835 = ( ~w1700 & w1833 ) | ( ~w1700 & w1834 ) | ( w1833 & w1834 ) ;
  assign w1836 = w1834 | w1835 ;
  assign w1837 = \pi080 ^ w1693 ;
  assign w1838 = w1694 & ~w1837 ;
  assign w1839 = ( w1836 & w1837 ) | ( w1836 & ~w1838 ) | ( w1837 & ~w1838 ) ;
  assign w1840 = ~\pi080 & w1693 ;
  assign w1841 = w1839 & ~w1840 ;
  assign w1842 = w331 | w1841 ;
  assign w1843 = w1688 & w1842 ;
  assign w1844 = ~w1700 & w1833 ;
  assign w1845 = w1834 ^ w1844 ;
  assign w1846 = ~w1842 & w1845 ;
  assign w1847 = w1843 | w1846 ;
  assign w1848 = ~\pi080 & w1847 ;
  assign w1849 = w1699 & w1842 ;
  assign w1850 = ~w1706 & w1830 ;
  assign w1851 = w1831 ^ w1850 ;
  assign w1852 = ~w1842 & w1851 ;
  assign w1853 = w1849 | w1852 ;
  assign w1854 = ~\pi079 & w1853 ;
  assign w1855 = w1705 & w1842 ;
  assign w1856 = ~w1712 & w1827 ;
  assign w1857 = w1828 ^ w1856 ;
  assign w1858 = ~w1842 & w1857 ;
  assign w1859 = w1855 | w1858 ;
  assign w1860 = ~\pi078 & w1859 ;
  assign w1861 = w1711 & w1842 ;
  assign w1862 = ~w1718 & w1824 ;
  assign w1863 = w1825 ^ w1862 ;
  assign w1864 = ~w1842 & w1863 ;
  assign w1865 = w1861 | w1864 ;
  assign w1866 = ~\pi077 & w1865 ;
  assign w1867 = w1717 & w1842 ;
  assign w1868 = ~w1724 & w1821 ;
  assign w1869 = w1822 ^ w1868 ;
  assign w1870 = ~w1842 & w1869 ;
  assign w1871 = w1867 | w1870 ;
  assign w1872 = ~\pi076 & w1871 ;
  assign w1873 = w1723 & w1842 ;
  assign w1874 = ~w1730 & w1818 ;
  assign w1875 = w1819 ^ w1874 ;
  assign w1876 = ~w1842 & w1875 ;
  assign w1877 = w1873 | w1876 ;
  assign w1878 = ~\pi075 & w1877 ;
  assign w1879 = w1729 & w1842 ;
  assign w1880 = ~w1736 & w1815 ;
  assign w1881 = w1816 ^ w1880 ;
  assign w1882 = ~w1842 & w1881 ;
  assign w1883 = w1879 | w1882 ;
  assign w1884 = ~\pi074 & w1883 ;
  assign w1885 = w1735 & w1842 ;
  assign w1886 = ~w1742 & w1812 ;
  assign w1887 = w1813 ^ w1886 ;
  assign w1888 = ~w1842 & w1887 ;
  assign w1889 = w1885 | w1888 ;
  assign w1890 = ~\pi073 & w1889 ;
  assign w1891 = w1741 & w1842 ;
  assign w1892 = ~w1748 & w1809 ;
  assign w1893 = w1810 ^ w1892 ;
  assign w1894 = ~w1842 & w1893 ;
  assign w1895 = w1891 | w1894 ;
  assign w1896 = ~\pi072 & w1895 ;
  assign w1897 = w1747 & w1842 ;
  assign w1898 = ~w1754 & w1806 ;
  assign w1899 = w1807 ^ w1898 ;
  assign w1900 = ~w1842 & w1899 ;
  assign w1901 = w1897 | w1900 ;
  assign w1902 = ~\pi071 & w1901 ;
  assign w1903 = w1753 & w1842 ;
  assign w1904 = ~w1760 & w1803 ;
  assign w1905 = w1804 ^ w1904 ;
  assign w1906 = ~w1842 & w1905 ;
  assign w1907 = w1903 | w1906 ;
  assign w1908 = ~\pi070 & w1907 ;
  assign w1909 = w1759 & w1842 ;
  assign w1910 = ~w1768 & w1800 ;
  assign w1911 = w1801 ^ w1910 ;
  assign w1912 = ~w1842 & w1911 ;
  assign w1913 = w1909 | w1912 ;
  assign w1914 = ~\pi069 & w1913 ;
  assign w1915 = w1767 & w1842 ;
  assign w1916 = ~w1779 & w1797 ;
  assign w1917 = w1798 ^ w1916 ;
  assign w1918 = ~w1842 & w1917 ;
  assign w1919 = w1915 | w1918 ;
  assign w1920 = ~\pi068 & w1919 ;
  assign w1921 = w1778 & w1842 ;
  assign w1922 = ~w1788 & w1791 ;
  assign w1923 = ( \pi065 & w1791 ) | ( \pi065 & w1922 ) | ( w1791 & w1922 ) ;
  assign w1924 = w1794 ^ w1923 ;
  assign w1925 = ~w1842 & w1924 ;
  assign w1926 = w1921 | w1925 ;
  assign w1927 = ~\pi067 & w1926 ;
  assign w1928 = w1788 & w1842 ;
  assign w1929 = ( ~w331 & w1784 ) | ( ~w331 & w1787 ) | ( w1784 & w1787 ) ;
  assign w1930 = \pi065 ^ w1929 ;
  assign w1931 = ( ~w331 & w1789 ) | ( ~w331 & w1930 ) | ( w1789 & w1930 ) ;
  assign w1932 = ( w1789 & w1841 ) | ( w1789 & w1930 ) | ( w1841 & w1930 ) ;
  assign w1933 = w1931 & ~w1932 ;
  assign w1934 = w1928 | w1933 ;
  assign w1935 = ~\pi066 & w1934 ;
  assign w1936 = ( \pi064 & ~\pi081 ) | ( \pi064 & \pi082 ) | ( ~\pi081 & \pi082 ) ;
  assign w1937 = w176 | w205 ;
  assign w1938 = ( \pi082 & \pi083 ) | ( \pi082 & ~w176 ) | ( \pi083 & ~w176 ) ;
  assign w1939 = w1937 | w1938 ;
  assign w1940 = w1936 & ~w1939 ;
  assign w1941 = ( ~w201 & w204 ) | ( ~w201 & w1940 ) | ( w204 & w1940 ) ;
  assign w1942 = ~w204 & w1941 ;
  assign w1943 = ( \pi047 & w1841 ) | ( \pi047 & ~w1942 ) | ( w1841 & ~w1942 ) ;
  assign w1944 = \pi047 & w1943 ;
  assign w1945 = ~w237 & w1789 ;
  assign w1946 = ~w452 & w1945 ;
  assign w1947 = ( w443 & ~w452 ) | ( w443 & w1841 ) | ( ~w452 & w1841 ) ;
  assign w1948 = w1946 & ~w1947 ;
  assign w1949 = w1944 | w1948 ;
  assign w1950 = ~\pi046 & \pi064 ;
  assign w1951 = ( w1944 & w1948 ) | ( w1944 & ~w1950 ) | ( w1948 & ~w1950 ) ;
  assign w1952 = \pi065 ^ w1951 ;
  assign w1953 = w1950 | w1952 ;
  assign w1954 = ~\pi065 & w1949 ;
  assign w1955 = \pi066 ^ w1934 ;
  assign w1956 = ( w1953 & ~w1954 ) | ( w1953 & w1955 ) | ( ~w1954 & w1955 ) ;
  assign w1957 = w1955 | w1956 ;
  assign w1958 = \pi067 ^ w1926 ;
  assign w1959 = ( ~w1935 & w1957 ) | ( ~w1935 & w1958 ) | ( w1957 & w1958 ) ;
  assign w1960 = w1958 | w1959 ;
  assign w1961 = \pi068 ^ w1919 ;
  assign w1962 = ( ~w1927 & w1960 ) | ( ~w1927 & w1961 ) | ( w1960 & w1961 ) ;
  assign w1963 = w1961 | w1962 ;
  assign w1964 = \pi069 ^ w1913 ;
  assign w1965 = ( ~w1920 & w1963 ) | ( ~w1920 & w1964 ) | ( w1963 & w1964 ) ;
  assign w1966 = w1964 | w1965 ;
  assign w1967 = \pi070 ^ w1907 ;
  assign w1968 = ( ~w1914 & w1966 ) | ( ~w1914 & w1967 ) | ( w1966 & w1967 ) ;
  assign w1969 = w1967 | w1968 ;
  assign w1970 = \pi071 ^ w1901 ;
  assign w1971 = ( ~w1908 & w1969 ) | ( ~w1908 & w1970 ) | ( w1969 & w1970 ) ;
  assign w1972 = w1970 | w1971 ;
  assign w1973 = \pi072 ^ w1895 ;
  assign w1974 = ( ~w1902 & w1972 ) | ( ~w1902 & w1973 ) | ( w1972 & w1973 ) ;
  assign w1975 = w1973 | w1974 ;
  assign w1976 = \pi073 ^ w1889 ;
  assign w1977 = ( ~w1896 & w1975 ) | ( ~w1896 & w1976 ) | ( w1975 & w1976 ) ;
  assign w1978 = w1976 | w1977 ;
  assign w1979 = \pi074 ^ w1883 ;
  assign w1980 = ( ~w1890 & w1978 ) | ( ~w1890 & w1979 ) | ( w1978 & w1979 ) ;
  assign w1981 = w1979 | w1980 ;
  assign w1982 = \pi075 ^ w1877 ;
  assign w1983 = ( ~w1884 & w1981 ) | ( ~w1884 & w1982 ) | ( w1981 & w1982 ) ;
  assign w1984 = w1982 | w1983 ;
  assign w1985 = \pi076 ^ w1871 ;
  assign w1986 = ( ~w1878 & w1984 ) | ( ~w1878 & w1985 ) | ( w1984 & w1985 ) ;
  assign w1987 = w1985 | w1986 ;
  assign w1988 = \pi077 ^ w1865 ;
  assign w1989 = ( ~w1872 & w1987 ) | ( ~w1872 & w1988 ) | ( w1987 & w1988 ) ;
  assign w1990 = w1988 | w1989 ;
  assign w1991 = \pi078 ^ w1859 ;
  assign w1992 = ( ~w1866 & w1990 ) | ( ~w1866 & w1991 ) | ( w1990 & w1991 ) ;
  assign w1993 = w1991 | w1992 ;
  assign w1994 = \pi079 ^ w1853 ;
  assign w1995 = ( ~w1860 & w1993 ) | ( ~w1860 & w1994 ) | ( w1993 & w1994 ) ;
  assign w1996 = w1994 | w1995 ;
  assign w1997 = \pi080 ^ w1847 ;
  assign w1998 = ( ~w1854 & w1996 ) | ( ~w1854 & w1997 ) | ( w1996 & w1997 ) ;
  assign w1999 = w1997 | w1998 ;
  assign w2000 = w1693 & w1842 ;
  assign w2001 = ~w1694 & w1836 ;
  assign w2002 = w1837 ^ w2001 ;
  assign w2003 = ~w1842 & w2002 ;
  assign w2004 = w2000 | w2003 ;
  assign w2005 = ~\pi081 & w2004 ;
  assign w2006 = ( \pi081 & ~w2000 ) | ( \pi081 & w2003 ) | ( ~w2000 & w2003 ) ;
  assign w2007 = ~w2003 & w2006 ;
  assign w2008 = ( ~\pi082 & w176 ) | ( ~\pi082 & w205 ) | ( w176 & w205 ) ;
  assign w2009 = ( \pi082 & \pi083 ) | ( \pi082 & ~w204 ) | ( \pi083 & ~w204 ) ;
  assign w2010 = w298 | w2009 ;
  assign w2011 = w2008 | w2010 ;
  assign w2012 = w2005 | w2007 ;
  assign w2013 = ( ~w1848 & w1999 ) | ( ~w1848 & w2012 ) | ( w1999 & w2012 ) ;
  assign w2014 = ( w2011 & ~w2012 ) | ( w2011 & w2013 ) | ( ~w2012 & w2013 ) ;
  assign w2015 = w2012 | w2014 ;
  assign w2016 = ~w331 & w2004 ;
  assign w2017 = w2015 & ~w2016 ;
  assign w2018 = ~w1854 & w1996 ;
  assign w2019 = w1997 ^ w2018 ;
  assign w2020 = ~w2017 & w2019 ;
  assign w2021 = ( w1847 & w2015 ) | ( w1847 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2022 = ~w2016 & w2021 ;
  assign w2023 = w2020 | w2022 ;
  assign w2024 = ( ~w1848 & w1999 ) | ( ~w1848 & w2017 ) | ( w1999 & w2017 ) ;
  assign w2025 = w2012 ^ w2024 ;
  assign w2026 = ~w2017 & w2025 ;
  assign w2027 = ( w331 & ~w2004 ) | ( w331 & w2015 ) | ( ~w2004 & w2015 ) ;
  assign w2028 = w2004 & w2027 ;
  assign w2029 = w2026 | w2028 ;
  assign w2030 = ~\pi081 & w2023 ;
  assign w2031 = ~w1860 & w1993 ;
  assign w2032 = w1994 ^ w2031 ;
  assign w2033 = ~w2017 & w2032 ;
  assign w2034 = ( w1853 & w2015 ) | ( w1853 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2035 = ~w2016 & w2034 ;
  assign w2036 = w2033 | w2035 ;
  assign w2037 = ~\pi080 & w2036 ;
  assign w2038 = ~w1866 & w1990 ;
  assign w2039 = w1991 ^ w2038 ;
  assign w2040 = ~w2017 & w2039 ;
  assign w2041 = ( w1859 & w2015 ) | ( w1859 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2042 = ~w2016 & w2041 ;
  assign w2043 = w2040 | w2042 ;
  assign w2044 = ~\pi079 & w2043 ;
  assign w2045 = ~w1872 & w1987 ;
  assign w2046 = w1988 ^ w2045 ;
  assign w2047 = ~w2017 & w2046 ;
  assign w2048 = ( w1865 & w2015 ) | ( w1865 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2049 = ~w2016 & w2048 ;
  assign w2050 = w2047 | w2049 ;
  assign w2051 = ~\pi078 & w2050 ;
  assign w2052 = ~w1878 & w1984 ;
  assign w2053 = w1985 ^ w2052 ;
  assign w2054 = ~w2017 & w2053 ;
  assign w2055 = ( w1871 & w2015 ) | ( w1871 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2056 = ~w2016 & w2055 ;
  assign w2057 = w2054 | w2056 ;
  assign w2058 = ~\pi077 & w2057 ;
  assign w2059 = ~w1884 & w1981 ;
  assign w2060 = w1982 ^ w2059 ;
  assign w2061 = ~w2017 & w2060 ;
  assign w2062 = ( w1877 & w2015 ) | ( w1877 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2063 = ~w2016 & w2062 ;
  assign w2064 = w2061 | w2063 ;
  assign w2065 = ~\pi076 & w2064 ;
  assign w2066 = ~w1890 & w1978 ;
  assign w2067 = w1979 ^ w2066 ;
  assign w2068 = ~w2017 & w2067 ;
  assign w2069 = ( w1883 & w2015 ) | ( w1883 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2070 = ~w2016 & w2069 ;
  assign w2071 = w2068 | w2070 ;
  assign w2072 = ~\pi075 & w2071 ;
  assign w2073 = ~w1896 & w1975 ;
  assign w2074 = w1976 ^ w2073 ;
  assign w2075 = ~w2017 & w2074 ;
  assign w2076 = ( w1889 & w2015 ) | ( w1889 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2077 = ~w2016 & w2076 ;
  assign w2078 = w2075 | w2077 ;
  assign w2079 = ~\pi074 & w2078 ;
  assign w2080 = ~w1902 & w1972 ;
  assign w2081 = w1973 ^ w2080 ;
  assign w2082 = ~w2017 & w2081 ;
  assign w2083 = ( w1895 & w2015 ) | ( w1895 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2084 = ~w2016 & w2083 ;
  assign w2085 = w2082 | w2084 ;
  assign w2086 = ~\pi073 & w2085 ;
  assign w2087 = ~w1908 & w1969 ;
  assign w2088 = w1970 ^ w2087 ;
  assign w2089 = ~w2017 & w2088 ;
  assign w2090 = ( w1901 & w2015 ) | ( w1901 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2091 = ~w2016 & w2090 ;
  assign w2092 = w2089 | w2091 ;
  assign w2093 = ~\pi072 & w2092 ;
  assign w2094 = ~w1914 & w1966 ;
  assign w2095 = w1967 ^ w2094 ;
  assign w2096 = ~w2017 & w2095 ;
  assign w2097 = ( w1907 & w2015 ) | ( w1907 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2098 = ~w2016 & w2097 ;
  assign w2099 = w2096 | w2098 ;
  assign w2100 = ~\pi071 & w2099 ;
  assign w2101 = ~w1920 & w1963 ;
  assign w2102 = w1964 ^ w2101 ;
  assign w2103 = ~w2017 & w2102 ;
  assign w2104 = ( w1913 & w2015 ) | ( w1913 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2105 = ~w2016 & w2104 ;
  assign w2106 = w2103 | w2105 ;
  assign w2107 = ~\pi070 & w2106 ;
  assign w2108 = ~w1927 & w1960 ;
  assign w2109 = w1961 ^ w2108 ;
  assign w2110 = ~w2017 & w2109 ;
  assign w2111 = ( w1919 & w2015 ) | ( w1919 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2112 = ~w2016 & w2111 ;
  assign w2113 = w2110 | w2112 ;
  assign w2114 = ~\pi069 & w2113 ;
  assign w2115 = ~w1935 & w1957 ;
  assign w2116 = w1958 ^ w2115 ;
  assign w2117 = ~w2017 & w2116 ;
  assign w2118 = ( w1926 & w2015 ) | ( w1926 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2119 = ~w2016 & w2118 ;
  assign w2120 = w2117 | w2119 ;
  assign w2121 = ~\pi068 & w2120 ;
  assign w2122 = w1953 & ~w1954 ;
  assign w2123 = w1955 ^ w2122 ;
  assign w2124 = ~w2017 & w2123 ;
  assign w2125 = ( w1934 & w2015 ) | ( w1934 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2126 = ~w2016 & w2125 ;
  assign w2127 = w2124 | w2126 ;
  assign w2128 = ~\pi067 & w2127 ;
  assign w2129 = ( w1944 & w1948 ) | ( w1944 & ~w2017 ) | ( w1948 & ~w2017 ) ;
  assign w2130 = ( ~\pi046 & \pi064 ) | ( ~\pi046 & w2017 ) | ( \pi064 & w2017 ) ;
  assign w2131 = w2129 ^ w2130 ;
  assign w2132 = \pi065 ^ w2131 ;
  assign w2133 = ~w2017 & w2132 ;
  assign w2134 = ( w1949 & w2015 ) | ( w1949 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2135 = ~w2016 & w2134 ;
  assign w2136 = w2133 | w2135 ;
  assign w2137 = ~\pi066 & w2136 ;
  assign w2138 = \pi066 ^ w2136 ;
  assign w2139 = \pi064 & ~w2017 ;
  assign w2140 = \pi046 ^ w2139 ;
  assign w2141 = ( ~\pi045 & \pi064 ) | ( ~\pi045 & w2138 ) | ( \pi064 & w2138 ) ;
  assign w2142 = ( \pi065 & ~w2140 ) | ( \pi065 & w2141 ) | ( ~w2140 & w2141 ) ;
  assign w2143 = w2138 | w2142 ;
  assign w2144 = \pi067 ^ w2127 ;
  assign w2145 = ( ~w2137 & w2143 ) | ( ~w2137 & w2144 ) | ( w2143 & w2144 ) ;
  assign w2146 = w2144 | w2145 ;
  assign w2147 = \pi068 ^ w2120 ;
  assign w2148 = ( ~w2128 & w2146 ) | ( ~w2128 & w2147 ) | ( w2146 & w2147 ) ;
  assign w2149 = w2147 | w2148 ;
  assign w2150 = \pi069 ^ w2113 ;
  assign w2151 = ( ~w2121 & w2149 ) | ( ~w2121 & w2150 ) | ( w2149 & w2150 ) ;
  assign w2152 = w2150 | w2151 ;
  assign w2153 = \pi070 ^ w2106 ;
  assign w2154 = ( ~w2114 & w2152 ) | ( ~w2114 & w2153 ) | ( w2152 & w2153 ) ;
  assign w2155 = w2153 | w2154 ;
  assign w2156 = \pi071 ^ w2099 ;
  assign w2157 = ( ~w2107 & w2155 ) | ( ~w2107 & w2156 ) | ( w2155 & w2156 ) ;
  assign w2158 = w2156 | w2157 ;
  assign w2159 = \pi072 ^ w2092 ;
  assign w2160 = ( ~w2100 & w2158 ) | ( ~w2100 & w2159 ) | ( w2158 & w2159 ) ;
  assign w2161 = w2159 | w2160 ;
  assign w2162 = \pi073 ^ w2085 ;
  assign w2163 = ( ~w2093 & w2161 ) | ( ~w2093 & w2162 ) | ( w2161 & w2162 ) ;
  assign w2164 = w2162 | w2163 ;
  assign w2165 = \pi074 ^ w2078 ;
  assign w2166 = ( ~w2086 & w2164 ) | ( ~w2086 & w2165 ) | ( w2164 & w2165 ) ;
  assign w2167 = w2165 | w2166 ;
  assign w2168 = \pi075 ^ w2071 ;
  assign w2169 = ( ~w2079 & w2167 ) | ( ~w2079 & w2168 ) | ( w2167 & w2168 ) ;
  assign w2170 = w2168 | w2169 ;
  assign w2171 = \pi076 ^ w2064 ;
  assign w2172 = ( ~w2072 & w2170 ) | ( ~w2072 & w2171 ) | ( w2170 & w2171 ) ;
  assign w2173 = w2171 | w2172 ;
  assign w2174 = \pi077 ^ w2057 ;
  assign w2175 = ( ~w2065 & w2173 ) | ( ~w2065 & w2174 ) | ( w2173 & w2174 ) ;
  assign w2176 = w2174 | w2175 ;
  assign w2177 = \pi078 ^ w2050 ;
  assign w2178 = ( ~w2058 & w2176 ) | ( ~w2058 & w2177 ) | ( w2176 & w2177 ) ;
  assign w2179 = w2177 | w2178 ;
  assign w2180 = \pi079 ^ w2043 ;
  assign w2181 = ( ~w2051 & w2179 ) | ( ~w2051 & w2180 ) | ( w2179 & w2180 ) ;
  assign w2182 = w2180 | w2181 ;
  assign w2183 = \pi080 ^ w2036 ;
  assign w2184 = ( ~w2044 & w2182 ) | ( ~w2044 & w2183 ) | ( w2182 & w2183 ) ;
  assign w2185 = w2183 | w2184 ;
  assign w2186 = \pi081 ^ w2023 ;
  assign w2187 = ( ~w2037 & w2185 ) | ( ~w2037 & w2186 ) | ( w2185 & w2186 ) ;
  assign w2188 = w2186 | w2187 ;
  assign w2189 = \pi082 ^ w2029 ;
  assign w2190 = w2030 & ~w2189 ;
  assign w2191 = ( w2188 & w2189 ) | ( w2188 & ~w2190 ) | ( w2189 & ~w2190 ) ;
  assign w2192 = ~\pi082 & w2029 ;
  assign w2193 = w2191 & ~w2192 ;
  assign w2194 = ( ~\pi083 & w234 ) | ( ~\pi083 & w244 ) | ( w234 & w244 ) ;
  assign w2195 = ( \pi083 & \pi084 ) | ( \pi083 & ~w290 ) | ( \pi084 & ~w290 ) ;
  assign w2196 = w291 | w2195 ;
  assign w2197 = w2194 | w2196 ;
  assign w2198 = w2193 | w2197 ;
  assign w2199 = w2023 & w2198 ;
  assign w2200 = ~w2037 & w2185 ;
  assign w2201 = w2186 ^ w2200 ;
  assign w2202 = ~w2198 & w2201 ;
  assign w2203 = w2199 | w2202 ;
  assign w2204 = w2029 & w2198 ;
  assign w2205 = ~w2030 & w2188 ;
  assign w2206 = w2189 ^ w2205 ;
  assign w2207 = ~w2198 & w2206 ;
  assign w2208 = w2204 | w2207 ;
  assign w2209 = ~\pi082 & w2203 ;
  assign w2210 = w2036 & w2198 ;
  assign w2211 = ~w2044 & w2182 ;
  assign w2212 = w2183 ^ w2211 ;
  assign w2213 = ~w2198 & w2212 ;
  assign w2214 = w2210 | w2213 ;
  assign w2215 = ~\pi081 & w2214 ;
  assign w2216 = w2043 & w2198 ;
  assign w2217 = ~w2051 & w2179 ;
  assign w2218 = w2180 ^ w2217 ;
  assign w2219 = ~w2198 & w2218 ;
  assign w2220 = w2216 | w2219 ;
  assign w2221 = ~\pi080 & w2220 ;
  assign w2222 = w2050 & w2198 ;
  assign w2223 = ~w2058 & w2176 ;
  assign w2224 = w2177 ^ w2223 ;
  assign w2225 = ~w2198 & w2224 ;
  assign w2226 = w2222 | w2225 ;
  assign w2227 = ~\pi079 & w2226 ;
  assign w2228 = w2057 & w2198 ;
  assign w2229 = ~w2065 & w2173 ;
  assign w2230 = w2174 ^ w2229 ;
  assign w2231 = ~w2198 & w2230 ;
  assign w2232 = w2228 | w2231 ;
  assign w2233 = ~\pi078 & w2232 ;
  assign w2234 = w2064 & w2198 ;
  assign w2235 = ~w2072 & w2170 ;
  assign w2236 = w2171 ^ w2235 ;
  assign w2237 = ~w2198 & w2236 ;
  assign w2238 = w2234 | w2237 ;
  assign w2239 = ~\pi077 & w2238 ;
  assign w2240 = w2071 & w2198 ;
  assign w2241 = ~w2079 & w2167 ;
  assign w2242 = w2168 ^ w2241 ;
  assign w2243 = ~w2198 & w2242 ;
  assign w2244 = w2240 | w2243 ;
  assign w2245 = ~\pi076 & w2244 ;
  assign w2246 = w2078 & w2198 ;
  assign w2247 = ~w2086 & w2164 ;
  assign w2248 = w2165 ^ w2247 ;
  assign w2249 = ~w2198 & w2248 ;
  assign w2250 = w2246 | w2249 ;
  assign w2251 = ~\pi075 & w2250 ;
  assign w2252 = w2085 & w2198 ;
  assign w2253 = ~w2093 & w2161 ;
  assign w2254 = w2162 ^ w2253 ;
  assign w2255 = ~w2198 & w2254 ;
  assign w2256 = w2252 | w2255 ;
  assign w2257 = ~\pi074 & w2256 ;
  assign w2258 = w2092 & w2198 ;
  assign w2259 = ~w2100 & w2158 ;
  assign w2260 = w2159 ^ w2259 ;
  assign w2261 = ~w2198 & w2260 ;
  assign w2262 = w2258 | w2261 ;
  assign w2263 = ~\pi073 & w2262 ;
  assign w2264 = w2099 & w2198 ;
  assign w2265 = ~w2107 & w2155 ;
  assign w2266 = w2156 ^ w2265 ;
  assign w2267 = ~w2198 & w2266 ;
  assign w2268 = w2264 | w2267 ;
  assign w2269 = ~\pi072 & w2268 ;
  assign w2270 = w2106 & w2198 ;
  assign w2271 = ~w2114 & w2152 ;
  assign w2272 = w2153 ^ w2271 ;
  assign w2273 = ~w2198 & w2272 ;
  assign w2274 = w2270 | w2273 ;
  assign w2275 = ~\pi071 & w2274 ;
  assign w2276 = w2113 & w2198 ;
  assign w2277 = ~w2121 & w2149 ;
  assign w2278 = w2150 ^ w2277 ;
  assign w2279 = ~w2198 & w2278 ;
  assign w2280 = w2276 | w2279 ;
  assign w2281 = ~\pi070 & w2280 ;
  assign w2282 = w2120 & w2198 ;
  assign w2283 = ~w2128 & w2146 ;
  assign w2284 = w2147 ^ w2283 ;
  assign w2285 = ~w2198 & w2284 ;
  assign w2286 = w2282 | w2285 ;
  assign w2287 = ~\pi069 & w2286 ;
  assign w2288 = w2127 & w2198 ;
  assign w2289 = ~w2137 & w2143 ;
  assign w2290 = w2144 ^ w2289 ;
  assign w2291 = ~w2198 & w2290 ;
  assign w2292 = w2288 | w2291 ;
  assign w2293 = ~\pi068 & w2292 ;
  assign w2294 = w2136 & w2198 ;
  assign w2295 = ~\pi045 & \pi064 ;
  assign w2296 = ( \pi065 & ~w2140 ) | ( \pi065 & w2295 ) | ( ~w2140 & w2295 ) ;
  assign w2297 = w2138 ^ w2296 ;
  assign w2298 = ( w2193 & w2197 ) | ( w2193 & w2297 ) | ( w2197 & w2297 ) ;
  assign w2299 = w2297 & ~w2298 ;
  assign w2300 = w2294 | w2299 ;
  assign w2301 = ~\pi067 & w2300 ;
  assign w2302 = \pi046 ^ \pi065 ;
  assign w2303 = \pi045 ^ w2017 ;
  assign w2304 = ( \pi064 & w2197 ) | ( \pi064 & w2303 ) | ( w2197 & w2303 ) ;
  assign w2305 = w2302 ^ w2304 ;
  assign w2306 = ~w2197 & w2305 ;
  assign w2307 = ~w2193 & w2306 ;
  assign w2308 = ( ~\pi064 & w2017 ) | ( ~\pi064 & w2198 ) | ( w2017 & w2198 ) ;
  assign w2309 = \pi046 ^ w2308 ;
  assign w2310 = w2198 & ~w2309 ;
  assign w2311 = w2307 | w2310 ;
  assign w2312 = ~\pi066 & w2311 ;
  assign w2313 = ( \pi064 & w176 ) | ( \pi064 & w205 ) | ( w176 & w205 ) ;
  assign w2314 = ( \pi064 & ~\pi083 ) | ( \pi064 & w204 ) | ( ~\pi083 & w204 ) ;
  assign w2315 = ~w298 & w2314 ;
  assign w2316 = ~w2313 & w2315 ;
  assign w2317 = ( \pi045 & w2193 ) | ( \pi045 & ~w2316 ) | ( w2193 & ~w2316 ) ;
  assign w2318 = \pi045 & w2317 ;
  assign w2319 = ( ~\pi045 & \pi064 ) | ( ~\pi045 & \pi083 ) | ( \pi064 & \pi083 ) ;
  assign w2320 = w234 | w244 ;
  assign w2321 = ( \pi083 & \pi084 ) | ( \pi083 & ~w234 ) | ( \pi084 & ~w234 ) ;
  assign w2322 = w2320 | w2321 ;
  assign w2323 = w2319 & ~w2322 ;
  assign w2324 = ( ~w275 & w290 ) | ( ~w275 & w2323 ) | ( w290 & w2323 ) ;
  assign w2325 = ~w290 & w2324 ;
  assign w2326 = ~w2193 & w2325 ;
  assign w2327 = w2318 | w2326 ;
  assign w2328 = ~\pi044 & \pi064 ;
  assign w2329 = \pi065 ^ w2327 ;
  assign w2330 = w2328 | w2329 ;
  assign w2331 = ~\pi065 & w2327 ;
  assign w2332 = w2198 | w2307 ;
  assign w2333 = ( w2140 & w2307 ) | ( w2140 & w2332 ) | ( w2307 & w2332 ) ;
  assign w2334 = \pi066 ^ w2333 ;
  assign w2335 = ( w2330 & ~w2331 ) | ( w2330 & w2334 ) | ( ~w2331 & w2334 ) ;
  assign w2336 = w2334 | w2335 ;
  assign w2337 = \pi067 ^ w2300 ;
  assign w2338 = ( ~w2312 & w2336 ) | ( ~w2312 & w2337 ) | ( w2336 & w2337 ) ;
  assign w2339 = w2337 | w2338 ;
  assign w2340 = \pi068 ^ w2292 ;
  assign w2341 = ( ~w2301 & w2339 ) | ( ~w2301 & w2340 ) | ( w2339 & w2340 ) ;
  assign w2342 = w2340 | w2341 ;
  assign w2343 = \pi069 ^ w2286 ;
  assign w2344 = ( ~w2293 & w2342 ) | ( ~w2293 & w2343 ) | ( w2342 & w2343 ) ;
  assign w2345 = w2343 | w2344 ;
  assign w2346 = \pi070 ^ w2280 ;
  assign w2347 = ( ~w2287 & w2345 ) | ( ~w2287 & w2346 ) | ( w2345 & w2346 ) ;
  assign w2348 = w2346 | w2347 ;
  assign w2349 = \pi071 ^ w2274 ;
  assign w2350 = ( ~w2281 & w2348 ) | ( ~w2281 & w2349 ) | ( w2348 & w2349 ) ;
  assign w2351 = w2349 | w2350 ;
  assign w2352 = \pi072 ^ w2268 ;
  assign w2353 = ( ~w2275 & w2351 ) | ( ~w2275 & w2352 ) | ( w2351 & w2352 ) ;
  assign w2354 = w2352 | w2353 ;
  assign w2355 = \pi073 ^ w2262 ;
  assign w2356 = ( ~w2269 & w2354 ) | ( ~w2269 & w2355 ) | ( w2354 & w2355 ) ;
  assign w2357 = w2355 | w2356 ;
  assign w2358 = \pi074 ^ w2256 ;
  assign w2359 = ( ~w2263 & w2357 ) | ( ~w2263 & w2358 ) | ( w2357 & w2358 ) ;
  assign w2360 = w2358 | w2359 ;
  assign w2361 = \pi075 ^ w2250 ;
  assign w2362 = ( ~w2257 & w2360 ) | ( ~w2257 & w2361 ) | ( w2360 & w2361 ) ;
  assign w2363 = w2361 | w2362 ;
  assign w2364 = \pi076 ^ w2244 ;
  assign w2365 = ( ~w2251 & w2363 ) | ( ~w2251 & w2364 ) | ( w2363 & w2364 ) ;
  assign w2366 = w2364 | w2365 ;
  assign w2367 = \pi077 ^ w2238 ;
  assign w2368 = ( ~w2245 & w2366 ) | ( ~w2245 & w2367 ) | ( w2366 & w2367 ) ;
  assign w2369 = w2367 | w2368 ;
  assign w2370 = \pi078 ^ w2232 ;
  assign w2371 = ( ~w2239 & w2369 ) | ( ~w2239 & w2370 ) | ( w2369 & w2370 ) ;
  assign w2372 = w2370 | w2371 ;
  assign w2373 = \pi079 ^ w2226 ;
  assign w2374 = ( ~w2233 & w2372 ) | ( ~w2233 & w2373 ) | ( w2372 & w2373 ) ;
  assign w2375 = w2373 | w2374 ;
  assign w2376 = \pi080 ^ w2220 ;
  assign w2377 = ( ~w2227 & w2375 ) | ( ~w2227 & w2376 ) | ( w2375 & w2376 ) ;
  assign w2378 = w2376 | w2377 ;
  assign w2379 = \pi081 ^ w2214 ;
  assign w2380 = ( ~w2221 & w2378 ) | ( ~w2221 & w2379 ) | ( w2378 & w2379 ) ;
  assign w2381 = w2379 | w2380 ;
  assign w2382 = \pi082 ^ w2203 ;
  assign w2383 = ( ~w2215 & w2381 ) | ( ~w2215 & w2382 ) | ( w2381 & w2382 ) ;
  assign w2384 = w2382 | w2383 ;
  assign w2385 = \pi083 ^ w2208 ;
  assign w2386 = w2209 & ~w2385 ;
  assign w2387 = ( w2384 & w2385 ) | ( w2384 & ~w2386 ) | ( w2385 & ~w2386 ) ;
  assign w2388 = ~\pi083 & w2208 ;
  assign w2389 = w2387 & ~w2388 ;
  assign w2390 = w187 | w2389 ;
  assign w2391 = w2203 & w2390 ;
  assign w2392 = ~w2215 & w2381 ;
  assign w2393 = w2382 ^ w2392 ;
  assign w2394 = ~w2390 & w2393 ;
  assign w2395 = w2391 | w2394 ;
  assign w2396 = ~\pi083 & w2395 ;
  assign w2397 = w2214 & w2390 ;
  assign w2398 = ~w2221 & w2378 ;
  assign w2399 = w2379 ^ w2398 ;
  assign w2400 = ~w2390 & w2399 ;
  assign w2401 = w2397 | w2400 ;
  assign w2402 = ~\pi082 & w2401 ;
  assign w2403 = w2220 & w2390 ;
  assign w2404 = ~w2227 & w2375 ;
  assign w2405 = w2376 ^ w2404 ;
  assign w2406 = ~w2390 & w2405 ;
  assign w2407 = w2403 | w2406 ;
  assign w2408 = ~\pi081 & w2407 ;
  assign w2409 = w2226 & w2390 ;
  assign w2410 = ~w2233 & w2372 ;
  assign w2411 = w2373 ^ w2410 ;
  assign w2412 = ~w2390 & w2411 ;
  assign w2413 = w2409 | w2412 ;
  assign w2414 = ~\pi080 & w2413 ;
  assign w2415 = w2232 & w2390 ;
  assign w2416 = ~w2239 & w2369 ;
  assign w2417 = w2370 ^ w2416 ;
  assign w2418 = ~w2390 & w2417 ;
  assign w2419 = w2415 | w2418 ;
  assign w2420 = ~\pi079 & w2419 ;
  assign w2421 = w2238 & w2390 ;
  assign w2422 = ~w2245 & w2366 ;
  assign w2423 = w2367 ^ w2422 ;
  assign w2424 = ~w2390 & w2423 ;
  assign w2425 = w2421 | w2424 ;
  assign w2426 = ~\pi078 & w2425 ;
  assign w2427 = w2244 & w2390 ;
  assign w2428 = ~w2251 & w2363 ;
  assign w2429 = w2364 ^ w2428 ;
  assign w2430 = ~w2390 & w2429 ;
  assign w2431 = w2427 | w2430 ;
  assign w2432 = ~\pi077 & w2431 ;
  assign w2433 = w2250 & w2390 ;
  assign w2434 = ~w2257 & w2360 ;
  assign w2435 = w2361 ^ w2434 ;
  assign w2436 = ~w2390 & w2435 ;
  assign w2437 = w2433 | w2436 ;
  assign w2438 = ~\pi076 & w2437 ;
  assign w2439 = w2256 & w2390 ;
  assign w2440 = ~w2263 & w2357 ;
  assign w2441 = w2358 ^ w2440 ;
  assign w2442 = ~w2390 & w2441 ;
  assign w2443 = w2439 | w2442 ;
  assign w2444 = ~\pi075 & w2443 ;
  assign w2445 = w2262 & w2390 ;
  assign w2446 = ~w2269 & w2354 ;
  assign w2447 = w2355 ^ w2446 ;
  assign w2448 = ~w2390 & w2447 ;
  assign w2449 = w2445 | w2448 ;
  assign w2450 = ~\pi074 & w2449 ;
  assign w2451 = w2268 & w2390 ;
  assign w2452 = ~w2275 & w2351 ;
  assign w2453 = w2352 ^ w2452 ;
  assign w2454 = ~w2390 & w2453 ;
  assign w2455 = w2451 | w2454 ;
  assign w2456 = ~\pi073 & w2455 ;
  assign w2457 = w2274 & w2390 ;
  assign w2458 = ~w2281 & w2348 ;
  assign w2459 = w2349 ^ w2458 ;
  assign w2460 = ~w2390 & w2459 ;
  assign w2461 = w2457 | w2460 ;
  assign w2462 = ~\pi072 & w2461 ;
  assign w2463 = w2280 & w2390 ;
  assign w2464 = ~w2287 & w2345 ;
  assign w2465 = w2346 ^ w2464 ;
  assign w2466 = ~w2390 & w2465 ;
  assign w2467 = w2463 | w2466 ;
  assign w2468 = ~\pi071 & w2467 ;
  assign w2469 = w2286 & w2390 ;
  assign w2470 = ~w2293 & w2342 ;
  assign w2471 = w2343 ^ w2470 ;
  assign w2472 = ~w2390 & w2471 ;
  assign w2473 = w2469 | w2472 ;
  assign w2474 = ~\pi070 & w2473 ;
  assign w2475 = w2292 & w2390 ;
  assign w2476 = ~w2301 & w2339 ;
  assign w2477 = w2340 ^ w2476 ;
  assign w2478 = ~w2390 & w2477 ;
  assign w2479 = w2475 | w2478 ;
  assign w2480 = ~\pi069 & w2479 ;
  assign w2481 = w2300 & w2390 ;
  assign w2482 = ~w2312 & w2336 ;
  assign w2483 = w2337 ^ w2482 ;
  assign w2484 = ~w2390 & w2483 ;
  assign w2485 = w2481 | w2484 ;
  assign w2486 = ~\pi068 & w2485 ;
  assign w2487 = w2311 & w2390 ;
  assign w2488 = w2330 & ~w2331 ;
  assign w2489 = w2334 ^ w2488 ;
  assign w2490 = ~w2390 & w2489 ;
  assign w2491 = w2487 | w2490 ;
  assign w2492 = ~\pi067 & w2491 ;
  assign w2493 = w2327 & w2390 ;
  assign w2494 = ( ~w187 & w2318 ) | ( ~w187 & w2326 ) | ( w2318 & w2326 ) ;
  assign w2495 = \pi065 ^ w2494 ;
  assign w2496 = ( ~w187 & w2328 ) | ( ~w187 & w2495 ) | ( w2328 & w2495 ) ;
  assign w2497 = ( w2328 & w2389 ) | ( w2328 & w2495 ) | ( w2389 & w2495 ) ;
  assign w2498 = w2496 & ~w2497 ;
  assign w2499 = w2493 | w2498 ;
  assign w2500 = ~\pi066 & w2499 ;
  assign w2501 = ( \pi064 & w234 ) | ( \pi064 & w244 ) | ( w234 & w244 ) ;
  assign w2502 = ( \pi064 & ~\pi084 ) | ( \pi064 & w290 ) | ( ~\pi084 & w290 ) ;
  assign w2503 = ~w291 & w2502 ;
  assign w2504 = ~w2501 & w2503 ;
  assign w2505 = ~w176 & w2328 ;
  assign w2506 = ~w204 & w2505 ;
  assign w2507 = ( w201 & ~w204 ) | ( w201 & w205 ) | ( ~w204 & w205 ) ;
  assign w2508 = w2506 & ~w2507 ;
  assign w2509 = ( \pi044 & w2389 ) | ( \pi044 & ~w2504 ) | ( w2389 & ~w2504 ) ;
  assign w2510 = \pi044 & w2509 ;
  assign w2511 = w2389 | w2508 ;
  assign w2512 = ( ~w2389 & w2510 ) | ( ~w2389 & w2511 ) | ( w2510 & w2511 ) ;
  assign w2513 = ~\pi043 & \pi064 ;
  assign w2514 = w2504 & ~w2511 ;
  assign w2515 = \pi044 & ~w2514 ;
  assign w2516 = ( ~w2389 & w2511 ) | ( ~w2389 & w2515 ) | ( w2511 & w2515 ) ;
  assign w2517 = \pi065 ^ w2516 ;
  assign w2518 = w2513 | w2517 ;
  assign w2519 = ~\pi065 & w2512 ;
  assign w2520 = \pi066 ^ w2499 ;
  assign w2521 = ( w2518 & ~w2519 ) | ( w2518 & w2520 ) | ( ~w2519 & w2520 ) ;
  assign w2522 = w2520 | w2521 ;
  assign w2523 = \pi067 ^ w2491 ;
  assign w2524 = ( ~w2500 & w2522 ) | ( ~w2500 & w2523 ) | ( w2522 & w2523 ) ;
  assign w2525 = w2523 | w2524 ;
  assign w2526 = \pi068 ^ w2485 ;
  assign w2527 = ( ~w2492 & w2525 ) | ( ~w2492 & w2526 ) | ( w2525 & w2526 ) ;
  assign w2528 = w2526 | w2527 ;
  assign w2529 = \pi069 ^ w2479 ;
  assign w2530 = ( ~w2486 & w2528 ) | ( ~w2486 & w2529 ) | ( w2528 & w2529 ) ;
  assign w2531 = w2529 | w2530 ;
  assign w2532 = \pi070 ^ w2473 ;
  assign w2533 = ( ~w2480 & w2531 ) | ( ~w2480 & w2532 ) | ( w2531 & w2532 ) ;
  assign w2534 = w2532 | w2533 ;
  assign w2535 = \pi071 ^ w2467 ;
  assign w2536 = ( ~w2474 & w2534 ) | ( ~w2474 & w2535 ) | ( w2534 & w2535 ) ;
  assign w2537 = w2535 | w2536 ;
  assign w2538 = \pi072 ^ w2461 ;
  assign w2539 = ( ~w2468 & w2537 ) | ( ~w2468 & w2538 ) | ( w2537 & w2538 ) ;
  assign w2540 = w2538 | w2539 ;
  assign w2541 = \pi073 ^ w2455 ;
  assign w2542 = ( ~w2462 & w2540 ) | ( ~w2462 & w2541 ) | ( w2540 & w2541 ) ;
  assign w2543 = w2541 | w2542 ;
  assign w2544 = \pi074 ^ w2449 ;
  assign w2545 = ( ~w2456 & w2543 ) | ( ~w2456 & w2544 ) | ( w2543 & w2544 ) ;
  assign w2546 = w2544 | w2545 ;
  assign w2547 = \pi075 ^ w2443 ;
  assign w2548 = ( ~w2450 & w2546 ) | ( ~w2450 & w2547 ) | ( w2546 & w2547 ) ;
  assign w2549 = w2547 | w2548 ;
  assign w2550 = \pi076 ^ w2437 ;
  assign w2551 = ( ~w2444 & w2549 ) | ( ~w2444 & w2550 ) | ( w2549 & w2550 ) ;
  assign w2552 = w2550 | w2551 ;
  assign w2553 = \pi077 ^ w2431 ;
  assign w2554 = ( ~w2438 & w2552 ) | ( ~w2438 & w2553 ) | ( w2552 & w2553 ) ;
  assign w2555 = w2553 | w2554 ;
  assign w2556 = \pi078 ^ w2425 ;
  assign w2557 = ( ~w2432 & w2555 ) | ( ~w2432 & w2556 ) | ( w2555 & w2556 ) ;
  assign w2558 = w2556 | w2557 ;
  assign w2559 = \pi079 ^ w2419 ;
  assign w2560 = ( ~w2426 & w2558 ) | ( ~w2426 & w2559 ) | ( w2558 & w2559 ) ;
  assign w2561 = w2559 | w2560 ;
  assign w2562 = \pi080 ^ w2413 ;
  assign w2563 = ( ~w2420 & w2561 ) | ( ~w2420 & w2562 ) | ( w2561 & w2562 ) ;
  assign w2564 = w2562 | w2563 ;
  assign w2565 = \pi081 ^ w2407 ;
  assign w2566 = ( ~w2414 & w2564 ) | ( ~w2414 & w2565 ) | ( w2564 & w2565 ) ;
  assign w2567 = w2565 | w2566 ;
  assign w2568 = \pi082 ^ w2401 ;
  assign w2569 = ( ~w2408 & w2567 ) | ( ~w2408 & w2568 ) | ( w2567 & w2568 ) ;
  assign w2570 = w2568 | w2569 ;
  assign w2571 = \pi083 ^ w2395 ;
  assign w2572 = ( ~w2402 & w2570 ) | ( ~w2402 & w2571 ) | ( w2570 & w2571 ) ;
  assign w2573 = w2571 | w2572 ;
  assign w2574 = w2208 & w2390 ;
  assign w2575 = ~w2209 & w2384 ;
  assign w2576 = w2385 ^ w2575 ;
  assign w2577 = ~w2390 & w2576 ;
  assign w2578 = w2574 | w2577 ;
  assign w2579 = ~\pi084 & w2578 ;
  assign w2580 = ( \pi084 & ~w2574 ) | ( \pi084 & w2577 ) | ( ~w2574 & w2577 ) ;
  assign w2581 = ~w2577 & w2580 ;
  assign w2582 = w2579 | w2581 ;
  assign w2583 = ( ~w2396 & w2573 ) | ( ~w2396 & w2582 ) | ( w2573 & w2582 ) ;
  assign w2584 = ( w491 & ~w2582 ) | ( w491 & w2583 ) | ( ~w2582 & w2583 ) ;
  assign w2585 = w2582 | w2584 ;
  assign w2586 = ~w187 & w2578 ;
  assign w2587 = w2585 & ~w2586 ;
  assign w2588 = ~w2402 & w2570 ;
  assign w2589 = w2571 ^ w2588 ;
  assign w2590 = ~w2587 & w2589 ;
  assign w2591 = ( w2395 & w2585 ) | ( w2395 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2592 = ~w2586 & w2591 ;
  assign w2593 = w2590 | w2592 ;
  assign w2594 = ( ~w2396 & w2573 ) | ( ~w2396 & w2587 ) | ( w2573 & w2587 ) ;
  assign w2595 = w2582 ^ w2594 ;
  assign w2596 = ~w2587 & w2595 ;
  assign w2597 = ( w187 & ~w2578 ) | ( w187 & w2585 ) | ( ~w2578 & w2585 ) ;
  assign w2598 = w2578 & w2597 ;
  assign w2599 = w2596 | w2598 ;
  assign w2600 = ~\pi084 & w2593 ;
  assign w2601 = ~w2408 & w2567 ;
  assign w2602 = w2568 ^ w2601 ;
  assign w2603 = ~w2587 & w2602 ;
  assign w2604 = ( w2401 & w2585 ) | ( w2401 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2605 = ~w2586 & w2604 ;
  assign w2606 = w2603 | w2605 ;
  assign w2607 = ~\pi083 & w2606 ;
  assign w2608 = ~w2414 & w2564 ;
  assign w2609 = w2565 ^ w2608 ;
  assign w2610 = ~w2587 & w2609 ;
  assign w2611 = ( w2407 & w2585 ) | ( w2407 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2612 = ~w2586 & w2611 ;
  assign w2613 = w2610 | w2612 ;
  assign w2614 = ~\pi082 & w2613 ;
  assign w2615 = ~w2420 & w2561 ;
  assign w2616 = w2562 ^ w2615 ;
  assign w2617 = ~w2587 & w2616 ;
  assign w2618 = ( w2413 & w2585 ) | ( w2413 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2619 = ~w2586 & w2618 ;
  assign w2620 = w2617 | w2619 ;
  assign w2621 = ~\pi081 & w2620 ;
  assign w2622 = ~w2426 & w2558 ;
  assign w2623 = w2559 ^ w2622 ;
  assign w2624 = ~w2587 & w2623 ;
  assign w2625 = ( w2419 & w2585 ) | ( w2419 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2626 = ~w2586 & w2625 ;
  assign w2627 = w2624 | w2626 ;
  assign w2628 = ~\pi080 & w2627 ;
  assign w2629 = ~w2432 & w2555 ;
  assign w2630 = w2556 ^ w2629 ;
  assign w2631 = ~w2587 & w2630 ;
  assign w2632 = ( w2425 & w2585 ) | ( w2425 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2633 = ~w2586 & w2632 ;
  assign w2634 = w2631 | w2633 ;
  assign w2635 = ~\pi079 & w2634 ;
  assign w2636 = ~w2438 & w2552 ;
  assign w2637 = w2553 ^ w2636 ;
  assign w2638 = ~w2587 & w2637 ;
  assign w2639 = ( w2431 & w2585 ) | ( w2431 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2640 = ~w2586 & w2639 ;
  assign w2641 = w2638 | w2640 ;
  assign w2642 = ~\pi078 & w2641 ;
  assign w2643 = ~w2444 & w2549 ;
  assign w2644 = w2550 ^ w2643 ;
  assign w2645 = ~w2587 & w2644 ;
  assign w2646 = ( w2437 & w2585 ) | ( w2437 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2647 = ~w2586 & w2646 ;
  assign w2648 = w2645 | w2647 ;
  assign w2649 = ~\pi077 & w2648 ;
  assign w2650 = ~w2450 & w2546 ;
  assign w2651 = w2547 ^ w2650 ;
  assign w2652 = ~w2587 & w2651 ;
  assign w2653 = ( w2443 & w2585 ) | ( w2443 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2654 = ~w2586 & w2653 ;
  assign w2655 = w2652 | w2654 ;
  assign w2656 = ~\pi076 & w2655 ;
  assign w2657 = ~w2456 & w2543 ;
  assign w2658 = w2544 ^ w2657 ;
  assign w2659 = ~w2587 & w2658 ;
  assign w2660 = ( w2449 & w2585 ) | ( w2449 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2661 = ~w2586 & w2660 ;
  assign w2662 = w2659 | w2661 ;
  assign w2663 = ~\pi075 & w2662 ;
  assign w2664 = ~w2462 & w2540 ;
  assign w2665 = w2541 ^ w2664 ;
  assign w2666 = ~w2587 & w2665 ;
  assign w2667 = ( w2455 & w2585 ) | ( w2455 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2668 = ~w2586 & w2667 ;
  assign w2669 = w2666 | w2668 ;
  assign w2670 = ~\pi074 & w2669 ;
  assign w2671 = ~w2468 & w2537 ;
  assign w2672 = w2538 ^ w2671 ;
  assign w2673 = ~w2587 & w2672 ;
  assign w2674 = ( w2461 & w2585 ) | ( w2461 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2675 = ~w2586 & w2674 ;
  assign w2676 = w2673 | w2675 ;
  assign w2677 = ~\pi073 & w2676 ;
  assign w2678 = ~w2474 & w2534 ;
  assign w2679 = w2535 ^ w2678 ;
  assign w2680 = ~w2587 & w2679 ;
  assign w2681 = ( w2467 & w2585 ) | ( w2467 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2682 = ~w2586 & w2681 ;
  assign w2683 = w2680 | w2682 ;
  assign w2684 = ~\pi072 & w2683 ;
  assign w2685 = ~w2480 & w2531 ;
  assign w2686 = w2532 ^ w2685 ;
  assign w2687 = ~w2587 & w2686 ;
  assign w2688 = ( w2473 & w2585 ) | ( w2473 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2689 = ~w2586 & w2688 ;
  assign w2690 = w2687 | w2689 ;
  assign w2691 = ~\pi071 & w2690 ;
  assign w2692 = ~w2486 & w2528 ;
  assign w2693 = w2529 ^ w2692 ;
  assign w2694 = ~w2587 & w2693 ;
  assign w2695 = ( w2479 & w2585 ) | ( w2479 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2696 = ~w2586 & w2695 ;
  assign w2697 = w2694 | w2696 ;
  assign w2698 = ~\pi070 & w2697 ;
  assign w2699 = ~w2492 & w2525 ;
  assign w2700 = w2526 ^ w2699 ;
  assign w2701 = ~w2587 & w2700 ;
  assign w2702 = ( w2485 & w2585 ) | ( w2485 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2703 = ~w2586 & w2702 ;
  assign w2704 = w2701 | w2703 ;
  assign w2705 = ~\pi069 & w2704 ;
  assign w2706 = ~w2500 & w2522 ;
  assign w2707 = w2523 ^ w2706 ;
  assign w2708 = ~w2587 & w2707 ;
  assign w2709 = ( w2491 & w2585 ) | ( w2491 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2710 = ~w2586 & w2709 ;
  assign w2711 = w2708 | w2710 ;
  assign w2712 = ~\pi068 & w2711 ;
  assign w2713 = w2518 & ~w2519 ;
  assign w2714 = w2520 ^ w2713 ;
  assign w2715 = ~w2587 & w2714 ;
  assign w2716 = ( w2499 & w2585 ) | ( w2499 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2717 = ~w2586 & w2716 ;
  assign w2718 = w2715 | w2717 ;
  assign w2719 = ~\pi067 & w2718 ;
  assign w2720 = w2504 & ~w2508 ;
  assign w2721 = w2389 ^ w2508 ;
  assign w2722 = ( \pi044 & ~w2720 ) | ( \pi044 & w2721 ) | ( ~w2720 & w2721 ) ;
  assign w2723 = ( \pi044 & w2508 ) | ( \pi044 & w2722 ) | ( w2508 & w2722 ) ;
  assign w2724 = w2513 ^ w2723 ;
  assign w2725 = \pi065 ^ w2724 ;
  assign w2726 = ~w2587 & w2725 ;
  assign w2727 = ( w2512 & w2585 ) | ( w2512 & w2586 ) | ( w2585 & w2586 ) ;
  assign w2728 = ~w2586 & w2727 ;
  assign w2729 = w2726 | w2728 ;
  assign w2730 = ~\pi066 & w2729 ;
  assign w2731 = \pi066 ^ w2729 ;
  assign w2732 = \pi064 & ~w2587 ;
  assign w2733 = \pi043 ^ w2732 ;
  assign w2734 = ( ~\pi042 & \pi064 ) | ( ~\pi042 & w2731 ) | ( \pi064 & w2731 ) ;
  assign w2735 = ( \pi065 & ~w2733 ) | ( \pi065 & w2734 ) | ( ~w2733 & w2734 ) ;
  assign w2736 = w2731 | w2735 ;
  assign w2737 = \pi067 ^ w2718 ;
  assign w2738 = ( ~w2730 & w2736 ) | ( ~w2730 & w2737 ) | ( w2736 & w2737 ) ;
  assign w2739 = w2737 | w2738 ;
  assign w2740 = \pi068 ^ w2711 ;
  assign w2741 = ( ~w2719 & w2739 ) | ( ~w2719 & w2740 ) | ( w2739 & w2740 ) ;
  assign w2742 = w2740 | w2741 ;
  assign w2743 = \pi069 ^ w2704 ;
  assign w2744 = ( ~w2712 & w2742 ) | ( ~w2712 & w2743 ) | ( w2742 & w2743 ) ;
  assign w2745 = w2743 | w2744 ;
  assign w2746 = \pi070 ^ w2697 ;
  assign w2747 = ( ~w2705 & w2745 ) | ( ~w2705 & w2746 ) | ( w2745 & w2746 ) ;
  assign w2748 = w2746 | w2747 ;
  assign w2749 = \pi071 ^ w2690 ;
  assign w2750 = ( ~w2698 & w2748 ) | ( ~w2698 & w2749 ) | ( w2748 & w2749 ) ;
  assign w2751 = w2749 | w2750 ;
  assign w2752 = \pi072 ^ w2683 ;
  assign w2753 = ( ~w2691 & w2751 ) | ( ~w2691 & w2752 ) | ( w2751 & w2752 ) ;
  assign w2754 = w2752 | w2753 ;
  assign w2755 = \pi073 ^ w2676 ;
  assign w2756 = ( ~w2684 & w2754 ) | ( ~w2684 & w2755 ) | ( w2754 & w2755 ) ;
  assign w2757 = w2755 | w2756 ;
  assign w2758 = \pi074 ^ w2669 ;
  assign w2759 = ( ~w2677 & w2757 ) | ( ~w2677 & w2758 ) | ( w2757 & w2758 ) ;
  assign w2760 = w2758 | w2759 ;
  assign w2761 = \pi075 ^ w2662 ;
  assign w2762 = ( ~w2670 & w2760 ) | ( ~w2670 & w2761 ) | ( w2760 & w2761 ) ;
  assign w2763 = w2761 | w2762 ;
  assign w2764 = \pi076 ^ w2655 ;
  assign w2765 = ( ~w2663 & w2763 ) | ( ~w2663 & w2764 ) | ( w2763 & w2764 ) ;
  assign w2766 = w2764 | w2765 ;
  assign w2767 = \pi077 ^ w2648 ;
  assign w2768 = ( ~w2656 & w2766 ) | ( ~w2656 & w2767 ) | ( w2766 & w2767 ) ;
  assign w2769 = w2767 | w2768 ;
  assign w2770 = \pi078 ^ w2641 ;
  assign w2771 = ( ~w2649 & w2769 ) | ( ~w2649 & w2770 ) | ( w2769 & w2770 ) ;
  assign w2772 = w2770 | w2771 ;
  assign w2773 = \pi079 ^ w2634 ;
  assign w2774 = ( ~w2642 & w2772 ) | ( ~w2642 & w2773 ) | ( w2772 & w2773 ) ;
  assign w2775 = w2773 | w2774 ;
  assign w2776 = \pi080 ^ w2627 ;
  assign w2777 = ( ~w2635 & w2775 ) | ( ~w2635 & w2776 ) | ( w2775 & w2776 ) ;
  assign w2778 = w2776 | w2777 ;
  assign w2779 = \pi081 ^ w2620 ;
  assign w2780 = ( ~w2628 & w2778 ) | ( ~w2628 & w2779 ) | ( w2778 & w2779 ) ;
  assign w2781 = w2779 | w2780 ;
  assign w2782 = \pi082 ^ w2613 ;
  assign w2783 = ( ~w2621 & w2781 ) | ( ~w2621 & w2782 ) | ( w2781 & w2782 ) ;
  assign w2784 = w2782 | w2783 ;
  assign w2785 = \pi083 ^ w2606 ;
  assign w2786 = ( ~w2614 & w2784 ) | ( ~w2614 & w2785 ) | ( w2784 & w2785 ) ;
  assign w2787 = w2785 | w2786 ;
  assign w2788 = \pi084 ^ w2593 ;
  assign w2789 = ( ~w2607 & w2787 ) | ( ~w2607 & w2788 ) | ( w2787 & w2788 ) ;
  assign w2790 = w2788 | w2789 ;
  assign w2791 = \pi085 ^ w2599 ;
  assign w2792 = w2600 & ~w2791 ;
  assign w2793 = ( w2790 & w2791 ) | ( w2790 & ~w2792 ) | ( w2791 & ~w2792 ) ;
  assign w2794 = ~\pi085 & w2599 ;
  assign w2795 = w2793 & ~w2794 ;
  assign w2796 = ( ~\pi086 & w173 ) | ( ~\pi086 & w183 ) | ( w173 & w183 ) ;
  assign w2797 = ( \pi086 & \pi087 ) | ( \pi086 & ~w155 ) | ( \pi087 & ~w155 ) ;
  assign w2798 = w368 | w2797 ;
  assign w2799 = w2796 | w2798 ;
  assign w2800 = w2795 | w2799 ;
  assign w2801 = w2593 & w2800 ;
  assign w2802 = ~w2607 & w2787 ;
  assign w2803 = w2788 ^ w2802 ;
  assign w2804 = ~w2800 & w2803 ;
  assign w2805 = w2801 | w2804 ;
  assign w2806 = w2599 & w2800 ;
  assign w2807 = ~w2600 & w2790 ;
  assign w2808 = w2791 ^ w2807 ;
  assign w2809 = ~w2800 & w2808 ;
  assign w2810 = w2806 | w2809 ;
  assign w2811 = ~\pi085 & w2805 ;
  assign w2812 = w2606 & w2800 ;
  assign w2813 = ~w2614 & w2784 ;
  assign w2814 = w2785 ^ w2813 ;
  assign w2815 = ~w2800 & w2814 ;
  assign w2816 = w2812 | w2815 ;
  assign w2817 = ~\pi084 & w2816 ;
  assign w2818 = w2613 & w2800 ;
  assign w2819 = ~w2621 & w2781 ;
  assign w2820 = w2782 ^ w2819 ;
  assign w2821 = ~w2800 & w2820 ;
  assign w2822 = w2818 | w2821 ;
  assign w2823 = ~\pi083 & w2822 ;
  assign w2824 = w2620 & w2800 ;
  assign w2825 = ~w2628 & w2778 ;
  assign w2826 = w2779 ^ w2825 ;
  assign w2827 = ~w2800 & w2826 ;
  assign w2828 = w2824 | w2827 ;
  assign w2829 = ~\pi082 & w2828 ;
  assign w2830 = w2627 & w2800 ;
  assign w2831 = ~w2635 & w2775 ;
  assign w2832 = w2776 ^ w2831 ;
  assign w2833 = ~w2800 & w2832 ;
  assign w2834 = w2830 | w2833 ;
  assign w2835 = ~\pi081 & w2834 ;
  assign w2836 = w2634 & w2800 ;
  assign w2837 = ~w2642 & w2772 ;
  assign w2838 = w2773 ^ w2837 ;
  assign w2839 = ~w2800 & w2838 ;
  assign w2840 = w2836 | w2839 ;
  assign w2841 = ~\pi080 & w2840 ;
  assign w2842 = w2641 & w2800 ;
  assign w2843 = ~w2649 & w2769 ;
  assign w2844 = w2770 ^ w2843 ;
  assign w2845 = ~w2800 & w2844 ;
  assign w2846 = w2842 | w2845 ;
  assign w2847 = ~\pi079 & w2846 ;
  assign w2848 = w2648 & w2800 ;
  assign w2849 = ~w2656 & w2766 ;
  assign w2850 = w2767 ^ w2849 ;
  assign w2851 = ~w2800 & w2850 ;
  assign w2852 = w2848 | w2851 ;
  assign w2853 = ~\pi078 & w2852 ;
  assign w2854 = w2655 & w2800 ;
  assign w2855 = ~w2663 & w2763 ;
  assign w2856 = w2764 ^ w2855 ;
  assign w2857 = ~w2800 & w2856 ;
  assign w2858 = w2854 | w2857 ;
  assign w2859 = ~\pi077 & w2858 ;
  assign w2860 = w2662 & w2800 ;
  assign w2861 = ~w2670 & w2760 ;
  assign w2862 = w2761 ^ w2861 ;
  assign w2863 = ~w2800 & w2862 ;
  assign w2864 = w2860 | w2863 ;
  assign w2865 = ~\pi076 & w2864 ;
  assign w2866 = w2669 & w2800 ;
  assign w2867 = ~w2677 & w2757 ;
  assign w2868 = w2758 ^ w2867 ;
  assign w2869 = ~w2800 & w2868 ;
  assign w2870 = w2866 | w2869 ;
  assign w2871 = ~\pi075 & w2870 ;
  assign w2872 = w2676 & w2800 ;
  assign w2873 = ~w2684 & w2754 ;
  assign w2874 = w2755 ^ w2873 ;
  assign w2875 = ~w2800 & w2874 ;
  assign w2876 = w2872 | w2875 ;
  assign w2877 = ~\pi074 & w2876 ;
  assign w2878 = w2683 & w2800 ;
  assign w2879 = ~w2691 & w2751 ;
  assign w2880 = w2752 ^ w2879 ;
  assign w2881 = ~w2800 & w2880 ;
  assign w2882 = w2878 | w2881 ;
  assign w2883 = ~\pi073 & w2882 ;
  assign w2884 = w2690 & w2800 ;
  assign w2885 = ~w2698 & w2748 ;
  assign w2886 = w2749 ^ w2885 ;
  assign w2887 = ~w2800 & w2886 ;
  assign w2888 = w2884 | w2887 ;
  assign w2889 = ~\pi072 & w2888 ;
  assign w2890 = w2697 & w2800 ;
  assign w2891 = ~w2705 & w2745 ;
  assign w2892 = w2746 ^ w2891 ;
  assign w2893 = ~w2800 & w2892 ;
  assign w2894 = w2890 | w2893 ;
  assign w2895 = ~\pi071 & w2894 ;
  assign w2896 = w2704 & w2800 ;
  assign w2897 = ~w2712 & w2742 ;
  assign w2898 = w2743 ^ w2897 ;
  assign w2899 = ~w2800 & w2898 ;
  assign w2900 = w2896 | w2899 ;
  assign w2901 = ~\pi070 & w2900 ;
  assign w2902 = w2711 & w2800 ;
  assign w2903 = ~w2719 & w2739 ;
  assign w2904 = w2740 ^ w2903 ;
  assign w2905 = ~w2800 & w2904 ;
  assign w2906 = w2902 | w2905 ;
  assign w2907 = ~\pi069 & w2906 ;
  assign w2908 = w2718 & w2800 ;
  assign w2909 = ~w2730 & w2736 ;
  assign w2910 = w2737 ^ w2909 ;
  assign w2911 = ~w2800 & w2910 ;
  assign w2912 = w2908 | w2911 ;
  assign w2913 = ~\pi068 & w2912 ;
  assign w2914 = w2729 & w2800 ;
  assign w2915 = ~\pi042 & \pi064 ;
  assign w2916 = ( \pi065 & ~w2733 ) | ( \pi065 & w2915 ) | ( ~w2733 & w2915 ) ;
  assign w2917 = w2731 ^ w2916 ;
  assign w2918 = ( w2795 & w2799 ) | ( w2795 & w2917 ) | ( w2799 & w2917 ) ;
  assign w2919 = w2917 & ~w2918 ;
  assign w2920 = w2914 | w2919 ;
  assign w2921 = ~\pi067 & w2920 ;
  assign w2922 = \pi043 ^ \pi065 ;
  assign w2923 = \pi042 ^ w2587 ;
  assign w2924 = ( \pi064 & w2799 ) | ( \pi064 & w2923 ) | ( w2799 & w2923 ) ;
  assign w2925 = w2922 ^ w2924 ;
  assign w2926 = ~w2799 & w2925 ;
  assign w2927 = ~w2795 & w2926 ;
  assign w2928 = ( ~\pi064 & w2587 ) | ( ~\pi064 & w2800 ) | ( w2587 & w2800 ) ;
  assign w2929 = \pi043 ^ w2928 ;
  assign w2930 = w2800 & ~w2929 ;
  assign w2931 = w2927 | w2930 ;
  assign w2932 = ~\pi066 & w2931 ;
  assign w2933 = ( \pi064 & ~\pi086 ) | ( \pi064 & \pi087 ) | ( ~\pi086 & \pi087 ) ;
  assign w2934 = w243 | w441 ;
  assign w2935 = ( \pi087 & \pi088 ) | ( \pi087 & ~w243 ) | ( \pi088 & ~w243 ) ;
  assign w2936 = w2934 | w2935 ;
  assign w2937 = w2933 & ~w2936 ;
  assign w2938 = ( ~w448 & w451 ) | ( ~w448 & w2937 ) | ( w451 & w2937 ) ;
  assign w2939 = ~w451 & w2938 ;
  assign w2940 = ( \pi042 & w2795 ) | ( \pi042 & ~w2939 ) | ( w2795 & ~w2939 ) ;
  assign w2941 = \pi042 & w2940 ;
  assign w2942 = ( ~\pi042 & \pi064 ) | ( ~\pi042 & \pi086 ) | ( \pi064 & \pi086 ) ;
  assign w2943 = w173 | w183 ;
  assign w2944 = ( \pi086 & \pi087 ) | ( \pi086 & ~w173 ) | ( \pi087 & ~w173 ) ;
  assign w2945 = w2943 | w2944 ;
  assign w2946 = w2942 & ~w2945 ;
  assign w2947 = ( w155 & w170 ) | ( w155 & w2946 ) | ( w170 & w2946 ) ;
  assign w2948 = w2946 & ~w2947 ;
  assign w2949 = ~w2795 & w2948 ;
  assign w2950 = w2941 | w2949 ;
  assign w2951 = ~\pi041 & \pi064 ;
  assign w2952 = \pi065 ^ w2950 ;
  assign w2953 = w2951 | w2952 ;
  assign w2954 = ~\pi065 & w2950 ;
  assign w2955 = w2800 | w2927 ;
  assign w2956 = ( w2733 & w2927 ) | ( w2733 & w2955 ) | ( w2927 & w2955 ) ;
  assign w2957 = \pi066 ^ w2956 ;
  assign w2958 = ( w2953 & ~w2954 ) | ( w2953 & w2957 ) | ( ~w2954 & w2957 ) ;
  assign w2959 = w2957 | w2958 ;
  assign w2960 = \pi067 ^ w2920 ;
  assign w2961 = ( ~w2932 & w2959 ) | ( ~w2932 & w2960 ) | ( w2959 & w2960 ) ;
  assign w2962 = w2960 | w2961 ;
  assign w2963 = \pi068 ^ w2912 ;
  assign w2964 = ( ~w2921 & w2962 ) | ( ~w2921 & w2963 ) | ( w2962 & w2963 ) ;
  assign w2965 = w2963 | w2964 ;
  assign w2966 = \pi069 ^ w2906 ;
  assign w2967 = ( ~w2913 & w2965 ) | ( ~w2913 & w2966 ) | ( w2965 & w2966 ) ;
  assign w2968 = w2966 | w2967 ;
  assign w2969 = \pi070 ^ w2900 ;
  assign w2970 = ( ~w2907 & w2968 ) | ( ~w2907 & w2969 ) | ( w2968 & w2969 ) ;
  assign w2971 = w2969 | w2970 ;
  assign w2972 = \pi071 ^ w2894 ;
  assign w2973 = ( ~w2901 & w2971 ) | ( ~w2901 & w2972 ) | ( w2971 & w2972 ) ;
  assign w2974 = w2972 | w2973 ;
  assign w2975 = \pi072 ^ w2888 ;
  assign w2976 = ( ~w2895 & w2974 ) | ( ~w2895 & w2975 ) | ( w2974 & w2975 ) ;
  assign w2977 = w2975 | w2976 ;
  assign w2978 = \pi073 ^ w2882 ;
  assign w2979 = ( ~w2889 & w2977 ) | ( ~w2889 & w2978 ) | ( w2977 & w2978 ) ;
  assign w2980 = w2978 | w2979 ;
  assign w2981 = \pi074 ^ w2876 ;
  assign w2982 = ( ~w2883 & w2980 ) | ( ~w2883 & w2981 ) | ( w2980 & w2981 ) ;
  assign w2983 = w2981 | w2982 ;
  assign w2984 = \pi075 ^ w2870 ;
  assign w2985 = ( ~w2877 & w2983 ) | ( ~w2877 & w2984 ) | ( w2983 & w2984 ) ;
  assign w2986 = w2984 | w2985 ;
  assign w2987 = \pi076 ^ w2864 ;
  assign w2988 = ( ~w2871 & w2986 ) | ( ~w2871 & w2987 ) | ( w2986 & w2987 ) ;
  assign w2989 = w2987 | w2988 ;
  assign w2990 = \pi077 ^ w2858 ;
  assign w2991 = ( ~w2865 & w2989 ) | ( ~w2865 & w2990 ) | ( w2989 & w2990 ) ;
  assign w2992 = w2990 | w2991 ;
  assign w2993 = \pi078 ^ w2852 ;
  assign w2994 = ( ~w2859 & w2992 ) | ( ~w2859 & w2993 ) | ( w2992 & w2993 ) ;
  assign w2995 = w2993 | w2994 ;
  assign w2996 = \pi079 ^ w2846 ;
  assign w2997 = ( ~w2853 & w2995 ) | ( ~w2853 & w2996 ) | ( w2995 & w2996 ) ;
  assign w2998 = w2996 | w2997 ;
  assign w2999 = \pi080 ^ w2840 ;
  assign w3000 = ( ~w2847 & w2998 ) | ( ~w2847 & w2999 ) | ( w2998 & w2999 ) ;
  assign w3001 = w2999 | w3000 ;
  assign w3002 = \pi081 ^ w2834 ;
  assign w3003 = ( ~w2841 & w3001 ) | ( ~w2841 & w3002 ) | ( w3001 & w3002 ) ;
  assign w3004 = w3002 | w3003 ;
  assign w3005 = \pi082 ^ w2828 ;
  assign w3006 = ( ~w2835 & w3004 ) | ( ~w2835 & w3005 ) | ( w3004 & w3005 ) ;
  assign w3007 = w3005 | w3006 ;
  assign w3008 = \pi083 ^ w2822 ;
  assign w3009 = ( ~w2829 & w3007 ) | ( ~w2829 & w3008 ) | ( w3007 & w3008 ) ;
  assign w3010 = w3008 | w3009 ;
  assign w3011 = \pi084 ^ w2816 ;
  assign w3012 = ( ~w2823 & w3010 ) | ( ~w2823 & w3011 ) | ( w3010 & w3011 ) ;
  assign w3013 = w3011 | w3012 ;
  assign w3014 = \pi085 ^ w2805 ;
  assign w3015 = ( ~w2817 & w3013 ) | ( ~w2817 & w3014 ) | ( w3013 & w3014 ) ;
  assign w3016 = w3014 | w3015 ;
  assign w3017 = \pi086 ^ w2810 ;
  assign w3018 = w2811 & ~w3017 ;
  assign w3019 = ( w3016 & w3017 ) | ( w3016 & ~w3018 ) | ( w3017 & ~w3018 ) ;
  assign w3020 = ~\pi086 & w2810 ;
  assign w3021 = w3019 & ~w3020 ;
  assign w3022 = ( ~\pi087 & w243 ) | ( ~\pi087 & w441 ) | ( w243 & w441 ) ;
  assign w3023 = ( \pi087 & \pi088 ) | ( \pi087 & ~w451 ) | ( \pi088 & ~w451 ) ;
  assign w3024 = w452 | w3023 ;
  assign w3025 = w3022 | w3024 ;
  assign w3026 = w3021 | w3025 ;
  assign w3027 = w2805 & w3026 ;
  assign w3028 = ~w2817 & w3013 ;
  assign w3029 = w3014 ^ w3028 ;
  assign w3030 = ~w3026 & w3029 ;
  assign w3031 = w3027 | w3030 ;
  assign w3032 = ~\pi086 & w3031 ;
  assign w3033 = w2816 & w3026 ;
  assign w3034 = ~w2823 & w3010 ;
  assign w3035 = w3011 ^ w3034 ;
  assign w3036 = ~w3026 & w3035 ;
  assign w3037 = w3033 | w3036 ;
  assign w3038 = ~\pi085 & w3037 ;
  assign w3039 = w2822 & w3026 ;
  assign w3040 = ~w2829 & w3007 ;
  assign w3041 = w3008 ^ w3040 ;
  assign w3042 = ~w3026 & w3041 ;
  assign w3043 = w3039 | w3042 ;
  assign w3044 = ~\pi084 & w3043 ;
  assign w3045 = w2828 & w3026 ;
  assign w3046 = ~w2835 & w3004 ;
  assign w3047 = w3005 ^ w3046 ;
  assign w3048 = ~w3026 & w3047 ;
  assign w3049 = w3045 | w3048 ;
  assign w3050 = ~\pi083 & w3049 ;
  assign w3051 = w2834 & w3026 ;
  assign w3052 = ~w2841 & w3001 ;
  assign w3053 = w3002 ^ w3052 ;
  assign w3054 = ~w3026 & w3053 ;
  assign w3055 = w3051 | w3054 ;
  assign w3056 = ~\pi082 & w3055 ;
  assign w3057 = w2840 & w3026 ;
  assign w3058 = ~w2847 & w2998 ;
  assign w3059 = w2999 ^ w3058 ;
  assign w3060 = ~w3026 & w3059 ;
  assign w3061 = w3057 | w3060 ;
  assign w3062 = ~\pi081 & w3061 ;
  assign w3063 = w2846 & w3026 ;
  assign w3064 = ~w2853 & w2995 ;
  assign w3065 = w2996 ^ w3064 ;
  assign w3066 = ~w3026 & w3065 ;
  assign w3067 = w3063 | w3066 ;
  assign w3068 = ~\pi080 & w3067 ;
  assign w3069 = w2852 & w3026 ;
  assign w3070 = ~w2859 & w2992 ;
  assign w3071 = w2993 ^ w3070 ;
  assign w3072 = ~w3026 & w3071 ;
  assign w3073 = w3069 | w3072 ;
  assign w3074 = ~\pi079 & w3073 ;
  assign w3075 = w2858 & w3026 ;
  assign w3076 = ~w2865 & w2989 ;
  assign w3077 = w2990 ^ w3076 ;
  assign w3078 = ~w3026 & w3077 ;
  assign w3079 = w3075 | w3078 ;
  assign w3080 = ~\pi078 & w3079 ;
  assign w3081 = w2864 & w3026 ;
  assign w3082 = ~w2871 & w2986 ;
  assign w3083 = w2987 ^ w3082 ;
  assign w3084 = ~w3026 & w3083 ;
  assign w3085 = w3081 | w3084 ;
  assign w3086 = ~\pi077 & w3085 ;
  assign w3087 = w2870 & w3026 ;
  assign w3088 = ~w2877 & w2983 ;
  assign w3089 = w2984 ^ w3088 ;
  assign w3090 = ~w3026 & w3089 ;
  assign w3091 = w3087 | w3090 ;
  assign w3092 = ~\pi076 & w3091 ;
  assign w3093 = w2876 & w3026 ;
  assign w3094 = ~w2883 & w2980 ;
  assign w3095 = w2981 ^ w3094 ;
  assign w3096 = ~w3026 & w3095 ;
  assign w3097 = w3093 | w3096 ;
  assign w3098 = ~\pi075 & w3097 ;
  assign w3099 = w2882 & w3026 ;
  assign w3100 = ~w2889 & w2977 ;
  assign w3101 = w2978 ^ w3100 ;
  assign w3102 = ~w3026 & w3101 ;
  assign w3103 = w3099 | w3102 ;
  assign w3104 = ~\pi074 & w3103 ;
  assign w3105 = w2888 & w3026 ;
  assign w3106 = ~w2895 & w2974 ;
  assign w3107 = w2975 ^ w3106 ;
  assign w3108 = ~w3026 & w3107 ;
  assign w3109 = w3105 | w3108 ;
  assign w3110 = ~\pi073 & w3109 ;
  assign w3111 = w2894 & w3026 ;
  assign w3112 = ~w2901 & w2971 ;
  assign w3113 = w2972 ^ w3112 ;
  assign w3114 = ~w3026 & w3113 ;
  assign w3115 = w3111 | w3114 ;
  assign w3116 = ~\pi072 & w3115 ;
  assign w3117 = w2900 & w3026 ;
  assign w3118 = ~w2907 & w2968 ;
  assign w3119 = w2969 ^ w3118 ;
  assign w3120 = ~w3026 & w3119 ;
  assign w3121 = w3117 | w3120 ;
  assign w3122 = ~\pi071 & w3121 ;
  assign w3123 = w2906 & w3026 ;
  assign w3124 = ~w2913 & w2965 ;
  assign w3125 = w2966 ^ w3124 ;
  assign w3126 = ~w3026 & w3125 ;
  assign w3127 = w3123 | w3126 ;
  assign w3128 = ~\pi070 & w3127 ;
  assign w3129 = w2912 & w3026 ;
  assign w3130 = ~w2921 & w2962 ;
  assign w3131 = w2963 ^ w3130 ;
  assign w3132 = ~w3026 & w3131 ;
  assign w3133 = w3129 | w3132 ;
  assign w3134 = ~\pi069 & w3133 ;
  assign w3135 = w2920 & w3026 ;
  assign w3136 = ~w2932 & w2959 ;
  assign w3137 = w2960 ^ w3136 ;
  assign w3138 = ~w3026 & w3137 ;
  assign w3139 = w3135 | w3138 ;
  assign w3140 = ~\pi068 & w3139 ;
  assign w3141 = w2931 & w3026 ;
  assign w3142 = w2953 & ~w2954 ;
  assign w3143 = w2957 ^ w3142 ;
  assign w3144 = ~w3026 & w3143 ;
  assign w3145 = w3141 | w3144 ;
  assign w3146 = ~\pi067 & w3145 ;
  assign w3147 = w2951 ^ w2952 ;
  assign w3148 = ~w3025 & w3147 ;
  assign w3149 = ( w2950 & w3021 ) | ( w2950 & w3025 ) | ( w3021 & w3025 ) ;
  assign w3150 = w2950 & w3149 ;
  assign w3151 = w3021 | w3148 ;
  assign w3152 = ( ~w3021 & w3150 ) | ( ~w3021 & w3151 ) | ( w3150 & w3151 ) ;
  assign w3153 = ~\pi066 & w3152 ;
  assign w3154 = ( \pi064 & w173 ) | ( \pi064 & w183 ) | ( w173 & w183 ) ;
  assign w3155 = ( \pi064 & ~\pi087 ) | ( \pi064 & w155 ) | ( ~\pi087 & w155 ) ;
  assign w3156 = ~w368 & w3155 ;
  assign w3157 = ~w3154 & w3156 ;
  assign w3158 = ( \pi041 & w3021 ) | ( \pi041 & ~w3157 ) | ( w3021 & ~w3157 ) ;
  assign w3159 = \pi041 & w3158 ;
  assign w3160 = \pi087 | \pi088 ;
  assign w3161 = w243 | w3160 ;
  assign w3162 = ( w243 & ~w441 ) | ( w243 & w2951 ) | ( ~w441 & w2951 ) ;
  assign w3163 = ~w3161 & w3162 ;
  assign w3164 = ( ~w448 & w451 ) | ( ~w448 & w3163 ) | ( w451 & w3163 ) ;
  assign w3165 = ~w451 & w3164 ;
  assign w3166 = ~w3021 & w3165 ;
  assign w3167 = w3159 | w3166 ;
  assign w3168 = ~\pi040 & \pi064 ;
  assign w3169 = ( w3159 & w3166 ) | ( w3159 & ~w3168 ) | ( w3166 & ~w3168 ) ;
  assign w3170 = \pi065 ^ w3169 ;
  assign w3171 = w3168 | w3170 ;
  assign w3172 = ~\pi065 & w3167 ;
  assign w3173 = ~w3021 & w3148 ;
  assign w3174 = ( ~w3021 & w3025 ) | ( ~w3021 & w3173 ) | ( w3025 & w3173 ) ;
  assign w3175 = w2950 | w3173 ;
  assign w3176 = ( w3021 & w3174 ) | ( w3021 & w3175 ) | ( w3174 & w3175 ) ;
  assign w3177 = \pi066 ^ w3176 ;
  assign w3178 = ( w3171 & ~w3172 ) | ( w3171 & w3177 ) | ( ~w3172 & w3177 ) ;
  assign w3179 = w3177 | w3178 ;
  assign w3180 = \pi067 ^ w3145 ;
  assign w3181 = ( ~w3153 & w3179 ) | ( ~w3153 & w3180 ) | ( w3179 & w3180 ) ;
  assign w3182 = w3180 | w3181 ;
  assign w3183 = \pi068 ^ w3139 ;
  assign w3184 = ( ~w3146 & w3182 ) | ( ~w3146 & w3183 ) | ( w3182 & w3183 ) ;
  assign w3185 = w3183 | w3184 ;
  assign w3186 = \pi069 ^ w3133 ;
  assign w3187 = ( ~w3140 & w3185 ) | ( ~w3140 & w3186 ) | ( w3185 & w3186 ) ;
  assign w3188 = w3186 | w3187 ;
  assign w3189 = \pi070 ^ w3127 ;
  assign w3190 = ( ~w3134 & w3188 ) | ( ~w3134 & w3189 ) | ( w3188 & w3189 ) ;
  assign w3191 = w3189 | w3190 ;
  assign w3192 = \pi071 ^ w3121 ;
  assign w3193 = ( ~w3128 & w3191 ) | ( ~w3128 & w3192 ) | ( w3191 & w3192 ) ;
  assign w3194 = w3192 | w3193 ;
  assign w3195 = \pi072 ^ w3115 ;
  assign w3196 = ( ~w3122 & w3194 ) | ( ~w3122 & w3195 ) | ( w3194 & w3195 ) ;
  assign w3197 = w3195 | w3196 ;
  assign w3198 = \pi073 ^ w3109 ;
  assign w3199 = ( ~w3116 & w3197 ) | ( ~w3116 & w3198 ) | ( w3197 & w3198 ) ;
  assign w3200 = w3198 | w3199 ;
  assign w3201 = \pi074 ^ w3103 ;
  assign w3202 = ( ~w3110 & w3200 ) | ( ~w3110 & w3201 ) | ( w3200 & w3201 ) ;
  assign w3203 = w3201 | w3202 ;
  assign w3204 = \pi075 ^ w3097 ;
  assign w3205 = ( ~w3104 & w3203 ) | ( ~w3104 & w3204 ) | ( w3203 & w3204 ) ;
  assign w3206 = w3204 | w3205 ;
  assign w3207 = \pi076 ^ w3091 ;
  assign w3208 = ( ~w3098 & w3206 ) | ( ~w3098 & w3207 ) | ( w3206 & w3207 ) ;
  assign w3209 = w3207 | w3208 ;
  assign w3210 = \pi077 ^ w3085 ;
  assign w3211 = ( ~w3092 & w3209 ) | ( ~w3092 & w3210 ) | ( w3209 & w3210 ) ;
  assign w3212 = w3210 | w3211 ;
  assign w3213 = \pi078 ^ w3079 ;
  assign w3214 = ( ~w3086 & w3212 ) | ( ~w3086 & w3213 ) | ( w3212 & w3213 ) ;
  assign w3215 = w3213 | w3214 ;
  assign w3216 = \pi079 ^ w3073 ;
  assign w3217 = ( ~w3080 & w3215 ) | ( ~w3080 & w3216 ) | ( w3215 & w3216 ) ;
  assign w3218 = w3216 | w3217 ;
  assign w3219 = \pi080 ^ w3067 ;
  assign w3220 = ( ~w3074 & w3218 ) | ( ~w3074 & w3219 ) | ( w3218 & w3219 ) ;
  assign w3221 = w3219 | w3220 ;
  assign w3222 = \pi081 ^ w3061 ;
  assign w3223 = ( ~w3068 & w3221 ) | ( ~w3068 & w3222 ) | ( w3221 & w3222 ) ;
  assign w3224 = w3222 | w3223 ;
  assign w3225 = \pi082 ^ w3055 ;
  assign w3226 = ( ~w3062 & w3224 ) | ( ~w3062 & w3225 ) | ( w3224 & w3225 ) ;
  assign w3227 = w3225 | w3226 ;
  assign w3228 = \pi083 ^ w3049 ;
  assign w3229 = ( ~w3056 & w3227 ) | ( ~w3056 & w3228 ) | ( w3227 & w3228 ) ;
  assign w3230 = w3228 | w3229 ;
  assign w3231 = \pi084 ^ w3043 ;
  assign w3232 = ( ~w3050 & w3230 ) | ( ~w3050 & w3231 ) | ( w3230 & w3231 ) ;
  assign w3233 = w3231 | w3232 ;
  assign w3234 = \pi085 ^ w3037 ;
  assign w3235 = ( ~w3044 & w3233 ) | ( ~w3044 & w3234 ) | ( w3233 & w3234 ) ;
  assign w3236 = w3234 | w3235 ;
  assign w3237 = \pi086 ^ w3031 ;
  assign w3238 = ( ~w3038 & w3236 ) | ( ~w3038 & w3237 ) | ( w3236 & w3237 ) ;
  assign w3239 = w3237 | w3238 ;
  assign w3240 = w2810 & w3026 ;
  assign w3241 = ~w2811 & w3016 ;
  assign w3242 = w3017 ^ w3241 ;
  assign w3243 = ~w3026 & w3242 ;
  assign w3244 = w3240 | w3243 ;
  assign w3245 = ~\pi087 & w3244 ;
  assign w3246 = ( \pi087 & ~w3240 ) | ( \pi087 & w3243 ) | ( ~w3240 & w3243 ) ;
  assign w3247 = ~w3243 & w3246 ;
  assign w3248 = w204 | w205 ;
  assign w3249 = w3247 | w3248 ;
  assign w3250 = ( w201 & w3245 ) | ( w201 & ~w3247 ) | ( w3245 & ~w3247 ) ;
  assign w3251 = w3249 | w3250 ;
  assign w3252 = ( ~w3032 & w3239 ) | ( ~w3032 & w3251 ) | ( w3239 & w3251 ) ;
  assign w3253 = w3251 | w3252 ;
  assign w3254 = ~w3025 & w3244 ;
  assign w3255 = w3253 & ~w3254 ;
  assign w3256 = ~w3038 & w3236 ;
  assign w3257 = w3237 ^ w3256 ;
  assign w3258 = ~w3255 & w3257 ;
  assign w3259 = ( w3031 & w3253 ) | ( w3031 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3260 = ~w3254 & w3259 ;
  assign w3261 = w3258 | w3260 ;
  assign w3262 = w3245 | w3247 ;
  assign w3263 = ( ~w3032 & w3239 ) | ( ~w3032 & w3255 ) | ( w3239 & w3255 ) ;
  assign w3264 = w3262 ^ w3263 ;
  assign w3265 = ~w3255 & w3264 ;
  assign w3266 = ( w3025 & ~w3244 ) | ( w3025 & w3253 ) | ( ~w3244 & w3253 ) ;
  assign w3267 = w3244 & w3266 ;
  assign w3268 = w3265 | w3267 ;
  assign w3269 = ~\pi087 & w3261 ;
  assign w3270 = ~w3044 & w3233 ;
  assign w3271 = w3234 ^ w3270 ;
  assign w3272 = ~w3255 & w3271 ;
  assign w3273 = ( w3037 & w3253 ) | ( w3037 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3274 = ~w3254 & w3273 ;
  assign w3275 = w3272 | w3274 ;
  assign w3276 = ~\pi086 & w3275 ;
  assign w3277 = ~w3050 & w3230 ;
  assign w3278 = w3231 ^ w3277 ;
  assign w3279 = ~w3255 & w3278 ;
  assign w3280 = ( w3043 & w3253 ) | ( w3043 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3281 = ~w3254 & w3280 ;
  assign w3282 = w3279 | w3281 ;
  assign w3283 = ~\pi085 & w3282 ;
  assign w3284 = ~w3056 & w3227 ;
  assign w3285 = w3228 ^ w3284 ;
  assign w3286 = ~w3255 & w3285 ;
  assign w3287 = ( w3049 & w3253 ) | ( w3049 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3288 = ~w3254 & w3287 ;
  assign w3289 = w3286 | w3288 ;
  assign w3290 = ~\pi084 & w3289 ;
  assign w3291 = ~w3062 & w3224 ;
  assign w3292 = w3225 ^ w3291 ;
  assign w3293 = ~w3255 & w3292 ;
  assign w3294 = ( w3055 & w3253 ) | ( w3055 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3295 = ~w3254 & w3294 ;
  assign w3296 = w3293 | w3295 ;
  assign w3297 = ~\pi083 & w3296 ;
  assign w3298 = ~w3068 & w3221 ;
  assign w3299 = w3222 ^ w3298 ;
  assign w3300 = ~w3255 & w3299 ;
  assign w3301 = ( w3061 & w3253 ) | ( w3061 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3302 = ~w3254 & w3301 ;
  assign w3303 = w3300 | w3302 ;
  assign w3304 = ~\pi082 & w3303 ;
  assign w3305 = ~w3074 & w3218 ;
  assign w3306 = w3219 ^ w3305 ;
  assign w3307 = ~w3255 & w3306 ;
  assign w3308 = ( w3067 & w3253 ) | ( w3067 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3309 = ~w3254 & w3308 ;
  assign w3310 = w3307 | w3309 ;
  assign w3311 = ~\pi081 & w3310 ;
  assign w3312 = ~w3080 & w3215 ;
  assign w3313 = w3216 ^ w3312 ;
  assign w3314 = ~w3255 & w3313 ;
  assign w3315 = ( w3073 & w3253 ) | ( w3073 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3316 = ~w3254 & w3315 ;
  assign w3317 = w3314 | w3316 ;
  assign w3318 = ~\pi080 & w3317 ;
  assign w3319 = ~w3086 & w3212 ;
  assign w3320 = w3213 ^ w3319 ;
  assign w3321 = ~w3255 & w3320 ;
  assign w3322 = ( w3079 & w3253 ) | ( w3079 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3323 = ~w3254 & w3322 ;
  assign w3324 = w3321 | w3323 ;
  assign w3325 = ~\pi079 & w3324 ;
  assign w3326 = ~w3092 & w3209 ;
  assign w3327 = w3210 ^ w3326 ;
  assign w3328 = ~w3255 & w3327 ;
  assign w3329 = ( w3085 & w3253 ) | ( w3085 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3330 = ~w3254 & w3329 ;
  assign w3331 = w3328 | w3330 ;
  assign w3332 = ~\pi078 & w3331 ;
  assign w3333 = ~w3098 & w3206 ;
  assign w3334 = w3207 ^ w3333 ;
  assign w3335 = ~w3255 & w3334 ;
  assign w3336 = ( w3091 & w3253 ) | ( w3091 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3337 = ~w3254 & w3336 ;
  assign w3338 = w3335 | w3337 ;
  assign w3339 = ~\pi077 & w3338 ;
  assign w3340 = ~w3104 & w3203 ;
  assign w3341 = w3204 ^ w3340 ;
  assign w3342 = ~w3255 & w3341 ;
  assign w3343 = ( w3097 & w3253 ) | ( w3097 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3344 = ~w3254 & w3343 ;
  assign w3345 = w3342 | w3344 ;
  assign w3346 = ~\pi076 & w3345 ;
  assign w3347 = ~w3110 & w3200 ;
  assign w3348 = w3201 ^ w3347 ;
  assign w3349 = ~w3255 & w3348 ;
  assign w3350 = ( w3103 & w3253 ) | ( w3103 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3351 = ~w3254 & w3350 ;
  assign w3352 = w3349 | w3351 ;
  assign w3353 = ~\pi075 & w3352 ;
  assign w3354 = ~w3116 & w3197 ;
  assign w3355 = w3198 ^ w3354 ;
  assign w3356 = ~w3255 & w3355 ;
  assign w3357 = ( w3109 & w3253 ) | ( w3109 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3358 = ~w3254 & w3357 ;
  assign w3359 = w3356 | w3358 ;
  assign w3360 = ~\pi074 & w3359 ;
  assign w3361 = ~w3122 & w3194 ;
  assign w3362 = w3195 ^ w3361 ;
  assign w3363 = ~w3255 & w3362 ;
  assign w3364 = ( w3115 & w3253 ) | ( w3115 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3365 = ~w3254 & w3364 ;
  assign w3366 = w3363 | w3365 ;
  assign w3367 = ~\pi073 & w3366 ;
  assign w3368 = ~w3128 & w3191 ;
  assign w3369 = w3192 ^ w3368 ;
  assign w3370 = ~w3255 & w3369 ;
  assign w3371 = ( w3121 & w3253 ) | ( w3121 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3372 = ~w3254 & w3371 ;
  assign w3373 = w3370 | w3372 ;
  assign w3374 = ~\pi072 & w3373 ;
  assign w3375 = ~w3134 & w3188 ;
  assign w3376 = w3189 ^ w3375 ;
  assign w3377 = ~w3255 & w3376 ;
  assign w3378 = ( w3127 & w3253 ) | ( w3127 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3379 = ~w3254 & w3378 ;
  assign w3380 = w3377 | w3379 ;
  assign w3381 = ~\pi071 & w3380 ;
  assign w3382 = ~w3140 & w3185 ;
  assign w3383 = w3186 ^ w3382 ;
  assign w3384 = ~w3255 & w3383 ;
  assign w3385 = ( w3133 & w3253 ) | ( w3133 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3386 = ~w3254 & w3385 ;
  assign w3387 = w3384 | w3386 ;
  assign w3388 = ~\pi070 & w3387 ;
  assign w3389 = ~w3146 & w3182 ;
  assign w3390 = w3183 ^ w3389 ;
  assign w3391 = ~w3255 & w3390 ;
  assign w3392 = ( w3139 & w3253 ) | ( w3139 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3393 = ~w3254 & w3392 ;
  assign w3394 = w3391 | w3393 ;
  assign w3395 = ~\pi069 & w3394 ;
  assign w3396 = ~w3153 & w3179 ;
  assign w3397 = w3180 ^ w3396 ;
  assign w3398 = ~w3255 & w3397 ;
  assign w3399 = ( w3145 & w3253 ) | ( w3145 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3400 = ~w3254 & w3399 ;
  assign w3401 = w3398 | w3400 ;
  assign w3402 = ~\pi068 & w3401 ;
  assign w3403 = w3171 & ~w3172 ;
  assign w3404 = w3177 ^ w3403 ;
  assign w3405 = ~w3255 & w3404 ;
  assign w3406 = ( w3152 & w3253 ) | ( w3152 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3407 = ~w3254 & w3406 ;
  assign w3408 = w3405 | w3407 ;
  assign w3409 = ~\pi067 & w3408 ;
  assign w3410 = ( w3159 & w3166 ) | ( w3159 & ~w3255 ) | ( w3166 & ~w3255 ) ;
  assign w3411 = ( ~\pi040 & \pi064 ) | ( ~\pi040 & w3255 ) | ( \pi064 & w3255 ) ;
  assign w3412 = w3410 ^ w3411 ;
  assign w3413 = \pi065 ^ w3412 ;
  assign w3414 = ~w3255 & w3413 ;
  assign w3415 = ( w3167 & w3253 ) | ( w3167 & w3254 ) | ( w3253 & w3254 ) ;
  assign w3416 = ~w3254 & w3415 ;
  assign w3417 = w3414 | w3416 ;
  assign w3418 = ~\pi066 & w3417 ;
  assign w3419 = \pi066 ^ w3417 ;
  assign w3420 = \pi064 & ~w3255 ;
  assign w3421 = \pi040 ^ w3420 ;
  assign w3422 = ( ~\pi039 & \pi064 ) | ( ~\pi039 & w3419 ) | ( \pi064 & w3419 ) ;
  assign w3423 = ( \pi065 & ~w3421 ) | ( \pi065 & w3422 ) | ( ~w3421 & w3422 ) ;
  assign w3424 = w3419 | w3423 ;
  assign w3425 = \pi067 ^ w3408 ;
  assign w3426 = ( ~w3418 & w3424 ) | ( ~w3418 & w3425 ) | ( w3424 & w3425 ) ;
  assign w3427 = w3425 | w3426 ;
  assign w3428 = \pi068 ^ w3401 ;
  assign w3429 = ( ~w3409 & w3427 ) | ( ~w3409 & w3428 ) | ( w3427 & w3428 ) ;
  assign w3430 = w3428 | w3429 ;
  assign w3431 = \pi069 ^ w3394 ;
  assign w3432 = ( ~w3402 & w3430 ) | ( ~w3402 & w3431 ) | ( w3430 & w3431 ) ;
  assign w3433 = w3431 | w3432 ;
  assign w3434 = \pi070 ^ w3387 ;
  assign w3435 = ( ~w3395 & w3433 ) | ( ~w3395 & w3434 ) | ( w3433 & w3434 ) ;
  assign w3436 = w3434 | w3435 ;
  assign w3437 = \pi071 ^ w3380 ;
  assign w3438 = ( ~w3388 & w3436 ) | ( ~w3388 & w3437 ) | ( w3436 & w3437 ) ;
  assign w3439 = w3437 | w3438 ;
  assign w3440 = \pi072 ^ w3373 ;
  assign w3441 = ( ~w3381 & w3439 ) | ( ~w3381 & w3440 ) | ( w3439 & w3440 ) ;
  assign w3442 = w3440 | w3441 ;
  assign w3443 = \pi073 ^ w3366 ;
  assign w3444 = ( ~w3374 & w3442 ) | ( ~w3374 & w3443 ) | ( w3442 & w3443 ) ;
  assign w3445 = w3443 | w3444 ;
  assign w3446 = \pi074 ^ w3359 ;
  assign w3447 = ( ~w3367 & w3445 ) | ( ~w3367 & w3446 ) | ( w3445 & w3446 ) ;
  assign w3448 = w3446 | w3447 ;
  assign w3449 = \pi075 ^ w3352 ;
  assign w3450 = ( ~w3360 & w3448 ) | ( ~w3360 & w3449 ) | ( w3448 & w3449 ) ;
  assign w3451 = w3449 | w3450 ;
  assign w3452 = \pi076 ^ w3345 ;
  assign w3453 = ( ~w3353 & w3451 ) | ( ~w3353 & w3452 ) | ( w3451 & w3452 ) ;
  assign w3454 = w3452 | w3453 ;
  assign w3455 = \pi077 ^ w3338 ;
  assign w3456 = ( ~w3346 & w3454 ) | ( ~w3346 & w3455 ) | ( w3454 & w3455 ) ;
  assign w3457 = w3455 | w3456 ;
  assign w3458 = \pi078 ^ w3331 ;
  assign w3459 = ( ~w3339 & w3457 ) | ( ~w3339 & w3458 ) | ( w3457 & w3458 ) ;
  assign w3460 = w3458 | w3459 ;
  assign w3461 = \pi079 ^ w3324 ;
  assign w3462 = ( ~w3332 & w3460 ) | ( ~w3332 & w3461 ) | ( w3460 & w3461 ) ;
  assign w3463 = w3461 | w3462 ;
  assign w3464 = \pi080 ^ w3317 ;
  assign w3465 = ( ~w3325 & w3463 ) | ( ~w3325 & w3464 ) | ( w3463 & w3464 ) ;
  assign w3466 = w3464 | w3465 ;
  assign w3467 = \pi081 ^ w3310 ;
  assign w3468 = ( ~w3318 & w3466 ) | ( ~w3318 & w3467 ) | ( w3466 & w3467 ) ;
  assign w3469 = w3467 | w3468 ;
  assign w3470 = \pi082 ^ w3303 ;
  assign w3471 = ( ~w3311 & w3469 ) | ( ~w3311 & w3470 ) | ( w3469 & w3470 ) ;
  assign w3472 = w3470 | w3471 ;
  assign w3473 = \pi083 ^ w3296 ;
  assign w3474 = ( ~w3304 & w3472 ) | ( ~w3304 & w3473 ) | ( w3472 & w3473 ) ;
  assign w3475 = w3473 | w3474 ;
  assign w3476 = \pi084 ^ w3289 ;
  assign w3477 = ( ~w3297 & w3475 ) | ( ~w3297 & w3476 ) | ( w3475 & w3476 ) ;
  assign w3478 = w3476 | w3477 ;
  assign w3479 = \pi085 ^ w3282 ;
  assign w3480 = ( ~w3290 & w3478 ) | ( ~w3290 & w3479 ) | ( w3478 & w3479 ) ;
  assign w3481 = w3479 | w3480 ;
  assign w3482 = \pi086 ^ w3275 ;
  assign w3483 = ( ~w3283 & w3481 ) | ( ~w3283 & w3482 ) | ( w3481 & w3482 ) ;
  assign w3484 = w3482 | w3483 ;
  assign w3485 = \pi087 ^ w3261 ;
  assign w3486 = ( ~w3276 & w3484 ) | ( ~w3276 & w3485 ) | ( w3484 & w3485 ) ;
  assign w3487 = w3485 | w3486 ;
  assign w3488 = \pi088 ^ w3268 ;
  assign w3489 = w3269 & ~w3488 ;
  assign w3490 = ( w3487 & w3488 ) | ( w3487 & ~w3489 ) | ( w3488 & ~w3489 ) ;
  assign w3491 = ~\pi088 & w3268 ;
  assign w3492 = w3490 & ~w3491 ;
  assign w3493 = ( w244 & w275 ) | ( w244 & ~w290 ) | ( w275 & ~w290 ) ;
  assign w3494 = w290 | w3493 ;
  assign w3495 = w3492 | w3494 ;
  assign w3496 = w3261 & w3495 ;
  assign w3497 = ~w3276 & w3484 ;
  assign w3498 = w3485 ^ w3497 ;
  assign w3499 = ~w3495 & w3498 ;
  assign w3500 = w3496 | w3499 ;
  assign w3501 = w3268 & w3495 ;
  assign w3502 = ~w3269 & w3487 ;
  assign w3503 = w3488 ^ w3502 ;
  assign w3504 = ~w3495 & w3503 ;
  assign w3505 = w3501 | w3504 ;
  assign w3506 = ~\pi088 & w3500 ;
  assign w3507 = w3275 & w3495 ;
  assign w3508 = ~w3283 & w3481 ;
  assign w3509 = w3482 ^ w3508 ;
  assign w3510 = ~w3495 & w3509 ;
  assign w3511 = w3507 | w3510 ;
  assign w3512 = ~\pi087 & w3511 ;
  assign w3513 = w3282 & w3495 ;
  assign w3514 = ~w3290 & w3478 ;
  assign w3515 = w3479 ^ w3514 ;
  assign w3516 = ~w3495 & w3515 ;
  assign w3517 = w3513 | w3516 ;
  assign w3518 = ~\pi086 & w3517 ;
  assign w3519 = w3289 & w3495 ;
  assign w3520 = ~w3297 & w3475 ;
  assign w3521 = w3476 ^ w3520 ;
  assign w3522 = ~w3495 & w3521 ;
  assign w3523 = w3519 | w3522 ;
  assign w3524 = ~\pi085 & w3523 ;
  assign w3525 = w3296 & w3495 ;
  assign w3526 = ~w3304 & w3472 ;
  assign w3527 = w3473 ^ w3526 ;
  assign w3528 = ~w3495 & w3527 ;
  assign w3529 = w3525 | w3528 ;
  assign w3530 = ~\pi084 & w3529 ;
  assign w3531 = w3303 & w3495 ;
  assign w3532 = ~w3311 & w3469 ;
  assign w3533 = w3470 ^ w3532 ;
  assign w3534 = ~w3495 & w3533 ;
  assign w3535 = w3531 | w3534 ;
  assign w3536 = ~\pi083 & w3535 ;
  assign w3537 = w3310 & w3495 ;
  assign w3538 = ~w3318 & w3466 ;
  assign w3539 = w3467 ^ w3538 ;
  assign w3540 = ~w3495 & w3539 ;
  assign w3541 = w3537 | w3540 ;
  assign w3542 = ~\pi082 & w3541 ;
  assign w3543 = w3317 & w3495 ;
  assign w3544 = ~w3325 & w3463 ;
  assign w3545 = w3464 ^ w3544 ;
  assign w3546 = ~w3495 & w3545 ;
  assign w3547 = w3543 | w3546 ;
  assign w3548 = ~\pi081 & w3547 ;
  assign w3549 = w3324 & w3495 ;
  assign w3550 = ~w3332 & w3460 ;
  assign w3551 = w3461 ^ w3550 ;
  assign w3552 = ~w3495 & w3551 ;
  assign w3553 = w3549 | w3552 ;
  assign w3554 = ~\pi080 & w3553 ;
  assign w3555 = w3331 & w3495 ;
  assign w3556 = ~w3339 & w3457 ;
  assign w3557 = w3458 ^ w3556 ;
  assign w3558 = ~w3495 & w3557 ;
  assign w3559 = w3555 | w3558 ;
  assign w3560 = ~\pi079 & w3559 ;
  assign w3561 = w3338 & w3495 ;
  assign w3562 = ~w3346 & w3454 ;
  assign w3563 = w3455 ^ w3562 ;
  assign w3564 = ~w3495 & w3563 ;
  assign w3565 = w3561 | w3564 ;
  assign w3566 = ~\pi078 & w3565 ;
  assign w3567 = w3345 & w3495 ;
  assign w3568 = ~w3353 & w3451 ;
  assign w3569 = w3452 ^ w3568 ;
  assign w3570 = ~w3495 & w3569 ;
  assign w3571 = w3567 | w3570 ;
  assign w3572 = ~\pi077 & w3571 ;
  assign w3573 = w3352 & w3495 ;
  assign w3574 = ~w3360 & w3448 ;
  assign w3575 = w3449 ^ w3574 ;
  assign w3576 = ~w3495 & w3575 ;
  assign w3577 = w3573 | w3576 ;
  assign w3578 = ~\pi076 & w3577 ;
  assign w3579 = w3359 & w3495 ;
  assign w3580 = ~w3367 & w3445 ;
  assign w3581 = w3446 ^ w3580 ;
  assign w3582 = ~w3495 & w3581 ;
  assign w3583 = w3579 | w3582 ;
  assign w3584 = ~\pi075 & w3583 ;
  assign w3585 = w3366 & w3495 ;
  assign w3586 = ~w3374 & w3442 ;
  assign w3587 = w3443 ^ w3586 ;
  assign w3588 = ~w3495 & w3587 ;
  assign w3589 = w3585 | w3588 ;
  assign w3590 = ~\pi074 & w3589 ;
  assign w3591 = w3373 & w3495 ;
  assign w3592 = ~w3381 & w3439 ;
  assign w3593 = w3440 ^ w3592 ;
  assign w3594 = ~w3495 & w3593 ;
  assign w3595 = w3591 | w3594 ;
  assign w3596 = ~\pi073 & w3595 ;
  assign w3597 = w3380 & w3495 ;
  assign w3598 = ~w3388 & w3436 ;
  assign w3599 = w3437 ^ w3598 ;
  assign w3600 = ~w3495 & w3599 ;
  assign w3601 = w3597 | w3600 ;
  assign w3602 = ~\pi072 & w3601 ;
  assign w3603 = w3387 & w3495 ;
  assign w3604 = ~w3395 & w3433 ;
  assign w3605 = w3434 ^ w3604 ;
  assign w3606 = ~w3495 & w3605 ;
  assign w3607 = w3603 | w3606 ;
  assign w3608 = ~\pi071 & w3607 ;
  assign w3609 = w3394 & w3495 ;
  assign w3610 = ~w3402 & w3430 ;
  assign w3611 = w3431 ^ w3610 ;
  assign w3612 = ~w3495 & w3611 ;
  assign w3613 = w3609 | w3612 ;
  assign w3614 = ~\pi070 & w3613 ;
  assign w3615 = w3401 & w3495 ;
  assign w3616 = ~w3409 & w3427 ;
  assign w3617 = w3428 ^ w3616 ;
  assign w3618 = ~w3495 & w3617 ;
  assign w3619 = w3615 | w3618 ;
  assign w3620 = ~\pi069 & w3619 ;
  assign w3621 = w3408 & w3495 ;
  assign w3622 = ~w3418 & w3424 ;
  assign w3623 = w3425 ^ w3622 ;
  assign w3624 = ~w3495 & w3623 ;
  assign w3625 = w3621 | w3624 ;
  assign w3626 = ~\pi068 & w3625 ;
  assign w3627 = w3417 & w3495 ;
  assign w3628 = ~\pi039 & \pi064 ;
  assign w3629 = ( \pi065 & ~w3421 ) | ( \pi065 & w3628 ) | ( ~w3421 & w3628 ) ;
  assign w3630 = w3419 ^ w3629 ;
  assign w3631 = ( w3492 & w3494 ) | ( w3492 & w3630 ) | ( w3494 & w3630 ) ;
  assign w3632 = w3630 & ~w3631 ;
  assign w3633 = w3627 | w3632 ;
  assign w3634 = ~\pi067 & w3633 ;
  assign w3635 = \pi040 ^ \pi065 ;
  assign w3636 = \pi039 ^ w3255 ;
  assign w3637 = ( \pi064 & w3494 ) | ( \pi064 & w3636 ) | ( w3494 & w3636 ) ;
  assign w3638 = w3635 ^ w3637 ;
  assign w3639 = ~w3494 & w3638 ;
  assign w3640 = ~w3492 & w3639 ;
  assign w3641 = ( ~\pi064 & w3255 ) | ( ~\pi064 & w3495 ) | ( w3255 & w3495 ) ;
  assign w3642 = \pi040 ^ w3641 ;
  assign w3643 = w3495 & ~w3642 ;
  assign w3644 = w3640 | w3643 ;
  assign w3645 = ~\pi066 & w3644 ;
  assign w3646 = ( \pi064 & ~\pi089 ) | ( \pi064 & \pi090 ) | ( ~\pi089 & \pi090 ) ;
  assign w3647 = w182 | w204 ;
  assign w3648 = ( \pi090 & \pi091 ) | ( \pi090 & ~w182 ) | ( \pi091 & ~w182 ) ;
  assign w3649 = w3647 | w3648 ;
  assign w3650 = w3646 & ~w3649 ;
  assign w3651 = ~w201 & w3650 ;
  assign w3652 = ( \pi039 & w3492 ) | ( \pi039 & ~w3651 ) | ( w3492 & ~w3651 ) ;
  assign w3653 = \pi039 & w3652 ;
  assign w3654 = ( ~\pi039 & w243 ) | ( ~\pi039 & w441 ) | ( w243 & w441 ) ;
  assign w3655 = ( ~\pi039 & \pi064 ) | ( ~\pi039 & w451 ) | ( \pi064 & w451 ) ;
  assign w3656 = ~w452 & w3655 ;
  assign w3657 = ~w3654 & w3656 ;
  assign w3658 = ~w3492 & w3657 ;
  assign w3659 = w3653 | w3658 ;
  assign w3660 = ~\pi038 & \pi064 ;
  assign w3661 = \pi065 ^ w3659 ;
  assign w3662 = w3660 | w3661 ;
  assign w3663 = w3495 | w3640 ;
  assign w3664 = ( w3421 & w3640 ) | ( w3421 & w3663 ) | ( w3640 & w3663 ) ;
  assign w3665 = \pi066 ^ w3664 ;
  assign w3666 = ~\pi065 & w3659 ;
  assign w3667 = w3662 | w3666 ;
  assign w3668 = ( w3665 & ~w3666 ) | ( w3665 & w3667 ) | ( ~w3666 & w3667 ) ;
  assign w3669 = \pi067 ^ w3633 ;
  assign w3670 = ( ~w3645 & w3668 ) | ( ~w3645 & w3669 ) | ( w3668 & w3669 ) ;
  assign w3671 = w3669 | w3670 ;
  assign w3672 = \pi068 ^ w3625 ;
  assign w3673 = ( ~w3634 & w3671 ) | ( ~w3634 & w3672 ) | ( w3671 & w3672 ) ;
  assign w3674 = w3672 | w3673 ;
  assign w3675 = \pi069 ^ w3619 ;
  assign w3676 = ( ~w3626 & w3674 ) | ( ~w3626 & w3675 ) | ( w3674 & w3675 ) ;
  assign w3677 = w3675 | w3676 ;
  assign w3678 = \pi070 ^ w3613 ;
  assign w3679 = ( ~w3620 & w3677 ) | ( ~w3620 & w3678 ) | ( w3677 & w3678 ) ;
  assign w3680 = w3678 | w3679 ;
  assign w3681 = \pi071 ^ w3607 ;
  assign w3682 = ( ~w3614 & w3680 ) | ( ~w3614 & w3681 ) | ( w3680 & w3681 ) ;
  assign w3683 = w3681 | w3682 ;
  assign w3684 = \pi072 ^ w3601 ;
  assign w3685 = ( ~w3608 & w3683 ) | ( ~w3608 & w3684 ) | ( w3683 & w3684 ) ;
  assign w3686 = w3684 | w3685 ;
  assign w3687 = \pi073 ^ w3595 ;
  assign w3688 = ( ~w3602 & w3686 ) | ( ~w3602 & w3687 ) | ( w3686 & w3687 ) ;
  assign w3689 = w3687 | w3688 ;
  assign w3690 = \pi074 ^ w3589 ;
  assign w3691 = ( ~w3596 & w3689 ) | ( ~w3596 & w3690 ) | ( w3689 & w3690 ) ;
  assign w3692 = w3690 | w3691 ;
  assign w3693 = \pi075 ^ w3583 ;
  assign w3694 = ( ~w3590 & w3692 ) | ( ~w3590 & w3693 ) | ( w3692 & w3693 ) ;
  assign w3695 = w3693 | w3694 ;
  assign w3696 = \pi076 ^ w3577 ;
  assign w3697 = ( ~w3584 & w3695 ) | ( ~w3584 & w3696 ) | ( w3695 & w3696 ) ;
  assign w3698 = w3696 | w3697 ;
  assign w3699 = \pi077 ^ w3571 ;
  assign w3700 = ( ~w3578 & w3698 ) | ( ~w3578 & w3699 ) | ( w3698 & w3699 ) ;
  assign w3701 = w3699 | w3700 ;
  assign w3702 = \pi078 ^ w3565 ;
  assign w3703 = ( ~w3572 & w3701 ) | ( ~w3572 & w3702 ) | ( w3701 & w3702 ) ;
  assign w3704 = w3702 | w3703 ;
  assign w3705 = \pi079 ^ w3559 ;
  assign w3706 = ( ~w3566 & w3704 ) | ( ~w3566 & w3705 ) | ( w3704 & w3705 ) ;
  assign w3707 = w3705 | w3706 ;
  assign w3708 = \pi080 ^ w3553 ;
  assign w3709 = ( ~w3560 & w3707 ) | ( ~w3560 & w3708 ) | ( w3707 & w3708 ) ;
  assign w3710 = w3708 | w3709 ;
  assign w3711 = \pi081 ^ w3547 ;
  assign w3712 = ( ~w3554 & w3710 ) | ( ~w3554 & w3711 ) | ( w3710 & w3711 ) ;
  assign w3713 = w3711 | w3712 ;
  assign w3714 = \pi082 ^ w3541 ;
  assign w3715 = ( ~w3548 & w3713 ) | ( ~w3548 & w3714 ) | ( w3713 & w3714 ) ;
  assign w3716 = w3714 | w3715 ;
  assign w3717 = \pi083 ^ w3535 ;
  assign w3718 = ( ~w3542 & w3716 ) | ( ~w3542 & w3717 ) | ( w3716 & w3717 ) ;
  assign w3719 = w3717 | w3718 ;
  assign w3720 = \pi084 ^ w3529 ;
  assign w3721 = ( ~w3536 & w3719 ) | ( ~w3536 & w3720 ) | ( w3719 & w3720 ) ;
  assign w3722 = w3720 | w3721 ;
  assign w3723 = \pi085 ^ w3523 ;
  assign w3724 = ( ~w3530 & w3722 ) | ( ~w3530 & w3723 ) | ( w3722 & w3723 ) ;
  assign w3725 = w3723 | w3724 ;
  assign w3726 = \pi086 ^ w3517 ;
  assign w3727 = ( ~w3524 & w3725 ) | ( ~w3524 & w3726 ) | ( w3725 & w3726 ) ;
  assign w3728 = w3726 | w3727 ;
  assign w3729 = \pi087 ^ w3511 ;
  assign w3730 = ( ~w3518 & w3728 ) | ( ~w3518 & w3729 ) | ( w3728 & w3729 ) ;
  assign w3731 = w3729 | w3730 ;
  assign w3732 = \pi088 ^ w3500 ;
  assign w3733 = ( ~w3512 & w3731 ) | ( ~w3512 & w3732 ) | ( w3731 & w3732 ) ;
  assign w3734 = w3732 | w3733 ;
  assign w3735 = \pi089 ^ w3505 ;
  assign w3736 = w3506 & ~w3735 ;
  assign w3737 = ( w3734 & w3735 ) | ( w3734 & ~w3736 ) | ( w3735 & ~w3736 ) ;
  assign w3738 = ~\pi089 & w3505 ;
  assign w3739 = w3737 & ~w3738 ;
  assign w3740 = \pi090 | \pi091 ;
  assign w3741 = w204 | w3740 ;
  assign w3742 = ( w182 & w201 ) | ( w182 & ~w204 ) | ( w201 & ~w204 ) ;
  assign w3743 = w3741 | w3742 ;
  assign w3744 = w3739 | w3743 ;
  assign w3745 = w3500 & w3744 ;
  assign w3746 = ~w3512 & w3731 ;
  assign w3747 = w3732 ^ w3746 ;
  assign w3748 = ~w3744 & w3747 ;
  assign w3749 = w3745 | w3748 ;
  assign w3750 = ~\pi089 & w3749 ;
  assign w3751 = w3511 & w3744 ;
  assign w3752 = ~w3518 & w3728 ;
  assign w3753 = w3729 ^ w3752 ;
  assign w3754 = ~w3744 & w3753 ;
  assign w3755 = w3751 | w3754 ;
  assign w3756 = ~\pi088 & w3755 ;
  assign w3757 = w3517 & w3744 ;
  assign w3758 = ~w3524 & w3725 ;
  assign w3759 = w3726 ^ w3758 ;
  assign w3760 = ~w3744 & w3759 ;
  assign w3761 = w3757 | w3760 ;
  assign w3762 = ~\pi087 & w3761 ;
  assign w3763 = w3523 & w3744 ;
  assign w3764 = ~w3530 & w3722 ;
  assign w3765 = w3723 ^ w3764 ;
  assign w3766 = ~w3744 & w3765 ;
  assign w3767 = w3763 | w3766 ;
  assign w3768 = ~\pi086 & w3767 ;
  assign w3769 = w3529 & w3744 ;
  assign w3770 = ~w3536 & w3719 ;
  assign w3771 = w3720 ^ w3770 ;
  assign w3772 = ~w3744 & w3771 ;
  assign w3773 = w3769 | w3772 ;
  assign w3774 = ~\pi085 & w3773 ;
  assign w3775 = w3535 & w3744 ;
  assign w3776 = ~w3542 & w3716 ;
  assign w3777 = w3717 ^ w3776 ;
  assign w3778 = ~w3744 & w3777 ;
  assign w3779 = w3775 | w3778 ;
  assign w3780 = ~\pi084 & w3779 ;
  assign w3781 = w3541 & w3744 ;
  assign w3782 = ~w3548 & w3713 ;
  assign w3783 = w3714 ^ w3782 ;
  assign w3784 = ~w3744 & w3783 ;
  assign w3785 = w3781 | w3784 ;
  assign w3786 = ~\pi083 & w3785 ;
  assign w3787 = w3547 & w3744 ;
  assign w3788 = ~w3554 & w3710 ;
  assign w3789 = w3711 ^ w3788 ;
  assign w3790 = ~w3744 & w3789 ;
  assign w3791 = w3787 | w3790 ;
  assign w3792 = ~\pi082 & w3791 ;
  assign w3793 = w3553 & w3744 ;
  assign w3794 = ~w3560 & w3707 ;
  assign w3795 = w3708 ^ w3794 ;
  assign w3796 = ~w3744 & w3795 ;
  assign w3797 = w3793 | w3796 ;
  assign w3798 = ~\pi081 & w3797 ;
  assign w3799 = w3559 & w3744 ;
  assign w3800 = ~w3566 & w3704 ;
  assign w3801 = w3705 ^ w3800 ;
  assign w3802 = ~w3744 & w3801 ;
  assign w3803 = w3799 | w3802 ;
  assign w3804 = ~\pi080 & w3803 ;
  assign w3805 = w3565 & w3744 ;
  assign w3806 = ~w3572 & w3701 ;
  assign w3807 = w3702 ^ w3806 ;
  assign w3808 = ~w3744 & w3807 ;
  assign w3809 = w3805 | w3808 ;
  assign w3810 = ~\pi079 & w3809 ;
  assign w3811 = w3571 & w3744 ;
  assign w3812 = ~w3578 & w3698 ;
  assign w3813 = w3699 ^ w3812 ;
  assign w3814 = ~w3744 & w3813 ;
  assign w3815 = w3811 | w3814 ;
  assign w3816 = ~\pi078 & w3815 ;
  assign w3817 = w3577 & w3744 ;
  assign w3818 = ~w3584 & w3695 ;
  assign w3819 = w3696 ^ w3818 ;
  assign w3820 = ~w3744 & w3819 ;
  assign w3821 = w3817 | w3820 ;
  assign w3822 = ~\pi077 & w3821 ;
  assign w3823 = w3583 & w3744 ;
  assign w3824 = ~w3590 & w3692 ;
  assign w3825 = w3693 ^ w3824 ;
  assign w3826 = ~w3744 & w3825 ;
  assign w3827 = w3823 | w3826 ;
  assign w3828 = ~\pi076 & w3827 ;
  assign w3829 = w3589 & w3744 ;
  assign w3830 = ~w3596 & w3689 ;
  assign w3831 = w3690 ^ w3830 ;
  assign w3832 = ~w3744 & w3831 ;
  assign w3833 = w3829 | w3832 ;
  assign w3834 = ~\pi075 & w3833 ;
  assign w3835 = w3595 & w3744 ;
  assign w3836 = ~w3602 & w3686 ;
  assign w3837 = w3687 ^ w3836 ;
  assign w3838 = ~w3744 & w3837 ;
  assign w3839 = w3835 | w3838 ;
  assign w3840 = ~\pi074 & w3839 ;
  assign w3841 = w3601 & w3744 ;
  assign w3842 = ~w3608 & w3683 ;
  assign w3843 = w3684 ^ w3842 ;
  assign w3844 = ~w3744 & w3843 ;
  assign w3845 = w3841 | w3844 ;
  assign w3846 = ~\pi073 & w3845 ;
  assign w3847 = w3607 & w3744 ;
  assign w3848 = ~w3614 & w3680 ;
  assign w3849 = w3681 ^ w3848 ;
  assign w3850 = ~w3744 & w3849 ;
  assign w3851 = w3847 | w3850 ;
  assign w3852 = ~\pi072 & w3851 ;
  assign w3853 = w3613 & w3744 ;
  assign w3854 = ~w3620 & w3677 ;
  assign w3855 = w3678 ^ w3854 ;
  assign w3856 = ~w3744 & w3855 ;
  assign w3857 = w3853 | w3856 ;
  assign w3858 = ~\pi071 & w3857 ;
  assign w3859 = w3619 & w3744 ;
  assign w3860 = ~w3626 & w3674 ;
  assign w3861 = w3675 ^ w3860 ;
  assign w3862 = ~w3744 & w3861 ;
  assign w3863 = w3859 | w3862 ;
  assign w3864 = ~\pi070 & w3863 ;
  assign w3865 = w3625 & w3744 ;
  assign w3866 = ~w3634 & w3671 ;
  assign w3867 = w3672 ^ w3866 ;
  assign w3868 = ~w3744 & w3867 ;
  assign w3869 = w3865 | w3868 ;
  assign w3870 = ~\pi069 & w3869 ;
  assign w3871 = w3633 & w3744 ;
  assign w3872 = ~w3645 & w3668 ;
  assign w3873 = w3669 ^ w3872 ;
  assign w3874 = ~w3744 & w3873 ;
  assign w3875 = w3871 | w3874 ;
  assign w3876 = ~\pi068 & w3875 ;
  assign w3877 = w3644 & w3744 ;
  assign w3878 = ~w3659 & w3662 ;
  assign w3879 = ( \pi065 & w3662 ) | ( \pi065 & w3878 ) | ( w3662 & w3878 ) ;
  assign w3880 = w3665 ^ w3879 ;
  assign w3881 = ~w3744 & w3880 ;
  assign w3882 = w3877 | w3881 ;
  assign w3883 = ~\pi067 & w3882 ;
  assign w3884 = w3659 & w3744 ;
  assign w3885 = ( w3653 & w3658 ) | ( w3653 & ~w3743 ) | ( w3658 & ~w3743 ) ;
  assign w3886 = \pi065 ^ w3885 ;
  assign w3887 = ( w3660 & ~w3743 ) | ( w3660 & w3886 ) | ( ~w3743 & w3886 ) ;
  assign w3888 = ( w3660 & w3739 ) | ( w3660 & w3886 ) | ( w3739 & w3886 ) ;
  assign w3889 = w3887 & ~w3888 ;
  assign w3890 = w3884 | w3889 ;
  assign w3891 = ~\pi066 & w3890 ;
  assign w3892 = ( \pi064 & ~\pi090 ) | ( \pi064 & \pi091 ) | ( ~\pi090 & \pi091 ) ;
  assign w3893 = w240 | w290 ;
  assign w3894 = ( \pi091 & \pi092 ) | ( \pi091 & ~w240 ) | ( \pi092 & ~w240 ) ;
  assign w3895 = w3893 | w3894 ;
  assign w3896 = w3892 & ~w3895 ;
  assign w3897 = ~w275 & w3896 ;
  assign w3898 = ( \pi038 & w3739 ) | ( \pi038 & ~w3897 ) | ( w3739 & ~w3897 ) ;
  assign w3899 = \pi038 & w3898 ;
  assign w3900 = ( \pi090 & ~w182 ) | ( \pi090 & w3660 ) | ( ~w182 & w3660 ) ;
  assign w3901 = ( \pi090 & \pi091 ) | ( \pi090 & ~w204 ) | ( \pi091 & ~w204 ) ;
  assign w3902 = w298 | w3901 ;
  assign w3903 = w3900 & ~w3902 ;
  assign w3904 = ~w3739 & w3903 ;
  assign w3905 = w3899 | w3904 ;
  assign w3906 = ~\pi037 & \pi064 ;
  assign w3907 = \pi065 ^ w3905 ;
  assign w3908 = w3906 | w3907 ;
  assign w3909 = \pi066 ^ w3890 ;
  assign w3910 = ~\pi065 & w3905 ;
  assign w3911 = w3908 | w3910 ;
  assign w3912 = ( w3909 & ~w3910 ) | ( w3909 & w3911 ) | ( ~w3910 & w3911 ) ;
  assign w3913 = \pi067 ^ w3882 ;
  assign w3914 = ( ~w3891 & w3912 ) | ( ~w3891 & w3913 ) | ( w3912 & w3913 ) ;
  assign w3915 = w3913 | w3914 ;
  assign w3916 = \pi068 ^ w3875 ;
  assign w3917 = ( ~w3883 & w3915 ) | ( ~w3883 & w3916 ) | ( w3915 & w3916 ) ;
  assign w3918 = w3916 | w3917 ;
  assign w3919 = \pi069 ^ w3869 ;
  assign w3920 = ( ~w3876 & w3918 ) | ( ~w3876 & w3919 ) | ( w3918 & w3919 ) ;
  assign w3921 = w3919 | w3920 ;
  assign w3922 = \pi070 ^ w3863 ;
  assign w3923 = ( ~w3870 & w3921 ) | ( ~w3870 & w3922 ) | ( w3921 & w3922 ) ;
  assign w3924 = w3922 | w3923 ;
  assign w3925 = \pi071 ^ w3857 ;
  assign w3926 = ( ~w3864 & w3924 ) | ( ~w3864 & w3925 ) | ( w3924 & w3925 ) ;
  assign w3927 = w3925 | w3926 ;
  assign w3928 = \pi072 ^ w3851 ;
  assign w3929 = ( ~w3858 & w3927 ) | ( ~w3858 & w3928 ) | ( w3927 & w3928 ) ;
  assign w3930 = w3928 | w3929 ;
  assign w3931 = \pi073 ^ w3845 ;
  assign w3932 = ( ~w3852 & w3930 ) | ( ~w3852 & w3931 ) | ( w3930 & w3931 ) ;
  assign w3933 = w3931 | w3932 ;
  assign w3934 = \pi074 ^ w3839 ;
  assign w3935 = ( ~w3846 & w3933 ) | ( ~w3846 & w3934 ) | ( w3933 & w3934 ) ;
  assign w3936 = w3934 | w3935 ;
  assign w3937 = \pi075 ^ w3833 ;
  assign w3938 = ( ~w3840 & w3936 ) | ( ~w3840 & w3937 ) | ( w3936 & w3937 ) ;
  assign w3939 = w3937 | w3938 ;
  assign w3940 = \pi076 ^ w3827 ;
  assign w3941 = ( ~w3834 & w3939 ) | ( ~w3834 & w3940 ) | ( w3939 & w3940 ) ;
  assign w3942 = w3940 | w3941 ;
  assign w3943 = \pi077 ^ w3821 ;
  assign w3944 = ( ~w3828 & w3942 ) | ( ~w3828 & w3943 ) | ( w3942 & w3943 ) ;
  assign w3945 = w3943 | w3944 ;
  assign w3946 = \pi078 ^ w3815 ;
  assign w3947 = ( ~w3822 & w3945 ) | ( ~w3822 & w3946 ) | ( w3945 & w3946 ) ;
  assign w3948 = w3946 | w3947 ;
  assign w3949 = \pi079 ^ w3809 ;
  assign w3950 = ( ~w3816 & w3948 ) | ( ~w3816 & w3949 ) | ( w3948 & w3949 ) ;
  assign w3951 = w3949 | w3950 ;
  assign w3952 = \pi080 ^ w3803 ;
  assign w3953 = ( ~w3810 & w3951 ) | ( ~w3810 & w3952 ) | ( w3951 & w3952 ) ;
  assign w3954 = w3952 | w3953 ;
  assign w3955 = \pi081 ^ w3797 ;
  assign w3956 = ( ~w3804 & w3954 ) | ( ~w3804 & w3955 ) | ( w3954 & w3955 ) ;
  assign w3957 = w3955 | w3956 ;
  assign w3958 = \pi082 ^ w3791 ;
  assign w3959 = ( ~w3798 & w3957 ) | ( ~w3798 & w3958 ) | ( w3957 & w3958 ) ;
  assign w3960 = w3958 | w3959 ;
  assign w3961 = \pi083 ^ w3785 ;
  assign w3962 = ( ~w3792 & w3960 ) | ( ~w3792 & w3961 ) | ( w3960 & w3961 ) ;
  assign w3963 = w3961 | w3962 ;
  assign w3964 = \pi084 ^ w3779 ;
  assign w3965 = ( ~w3786 & w3963 ) | ( ~w3786 & w3964 ) | ( w3963 & w3964 ) ;
  assign w3966 = w3964 | w3965 ;
  assign w3967 = \pi085 ^ w3773 ;
  assign w3968 = ( ~w3780 & w3966 ) | ( ~w3780 & w3967 ) | ( w3966 & w3967 ) ;
  assign w3969 = w3967 | w3968 ;
  assign w3970 = \pi086 ^ w3767 ;
  assign w3971 = ( ~w3774 & w3969 ) | ( ~w3774 & w3970 ) | ( w3969 & w3970 ) ;
  assign w3972 = w3970 | w3971 ;
  assign w3973 = \pi087 ^ w3761 ;
  assign w3974 = ( ~w3768 & w3972 ) | ( ~w3768 & w3973 ) | ( w3972 & w3973 ) ;
  assign w3975 = w3973 | w3974 ;
  assign w3976 = \pi088 ^ w3755 ;
  assign w3977 = ( ~w3762 & w3975 ) | ( ~w3762 & w3976 ) | ( w3975 & w3976 ) ;
  assign w3978 = w3976 | w3977 ;
  assign w3979 = \pi089 ^ w3749 ;
  assign w3980 = ( ~w3756 & w3978 ) | ( ~w3756 & w3979 ) | ( w3978 & w3979 ) ;
  assign w3981 = w3979 | w3980 ;
  assign w3982 = w3505 & w3744 ;
  assign w3983 = ~w3506 & w3734 ;
  assign w3984 = w3735 ^ w3983 ;
  assign w3985 = ~w3744 & w3984 ;
  assign w3986 = w3982 | w3985 ;
  assign w3987 = ~\pi090 & w3986 ;
  assign w3988 = ( \pi090 & ~w3982 ) | ( \pi090 & w3985 ) | ( ~w3982 & w3985 ) ;
  assign w3989 = ~w3985 & w3988 ;
  assign w3990 = \pi091 | \pi092 ;
  assign w3991 = w290 | w3990 ;
  assign w3992 = ( w240 & w275 ) | ( w240 & ~w290 ) | ( w275 & ~w290 ) ;
  assign w3993 = w3991 | w3992 ;
  assign w3994 = w3987 | w3989 ;
  assign w3995 = ( ~w3750 & w3981 ) | ( ~w3750 & w3994 ) | ( w3981 & w3994 ) ;
  assign w3996 = ( w3993 & ~w3994 ) | ( w3993 & w3995 ) | ( ~w3994 & w3995 ) ;
  assign w3997 = w3994 | w3996 ;
  assign w3998 = ~w3743 & w3986 ;
  assign w3999 = w3997 & ~w3998 ;
  assign w4000 = ~w3756 & w3978 ;
  assign w4001 = w3979 ^ w4000 ;
  assign w4002 = ~w3999 & w4001 ;
  assign w4003 = ( w3749 & w3997 ) | ( w3749 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4004 = ~w3998 & w4003 ;
  assign w4005 = w4002 | w4004 ;
  assign w4006 = ( ~w3750 & w3981 ) | ( ~w3750 & w3999 ) | ( w3981 & w3999 ) ;
  assign w4007 = w3994 ^ w4006 ;
  assign w4008 = ~w3999 & w4007 ;
  assign w4009 = ( w3743 & ~w3986 ) | ( w3743 & w3997 ) | ( ~w3986 & w3997 ) ;
  assign w4010 = w3986 & w4009 ;
  assign w4011 = w4008 | w4010 ;
  assign w4012 = ~\pi090 & w4005 ;
  assign w4013 = ~w3762 & w3975 ;
  assign w4014 = w3976 ^ w4013 ;
  assign w4015 = ~w3999 & w4014 ;
  assign w4016 = ( w3755 & w3997 ) | ( w3755 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4017 = ~w3998 & w4016 ;
  assign w4018 = w4015 | w4017 ;
  assign w4019 = ~\pi089 & w4018 ;
  assign w4020 = ~w3768 & w3972 ;
  assign w4021 = w3973 ^ w4020 ;
  assign w4022 = ~w3999 & w4021 ;
  assign w4023 = ( w3761 & w3997 ) | ( w3761 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4024 = ~w3998 & w4023 ;
  assign w4025 = w4022 | w4024 ;
  assign w4026 = ~\pi088 & w4025 ;
  assign w4027 = ~w3774 & w3969 ;
  assign w4028 = w3970 ^ w4027 ;
  assign w4029 = ~w3999 & w4028 ;
  assign w4030 = ( w3767 & w3997 ) | ( w3767 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4031 = ~w3998 & w4030 ;
  assign w4032 = w4029 | w4031 ;
  assign w4033 = ~\pi087 & w4032 ;
  assign w4034 = ~w3780 & w3966 ;
  assign w4035 = w3967 ^ w4034 ;
  assign w4036 = ~w3999 & w4035 ;
  assign w4037 = ( w3773 & w3997 ) | ( w3773 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4038 = ~w3998 & w4037 ;
  assign w4039 = w4036 | w4038 ;
  assign w4040 = ~\pi086 & w4039 ;
  assign w4041 = ~w3786 & w3963 ;
  assign w4042 = w3964 ^ w4041 ;
  assign w4043 = ~w3999 & w4042 ;
  assign w4044 = ( w3779 & w3997 ) | ( w3779 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4045 = ~w3998 & w4044 ;
  assign w4046 = w4043 | w4045 ;
  assign w4047 = ~\pi085 & w4046 ;
  assign w4048 = ~w3792 & w3960 ;
  assign w4049 = w3961 ^ w4048 ;
  assign w4050 = ~w3999 & w4049 ;
  assign w4051 = ( w3785 & w3997 ) | ( w3785 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4052 = ~w3998 & w4051 ;
  assign w4053 = w4050 | w4052 ;
  assign w4054 = ~\pi084 & w4053 ;
  assign w4055 = ~w3798 & w3957 ;
  assign w4056 = w3958 ^ w4055 ;
  assign w4057 = ~w3999 & w4056 ;
  assign w4058 = ( w3791 & w3997 ) | ( w3791 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4059 = ~w3998 & w4058 ;
  assign w4060 = w4057 | w4059 ;
  assign w4061 = ~\pi083 & w4060 ;
  assign w4062 = ~w3804 & w3954 ;
  assign w4063 = w3955 ^ w4062 ;
  assign w4064 = ~w3999 & w4063 ;
  assign w4065 = ( w3797 & w3997 ) | ( w3797 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4066 = ~w3998 & w4065 ;
  assign w4067 = w4064 | w4066 ;
  assign w4068 = ~\pi082 & w4067 ;
  assign w4069 = ~w3810 & w3951 ;
  assign w4070 = w3952 ^ w4069 ;
  assign w4071 = ~w3999 & w4070 ;
  assign w4072 = ( w3803 & w3997 ) | ( w3803 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4073 = ~w3998 & w4072 ;
  assign w4074 = w4071 | w4073 ;
  assign w4075 = ~\pi081 & w4074 ;
  assign w4076 = ~w3816 & w3948 ;
  assign w4077 = w3949 ^ w4076 ;
  assign w4078 = ~w3999 & w4077 ;
  assign w4079 = ( w3809 & w3997 ) | ( w3809 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4080 = ~w3998 & w4079 ;
  assign w4081 = w4078 | w4080 ;
  assign w4082 = ~\pi080 & w4081 ;
  assign w4083 = ~w3822 & w3945 ;
  assign w4084 = w3946 ^ w4083 ;
  assign w4085 = ~w3999 & w4084 ;
  assign w4086 = ( w3815 & w3997 ) | ( w3815 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4087 = ~w3998 & w4086 ;
  assign w4088 = w4085 | w4087 ;
  assign w4089 = ~\pi079 & w4088 ;
  assign w4090 = ~w3828 & w3942 ;
  assign w4091 = w3943 ^ w4090 ;
  assign w4092 = ~w3999 & w4091 ;
  assign w4093 = ( w3821 & w3997 ) | ( w3821 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4094 = ~w3998 & w4093 ;
  assign w4095 = w4092 | w4094 ;
  assign w4096 = ~\pi078 & w4095 ;
  assign w4097 = ~w3834 & w3939 ;
  assign w4098 = w3940 ^ w4097 ;
  assign w4099 = ~w3999 & w4098 ;
  assign w4100 = ( w3827 & w3997 ) | ( w3827 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4101 = ~w3998 & w4100 ;
  assign w4102 = w4099 | w4101 ;
  assign w4103 = ~\pi077 & w4102 ;
  assign w4104 = ~w3840 & w3936 ;
  assign w4105 = w3937 ^ w4104 ;
  assign w4106 = ~w3999 & w4105 ;
  assign w4107 = ( w3833 & w3997 ) | ( w3833 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4108 = ~w3998 & w4107 ;
  assign w4109 = w4106 | w4108 ;
  assign w4110 = ~\pi076 & w4109 ;
  assign w4111 = ~w3846 & w3933 ;
  assign w4112 = w3934 ^ w4111 ;
  assign w4113 = ~w3999 & w4112 ;
  assign w4114 = ( w3839 & w3997 ) | ( w3839 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4115 = ~w3998 & w4114 ;
  assign w4116 = w4113 | w4115 ;
  assign w4117 = ~\pi075 & w4116 ;
  assign w4118 = ~w3852 & w3930 ;
  assign w4119 = w3931 ^ w4118 ;
  assign w4120 = ~w3999 & w4119 ;
  assign w4121 = ( w3845 & w3997 ) | ( w3845 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4122 = ~w3998 & w4121 ;
  assign w4123 = w4120 | w4122 ;
  assign w4124 = ~\pi074 & w4123 ;
  assign w4125 = ~w3858 & w3927 ;
  assign w4126 = w3928 ^ w4125 ;
  assign w4127 = ~w3999 & w4126 ;
  assign w4128 = ( w3851 & w3997 ) | ( w3851 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4129 = ~w3998 & w4128 ;
  assign w4130 = w4127 | w4129 ;
  assign w4131 = ~\pi073 & w4130 ;
  assign w4132 = ~w3864 & w3924 ;
  assign w4133 = w3925 ^ w4132 ;
  assign w4134 = ~w3999 & w4133 ;
  assign w4135 = ( w3857 & w3997 ) | ( w3857 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4136 = ~w3998 & w4135 ;
  assign w4137 = w4134 | w4136 ;
  assign w4138 = ~\pi072 & w4137 ;
  assign w4139 = ~w3870 & w3921 ;
  assign w4140 = w3922 ^ w4139 ;
  assign w4141 = ~w3999 & w4140 ;
  assign w4142 = ( w3863 & w3997 ) | ( w3863 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4143 = ~w3998 & w4142 ;
  assign w4144 = w4141 | w4143 ;
  assign w4145 = ~\pi071 & w4144 ;
  assign w4146 = ~w3876 & w3918 ;
  assign w4147 = w3919 ^ w4146 ;
  assign w4148 = ~w3999 & w4147 ;
  assign w4149 = ( w3869 & w3997 ) | ( w3869 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4150 = ~w3998 & w4149 ;
  assign w4151 = w4148 | w4150 ;
  assign w4152 = ~\pi070 & w4151 ;
  assign w4153 = ~w3883 & w3915 ;
  assign w4154 = w3916 ^ w4153 ;
  assign w4155 = ~w3999 & w4154 ;
  assign w4156 = ( w3875 & w3997 ) | ( w3875 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4157 = ~w3998 & w4156 ;
  assign w4158 = w4155 | w4157 ;
  assign w4159 = ~\pi069 & w4158 ;
  assign w4160 = ~w3891 & w3912 ;
  assign w4161 = w3913 ^ w4160 ;
  assign w4162 = ~w3999 & w4161 ;
  assign w4163 = ( w3882 & w3997 ) | ( w3882 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4164 = ~w3998 & w4163 ;
  assign w4165 = w4162 | w4164 ;
  assign w4166 = ~\pi068 & w4165 ;
  assign w4167 = ( \pi065 & w3905 ) | ( \pi065 & ~w3999 ) | ( w3905 & ~w3999 ) ;
  assign w4168 = ( \pi065 & w3908 ) | ( \pi065 & ~w4167 ) | ( w3908 & ~w4167 ) ;
  assign w4169 = w3909 ^ w4168 ;
  assign w4170 = ~w3999 & w4169 ;
  assign w4171 = ( w3890 & w3997 ) | ( w3890 & w3998 ) | ( w3997 & w3998 ) ;
  assign w4172 = ~w3998 & w4171 ;
  assign w4173 = w4170 | w4172 ;
  assign w4174 = ~\pi067 & w4173 ;
  assign w4175 = w3905 ^ w3906 ;
  assign w4176 = \pi065 ^ w4175 ;
  assign w4177 = w3999 ^ w4176 ;
  assign w4178 = ( w3905 & w4176 ) | ( w3905 & w4177 ) | ( w4176 & w4177 ) ;
  assign w4179 = ~\pi066 & w4178 ;
  assign w4180 = w3905 ^ w3999 ;
  assign w4181 = ( w3905 & w4176 ) | ( w3905 & ~w4180 ) | ( w4176 & ~w4180 ) ;
  assign w4182 = \pi066 ^ w4181 ;
  assign w4183 = \pi064 & ~w3999 ;
  assign w4184 = \pi037 ^ w4183 ;
  assign w4185 = ( ~\pi036 & \pi064 ) | ( ~\pi036 & w4182 ) | ( \pi064 & w4182 ) ;
  assign w4186 = ( \pi065 & ~w4184 ) | ( \pi065 & w4185 ) | ( ~w4184 & w4185 ) ;
  assign w4187 = w4182 | w4186 ;
  assign w4188 = \pi067 ^ w4173 ;
  assign w4189 = ( ~w4179 & w4187 ) | ( ~w4179 & w4188 ) | ( w4187 & w4188 ) ;
  assign w4190 = w4188 | w4189 ;
  assign w4191 = \pi068 ^ w4165 ;
  assign w4192 = ( ~w4174 & w4190 ) | ( ~w4174 & w4191 ) | ( w4190 & w4191 ) ;
  assign w4193 = w4191 | w4192 ;
  assign w4194 = \pi069 ^ w4158 ;
  assign w4195 = ( ~w4166 & w4193 ) | ( ~w4166 & w4194 ) | ( w4193 & w4194 ) ;
  assign w4196 = w4194 | w4195 ;
  assign w4197 = \pi070 ^ w4151 ;
  assign w4198 = ( ~w4159 & w4196 ) | ( ~w4159 & w4197 ) | ( w4196 & w4197 ) ;
  assign w4199 = w4197 | w4198 ;
  assign w4200 = \pi071 ^ w4144 ;
  assign w4201 = ( ~w4152 & w4199 ) | ( ~w4152 & w4200 ) | ( w4199 & w4200 ) ;
  assign w4202 = w4200 | w4201 ;
  assign w4203 = \pi072 ^ w4137 ;
  assign w4204 = ( ~w4145 & w4202 ) | ( ~w4145 & w4203 ) | ( w4202 & w4203 ) ;
  assign w4205 = w4203 | w4204 ;
  assign w4206 = \pi073 ^ w4130 ;
  assign w4207 = ( ~w4138 & w4205 ) | ( ~w4138 & w4206 ) | ( w4205 & w4206 ) ;
  assign w4208 = w4206 | w4207 ;
  assign w4209 = \pi074 ^ w4123 ;
  assign w4210 = ( ~w4131 & w4208 ) | ( ~w4131 & w4209 ) | ( w4208 & w4209 ) ;
  assign w4211 = w4209 | w4210 ;
  assign w4212 = \pi075 ^ w4116 ;
  assign w4213 = ( ~w4124 & w4211 ) | ( ~w4124 & w4212 ) | ( w4211 & w4212 ) ;
  assign w4214 = w4212 | w4213 ;
  assign w4215 = \pi076 ^ w4109 ;
  assign w4216 = ( ~w4117 & w4214 ) | ( ~w4117 & w4215 ) | ( w4214 & w4215 ) ;
  assign w4217 = w4215 | w4216 ;
  assign w4218 = \pi077 ^ w4102 ;
  assign w4219 = ( ~w4110 & w4217 ) | ( ~w4110 & w4218 ) | ( w4217 & w4218 ) ;
  assign w4220 = w4218 | w4219 ;
  assign w4221 = \pi078 ^ w4095 ;
  assign w4222 = ( ~w4103 & w4220 ) | ( ~w4103 & w4221 ) | ( w4220 & w4221 ) ;
  assign w4223 = w4221 | w4222 ;
  assign w4224 = \pi079 ^ w4088 ;
  assign w4225 = ( ~w4096 & w4223 ) | ( ~w4096 & w4224 ) | ( w4223 & w4224 ) ;
  assign w4226 = w4224 | w4225 ;
  assign w4227 = \pi080 ^ w4081 ;
  assign w4228 = ( ~w4089 & w4226 ) | ( ~w4089 & w4227 ) | ( w4226 & w4227 ) ;
  assign w4229 = w4227 | w4228 ;
  assign w4230 = \pi081 ^ w4074 ;
  assign w4231 = ( ~w4082 & w4229 ) | ( ~w4082 & w4230 ) | ( w4229 & w4230 ) ;
  assign w4232 = w4230 | w4231 ;
  assign w4233 = \pi082 ^ w4067 ;
  assign w4234 = ( ~w4075 & w4232 ) | ( ~w4075 & w4233 ) | ( w4232 & w4233 ) ;
  assign w4235 = w4233 | w4234 ;
  assign w4236 = \pi083 ^ w4060 ;
  assign w4237 = ( ~w4068 & w4235 ) | ( ~w4068 & w4236 ) | ( w4235 & w4236 ) ;
  assign w4238 = w4236 | w4237 ;
  assign w4239 = \pi084 ^ w4053 ;
  assign w4240 = ( ~w4061 & w4238 ) | ( ~w4061 & w4239 ) | ( w4238 & w4239 ) ;
  assign w4241 = w4239 | w4240 ;
  assign w4242 = \pi085 ^ w4046 ;
  assign w4243 = ( ~w4054 & w4241 ) | ( ~w4054 & w4242 ) | ( w4241 & w4242 ) ;
  assign w4244 = w4242 | w4243 ;
  assign w4245 = \pi086 ^ w4039 ;
  assign w4246 = ( ~w4047 & w4244 ) | ( ~w4047 & w4245 ) | ( w4244 & w4245 ) ;
  assign w4247 = w4245 | w4246 ;
  assign w4248 = \pi087 ^ w4032 ;
  assign w4249 = ( ~w4040 & w4247 ) | ( ~w4040 & w4248 ) | ( w4247 & w4248 ) ;
  assign w4250 = w4248 | w4249 ;
  assign w4251 = \pi088 ^ w4025 ;
  assign w4252 = ( ~w4033 & w4250 ) | ( ~w4033 & w4251 ) | ( w4250 & w4251 ) ;
  assign w4253 = w4251 | w4252 ;
  assign w4254 = \pi089 ^ w4018 ;
  assign w4255 = ( ~w4026 & w4253 ) | ( ~w4026 & w4254 ) | ( w4253 & w4254 ) ;
  assign w4256 = w4254 | w4255 ;
  assign w4257 = \pi090 ^ w4005 ;
  assign w4258 = ( ~w4019 & w4256 ) | ( ~w4019 & w4257 ) | ( w4256 & w4257 ) ;
  assign w4259 = w4257 | w4258 ;
  assign w4260 = \pi091 ^ w4011 ;
  assign w4261 = w4012 & ~w4260 ;
  assign w4262 = ( w4259 & w4260 ) | ( w4259 & ~w4261 ) | ( w4260 & ~w4261 ) ;
  assign w4263 = ~\pi091 & w4011 ;
  assign w4264 = w4262 & ~w4263 ;
  assign w4265 = ( ~w155 & w170 ) | ( ~w155 & w183 ) | ( w170 & w183 ) ;
  assign w4266 = w155 | w4265 ;
  assign w4267 = w4264 | w4266 ;
  assign w4268 = w4005 & w4267 ;
  assign w4269 = ~w4019 & w4256 ;
  assign w4270 = w4257 ^ w4269 ;
  assign w4271 = ~w4267 & w4270 ;
  assign w4272 = w4268 | w4271 ;
  assign w4273 = w4011 & w4267 ;
  assign w4274 = ~w4012 & w4259 ;
  assign w4275 = w4260 ^ w4274 ;
  assign w4276 = ~w4267 & w4275 ;
  assign w4277 = w4273 | w4276 ;
  assign w4278 = ~\pi091 & w4272 ;
  assign w4279 = w4018 & w4267 ;
  assign w4280 = ~w4026 & w4253 ;
  assign w4281 = w4254 ^ w4280 ;
  assign w4282 = ~w4267 & w4281 ;
  assign w4283 = w4279 | w4282 ;
  assign w4284 = ~\pi090 & w4283 ;
  assign w4285 = w4025 & w4267 ;
  assign w4286 = ~w4033 & w4250 ;
  assign w4287 = w4251 ^ w4286 ;
  assign w4288 = ~w4267 & w4287 ;
  assign w4289 = w4285 | w4288 ;
  assign w4290 = ~\pi089 & w4289 ;
  assign w4291 = w4032 & w4267 ;
  assign w4292 = ~w4040 & w4247 ;
  assign w4293 = w4248 ^ w4292 ;
  assign w4294 = ~w4267 & w4293 ;
  assign w4295 = w4291 | w4294 ;
  assign w4296 = ~\pi088 & w4295 ;
  assign w4297 = w4039 & w4267 ;
  assign w4298 = ~w4047 & w4244 ;
  assign w4299 = w4245 ^ w4298 ;
  assign w4300 = ~w4267 & w4299 ;
  assign w4301 = w4297 | w4300 ;
  assign w4302 = ~\pi087 & w4301 ;
  assign w4303 = w4046 & w4267 ;
  assign w4304 = ~w4054 & w4241 ;
  assign w4305 = w4242 ^ w4304 ;
  assign w4306 = ~w4267 & w4305 ;
  assign w4307 = w4303 | w4306 ;
  assign w4308 = ~\pi086 & w4307 ;
  assign w4309 = w4053 & w4267 ;
  assign w4310 = ~w4061 & w4238 ;
  assign w4311 = w4239 ^ w4310 ;
  assign w4312 = ~w4267 & w4311 ;
  assign w4313 = w4309 | w4312 ;
  assign w4314 = ~\pi085 & w4313 ;
  assign w4315 = w4060 & w4267 ;
  assign w4316 = ~w4068 & w4235 ;
  assign w4317 = w4236 ^ w4316 ;
  assign w4318 = ~w4267 & w4317 ;
  assign w4319 = w4315 | w4318 ;
  assign w4320 = ~\pi084 & w4319 ;
  assign w4321 = w4067 & w4267 ;
  assign w4322 = ~w4075 & w4232 ;
  assign w4323 = w4233 ^ w4322 ;
  assign w4324 = ~w4267 & w4323 ;
  assign w4325 = w4321 | w4324 ;
  assign w4326 = ~\pi083 & w4325 ;
  assign w4327 = w4074 & w4267 ;
  assign w4328 = ~w4082 & w4229 ;
  assign w4329 = w4230 ^ w4328 ;
  assign w4330 = ~w4267 & w4329 ;
  assign w4331 = w4327 | w4330 ;
  assign w4332 = ~\pi082 & w4331 ;
  assign w4333 = w4081 & w4267 ;
  assign w4334 = ~w4089 & w4226 ;
  assign w4335 = w4227 ^ w4334 ;
  assign w4336 = ~w4267 & w4335 ;
  assign w4337 = w4333 | w4336 ;
  assign w4338 = ~\pi081 & w4337 ;
  assign w4339 = w4088 & w4267 ;
  assign w4340 = ~w4096 & w4223 ;
  assign w4341 = w4224 ^ w4340 ;
  assign w4342 = ~w4267 & w4341 ;
  assign w4343 = w4339 | w4342 ;
  assign w4344 = ~\pi080 & w4343 ;
  assign w4345 = w4095 & w4267 ;
  assign w4346 = ~w4103 & w4220 ;
  assign w4347 = w4221 ^ w4346 ;
  assign w4348 = ~w4267 & w4347 ;
  assign w4349 = w4345 | w4348 ;
  assign w4350 = ~\pi079 & w4349 ;
  assign w4351 = w4102 & w4267 ;
  assign w4352 = ~w4110 & w4217 ;
  assign w4353 = w4218 ^ w4352 ;
  assign w4354 = ~w4267 & w4353 ;
  assign w4355 = w4351 | w4354 ;
  assign w4356 = ~\pi078 & w4355 ;
  assign w4357 = w4109 & w4267 ;
  assign w4358 = ~w4117 & w4214 ;
  assign w4359 = w4215 ^ w4358 ;
  assign w4360 = ~w4267 & w4359 ;
  assign w4361 = w4357 | w4360 ;
  assign w4362 = ~\pi077 & w4361 ;
  assign w4363 = w4116 & w4267 ;
  assign w4364 = ~w4124 & w4211 ;
  assign w4365 = w4212 ^ w4364 ;
  assign w4366 = ~w4267 & w4365 ;
  assign w4367 = w4363 | w4366 ;
  assign w4368 = ~\pi076 & w4367 ;
  assign w4369 = w4123 & w4267 ;
  assign w4370 = ~w4131 & w4208 ;
  assign w4371 = w4209 ^ w4370 ;
  assign w4372 = ~w4267 & w4371 ;
  assign w4373 = w4369 | w4372 ;
  assign w4374 = ~\pi075 & w4373 ;
  assign w4375 = w4130 & w4267 ;
  assign w4376 = ~w4138 & w4205 ;
  assign w4377 = w4206 ^ w4376 ;
  assign w4378 = ~w4267 & w4377 ;
  assign w4379 = w4375 | w4378 ;
  assign w4380 = ~\pi074 & w4379 ;
  assign w4381 = w4137 & w4267 ;
  assign w4382 = ~w4145 & w4202 ;
  assign w4383 = w4203 ^ w4382 ;
  assign w4384 = ~w4267 & w4383 ;
  assign w4385 = w4381 | w4384 ;
  assign w4386 = ~\pi073 & w4385 ;
  assign w4387 = w4144 & w4267 ;
  assign w4388 = ~w4152 & w4199 ;
  assign w4389 = w4200 ^ w4388 ;
  assign w4390 = ~w4267 & w4389 ;
  assign w4391 = w4387 | w4390 ;
  assign w4392 = ~\pi072 & w4391 ;
  assign w4393 = w4151 & w4267 ;
  assign w4394 = ~w4159 & w4196 ;
  assign w4395 = w4197 ^ w4394 ;
  assign w4396 = ~w4267 & w4395 ;
  assign w4397 = w4393 | w4396 ;
  assign w4398 = ~\pi071 & w4397 ;
  assign w4399 = w4158 & w4267 ;
  assign w4400 = ~w4166 & w4193 ;
  assign w4401 = w4194 ^ w4400 ;
  assign w4402 = ~w4267 & w4401 ;
  assign w4403 = w4399 | w4402 ;
  assign w4404 = ~\pi070 & w4403 ;
  assign w4405 = w4165 & w4267 ;
  assign w4406 = ~w4174 & w4190 ;
  assign w4407 = w4191 ^ w4406 ;
  assign w4408 = ~w4267 & w4407 ;
  assign w4409 = w4405 | w4408 ;
  assign w4410 = ~\pi069 & w4409 ;
  assign w4411 = w4173 & w4267 ;
  assign w4412 = ~w4179 & w4187 ;
  assign w4413 = w4188 ^ w4412 ;
  assign w4414 = ~w4267 & w4413 ;
  assign w4415 = w4411 | w4414 ;
  assign w4416 = ~\pi068 & w4415 ;
  assign w4417 = w4178 & w4267 ;
  assign w4418 = ~\pi036 & \pi064 ;
  assign w4419 = ( \pi065 & ~w4184 ) | ( \pi065 & w4418 ) | ( ~w4184 & w4418 ) ;
  assign w4420 = w4182 ^ w4419 ;
  assign w4421 = ( w4264 & w4266 ) | ( w4264 & w4420 ) | ( w4266 & w4420 ) ;
  assign w4422 = w4420 & ~w4421 ;
  assign w4423 = w4417 | w4422 ;
  assign w4424 = ~\pi067 & w4423 ;
  assign w4425 = \pi037 ^ \pi065 ;
  assign w4426 = \pi036 ^ w3999 ;
  assign w4427 = ( \pi064 & w4266 ) | ( \pi064 & w4426 ) | ( w4266 & w4426 ) ;
  assign w4428 = w4425 ^ w4427 ;
  assign w4429 = ~w4266 & w4428 ;
  assign w4430 = ~w4264 & w4429 ;
  assign w4431 = ( ~\pi064 & w3999 ) | ( ~\pi064 & w4267 ) | ( w3999 & w4267 ) ;
  assign w4432 = \pi037 ^ w4431 ;
  assign w4433 = w4267 & ~w4432 ;
  assign w4434 = w4430 | w4433 ;
  assign w4435 = ~\pi066 & w4434 ;
  assign w4436 = \pi064 & ~\pi092 ;
  assign w4437 = ~w290 & w4436 ;
  assign w4438 = ~w3992 & w4437 ;
  assign w4439 = ( \pi036 & w4264 ) | ( \pi036 & ~w4438 ) | ( w4264 & ~w4438 ) ;
  assign w4440 = \pi036 & w4439 ;
  assign w4441 = ~w204 & w4418 ;
  assign w4442 = ~w3742 & w4441 ;
  assign w4443 = ~w4264 & w4442 ;
  assign w4444 = w4440 | w4443 ;
  assign w4445 = ~\pi035 & \pi064 ;
  assign w4446 = \pi065 ^ w4444 ;
  assign w4447 = w4445 | w4446 ;
  assign w4448 = w4267 | w4430 ;
  assign w4449 = ( w4184 & w4430 ) | ( w4184 & w4448 ) | ( w4430 & w4448 ) ;
  assign w4450 = \pi066 ^ w4449 ;
  assign w4451 = ~\pi065 & w4444 ;
  assign w4452 = w4447 | w4451 ;
  assign w4453 = ( w4450 & ~w4451 ) | ( w4450 & w4452 ) | ( ~w4451 & w4452 ) ;
  assign w4454 = \pi067 ^ w4423 ;
  assign w4455 = ( ~w4435 & w4453 ) | ( ~w4435 & w4454 ) | ( w4453 & w4454 ) ;
  assign w4456 = w4454 | w4455 ;
  assign w4457 = \pi068 ^ w4415 ;
  assign w4458 = ( ~w4424 & w4456 ) | ( ~w4424 & w4457 ) | ( w4456 & w4457 ) ;
  assign w4459 = w4457 | w4458 ;
  assign w4460 = \pi069 ^ w4409 ;
  assign w4461 = ( ~w4416 & w4459 ) | ( ~w4416 & w4460 ) | ( w4459 & w4460 ) ;
  assign w4462 = w4460 | w4461 ;
  assign w4463 = \pi070 ^ w4403 ;
  assign w4464 = ( ~w4410 & w4462 ) | ( ~w4410 & w4463 ) | ( w4462 & w4463 ) ;
  assign w4465 = w4463 | w4464 ;
  assign w4466 = \pi071 ^ w4397 ;
  assign w4467 = ( ~w4404 & w4465 ) | ( ~w4404 & w4466 ) | ( w4465 & w4466 ) ;
  assign w4468 = w4466 | w4467 ;
  assign w4469 = \pi072 ^ w4391 ;
  assign w4470 = ( ~w4398 & w4468 ) | ( ~w4398 & w4469 ) | ( w4468 & w4469 ) ;
  assign w4471 = w4469 | w4470 ;
  assign w4472 = \pi073 ^ w4385 ;
  assign w4473 = ( ~w4392 & w4471 ) | ( ~w4392 & w4472 ) | ( w4471 & w4472 ) ;
  assign w4474 = w4472 | w4473 ;
  assign w4475 = \pi074 ^ w4379 ;
  assign w4476 = ( ~w4386 & w4474 ) | ( ~w4386 & w4475 ) | ( w4474 & w4475 ) ;
  assign w4477 = w4475 | w4476 ;
  assign w4478 = \pi075 ^ w4373 ;
  assign w4479 = ( ~w4380 & w4477 ) | ( ~w4380 & w4478 ) | ( w4477 & w4478 ) ;
  assign w4480 = w4478 | w4479 ;
  assign w4481 = \pi076 ^ w4367 ;
  assign w4482 = ( ~w4374 & w4480 ) | ( ~w4374 & w4481 ) | ( w4480 & w4481 ) ;
  assign w4483 = w4481 | w4482 ;
  assign w4484 = \pi077 ^ w4361 ;
  assign w4485 = ( ~w4368 & w4483 ) | ( ~w4368 & w4484 ) | ( w4483 & w4484 ) ;
  assign w4486 = w4484 | w4485 ;
  assign w4487 = \pi078 ^ w4355 ;
  assign w4488 = ( ~w4362 & w4486 ) | ( ~w4362 & w4487 ) | ( w4486 & w4487 ) ;
  assign w4489 = w4487 | w4488 ;
  assign w4490 = \pi079 ^ w4349 ;
  assign w4491 = ( ~w4356 & w4489 ) | ( ~w4356 & w4490 ) | ( w4489 & w4490 ) ;
  assign w4492 = w4490 | w4491 ;
  assign w4493 = \pi080 ^ w4343 ;
  assign w4494 = ( ~w4350 & w4492 ) | ( ~w4350 & w4493 ) | ( w4492 & w4493 ) ;
  assign w4495 = w4493 | w4494 ;
  assign w4496 = \pi081 ^ w4337 ;
  assign w4497 = ( ~w4344 & w4495 ) | ( ~w4344 & w4496 ) | ( w4495 & w4496 ) ;
  assign w4498 = w4496 | w4497 ;
  assign w4499 = \pi082 ^ w4331 ;
  assign w4500 = ( ~w4338 & w4498 ) | ( ~w4338 & w4499 ) | ( w4498 & w4499 ) ;
  assign w4501 = w4499 | w4500 ;
  assign w4502 = \pi083 ^ w4325 ;
  assign w4503 = ( ~w4332 & w4501 ) | ( ~w4332 & w4502 ) | ( w4501 & w4502 ) ;
  assign w4504 = w4502 | w4503 ;
  assign w4505 = \pi084 ^ w4319 ;
  assign w4506 = ( ~w4326 & w4504 ) | ( ~w4326 & w4505 ) | ( w4504 & w4505 ) ;
  assign w4507 = w4505 | w4506 ;
  assign w4508 = \pi085 ^ w4313 ;
  assign w4509 = ( ~w4320 & w4507 ) | ( ~w4320 & w4508 ) | ( w4507 & w4508 ) ;
  assign w4510 = w4508 | w4509 ;
  assign w4511 = \pi086 ^ w4307 ;
  assign w4512 = ( ~w4314 & w4510 ) | ( ~w4314 & w4511 ) | ( w4510 & w4511 ) ;
  assign w4513 = w4511 | w4512 ;
  assign w4514 = \pi087 ^ w4301 ;
  assign w4515 = ( ~w4308 & w4513 ) | ( ~w4308 & w4514 ) | ( w4513 & w4514 ) ;
  assign w4516 = w4514 | w4515 ;
  assign w4517 = \pi088 ^ w4295 ;
  assign w4518 = ( ~w4302 & w4516 ) | ( ~w4302 & w4517 ) | ( w4516 & w4517 ) ;
  assign w4519 = w4517 | w4518 ;
  assign w4520 = \pi089 ^ w4289 ;
  assign w4521 = ( ~w4296 & w4519 ) | ( ~w4296 & w4520 ) | ( w4519 & w4520 ) ;
  assign w4522 = w4520 | w4521 ;
  assign w4523 = \pi090 ^ w4283 ;
  assign w4524 = ( ~w4290 & w4522 ) | ( ~w4290 & w4523 ) | ( w4522 & w4523 ) ;
  assign w4525 = w4523 | w4524 ;
  assign w4526 = \pi091 ^ w4272 ;
  assign w4527 = ( ~w4284 & w4525 ) | ( ~w4284 & w4526 ) | ( w4525 & w4526 ) ;
  assign w4528 = w4526 | w4527 ;
  assign w4529 = \pi092 ^ w4277 ;
  assign w4530 = w4278 & ~w4529 ;
  assign w4531 = ( w4528 & w4529 ) | ( w4528 & ~w4530 ) | ( w4529 & ~w4530 ) ;
  assign w4532 = ~\pi092 & w4277 ;
  assign w4533 = w4531 & ~w4532 ;
  assign w4534 = ( w441 & w448 ) | ( w441 & ~w451 ) | ( w448 & ~w451 ) ;
  assign w4535 = w451 | w4534 ;
  assign w4536 = w4533 | w4535 ;
  assign w4537 = w4272 & w4536 ;
  assign w4538 = ~w4284 & w4525 ;
  assign w4539 = w4526 ^ w4538 ;
  assign w4540 = ~w4536 & w4539 ;
  assign w4541 = w4537 | w4540 ;
  assign w4542 = ~\pi092 & w4541 ;
  assign w4543 = w4283 & w4536 ;
  assign w4544 = ~w4290 & w4522 ;
  assign w4545 = w4523 ^ w4544 ;
  assign w4546 = ~w4536 & w4545 ;
  assign w4547 = w4543 | w4546 ;
  assign w4548 = ~\pi091 & w4547 ;
  assign w4549 = w4289 & w4536 ;
  assign w4550 = ~w4296 & w4519 ;
  assign w4551 = w4520 ^ w4550 ;
  assign w4552 = ~w4536 & w4551 ;
  assign w4553 = w4549 | w4552 ;
  assign w4554 = ~\pi090 & w4553 ;
  assign w4555 = w4295 & w4536 ;
  assign w4556 = ~w4302 & w4516 ;
  assign w4557 = w4517 ^ w4556 ;
  assign w4558 = ~w4536 & w4557 ;
  assign w4559 = w4555 | w4558 ;
  assign w4560 = ~\pi089 & w4559 ;
  assign w4561 = w4301 & w4536 ;
  assign w4562 = ~w4308 & w4513 ;
  assign w4563 = w4514 ^ w4562 ;
  assign w4564 = ~w4536 & w4563 ;
  assign w4565 = w4561 | w4564 ;
  assign w4566 = ~\pi088 & w4565 ;
  assign w4567 = w4307 & w4536 ;
  assign w4568 = ~w4314 & w4510 ;
  assign w4569 = w4511 ^ w4568 ;
  assign w4570 = ~w4536 & w4569 ;
  assign w4571 = w4567 | w4570 ;
  assign w4572 = ~\pi087 & w4571 ;
  assign w4573 = w4313 & w4536 ;
  assign w4574 = ~w4320 & w4507 ;
  assign w4575 = w4508 ^ w4574 ;
  assign w4576 = ~w4536 & w4575 ;
  assign w4577 = w4573 | w4576 ;
  assign w4578 = ~\pi086 & w4577 ;
  assign w4579 = w4319 & w4536 ;
  assign w4580 = ~w4326 & w4504 ;
  assign w4581 = w4505 ^ w4580 ;
  assign w4582 = ~w4536 & w4581 ;
  assign w4583 = w4579 | w4582 ;
  assign w4584 = ~\pi085 & w4583 ;
  assign w4585 = w4325 & w4536 ;
  assign w4586 = ~w4332 & w4501 ;
  assign w4587 = w4502 ^ w4586 ;
  assign w4588 = ~w4536 & w4587 ;
  assign w4589 = w4585 | w4588 ;
  assign w4590 = ~\pi084 & w4589 ;
  assign w4591 = w4331 & w4536 ;
  assign w4592 = ~w4338 & w4498 ;
  assign w4593 = w4499 ^ w4592 ;
  assign w4594 = ~w4536 & w4593 ;
  assign w4595 = w4591 | w4594 ;
  assign w4596 = ~\pi083 & w4595 ;
  assign w4597 = w4337 & w4536 ;
  assign w4598 = ~w4344 & w4495 ;
  assign w4599 = w4496 ^ w4598 ;
  assign w4600 = ~w4536 & w4599 ;
  assign w4601 = w4597 | w4600 ;
  assign w4602 = ~\pi082 & w4601 ;
  assign w4603 = w4343 & w4536 ;
  assign w4604 = ~w4350 & w4492 ;
  assign w4605 = w4493 ^ w4604 ;
  assign w4606 = ~w4536 & w4605 ;
  assign w4607 = w4603 | w4606 ;
  assign w4608 = ~\pi081 & w4607 ;
  assign w4609 = w4349 & w4536 ;
  assign w4610 = ~w4356 & w4489 ;
  assign w4611 = w4490 ^ w4610 ;
  assign w4612 = ~w4536 & w4611 ;
  assign w4613 = w4609 | w4612 ;
  assign w4614 = ~\pi080 & w4613 ;
  assign w4615 = w4355 & w4536 ;
  assign w4616 = ~w4362 & w4486 ;
  assign w4617 = w4487 ^ w4616 ;
  assign w4618 = ~w4536 & w4617 ;
  assign w4619 = w4615 | w4618 ;
  assign w4620 = ~\pi079 & w4619 ;
  assign w4621 = w4361 & w4536 ;
  assign w4622 = ~w4368 & w4483 ;
  assign w4623 = w4484 ^ w4622 ;
  assign w4624 = ~w4536 & w4623 ;
  assign w4625 = w4621 | w4624 ;
  assign w4626 = ~\pi078 & w4625 ;
  assign w4627 = w4367 & w4536 ;
  assign w4628 = ~w4374 & w4480 ;
  assign w4629 = w4481 ^ w4628 ;
  assign w4630 = ~w4536 & w4629 ;
  assign w4631 = w4627 | w4630 ;
  assign w4632 = ~\pi077 & w4631 ;
  assign w4633 = w4373 & w4536 ;
  assign w4634 = ~w4380 & w4477 ;
  assign w4635 = w4478 ^ w4634 ;
  assign w4636 = ~w4536 & w4635 ;
  assign w4637 = w4633 | w4636 ;
  assign w4638 = ~\pi076 & w4637 ;
  assign w4639 = w4379 & w4536 ;
  assign w4640 = ~w4386 & w4474 ;
  assign w4641 = w4475 ^ w4640 ;
  assign w4642 = ~w4536 & w4641 ;
  assign w4643 = w4639 | w4642 ;
  assign w4644 = ~\pi075 & w4643 ;
  assign w4645 = w4385 & w4536 ;
  assign w4646 = ~w4392 & w4471 ;
  assign w4647 = w4472 ^ w4646 ;
  assign w4648 = ~w4536 & w4647 ;
  assign w4649 = w4645 | w4648 ;
  assign w4650 = ~\pi074 & w4649 ;
  assign w4651 = w4391 & w4536 ;
  assign w4652 = ~w4398 & w4468 ;
  assign w4653 = w4469 ^ w4652 ;
  assign w4654 = ~w4536 & w4653 ;
  assign w4655 = w4651 | w4654 ;
  assign w4656 = ~\pi073 & w4655 ;
  assign w4657 = w4397 & w4536 ;
  assign w4658 = ~w4404 & w4465 ;
  assign w4659 = w4466 ^ w4658 ;
  assign w4660 = ~w4536 & w4659 ;
  assign w4661 = w4657 | w4660 ;
  assign w4662 = ~\pi072 & w4661 ;
  assign w4663 = w4403 & w4536 ;
  assign w4664 = ~w4410 & w4462 ;
  assign w4665 = w4463 ^ w4664 ;
  assign w4666 = ~w4536 & w4665 ;
  assign w4667 = w4663 | w4666 ;
  assign w4668 = ~\pi071 & w4667 ;
  assign w4669 = w4409 & w4536 ;
  assign w4670 = ~w4416 & w4459 ;
  assign w4671 = w4460 ^ w4670 ;
  assign w4672 = ~w4536 & w4671 ;
  assign w4673 = w4669 | w4672 ;
  assign w4674 = ~\pi070 & w4673 ;
  assign w4675 = w4415 & w4536 ;
  assign w4676 = ~w4424 & w4456 ;
  assign w4677 = w4457 ^ w4676 ;
  assign w4678 = ~w4536 & w4677 ;
  assign w4679 = w4675 | w4678 ;
  assign w4680 = ~\pi069 & w4679 ;
  assign w4681 = w4423 & w4536 ;
  assign w4682 = ~w4435 & w4453 ;
  assign w4683 = w4454 ^ w4682 ;
  assign w4684 = ~w4536 & w4683 ;
  assign w4685 = w4681 | w4684 ;
  assign w4686 = ~\pi068 & w4685 ;
  assign w4687 = w4434 & w4536 ;
  assign w4688 = ~w4444 & w4447 ;
  assign w4689 = ( \pi065 & w4447 ) | ( \pi065 & w4688 ) | ( w4447 & w4688 ) ;
  assign w4690 = w4450 ^ w4689 ;
  assign w4691 = ~w4536 & w4690 ;
  assign w4692 = w4687 | w4691 ;
  assign w4693 = ~\pi067 & w4692 ;
  assign w4694 = ( w4440 & w4443 ) | ( w4440 & ~w4535 ) | ( w4443 & ~w4535 ) ;
  assign w4695 = \pi065 ^ w4694 ;
  assign w4696 = ( w4445 & ~w4535 ) | ( w4445 & w4695 ) | ( ~w4535 & w4695 ) ;
  assign w4697 = ( w4445 & w4533 ) | ( w4445 & w4695 ) | ( w4533 & w4695 ) ;
  assign w4698 = w4696 & ~w4697 ;
  assign w4699 = ( w4444 & w4536 ) | ( w4444 & w4698 ) | ( w4536 & w4698 ) ;
  assign w4700 = w4698 | w4699 ;
  assign w4701 = ~\pi066 & w4700 ;
  assign w4702 = ( \pi064 & ~\pi093 ) | ( \pi064 & \pi094 ) | ( ~\pi093 & \pi094 ) ;
  assign w4703 = w170 | w179 ;
  assign w4704 = ( \pi094 & \pi095 ) | ( \pi094 & ~w179 ) | ( \pi095 & ~w179 ) ;
  assign w4705 = w4703 | w4704 ;
  assign w4706 = w4702 & ~w4705 ;
  assign w4707 = ~w155 & w4706 ;
  assign w4708 = ( \pi035 & w4533 ) | ( \pi035 & ~w4707 ) | ( w4533 & ~w4707 ) ;
  assign w4709 = \pi035 & w4708 ;
  assign w4710 = ~w240 & w4445 ;
  assign w4711 = ~w275 & w4710 ;
  assign w4712 = ( ~w275 & w290 ) | ( ~w275 & w4533 ) | ( w290 & w4533 ) ;
  assign w4713 = w4711 & ~w4712 ;
  assign w4714 = ~\pi034 & \pi064 ;
  assign w4715 = ~w4444 & w4536 ;
  assign w4716 = ( w4536 & w4698 ) | ( w4536 & ~w4715 ) | ( w4698 & ~w4715 ) ;
  assign w4717 = \pi066 ^ w4716 ;
  assign w4718 = w4709 | w4713 ;
  assign w4719 = ( \pi065 & w4714 ) | ( \pi065 & ~w4718 ) | ( w4714 & ~w4718 ) ;
  assign w4720 = w4717 | w4719 ;
  assign w4721 = \pi067 ^ w4692 ;
  assign w4722 = ( ~w4701 & w4720 ) | ( ~w4701 & w4721 ) | ( w4720 & w4721 ) ;
  assign w4723 = w4721 | w4722 ;
  assign w4724 = \pi068 ^ w4685 ;
  assign w4725 = ( ~w4693 & w4723 ) | ( ~w4693 & w4724 ) | ( w4723 & w4724 ) ;
  assign w4726 = w4724 | w4725 ;
  assign w4727 = \pi069 ^ w4679 ;
  assign w4728 = ( ~w4686 & w4726 ) | ( ~w4686 & w4727 ) | ( w4726 & w4727 ) ;
  assign w4729 = w4727 | w4728 ;
  assign w4730 = \pi070 ^ w4673 ;
  assign w4731 = ( ~w4680 & w4729 ) | ( ~w4680 & w4730 ) | ( w4729 & w4730 ) ;
  assign w4732 = w4730 | w4731 ;
  assign w4733 = \pi071 ^ w4667 ;
  assign w4734 = ( ~w4674 & w4732 ) | ( ~w4674 & w4733 ) | ( w4732 & w4733 ) ;
  assign w4735 = w4733 | w4734 ;
  assign w4736 = \pi072 ^ w4661 ;
  assign w4737 = ( ~w4668 & w4735 ) | ( ~w4668 & w4736 ) | ( w4735 & w4736 ) ;
  assign w4738 = w4736 | w4737 ;
  assign w4739 = \pi073 ^ w4655 ;
  assign w4740 = ( ~w4662 & w4738 ) | ( ~w4662 & w4739 ) | ( w4738 & w4739 ) ;
  assign w4741 = w4739 | w4740 ;
  assign w4742 = \pi074 ^ w4649 ;
  assign w4743 = ( ~w4656 & w4741 ) | ( ~w4656 & w4742 ) | ( w4741 & w4742 ) ;
  assign w4744 = w4742 | w4743 ;
  assign w4745 = \pi075 ^ w4643 ;
  assign w4746 = ( ~w4650 & w4744 ) | ( ~w4650 & w4745 ) | ( w4744 & w4745 ) ;
  assign w4747 = w4745 | w4746 ;
  assign w4748 = \pi076 ^ w4637 ;
  assign w4749 = ( ~w4644 & w4747 ) | ( ~w4644 & w4748 ) | ( w4747 & w4748 ) ;
  assign w4750 = w4748 | w4749 ;
  assign w4751 = \pi077 ^ w4631 ;
  assign w4752 = ( ~w4638 & w4750 ) | ( ~w4638 & w4751 ) | ( w4750 & w4751 ) ;
  assign w4753 = w4751 | w4752 ;
  assign w4754 = \pi078 ^ w4625 ;
  assign w4755 = ( ~w4632 & w4753 ) | ( ~w4632 & w4754 ) | ( w4753 & w4754 ) ;
  assign w4756 = w4754 | w4755 ;
  assign w4757 = \pi079 ^ w4619 ;
  assign w4758 = ( ~w4626 & w4756 ) | ( ~w4626 & w4757 ) | ( w4756 & w4757 ) ;
  assign w4759 = w4757 | w4758 ;
  assign w4760 = \pi080 ^ w4613 ;
  assign w4761 = ( ~w4620 & w4759 ) | ( ~w4620 & w4760 ) | ( w4759 & w4760 ) ;
  assign w4762 = w4760 | w4761 ;
  assign w4763 = \pi081 ^ w4607 ;
  assign w4764 = ( ~w4614 & w4762 ) | ( ~w4614 & w4763 ) | ( w4762 & w4763 ) ;
  assign w4765 = w4763 | w4764 ;
  assign w4766 = \pi082 ^ w4601 ;
  assign w4767 = ( ~w4608 & w4765 ) | ( ~w4608 & w4766 ) | ( w4765 & w4766 ) ;
  assign w4768 = w4766 | w4767 ;
  assign w4769 = \pi083 ^ w4595 ;
  assign w4770 = ( ~w4602 & w4768 ) | ( ~w4602 & w4769 ) | ( w4768 & w4769 ) ;
  assign w4771 = w4769 | w4770 ;
  assign w4772 = \pi084 ^ w4589 ;
  assign w4773 = ( ~w4596 & w4771 ) | ( ~w4596 & w4772 ) | ( w4771 & w4772 ) ;
  assign w4774 = w4772 | w4773 ;
  assign w4775 = \pi085 ^ w4583 ;
  assign w4776 = ( ~w4590 & w4774 ) | ( ~w4590 & w4775 ) | ( w4774 & w4775 ) ;
  assign w4777 = w4775 | w4776 ;
  assign w4778 = \pi086 ^ w4577 ;
  assign w4779 = ( ~w4584 & w4777 ) | ( ~w4584 & w4778 ) | ( w4777 & w4778 ) ;
  assign w4780 = w4778 | w4779 ;
  assign w4781 = \pi087 ^ w4571 ;
  assign w4782 = ( ~w4578 & w4780 ) | ( ~w4578 & w4781 ) | ( w4780 & w4781 ) ;
  assign w4783 = w4781 | w4782 ;
  assign w4784 = \pi088 ^ w4565 ;
  assign w4785 = ( ~w4572 & w4783 ) | ( ~w4572 & w4784 ) | ( w4783 & w4784 ) ;
  assign w4786 = w4784 | w4785 ;
  assign w4787 = \pi089 ^ w4559 ;
  assign w4788 = ( ~w4566 & w4786 ) | ( ~w4566 & w4787 ) | ( w4786 & w4787 ) ;
  assign w4789 = w4787 | w4788 ;
  assign w4790 = \pi090 ^ w4553 ;
  assign w4791 = ( ~w4560 & w4789 ) | ( ~w4560 & w4790 ) | ( w4789 & w4790 ) ;
  assign w4792 = w4790 | w4791 ;
  assign w4793 = \pi091 ^ w4547 ;
  assign w4794 = ( ~w4554 & w4792 ) | ( ~w4554 & w4793 ) | ( w4792 & w4793 ) ;
  assign w4795 = w4793 | w4794 ;
  assign w4796 = \pi092 ^ w4541 ;
  assign w4797 = ( ~w4548 & w4795 ) | ( ~w4548 & w4796 ) | ( w4795 & w4796 ) ;
  assign w4798 = w4796 | w4797 ;
  assign w4799 = w4277 & w4536 ;
  assign w4800 = ~w4278 & w4528 ;
  assign w4801 = w4529 ^ w4800 ;
  assign w4802 = ~w4536 & w4801 ;
  assign w4803 = w4799 | w4802 ;
  assign w4804 = ~\pi093 & w4803 ;
  assign w4805 = ( \pi093 & ~w4799 ) | ( \pi093 & w4802 ) | ( ~w4799 & w4802 ) ;
  assign w4806 = ~w4802 & w4805 ;
  assign w4807 = \pi094 | \pi095 ;
  assign w4808 = w155 | w4807 ;
  assign w4809 = ( ~w155 & w170 ) | ( ~w155 & w179 ) | ( w170 & w179 ) ;
  assign w4810 = w4808 | w4809 ;
  assign w4811 = w4804 | w4806 ;
  assign w4812 = ( ~w4542 & w4798 ) | ( ~w4542 & w4811 ) | ( w4798 & w4811 ) ;
  assign w4813 = ( w4810 & ~w4811 ) | ( w4810 & w4812 ) | ( ~w4811 & w4812 ) ;
  assign w4814 = w4811 | w4813 ;
  assign w4815 = ~w4535 & w4803 ;
  assign w4816 = w4814 & ~w4815 ;
  assign w4817 = ~w4548 & w4795 ;
  assign w4818 = w4796 ^ w4817 ;
  assign w4819 = ~w4816 & w4818 ;
  assign w4820 = ( w4541 & w4814 ) | ( w4541 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4821 = ~w4815 & w4820 ;
  assign w4822 = w4819 | w4821 ;
  assign w4823 = ( ~w4542 & w4798 ) | ( ~w4542 & w4816 ) | ( w4798 & w4816 ) ;
  assign w4824 = w4811 ^ w4823 ;
  assign w4825 = ~w4816 & w4824 ;
  assign w4826 = ( w4535 & ~w4803 ) | ( w4535 & w4814 ) | ( ~w4803 & w4814 ) ;
  assign w4827 = w4803 & w4826 ;
  assign w4828 = w4825 | w4827 ;
  assign w4829 = ~\pi093 & w4822 ;
  assign w4830 = ~w4554 & w4792 ;
  assign w4831 = w4793 ^ w4830 ;
  assign w4832 = ~w4816 & w4831 ;
  assign w4833 = ( w4547 & w4814 ) | ( w4547 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4834 = ~w4815 & w4833 ;
  assign w4835 = w4832 | w4834 ;
  assign w4836 = ~\pi092 & w4835 ;
  assign w4837 = ~w4560 & w4789 ;
  assign w4838 = w4790 ^ w4837 ;
  assign w4839 = ~w4816 & w4838 ;
  assign w4840 = ( w4553 & w4814 ) | ( w4553 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4841 = ~w4815 & w4840 ;
  assign w4842 = w4839 | w4841 ;
  assign w4843 = ~\pi091 & w4842 ;
  assign w4844 = ~w4566 & w4786 ;
  assign w4845 = w4787 ^ w4844 ;
  assign w4846 = ~w4816 & w4845 ;
  assign w4847 = ( w4559 & w4814 ) | ( w4559 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4848 = ~w4815 & w4847 ;
  assign w4849 = w4846 | w4848 ;
  assign w4850 = ~\pi090 & w4849 ;
  assign w4851 = ~w4572 & w4783 ;
  assign w4852 = w4784 ^ w4851 ;
  assign w4853 = ~w4816 & w4852 ;
  assign w4854 = ( w4565 & w4814 ) | ( w4565 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4855 = ~w4815 & w4854 ;
  assign w4856 = w4853 | w4855 ;
  assign w4857 = ~\pi089 & w4856 ;
  assign w4858 = ~w4578 & w4780 ;
  assign w4859 = w4781 ^ w4858 ;
  assign w4860 = ~w4816 & w4859 ;
  assign w4861 = ( w4571 & w4814 ) | ( w4571 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4862 = ~w4815 & w4861 ;
  assign w4863 = w4860 | w4862 ;
  assign w4864 = ~\pi088 & w4863 ;
  assign w4865 = ~w4584 & w4777 ;
  assign w4866 = w4778 ^ w4865 ;
  assign w4867 = ~w4816 & w4866 ;
  assign w4868 = ( w4577 & w4814 ) | ( w4577 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4869 = ~w4815 & w4868 ;
  assign w4870 = w4867 | w4869 ;
  assign w4871 = ~\pi087 & w4870 ;
  assign w4872 = ~w4590 & w4774 ;
  assign w4873 = w4775 ^ w4872 ;
  assign w4874 = ~w4816 & w4873 ;
  assign w4875 = ( w4583 & w4814 ) | ( w4583 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4876 = ~w4815 & w4875 ;
  assign w4877 = w4874 | w4876 ;
  assign w4878 = ~\pi086 & w4877 ;
  assign w4879 = ~w4596 & w4771 ;
  assign w4880 = w4772 ^ w4879 ;
  assign w4881 = ~w4816 & w4880 ;
  assign w4882 = ( w4589 & w4814 ) | ( w4589 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4883 = ~w4815 & w4882 ;
  assign w4884 = w4881 | w4883 ;
  assign w4885 = ~\pi085 & w4884 ;
  assign w4886 = ~w4602 & w4768 ;
  assign w4887 = w4769 ^ w4886 ;
  assign w4888 = ~w4816 & w4887 ;
  assign w4889 = ( w4595 & w4814 ) | ( w4595 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4890 = ~w4815 & w4889 ;
  assign w4891 = w4888 | w4890 ;
  assign w4892 = ~\pi084 & w4891 ;
  assign w4893 = ~w4608 & w4765 ;
  assign w4894 = w4766 ^ w4893 ;
  assign w4895 = ~w4816 & w4894 ;
  assign w4896 = ( w4601 & w4814 ) | ( w4601 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4897 = ~w4815 & w4896 ;
  assign w4898 = w4895 | w4897 ;
  assign w4899 = ~\pi083 & w4898 ;
  assign w4900 = ~w4614 & w4762 ;
  assign w4901 = w4763 ^ w4900 ;
  assign w4902 = ~w4816 & w4901 ;
  assign w4903 = ( w4607 & w4814 ) | ( w4607 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4904 = ~w4815 & w4903 ;
  assign w4905 = w4902 | w4904 ;
  assign w4906 = ~\pi082 & w4905 ;
  assign w4907 = ~w4620 & w4759 ;
  assign w4908 = w4760 ^ w4907 ;
  assign w4909 = ~w4816 & w4908 ;
  assign w4910 = ( w4613 & w4814 ) | ( w4613 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4911 = ~w4815 & w4910 ;
  assign w4912 = w4909 | w4911 ;
  assign w4913 = ~\pi081 & w4912 ;
  assign w4914 = ~w4626 & w4756 ;
  assign w4915 = w4757 ^ w4914 ;
  assign w4916 = ~w4816 & w4915 ;
  assign w4917 = ( w4619 & w4814 ) | ( w4619 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4918 = ~w4815 & w4917 ;
  assign w4919 = w4916 | w4918 ;
  assign w4920 = ~\pi080 & w4919 ;
  assign w4921 = ~w4632 & w4753 ;
  assign w4922 = w4754 ^ w4921 ;
  assign w4923 = ~w4816 & w4922 ;
  assign w4924 = ( w4625 & w4814 ) | ( w4625 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4925 = ~w4815 & w4924 ;
  assign w4926 = w4923 | w4925 ;
  assign w4927 = ~\pi079 & w4926 ;
  assign w4928 = ~w4638 & w4750 ;
  assign w4929 = w4751 ^ w4928 ;
  assign w4930 = ~w4816 & w4929 ;
  assign w4931 = ( w4631 & w4814 ) | ( w4631 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4932 = ~w4815 & w4931 ;
  assign w4933 = w4930 | w4932 ;
  assign w4934 = ~\pi078 & w4933 ;
  assign w4935 = ~w4644 & w4747 ;
  assign w4936 = w4748 ^ w4935 ;
  assign w4937 = ~w4816 & w4936 ;
  assign w4938 = ( w4637 & w4814 ) | ( w4637 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4939 = ~w4815 & w4938 ;
  assign w4940 = w4937 | w4939 ;
  assign w4941 = ~\pi077 & w4940 ;
  assign w4942 = ~w4650 & w4744 ;
  assign w4943 = w4745 ^ w4942 ;
  assign w4944 = ~w4816 & w4943 ;
  assign w4945 = ( w4643 & w4814 ) | ( w4643 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4946 = ~w4815 & w4945 ;
  assign w4947 = w4944 | w4946 ;
  assign w4948 = ~\pi076 & w4947 ;
  assign w4949 = ~w4656 & w4741 ;
  assign w4950 = w4742 ^ w4949 ;
  assign w4951 = ~w4816 & w4950 ;
  assign w4952 = ( w4649 & w4814 ) | ( w4649 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4953 = ~w4815 & w4952 ;
  assign w4954 = w4951 | w4953 ;
  assign w4955 = ~\pi075 & w4954 ;
  assign w4956 = ~w4662 & w4738 ;
  assign w4957 = w4739 ^ w4956 ;
  assign w4958 = ~w4816 & w4957 ;
  assign w4959 = ( w4655 & w4814 ) | ( w4655 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4960 = ~w4815 & w4959 ;
  assign w4961 = w4958 | w4960 ;
  assign w4962 = ~\pi074 & w4961 ;
  assign w4963 = ~w4668 & w4735 ;
  assign w4964 = w4736 ^ w4963 ;
  assign w4965 = ~w4816 & w4964 ;
  assign w4966 = ( w4661 & w4814 ) | ( w4661 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4967 = ~w4815 & w4966 ;
  assign w4968 = w4965 | w4967 ;
  assign w4969 = ~\pi073 & w4968 ;
  assign w4970 = ~w4674 & w4732 ;
  assign w4971 = w4733 ^ w4970 ;
  assign w4972 = ~w4816 & w4971 ;
  assign w4973 = ( w4667 & w4814 ) | ( w4667 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4974 = ~w4815 & w4973 ;
  assign w4975 = w4972 | w4974 ;
  assign w4976 = ~\pi072 & w4975 ;
  assign w4977 = ~w4680 & w4729 ;
  assign w4978 = w4730 ^ w4977 ;
  assign w4979 = ~w4816 & w4978 ;
  assign w4980 = ( w4673 & w4814 ) | ( w4673 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4981 = ~w4815 & w4980 ;
  assign w4982 = w4979 | w4981 ;
  assign w4983 = ~\pi071 & w4982 ;
  assign w4984 = ~w4686 & w4726 ;
  assign w4985 = w4727 ^ w4984 ;
  assign w4986 = ~w4816 & w4985 ;
  assign w4987 = ( w4679 & w4814 ) | ( w4679 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4988 = ~w4815 & w4987 ;
  assign w4989 = w4986 | w4988 ;
  assign w4990 = ~\pi070 & w4989 ;
  assign w4991 = ~w4693 & w4723 ;
  assign w4992 = w4724 ^ w4991 ;
  assign w4993 = ~w4816 & w4992 ;
  assign w4994 = ( w4685 & w4814 ) | ( w4685 & w4815 ) | ( w4814 & w4815 ) ;
  assign w4995 = ~w4815 & w4994 ;
  assign w4996 = w4993 | w4995 ;
  assign w4997 = ~\pi069 & w4996 ;
  assign w4998 = ~w4701 & w4720 ;
  assign w4999 = w4721 ^ w4998 ;
  assign w5000 = ~w4816 & w4999 ;
  assign w5001 = ( w4692 & w4814 ) | ( w4692 & w4815 ) | ( w4814 & w4815 ) ;
  assign w5002 = ~w4815 & w5001 ;
  assign w5003 = w5000 | w5002 ;
  assign w5004 = ~\pi068 & w5003 ;
  assign w5005 = w4717 ^ w4719 ;
  assign w5006 = ~w4816 & w5005 ;
  assign w5007 = ( w4700 & w4814 ) | ( w4700 & w4815 ) | ( w4814 & w4815 ) ;
  assign w5008 = ~w4815 & w5007 ;
  assign w5009 = w5006 | w5008 ;
  assign w5010 = ~\pi067 & w5009 ;
  assign w5011 = w4714 ^ w4718 ;
  assign w5012 = \pi065 ^ w5011 ;
  assign w5013 = ~w4816 & w5012 ;
  assign w5014 = ( w4709 & w4713 ) | ( w4709 & ~w4815 ) | ( w4713 & ~w4815 ) ;
  assign w5015 = w4815 & w5014 ;
  assign w5016 = ( ~w4814 & w5014 ) | ( ~w4814 & w5015 ) | ( w5014 & w5015 ) ;
  assign w5017 = ( w5013 & w5014 ) | ( w5013 & ~w5016 ) | ( w5014 & ~w5016 ) ;
  assign w5018 = ~\pi066 & w5017 ;
  assign w5019 = w4814 | w4815 ;
  assign w5020 = ( w5013 & w5014 ) | ( w5013 & w5019 ) | ( w5014 & w5019 ) ;
  assign w5021 = ( ~w4815 & w5013 ) | ( ~w4815 & w5020 ) | ( w5013 & w5020 ) ;
  assign w5022 = \pi066 ^ w5021 ;
  assign w5023 = \pi064 & ~w4816 ;
  assign w5024 = \pi034 ^ w5023 ;
  assign w5025 = ( ~\pi033 & \pi064 ) | ( ~\pi033 & w5022 ) | ( \pi064 & w5022 ) ;
  assign w5026 = ( \pi065 & ~w5024 ) | ( \pi065 & w5025 ) | ( ~w5024 & w5025 ) ;
  assign w5027 = w5022 | w5026 ;
  assign w5028 = \pi067 ^ w5009 ;
  assign w5029 = ( ~w5018 & w5027 ) | ( ~w5018 & w5028 ) | ( w5027 & w5028 ) ;
  assign w5030 = w5028 | w5029 ;
  assign w5031 = \pi068 ^ w5003 ;
  assign w5032 = ( ~w5010 & w5030 ) | ( ~w5010 & w5031 ) | ( w5030 & w5031 ) ;
  assign w5033 = w5031 | w5032 ;
  assign w5034 = \pi069 ^ w4996 ;
  assign w5035 = ( ~w5004 & w5033 ) | ( ~w5004 & w5034 ) | ( w5033 & w5034 ) ;
  assign w5036 = w5034 | w5035 ;
  assign w5037 = \pi070 ^ w4989 ;
  assign w5038 = ( ~w4997 & w5036 ) | ( ~w4997 & w5037 ) | ( w5036 & w5037 ) ;
  assign w5039 = w5037 | w5038 ;
  assign w5040 = \pi071 ^ w4982 ;
  assign w5041 = ( ~w4990 & w5039 ) | ( ~w4990 & w5040 ) | ( w5039 & w5040 ) ;
  assign w5042 = w5040 | w5041 ;
  assign w5043 = \pi072 ^ w4975 ;
  assign w5044 = ( ~w4983 & w5042 ) | ( ~w4983 & w5043 ) | ( w5042 & w5043 ) ;
  assign w5045 = w5043 | w5044 ;
  assign w5046 = \pi073 ^ w4968 ;
  assign w5047 = ( ~w4976 & w5045 ) | ( ~w4976 & w5046 ) | ( w5045 & w5046 ) ;
  assign w5048 = w5046 | w5047 ;
  assign w5049 = \pi074 ^ w4961 ;
  assign w5050 = ( ~w4969 & w5048 ) | ( ~w4969 & w5049 ) | ( w5048 & w5049 ) ;
  assign w5051 = w5049 | w5050 ;
  assign w5052 = \pi075 ^ w4954 ;
  assign w5053 = ( ~w4962 & w5051 ) | ( ~w4962 & w5052 ) | ( w5051 & w5052 ) ;
  assign w5054 = w5052 | w5053 ;
  assign w5055 = \pi076 ^ w4947 ;
  assign w5056 = ( ~w4955 & w5054 ) | ( ~w4955 & w5055 ) | ( w5054 & w5055 ) ;
  assign w5057 = w5055 | w5056 ;
  assign w5058 = \pi077 ^ w4940 ;
  assign w5059 = ( ~w4948 & w5057 ) | ( ~w4948 & w5058 ) | ( w5057 & w5058 ) ;
  assign w5060 = w5058 | w5059 ;
  assign w5061 = \pi078 ^ w4933 ;
  assign w5062 = ( ~w4941 & w5060 ) | ( ~w4941 & w5061 ) | ( w5060 & w5061 ) ;
  assign w5063 = w5061 | w5062 ;
  assign w5064 = \pi079 ^ w4926 ;
  assign w5065 = ( ~w4934 & w5063 ) | ( ~w4934 & w5064 ) | ( w5063 & w5064 ) ;
  assign w5066 = w5064 | w5065 ;
  assign w5067 = \pi080 ^ w4919 ;
  assign w5068 = ( ~w4927 & w5066 ) | ( ~w4927 & w5067 ) | ( w5066 & w5067 ) ;
  assign w5069 = w5067 | w5068 ;
  assign w5070 = \pi081 ^ w4912 ;
  assign w5071 = ( ~w4920 & w5069 ) | ( ~w4920 & w5070 ) | ( w5069 & w5070 ) ;
  assign w5072 = w5070 | w5071 ;
  assign w5073 = \pi082 ^ w4905 ;
  assign w5074 = ( ~w4913 & w5072 ) | ( ~w4913 & w5073 ) | ( w5072 & w5073 ) ;
  assign w5075 = w5073 | w5074 ;
  assign w5076 = \pi083 ^ w4898 ;
  assign w5077 = ( ~w4906 & w5075 ) | ( ~w4906 & w5076 ) | ( w5075 & w5076 ) ;
  assign w5078 = w5076 | w5077 ;
  assign w5079 = \pi084 ^ w4891 ;
  assign w5080 = ( ~w4899 & w5078 ) | ( ~w4899 & w5079 ) | ( w5078 & w5079 ) ;
  assign w5081 = w5079 | w5080 ;
  assign w5082 = \pi085 ^ w4884 ;
  assign w5083 = ( ~w4892 & w5081 ) | ( ~w4892 & w5082 ) | ( w5081 & w5082 ) ;
  assign w5084 = w5082 | w5083 ;
  assign w5085 = \pi086 ^ w4877 ;
  assign w5086 = ( ~w4885 & w5084 ) | ( ~w4885 & w5085 ) | ( w5084 & w5085 ) ;
  assign w5087 = w5085 | w5086 ;
  assign w5088 = \pi087 ^ w4870 ;
  assign w5089 = ( ~w4878 & w5087 ) | ( ~w4878 & w5088 ) | ( w5087 & w5088 ) ;
  assign w5090 = w5088 | w5089 ;
  assign w5091 = \pi088 ^ w4863 ;
  assign w5092 = ( ~w4871 & w5090 ) | ( ~w4871 & w5091 ) | ( w5090 & w5091 ) ;
  assign w5093 = w5091 | w5092 ;
  assign w5094 = \pi089 ^ w4856 ;
  assign w5095 = ( ~w4864 & w5093 ) | ( ~w4864 & w5094 ) | ( w5093 & w5094 ) ;
  assign w5096 = w5094 | w5095 ;
  assign w5097 = \pi090 ^ w4849 ;
  assign w5098 = ( ~w4857 & w5096 ) | ( ~w4857 & w5097 ) | ( w5096 & w5097 ) ;
  assign w5099 = w5097 | w5098 ;
  assign w5100 = \pi091 ^ w4842 ;
  assign w5101 = ( ~w4850 & w5099 ) | ( ~w4850 & w5100 ) | ( w5099 & w5100 ) ;
  assign w5102 = w5100 | w5101 ;
  assign w5103 = \pi092 ^ w4835 ;
  assign w5104 = ( ~w4843 & w5102 ) | ( ~w4843 & w5103 ) | ( w5102 & w5103 ) ;
  assign w5105 = w5103 | w5104 ;
  assign w5106 = \pi093 ^ w4822 ;
  assign w5107 = ( ~w4836 & w5105 ) | ( ~w4836 & w5106 ) | ( w5105 & w5106 ) ;
  assign w5108 = w5106 | w5107 ;
  assign w5109 = \pi094 ^ w4828 ;
  assign w5110 = w4829 & ~w5109 ;
  assign w5111 = ( w5108 & w5109 ) | ( w5108 & ~w5110 ) | ( w5109 & ~w5110 ) ;
  assign w5112 = ~\pi094 & w4828 ;
  assign w5113 = w5111 & ~w5112 ;
  assign w5114 = \pi095 | \pi096 ;
  assign w5115 = w451 | w5114 ;
  assign w5116 = ( w281 & w448 ) | ( w281 & ~w451 ) | ( w448 & ~w451 ) ;
  assign w5117 = w5115 | w5116 ;
  assign w5118 = w5113 | w5117 ;
  assign w5119 = w4822 & w5118 ;
  assign w5120 = ~w4836 & w5105 ;
  assign w5121 = w5106 ^ w5120 ;
  assign w5122 = ~w5118 & w5121 ;
  assign w5123 = w5119 | w5122 ;
  assign w5124 = w4828 & w5118 ;
  assign w5125 = ~w4829 & w5108 ;
  assign w5126 = w5109 ^ w5125 ;
  assign w5127 = ~w5118 & w5126 ;
  assign w5128 = w5124 | w5127 ;
  assign w5129 = ~\pi094 & w5123 ;
  assign w5130 = w4835 & w5118 ;
  assign w5131 = ~w4843 & w5102 ;
  assign w5132 = w5103 ^ w5131 ;
  assign w5133 = ~w5118 & w5132 ;
  assign w5134 = w5130 | w5133 ;
  assign w5135 = ~\pi093 & w5134 ;
  assign w5136 = w4842 & w5118 ;
  assign w5137 = ~w4850 & w5099 ;
  assign w5138 = w5100 ^ w5137 ;
  assign w5139 = ~w5118 & w5138 ;
  assign w5140 = w5136 | w5139 ;
  assign w5141 = ~\pi092 & w5140 ;
  assign w5142 = w4849 & w5118 ;
  assign w5143 = ~w4857 & w5096 ;
  assign w5144 = w5097 ^ w5143 ;
  assign w5145 = ~w5118 & w5144 ;
  assign w5146 = w5142 | w5145 ;
  assign w5147 = ~\pi091 & w5146 ;
  assign w5148 = w4856 & w5118 ;
  assign w5149 = ~w4864 & w5093 ;
  assign w5150 = w5094 ^ w5149 ;
  assign w5151 = ~w5118 & w5150 ;
  assign w5152 = w5148 | w5151 ;
  assign w5153 = ~\pi090 & w5152 ;
  assign w5154 = w4863 & w5118 ;
  assign w5155 = ~w4871 & w5090 ;
  assign w5156 = w5091 ^ w5155 ;
  assign w5157 = ~w5118 & w5156 ;
  assign w5158 = w5154 | w5157 ;
  assign w5159 = ~\pi089 & w5158 ;
  assign w5160 = w4870 & w5118 ;
  assign w5161 = ~w4878 & w5087 ;
  assign w5162 = w5088 ^ w5161 ;
  assign w5163 = ~w5118 & w5162 ;
  assign w5164 = w5160 | w5163 ;
  assign w5165 = ~\pi088 & w5164 ;
  assign w5166 = w4877 & w5118 ;
  assign w5167 = ~w4885 & w5084 ;
  assign w5168 = w5085 ^ w5167 ;
  assign w5169 = ~w5118 & w5168 ;
  assign w5170 = w5166 | w5169 ;
  assign w5171 = ~\pi087 & w5170 ;
  assign w5172 = w4884 & w5118 ;
  assign w5173 = ~w4892 & w5081 ;
  assign w5174 = w5082 ^ w5173 ;
  assign w5175 = ~w5118 & w5174 ;
  assign w5176 = w5172 | w5175 ;
  assign w5177 = ~\pi086 & w5176 ;
  assign w5178 = w4891 & w5118 ;
  assign w5179 = ~w4899 & w5078 ;
  assign w5180 = w5079 ^ w5179 ;
  assign w5181 = ~w5118 & w5180 ;
  assign w5182 = w5178 | w5181 ;
  assign w5183 = ~\pi085 & w5182 ;
  assign w5184 = w4898 & w5118 ;
  assign w5185 = ~w4906 & w5075 ;
  assign w5186 = w5076 ^ w5185 ;
  assign w5187 = ~w5118 & w5186 ;
  assign w5188 = w5184 | w5187 ;
  assign w5189 = ~\pi084 & w5188 ;
  assign w5190 = w4905 & w5118 ;
  assign w5191 = ~w4913 & w5072 ;
  assign w5192 = w5073 ^ w5191 ;
  assign w5193 = ~w5118 & w5192 ;
  assign w5194 = w5190 | w5193 ;
  assign w5195 = ~\pi083 & w5194 ;
  assign w5196 = w4912 & w5118 ;
  assign w5197 = ~w4920 & w5069 ;
  assign w5198 = w5070 ^ w5197 ;
  assign w5199 = ~w5118 & w5198 ;
  assign w5200 = w5196 | w5199 ;
  assign w5201 = ~\pi082 & w5200 ;
  assign w5202 = w4919 & w5118 ;
  assign w5203 = ~w4927 & w5066 ;
  assign w5204 = w5067 ^ w5203 ;
  assign w5205 = ~w5118 & w5204 ;
  assign w5206 = w5202 | w5205 ;
  assign w5207 = ~\pi081 & w5206 ;
  assign w5208 = w4926 & w5118 ;
  assign w5209 = ~w4934 & w5063 ;
  assign w5210 = w5064 ^ w5209 ;
  assign w5211 = ~w5118 & w5210 ;
  assign w5212 = w5208 | w5211 ;
  assign w5213 = ~\pi080 & w5212 ;
  assign w5214 = w4933 & w5118 ;
  assign w5215 = ~w4941 & w5060 ;
  assign w5216 = w5061 ^ w5215 ;
  assign w5217 = ~w5118 & w5216 ;
  assign w5218 = w5214 | w5217 ;
  assign w5219 = ~\pi079 & w5218 ;
  assign w5220 = w4940 & w5118 ;
  assign w5221 = ~w4948 & w5057 ;
  assign w5222 = w5058 ^ w5221 ;
  assign w5223 = ~w5118 & w5222 ;
  assign w5224 = w5220 | w5223 ;
  assign w5225 = ~\pi078 & w5224 ;
  assign w5226 = w4947 & w5118 ;
  assign w5227 = ~w4955 & w5054 ;
  assign w5228 = w5055 ^ w5227 ;
  assign w5229 = ~w5118 & w5228 ;
  assign w5230 = w5226 | w5229 ;
  assign w5231 = ~\pi077 & w5230 ;
  assign w5232 = w4954 & w5118 ;
  assign w5233 = ~w4962 & w5051 ;
  assign w5234 = w5052 ^ w5233 ;
  assign w5235 = ~w5118 & w5234 ;
  assign w5236 = w5232 | w5235 ;
  assign w5237 = ~\pi076 & w5236 ;
  assign w5238 = w4961 & w5118 ;
  assign w5239 = ~w4969 & w5048 ;
  assign w5240 = w5049 ^ w5239 ;
  assign w5241 = ~w5118 & w5240 ;
  assign w5242 = w5238 | w5241 ;
  assign w5243 = ~\pi075 & w5242 ;
  assign w5244 = w4968 & w5118 ;
  assign w5245 = ~w4976 & w5045 ;
  assign w5246 = w5046 ^ w5245 ;
  assign w5247 = ~w5118 & w5246 ;
  assign w5248 = w5244 | w5247 ;
  assign w5249 = ~\pi074 & w5248 ;
  assign w5250 = w4975 & w5118 ;
  assign w5251 = ~w4983 & w5042 ;
  assign w5252 = w5043 ^ w5251 ;
  assign w5253 = ~w5118 & w5252 ;
  assign w5254 = w5250 | w5253 ;
  assign w5255 = ~\pi073 & w5254 ;
  assign w5256 = w4982 & w5118 ;
  assign w5257 = ~w4990 & w5039 ;
  assign w5258 = w5040 ^ w5257 ;
  assign w5259 = ~w5118 & w5258 ;
  assign w5260 = w5256 | w5259 ;
  assign w5261 = ~\pi072 & w5260 ;
  assign w5262 = w4989 & w5118 ;
  assign w5263 = ~w4997 & w5036 ;
  assign w5264 = w5037 ^ w5263 ;
  assign w5265 = ~w5118 & w5264 ;
  assign w5266 = w5262 | w5265 ;
  assign w5267 = ~\pi071 & w5266 ;
  assign w5268 = w4996 & w5118 ;
  assign w5269 = ~w5004 & w5033 ;
  assign w5270 = w5034 ^ w5269 ;
  assign w5271 = ~w5118 & w5270 ;
  assign w5272 = w5268 | w5271 ;
  assign w5273 = ~\pi070 & w5272 ;
  assign w5274 = w5003 & w5118 ;
  assign w5275 = ~w5010 & w5030 ;
  assign w5276 = w5031 ^ w5275 ;
  assign w5277 = ~w5118 & w5276 ;
  assign w5278 = w5274 | w5277 ;
  assign w5279 = ~\pi069 & w5278 ;
  assign w5280 = w5009 & w5118 ;
  assign w5281 = ~w5018 & w5027 ;
  assign w5282 = w5028 ^ w5281 ;
  assign w5283 = ~w5118 & w5282 ;
  assign w5284 = w5280 | w5283 ;
  assign w5285 = ~\pi068 & w5284 ;
  assign w5286 = w5017 & w5118 ;
  assign w5287 = ~\pi033 & \pi064 ;
  assign w5288 = ( \pi065 & ~w5024 ) | ( \pi065 & w5287 ) | ( ~w5024 & w5287 ) ;
  assign w5289 = w5022 ^ w5288 ;
  assign w5290 = ( w5113 & w5117 ) | ( w5113 & w5289 ) | ( w5117 & w5289 ) ;
  assign w5291 = w5289 & ~w5290 ;
  assign w5292 = w5286 | w5291 ;
  assign w5293 = ~\pi067 & w5292 ;
  assign w5294 = \pi034 ^ \pi065 ;
  assign w5295 = \pi033 ^ w4816 ;
  assign w5296 = ( \pi064 & w5117 ) | ( \pi064 & w5295 ) | ( w5117 & w5295 ) ;
  assign w5297 = w5294 ^ w5296 ;
  assign w5298 = ~w5117 & w5297 ;
  assign w5299 = ~w5113 & w5298 ;
  assign w5300 = ( ~\pi064 & w4816 ) | ( ~\pi064 & w5118 ) | ( w4816 & w5118 ) ;
  assign w5301 = \pi034 ^ w5300 ;
  assign w5302 = w5118 & ~w5301 ;
  assign w5303 = w5299 | w5302 ;
  assign w5304 = ~\pi066 & w5303 ;
  assign w5305 = \pi064 & ~\pi095 ;
  assign w5306 = ~w155 & w5305 ;
  assign w5307 = ~w4809 & w5306 ;
  assign w5308 = ( \pi033 & w5113 ) | ( \pi033 & ~w5307 ) | ( w5113 & ~w5307 ) ;
  assign w5309 = \pi033 & w5308 ;
  assign w5310 = ( ~\pi033 & \pi064 ) | ( ~\pi033 & \pi095 ) | ( \pi064 & \pi095 ) ;
  assign w5311 = w281 | w451 ;
  assign w5312 = ( \pi095 & \pi096 ) | ( \pi095 & ~w281 ) | ( \pi096 & ~w281 ) ;
  assign w5313 = w5311 | w5312 ;
  assign w5314 = w5310 & ~w5313 ;
  assign w5315 = ~w448 & w5314 ;
  assign w5316 = ~w5113 & w5315 ;
  assign w5317 = w5309 | w5316 ;
  assign w5318 = ~\pi032 & \pi064 ;
  assign w5319 = \pi065 ^ w5317 ;
  assign w5320 = w5318 | w5319 ;
  assign w5321 = w5118 | w5299 ;
  assign w5322 = ( w5024 & w5299 ) | ( w5024 & w5321 ) | ( w5299 & w5321 ) ;
  assign w5323 = \pi066 ^ w5322 ;
  assign w5324 = ~\pi065 & w5317 ;
  assign w5325 = w5320 | w5324 ;
  assign w5326 = ( w5323 & ~w5324 ) | ( w5323 & w5325 ) | ( ~w5324 & w5325 ) ;
  assign w5327 = \pi067 ^ w5292 ;
  assign w5328 = ( ~w5304 & w5326 ) | ( ~w5304 & w5327 ) | ( w5326 & w5327 ) ;
  assign w5329 = w5327 | w5328 ;
  assign w5330 = \pi068 ^ w5284 ;
  assign w5331 = ( ~w5293 & w5329 ) | ( ~w5293 & w5330 ) | ( w5329 & w5330 ) ;
  assign w5332 = w5330 | w5331 ;
  assign w5333 = \pi069 ^ w5278 ;
  assign w5334 = ( ~w5285 & w5332 ) | ( ~w5285 & w5333 ) | ( w5332 & w5333 ) ;
  assign w5335 = w5333 | w5334 ;
  assign w5336 = \pi070 ^ w5272 ;
  assign w5337 = ( ~w5279 & w5335 ) | ( ~w5279 & w5336 ) | ( w5335 & w5336 ) ;
  assign w5338 = w5336 | w5337 ;
  assign w5339 = \pi071 ^ w5266 ;
  assign w5340 = ( ~w5273 & w5338 ) | ( ~w5273 & w5339 ) | ( w5338 & w5339 ) ;
  assign w5341 = w5339 | w5340 ;
  assign w5342 = \pi072 ^ w5260 ;
  assign w5343 = ( ~w5267 & w5341 ) | ( ~w5267 & w5342 ) | ( w5341 & w5342 ) ;
  assign w5344 = w5342 | w5343 ;
  assign w5345 = \pi073 ^ w5254 ;
  assign w5346 = ( ~w5261 & w5344 ) | ( ~w5261 & w5345 ) | ( w5344 & w5345 ) ;
  assign w5347 = w5345 | w5346 ;
  assign w5348 = \pi074 ^ w5248 ;
  assign w5349 = ( ~w5255 & w5347 ) | ( ~w5255 & w5348 ) | ( w5347 & w5348 ) ;
  assign w5350 = w5348 | w5349 ;
  assign w5351 = \pi075 ^ w5242 ;
  assign w5352 = ( ~w5249 & w5350 ) | ( ~w5249 & w5351 ) | ( w5350 & w5351 ) ;
  assign w5353 = w5351 | w5352 ;
  assign w5354 = \pi076 ^ w5236 ;
  assign w5355 = ( ~w5243 & w5353 ) | ( ~w5243 & w5354 ) | ( w5353 & w5354 ) ;
  assign w5356 = w5354 | w5355 ;
  assign w5357 = \pi077 ^ w5230 ;
  assign w5358 = ( ~w5237 & w5356 ) | ( ~w5237 & w5357 ) | ( w5356 & w5357 ) ;
  assign w5359 = w5357 | w5358 ;
  assign w5360 = \pi078 ^ w5224 ;
  assign w5361 = ( ~w5231 & w5359 ) | ( ~w5231 & w5360 ) | ( w5359 & w5360 ) ;
  assign w5362 = w5360 | w5361 ;
  assign w5363 = \pi079 ^ w5218 ;
  assign w5364 = ( ~w5225 & w5362 ) | ( ~w5225 & w5363 ) | ( w5362 & w5363 ) ;
  assign w5365 = w5363 | w5364 ;
  assign w5366 = \pi080 ^ w5212 ;
  assign w5367 = ( ~w5219 & w5365 ) | ( ~w5219 & w5366 ) | ( w5365 & w5366 ) ;
  assign w5368 = w5366 | w5367 ;
  assign w5369 = \pi081 ^ w5206 ;
  assign w5370 = ( ~w5213 & w5368 ) | ( ~w5213 & w5369 ) | ( w5368 & w5369 ) ;
  assign w5371 = w5369 | w5370 ;
  assign w5372 = \pi082 ^ w5200 ;
  assign w5373 = ( ~w5207 & w5371 ) | ( ~w5207 & w5372 ) | ( w5371 & w5372 ) ;
  assign w5374 = w5372 | w5373 ;
  assign w5375 = \pi083 ^ w5194 ;
  assign w5376 = ( ~w5201 & w5374 ) | ( ~w5201 & w5375 ) | ( w5374 & w5375 ) ;
  assign w5377 = w5375 | w5376 ;
  assign w5378 = \pi084 ^ w5188 ;
  assign w5379 = ( ~w5195 & w5377 ) | ( ~w5195 & w5378 ) | ( w5377 & w5378 ) ;
  assign w5380 = w5378 | w5379 ;
  assign w5381 = \pi085 ^ w5182 ;
  assign w5382 = ( ~w5189 & w5380 ) | ( ~w5189 & w5381 ) | ( w5380 & w5381 ) ;
  assign w5383 = w5381 | w5382 ;
  assign w5384 = \pi086 ^ w5176 ;
  assign w5385 = ( ~w5183 & w5383 ) | ( ~w5183 & w5384 ) | ( w5383 & w5384 ) ;
  assign w5386 = w5384 | w5385 ;
  assign w5387 = \pi087 ^ w5170 ;
  assign w5388 = ( ~w5177 & w5386 ) | ( ~w5177 & w5387 ) | ( w5386 & w5387 ) ;
  assign w5389 = w5387 | w5388 ;
  assign w5390 = \pi088 ^ w5164 ;
  assign w5391 = ( ~w5171 & w5389 ) | ( ~w5171 & w5390 ) | ( w5389 & w5390 ) ;
  assign w5392 = w5390 | w5391 ;
  assign w5393 = \pi089 ^ w5158 ;
  assign w5394 = ( ~w5165 & w5392 ) | ( ~w5165 & w5393 ) | ( w5392 & w5393 ) ;
  assign w5395 = w5393 | w5394 ;
  assign w5396 = \pi090 ^ w5152 ;
  assign w5397 = ( ~w5159 & w5395 ) | ( ~w5159 & w5396 ) | ( w5395 & w5396 ) ;
  assign w5398 = w5396 | w5397 ;
  assign w5399 = \pi091 ^ w5146 ;
  assign w5400 = ( ~w5153 & w5398 ) | ( ~w5153 & w5399 ) | ( w5398 & w5399 ) ;
  assign w5401 = w5399 | w5400 ;
  assign w5402 = \pi092 ^ w5140 ;
  assign w5403 = ( ~w5147 & w5401 ) | ( ~w5147 & w5402 ) | ( w5401 & w5402 ) ;
  assign w5404 = w5402 | w5403 ;
  assign w5405 = \pi093 ^ w5134 ;
  assign w5406 = ( ~w5141 & w5404 ) | ( ~w5141 & w5405 ) | ( w5404 & w5405 ) ;
  assign w5407 = w5405 | w5406 ;
  assign w5408 = \pi094 ^ w5123 ;
  assign w5409 = ( ~w5135 & w5407 ) | ( ~w5135 & w5408 ) | ( w5407 & w5408 ) ;
  assign w5410 = w5408 | w5409 ;
  assign w5411 = \pi095 ^ w5128 ;
  assign w5412 = w5129 & ~w5411 ;
  assign w5413 = ( w5410 & w5411 ) | ( w5410 & ~w5412 ) | ( w5411 & ~w5412 ) ;
  assign w5414 = ~\pi095 & w5128 ;
  assign w5415 = w5413 & ~w5414 ;
  assign w5416 = w298 | w5415 ;
  assign w5417 = w5123 & w5416 ;
  assign w5418 = ~w5135 & w5407 ;
  assign w5419 = w5408 ^ w5418 ;
  assign w5420 = ~w5416 & w5419 ;
  assign w5421 = w5417 | w5420 ;
  assign w5422 = ~\pi095 & w5421 ;
  assign w5423 = w5134 & w5416 ;
  assign w5424 = ~w5141 & w5404 ;
  assign w5425 = w5405 ^ w5424 ;
  assign w5426 = ~w5416 & w5425 ;
  assign w5427 = w5423 | w5426 ;
  assign w5428 = ~\pi094 & w5427 ;
  assign w5429 = w5140 & w5416 ;
  assign w5430 = ~w5147 & w5401 ;
  assign w5431 = w5402 ^ w5430 ;
  assign w5432 = ~w5416 & w5431 ;
  assign w5433 = w5429 | w5432 ;
  assign w5434 = ~\pi093 & w5433 ;
  assign w5435 = w5146 & w5416 ;
  assign w5436 = ~w5153 & w5398 ;
  assign w5437 = w5399 ^ w5436 ;
  assign w5438 = ~w5416 & w5437 ;
  assign w5439 = w5435 | w5438 ;
  assign w5440 = ~\pi092 & w5439 ;
  assign w5441 = w5152 & w5416 ;
  assign w5442 = ~w5159 & w5395 ;
  assign w5443 = w5396 ^ w5442 ;
  assign w5444 = ~w5416 & w5443 ;
  assign w5445 = w5441 | w5444 ;
  assign w5446 = ~\pi091 & w5445 ;
  assign w5447 = w5158 & w5416 ;
  assign w5448 = ~w5165 & w5392 ;
  assign w5449 = w5393 ^ w5448 ;
  assign w5450 = ~w5416 & w5449 ;
  assign w5451 = w5447 | w5450 ;
  assign w5452 = ~\pi090 & w5451 ;
  assign w5453 = w5164 & w5416 ;
  assign w5454 = ~w5171 & w5389 ;
  assign w5455 = w5390 ^ w5454 ;
  assign w5456 = ~w5416 & w5455 ;
  assign w5457 = w5453 | w5456 ;
  assign w5458 = ~\pi089 & w5457 ;
  assign w5459 = w5170 & w5416 ;
  assign w5460 = ~w5177 & w5386 ;
  assign w5461 = w5387 ^ w5460 ;
  assign w5462 = ~w5416 & w5461 ;
  assign w5463 = w5459 | w5462 ;
  assign w5464 = ~\pi088 & w5463 ;
  assign w5465 = w5176 & w5416 ;
  assign w5466 = ~w5183 & w5383 ;
  assign w5467 = w5384 ^ w5466 ;
  assign w5468 = ~w5416 & w5467 ;
  assign w5469 = w5465 | w5468 ;
  assign w5470 = ~\pi087 & w5469 ;
  assign w5471 = w5182 & w5416 ;
  assign w5472 = ~w5189 & w5380 ;
  assign w5473 = w5381 ^ w5472 ;
  assign w5474 = ~w5416 & w5473 ;
  assign w5475 = w5471 | w5474 ;
  assign w5476 = ~\pi086 & w5475 ;
  assign w5477 = w5188 & w5416 ;
  assign w5478 = ~w5195 & w5377 ;
  assign w5479 = w5378 ^ w5478 ;
  assign w5480 = ~w5416 & w5479 ;
  assign w5481 = w5477 | w5480 ;
  assign w5482 = ~\pi085 & w5481 ;
  assign w5483 = w5194 & w5416 ;
  assign w5484 = ~w5201 & w5374 ;
  assign w5485 = w5375 ^ w5484 ;
  assign w5486 = ~w5416 & w5485 ;
  assign w5487 = w5483 | w5486 ;
  assign w5488 = ~\pi084 & w5487 ;
  assign w5489 = w5200 & w5416 ;
  assign w5490 = ~w5207 & w5371 ;
  assign w5491 = w5372 ^ w5490 ;
  assign w5492 = ~w5416 & w5491 ;
  assign w5493 = w5489 | w5492 ;
  assign w5494 = ~\pi083 & w5493 ;
  assign w5495 = w5206 & w5416 ;
  assign w5496 = ~w5213 & w5368 ;
  assign w5497 = w5369 ^ w5496 ;
  assign w5498 = ~w5416 & w5497 ;
  assign w5499 = w5495 | w5498 ;
  assign w5500 = ~\pi082 & w5499 ;
  assign w5501 = w5212 & w5416 ;
  assign w5502 = ~w5219 & w5365 ;
  assign w5503 = w5366 ^ w5502 ;
  assign w5504 = ~w5416 & w5503 ;
  assign w5505 = w5501 | w5504 ;
  assign w5506 = ~\pi081 & w5505 ;
  assign w5507 = w5218 & w5416 ;
  assign w5508 = ~w5225 & w5362 ;
  assign w5509 = w5363 ^ w5508 ;
  assign w5510 = ~w5416 & w5509 ;
  assign w5511 = w5507 | w5510 ;
  assign w5512 = ~\pi080 & w5511 ;
  assign w5513 = w5224 & w5416 ;
  assign w5514 = ~w5231 & w5359 ;
  assign w5515 = w5360 ^ w5514 ;
  assign w5516 = ~w5416 & w5515 ;
  assign w5517 = w5513 | w5516 ;
  assign w5518 = ~\pi079 & w5517 ;
  assign w5519 = w5230 & w5416 ;
  assign w5520 = ~w5237 & w5356 ;
  assign w5521 = w5357 ^ w5520 ;
  assign w5522 = ~w5416 & w5521 ;
  assign w5523 = w5519 | w5522 ;
  assign w5524 = ~\pi078 & w5523 ;
  assign w5525 = w5236 & w5416 ;
  assign w5526 = ~w5243 & w5353 ;
  assign w5527 = w5354 ^ w5526 ;
  assign w5528 = ~w5416 & w5527 ;
  assign w5529 = w5525 | w5528 ;
  assign w5530 = ~\pi077 & w5529 ;
  assign w5531 = w5242 & w5416 ;
  assign w5532 = ~w5249 & w5350 ;
  assign w5533 = w5351 ^ w5532 ;
  assign w5534 = ~w5416 & w5533 ;
  assign w5535 = w5531 | w5534 ;
  assign w5536 = ~\pi076 & w5535 ;
  assign w5537 = w5248 & w5416 ;
  assign w5538 = ~w5255 & w5347 ;
  assign w5539 = w5348 ^ w5538 ;
  assign w5540 = ~w5416 & w5539 ;
  assign w5541 = w5537 | w5540 ;
  assign w5542 = ~\pi075 & w5541 ;
  assign w5543 = w5254 & w5416 ;
  assign w5544 = ~w5261 & w5344 ;
  assign w5545 = w5345 ^ w5544 ;
  assign w5546 = ~w5416 & w5545 ;
  assign w5547 = w5543 | w5546 ;
  assign w5548 = ~\pi074 & w5547 ;
  assign w5549 = w5260 & w5416 ;
  assign w5550 = ~w5267 & w5341 ;
  assign w5551 = w5342 ^ w5550 ;
  assign w5552 = ~w5416 & w5551 ;
  assign w5553 = w5549 | w5552 ;
  assign w5554 = ~\pi073 & w5553 ;
  assign w5555 = w5266 & w5416 ;
  assign w5556 = ~w5273 & w5338 ;
  assign w5557 = w5339 ^ w5556 ;
  assign w5558 = ~w5416 & w5557 ;
  assign w5559 = w5555 | w5558 ;
  assign w5560 = ~\pi072 & w5559 ;
  assign w5561 = w5272 & w5416 ;
  assign w5562 = ~w5279 & w5335 ;
  assign w5563 = w5336 ^ w5562 ;
  assign w5564 = ~w5416 & w5563 ;
  assign w5565 = w5561 | w5564 ;
  assign w5566 = ~\pi071 & w5565 ;
  assign w5567 = w5278 & w5416 ;
  assign w5568 = ~w5285 & w5332 ;
  assign w5569 = w5333 ^ w5568 ;
  assign w5570 = ~w5416 & w5569 ;
  assign w5571 = w5567 | w5570 ;
  assign w5572 = ~\pi070 & w5571 ;
  assign w5573 = w5284 & w5416 ;
  assign w5574 = ~w5293 & w5329 ;
  assign w5575 = w5330 ^ w5574 ;
  assign w5576 = ~w5416 & w5575 ;
  assign w5577 = w5573 | w5576 ;
  assign w5578 = ~\pi069 & w5577 ;
  assign w5579 = w5292 & w5416 ;
  assign w5580 = ~w5304 & w5326 ;
  assign w5581 = w5327 ^ w5580 ;
  assign w5582 = ~w5416 & w5581 ;
  assign w5583 = w5579 | w5582 ;
  assign w5584 = ~\pi068 & w5583 ;
  assign w5585 = w5303 & w5416 ;
  assign w5586 = ~w5317 & w5320 ;
  assign w5587 = ( \pi065 & w5320 ) | ( \pi065 & w5586 ) | ( w5320 & w5586 ) ;
  assign w5588 = w5323 ^ w5587 ;
  assign w5589 = ~w5416 & w5588 ;
  assign w5590 = w5585 | w5589 ;
  assign w5591 = ~\pi067 & w5590 ;
  assign w5592 = ( ~w298 & w5309 ) | ( ~w298 & w5316 ) | ( w5309 & w5316 ) ;
  assign w5593 = \pi065 ^ w5592 ;
  assign w5594 = ( ~w298 & w5318 ) | ( ~w298 & w5593 ) | ( w5318 & w5593 ) ;
  assign w5595 = ( w5318 & w5415 ) | ( w5318 & w5593 ) | ( w5415 & w5593 ) ;
  assign w5596 = w5594 & ~w5595 ;
  assign w5597 = ( w5317 & w5416 ) | ( w5317 & w5596 ) | ( w5416 & w5596 ) ;
  assign w5598 = w5596 | w5597 ;
  assign w5599 = ~\pi066 & w5598 ;
  assign w5600 = \pi064 & ~\pi096 ;
  assign w5601 = ~w451 & w5600 ;
  assign w5602 = ~w5116 & w5601 ;
  assign w5603 = ( \pi032 & w5415 ) | ( \pi032 & ~w5602 ) | ( w5415 & ~w5602 ) ;
  assign w5604 = \pi032 & w5603 ;
  assign w5605 = ~w179 & w5318 ;
  assign w5606 = ~w170 & w5605 ;
  assign w5607 = ( w155 & ~w170 ) | ( w155 & w5415 ) | ( ~w170 & w5415 ) ;
  assign w5608 = w5606 & ~w5607 ;
  assign w5609 = ~\pi031 & \pi064 ;
  assign w5610 = ~w5317 & w5416 ;
  assign w5611 = ( w5416 & w5596 ) | ( w5416 & ~w5610 ) | ( w5596 & ~w5610 ) ;
  assign w5612 = \pi066 ^ w5611 ;
  assign w5613 = w5604 | w5608 ;
  assign w5614 = ( \pi065 & w5609 ) | ( \pi065 & ~w5613 ) | ( w5609 & ~w5613 ) ;
  assign w5615 = w5612 | w5614 ;
  assign w5616 = \pi067 ^ w5590 ;
  assign w5617 = ( ~w5599 & w5615 ) | ( ~w5599 & w5616 ) | ( w5615 & w5616 ) ;
  assign w5618 = w5616 | w5617 ;
  assign w5619 = \pi068 ^ w5583 ;
  assign w5620 = ( ~w5591 & w5618 ) | ( ~w5591 & w5619 ) | ( w5618 & w5619 ) ;
  assign w5621 = w5619 | w5620 ;
  assign w5622 = \pi069 ^ w5577 ;
  assign w5623 = ( ~w5584 & w5621 ) | ( ~w5584 & w5622 ) | ( w5621 & w5622 ) ;
  assign w5624 = w5622 | w5623 ;
  assign w5625 = \pi070 ^ w5571 ;
  assign w5626 = ( ~w5578 & w5624 ) | ( ~w5578 & w5625 ) | ( w5624 & w5625 ) ;
  assign w5627 = w5625 | w5626 ;
  assign w5628 = \pi071 ^ w5565 ;
  assign w5629 = ( ~w5572 & w5627 ) | ( ~w5572 & w5628 ) | ( w5627 & w5628 ) ;
  assign w5630 = w5628 | w5629 ;
  assign w5631 = \pi072 ^ w5559 ;
  assign w5632 = ( ~w5566 & w5630 ) | ( ~w5566 & w5631 ) | ( w5630 & w5631 ) ;
  assign w5633 = w5631 | w5632 ;
  assign w5634 = \pi073 ^ w5553 ;
  assign w5635 = ( ~w5560 & w5633 ) | ( ~w5560 & w5634 ) | ( w5633 & w5634 ) ;
  assign w5636 = w5634 | w5635 ;
  assign w5637 = \pi074 ^ w5547 ;
  assign w5638 = ( ~w5554 & w5636 ) | ( ~w5554 & w5637 ) | ( w5636 & w5637 ) ;
  assign w5639 = w5637 | w5638 ;
  assign w5640 = \pi075 ^ w5541 ;
  assign w5641 = ( ~w5548 & w5639 ) | ( ~w5548 & w5640 ) | ( w5639 & w5640 ) ;
  assign w5642 = w5640 | w5641 ;
  assign w5643 = \pi076 ^ w5535 ;
  assign w5644 = ( ~w5542 & w5642 ) | ( ~w5542 & w5643 ) | ( w5642 & w5643 ) ;
  assign w5645 = w5643 | w5644 ;
  assign w5646 = \pi077 ^ w5529 ;
  assign w5647 = ( ~w5536 & w5645 ) | ( ~w5536 & w5646 ) | ( w5645 & w5646 ) ;
  assign w5648 = w5646 | w5647 ;
  assign w5649 = \pi078 ^ w5523 ;
  assign w5650 = ( ~w5530 & w5648 ) | ( ~w5530 & w5649 ) | ( w5648 & w5649 ) ;
  assign w5651 = w5649 | w5650 ;
  assign w5652 = \pi079 ^ w5517 ;
  assign w5653 = ( ~w5524 & w5651 ) | ( ~w5524 & w5652 ) | ( w5651 & w5652 ) ;
  assign w5654 = w5652 | w5653 ;
  assign w5655 = \pi080 ^ w5511 ;
  assign w5656 = ( ~w5518 & w5654 ) | ( ~w5518 & w5655 ) | ( w5654 & w5655 ) ;
  assign w5657 = w5655 | w5656 ;
  assign w5658 = \pi081 ^ w5505 ;
  assign w5659 = ( ~w5512 & w5657 ) | ( ~w5512 & w5658 ) | ( w5657 & w5658 ) ;
  assign w5660 = w5658 | w5659 ;
  assign w5661 = \pi082 ^ w5499 ;
  assign w5662 = ( ~w5506 & w5660 ) | ( ~w5506 & w5661 ) | ( w5660 & w5661 ) ;
  assign w5663 = w5661 | w5662 ;
  assign w5664 = \pi083 ^ w5493 ;
  assign w5665 = ( ~w5500 & w5663 ) | ( ~w5500 & w5664 ) | ( w5663 & w5664 ) ;
  assign w5666 = w5664 | w5665 ;
  assign w5667 = \pi084 ^ w5487 ;
  assign w5668 = ( ~w5494 & w5666 ) | ( ~w5494 & w5667 ) | ( w5666 & w5667 ) ;
  assign w5669 = w5667 | w5668 ;
  assign w5670 = \pi085 ^ w5481 ;
  assign w5671 = ( ~w5488 & w5669 ) | ( ~w5488 & w5670 ) | ( w5669 & w5670 ) ;
  assign w5672 = w5670 | w5671 ;
  assign w5673 = \pi086 ^ w5475 ;
  assign w5674 = ( ~w5482 & w5672 ) | ( ~w5482 & w5673 ) | ( w5672 & w5673 ) ;
  assign w5675 = w5673 | w5674 ;
  assign w5676 = \pi087 ^ w5469 ;
  assign w5677 = ( ~w5476 & w5675 ) | ( ~w5476 & w5676 ) | ( w5675 & w5676 ) ;
  assign w5678 = w5676 | w5677 ;
  assign w5679 = \pi088 ^ w5463 ;
  assign w5680 = ( ~w5470 & w5678 ) | ( ~w5470 & w5679 ) | ( w5678 & w5679 ) ;
  assign w5681 = w5679 | w5680 ;
  assign w5682 = \pi089 ^ w5457 ;
  assign w5683 = ( ~w5464 & w5681 ) | ( ~w5464 & w5682 ) | ( w5681 & w5682 ) ;
  assign w5684 = w5682 | w5683 ;
  assign w5685 = \pi090 ^ w5451 ;
  assign w5686 = ( ~w5458 & w5684 ) | ( ~w5458 & w5685 ) | ( w5684 & w5685 ) ;
  assign w5687 = w5685 | w5686 ;
  assign w5688 = \pi091 ^ w5445 ;
  assign w5689 = ( ~w5452 & w5687 ) | ( ~w5452 & w5688 ) | ( w5687 & w5688 ) ;
  assign w5690 = w5688 | w5689 ;
  assign w5691 = \pi092 ^ w5439 ;
  assign w5692 = ( ~w5446 & w5690 ) | ( ~w5446 & w5691 ) | ( w5690 & w5691 ) ;
  assign w5693 = w5691 | w5692 ;
  assign w5694 = \pi093 ^ w5433 ;
  assign w5695 = ( ~w5440 & w5693 ) | ( ~w5440 & w5694 ) | ( w5693 & w5694 ) ;
  assign w5696 = w5694 | w5695 ;
  assign w5697 = \pi094 ^ w5427 ;
  assign w5698 = ( ~w5434 & w5696 ) | ( ~w5434 & w5697 ) | ( w5696 & w5697 ) ;
  assign w5699 = w5697 | w5698 ;
  assign w5700 = \pi095 ^ w5421 ;
  assign w5701 = ( ~w5428 & w5699 ) | ( ~w5428 & w5700 ) | ( w5699 & w5700 ) ;
  assign w5702 = w5700 | w5701 ;
  assign w5703 = w5128 & w5416 ;
  assign w5704 = ~w5129 & w5410 ;
  assign w5705 = w5411 ^ w5704 ;
  assign w5706 = ~w5416 & w5705 ;
  assign w5707 = w5703 | w5706 ;
  assign w5708 = ~\pi096 & w5707 ;
  assign w5709 = ( \pi096 & ~w5703 ) | ( \pi096 & w5706 ) | ( ~w5703 & w5706 ) ;
  assign w5710 = ~w5706 & w5709 ;
  assign w5711 = w5708 | w5710 ;
  assign w5712 = ( ~w5422 & w5702 ) | ( ~w5422 & w5711 ) | ( w5702 & w5711 ) ;
  assign w5713 = ( w291 & ~w5711 ) | ( w291 & w5712 ) | ( ~w5711 & w5712 ) ;
  assign w5714 = w5711 | w5713 ;
  assign w5715 = ~w298 & w5707 ;
  assign w5716 = w5714 & ~w5715 ;
  assign w5717 = ~w5428 & w5699 ;
  assign w5718 = w5700 ^ w5717 ;
  assign w5719 = ~w5716 & w5718 ;
  assign w5720 = ( w5421 & w5714 ) | ( w5421 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5721 = ~w5715 & w5720 ;
  assign w5722 = w5719 | w5721 ;
  assign w5723 = ( ~w5422 & w5702 ) | ( ~w5422 & w5716 ) | ( w5702 & w5716 ) ;
  assign w5724 = w5711 ^ w5723 ;
  assign w5725 = ~w5716 & w5724 ;
  assign w5726 = ( w298 & ~w5707 ) | ( w298 & w5714 ) | ( ~w5707 & w5714 ) ;
  assign w5727 = w5707 & w5726 ;
  assign w5728 = w5725 | w5727 ;
  assign w5729 = ~\pi096 & w5722 ;
  assign w5730 = ~w5434 & w5696 ;
  assign w5731 = w5697 ^ w5730 ;
  assign w5732 = ~w5716 & w5731 ;
  assign w5733 = ( w5427 & w5714 ) | ( w5427 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5734 = ~w5715 & w5733 ;
  assign w5735 = w5732 | w5734 ;
  assign w5736 = ~\pi095 & w5735 ;
  assign w5737 = ~w5440 & w5693 ;
  assign w5738 = w5694 ^ w5737 ;
  assign w5739 = ~w5716 & w5738 ;
  assign w5740 = ( w5433 & w5714 ) | ( w5433 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5741 = ~w5715 & w5740 ;
  assign w5742 = w5739 | w5741 ;
  assign w5743 = ~\pi094 & w5742 ;
  assign w5744 = ~w5446 & w5690 ;
  assign w5745 = w5691 ^ w5744 ;
  assign w5746 = ~w5716 & w5745 ;
  assign w5747 = ( w5439 & w5714 ) | ( w5439 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5748 = ~w5715 & w5747 ;
  assign w5749 = w5746 | w5748 ;
  assign w5750 = ~\pi093 & w5749 ;
  assign w5751 = ~w5452 & w5687 ;
  assign w5752 = w5688 ^ w5751 ;
  assign w5753 = ~w5716 & w5752 ;
  assign w5754 = ( w5445 & w5714 ) | ( w5445 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5755 = ~w5715 & w5754 ;
  assign w5756 = w5753 | w5755 ;
  assign w5757 = ~\pi092 & w5756 ;
  assign w5758 = ~w5458 & w5684 ;
  assign w5759 = w5685 ^ w5758 ;
  assign w5760 = ~w5716 & w5759 ;
  assign w5761 = ( w5451 & w5714 ) | ( w5451 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5762 = ~w5715 & w5761 ;
  assign w5763 = w5760 | w5762 ;
  assign w5764 = ~\pi091 & w5763 ;
  assign w5765 = ~w5464 & w5681 ;
  assign w5766 = w5682 ^ w5765 ;
  assign w5767 = ~w5716 & w5766 ;
  assign w5768 = ( w5457 & w5714 ) | ( w5457 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5769 = ~w5715 & w5768 ;
  assign w5770 = w5767 | w5769 ;
  assign w5771 = ~\pi090 & w5770 ;
  assign w5772 = ~w5470 & w5678 ;
  assign w5773 = w5679 ^ w5772 ;
  assign w5774 = ~w5716 & w5773 ;
  assign w5775 = ( w5463 & w5714 ) | ( w5463 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5776 = ~w5715 & w5775 ;
  assign w5777 = w5774 | w5776 ;
  assign w5778 = ~\pi089 & w5777 ;
  assign w5779 = ~w5476 & w5675 ;
  assign w5780 = w5676 ^ w5779 ;
  assign w5781 = ~w5716 & w5780 ;
  assign w5782 = ( w5469 & w5714 ) | ( w5469 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5783 = ~w5715 & w5782 ;
  assign w5784 = w5781 | w5783 ;
  assign w5785 = ~\pi088 & w5784 ;
  assign w5786 = ~w5482 & w5672 ;
  assign w5787 = w5673 ^ w5786 ;
  assign w5788 = ~w5716 & w5787 ;
  assign w5789 = ( w5475 & w5714 ) | ( w5475 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5790 = ~w5715 & w5789 ;
  assign w5791 = w5788 | w5790 ;
  assign w5792 = ~\pi087 & w5791 ;
  assign w5793 = ~w5488 & w5669 ;
  assign w5794 = w5670 ^ w5793 ;
  assign w5795 = ~w5716 & w5794 ;
  assign w5796 = ( w5481 & w5714 ) | ( w5481 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5797 = ~w5715 & w5796 ;
  assign w5798 = w5795 | w5797 ;
  assign w5799 = ~\pi086 & w5798 ;
  assign w5800 = ~w5494 & w5666 ;
  assign w5801 = w5667 ^ w5800 ;
  assign w5802 = ~w5716 & w5801 ;
  assign w5803 = ( w5487 & w5714 ) | ( w5487 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5804 = ~w5715 & w5803 ;
  assign w5805 = w5802 | w5804 ;
  assign w5806 = ~\pi085 & w5805 ;
  assign w5807 = ~w5500 & w5663 ;
  assign w5808 = w5664 ^ w5807 ;
  assign w5809 = ~w5716 & w5808 ;
  assign w5810 = ( w5493 & w5714 ) | ( w5493 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5811 = ~w5715 & w5810 ;
  assign w5812 = w5809 | w5811 ;
  assign w5813 = ~\pi084 & w5812 ;
  assign w5814 = ~w5506 & w5660 ;
  assign w5815 = w5661 ^ w5814 ;
  assign w5816 = ~w5716 & w5815 ;
  assign w5817 = ( w5499 & w5714 ) | ( w5499 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5818 = ~w5715 & w5817 ;
  assign w5819 = w5816 | w5818 ;
  assign w5820 = ~\pi083 & w5819 ;
  assign w5821 = ~w5512 & w5657 ;
  assign w5822 = w5658 ^ w5821 ;
  assign w5823 = ~w5716 & w5822 ;
  assign w5824 = ( w5505 & w5714 ) | ( w5505 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5825 = ~w5715 & w5824 ;
  assign w5826 = w5823 | w5825 ;
  assign w5827 = ~\pi082 & w5826 ;
  assign w5828 = ~w5518 & w5654 ;
  assign w5829 = w5655 ^ w5828 ;
  assign w5830 = ~w5716 & w5829 ;
  assign w5831 = ( w5511 & w5714 ) | ( w5511 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5832 = ~w5715 & w5831 ;
  assign w5833 = w5830 | w5832 ;
  assign w5834 = ~\pi081 & w5833 ;
  assign w5835 = ~w5524 & w5651 ;
  assign w5836 = w5652 ^ w5835 ;
  assign w5837 = ~w5716 & w5836 ;
  assign w5838 = ( w5517 & w5714 ) | ( w5517 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5839 = ~w5715 & w5838 ;
  assign w5840 = w5837 | w5839 ;
  assign w5841 = ~\pi080 & w5840 ;
  assign w5842 = ~w5530 & w5648 ;
  assign w5843 = w5649 ^ w5842 ;
  assign w5844 = ~w5716 & w5843 ;
  assign w5845 = ( w5523 & w5714 ) | ( w5523 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5846 = ~w5715 & w5845 ;
  assign w5847 = w5844 | w5846 ;
  assign w5848 = ~\pi079 & w5847 ;
  assign w5849 = ~w5536 & w5645 ;
  assign w5850 = w5646 ^ w5849 ;
  assign w5851 = ~w5716 & w5850 ;
  assign w5852 = ( w5529 & w5714 ) | ( w5529 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5853 = ~w5715 & w5852 ;
  assign w5854 = w5851 | w5853 ;
  assign w5855 = ~\pi078 & w5854 ;
  assign w5856 = ~w5542 & w5642 ;
  assign w5857 = w5643 ^ w5856 ;
  assign w5858 = ~w5716 & w5857 ;
  assign w5859 = ( w5535 & w5714 ) | ( w5535 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5860 = ~w5715 & w5859 ;
  assign w5861 = w5858 | w5860 ;
  assign w5862 = ~\pi077 & w5861 ;
  assign w5863 = ~w5548 & w5639 ;
  assign w5864 = w5640 ^ w5863 ;
  assign w5865 = ~w5716 & w5864 ;
  assign w5866 = ( w5541 & w5714 ) | ( w5541 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5867 = ~w5715 & w5866 ;
  assign w5868 = w5865 | w5867 ;
  assign w5869 = ~\pi076 & w5868 ;
  assign w5870 = ~w5554 & w5636 ;
  assign w5871 = w5637 ^ w5870 ;
  assign w5872 = ~w5716 & w5871 ;
  assign w5873 = ( w5547 & w5714 ) | ( w5547 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5874 = ~w5715 & w5873 ;
  assign w5875 = w5872 | w5874 ;
  assign w5876 = ~\pi075 & w5875 ;
  assign w5877 = ~w5560 & w5633 ;
  assign w5878 = w5634 ^ w5877 ;
  assign w5879 = ~w5716 & w5878 ;
  assign w5880 = ( w5553 & w5714 ) | ( w5553 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5881 = ~w5715 & w5880 ;
  assign w5882 = w5879 | w5881 ;
  assign w5883 = ~\pi074 & w5882 ;
  assign w5884 = ~w5566 & w5630 ;
  assign w5885 = w5631 ^ w5884 ;
  assign w5886 = ~w5716 & w5885 ;
  assign w5887 = ( w5559 & w5714 ) | ( w5559 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5888 = ~w5715 & w5887 ;
  assign w5889 = w5886 | w5888 ;
  assign w5890 = ~\pi073 & w5889 ;
  assign w5891 = ~w5572 & w5627 ;
  assign w5892 = w5628 ^ w5891 ;
  assign w5893 = ~w5716 & w5892 ;
  assign w5894 = ( w5565 & w5714 ) | ( w5565 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5895 = ~w5715 & w5894 ;
  assign w5896 = w5893 | w5895 ;
  assign w5897 = ~\pi072 & w5896 ;
  assign w5898 = ~w5578 & w5624 ;
  assign w5899 = w5625 ^ w5898 ;
  assign w5900 = ~w5716 & w5899 ;
  assign w5901 = ( w5571 & w5714 ) | ( w5571 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5902 = ~w5715 & w5901 ;
  assign w5903 = w5900 | w5902 ;
  assign w5904 = ~\pi071 & w5903 ;
  assign w5905 = ~w5584 & w5621 ;
  assign w5906 = w5622 ^ w5905 ;
  assign w5907 = ~w5716 & w5906 ;
  assign w5908 = ( w5577 & w5714 ) | ( w5577 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5909 = ~w5715 & w5908 ;
  assign w5910 = w5907 | w5909 ;
  assign w5911 = ~\pi070 & w5910 ;
  assign w5912 = ~w5591 & w5618 ;
  assign w5913 = w5619 ^ w5912 ;
  assign w5914 = ~w5716 & w5913 ;
  assign w5915 = ( w5583 & w5714 ) | ( w5583 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5916 = ~w5715 & w5915 ;
  assign w5917 = w5914 | w5916 ;
  assign w5918 = ~\pi069 & w5917 ;
  assign w5919 = ~w5599 & w5615 ;
  assign w5920 = w5616 ^ w5919 ;
  assign w5921 = ~w5716 & w5920 ;
  assign w5922 = ( w5590 & w5714 ) | ( w5590 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5923 = ~w5715 & w5922 ;
  assign w5924 = w5921 | w5923 ;
  assign w5925 = ~\pi068 & w5924 ;
  assign w5926 = w5612 ^ w5614 ;
  assign w5927 = ~w5716 & w5926 ;
  assign w5928 = ( w5598 & w5714 ) | ( w5598 & w5715 ) | ( w5714 & w5715 ) ;
  assign w5929 = ~w5715 & w5928 ;
  assign w5930 = w5927 | w5929 ;
  assign w5931 = ~\pi067 & w5930 ;
  assign w5932 = w5609 ^ w5613 ;
  assign w5933 = \pi065 ^ w5932 ;
  assign w5934 = ~w5716 & w5933 ;
  assign w5935 = ( w5604 & w5608 ) | ( w5604 & ~w5715 ) | ( w5608 & ~w5715 ) ;
  assign w5936 = w5715 & w5935 ;
  assign w5937 = ( ~w5714 & w5935 ) | ( ~w5714 & w5936 ) | ( w5935 & w5936 ) ;
  assign w5938 = ( w5934 & w5935 ) | ( w5934 & ~w5937 ) | ( w5935 & ~w5937 ) ;
  assign w5939 = ~\pi066 & w5938 ;
  assign w5940 = w5714 | w5715 ;
  assign w5941 = ( w5934 & w5935 ) | ( w5934 & w5940 ) | ( w5935 & w5940 ) ;
  assign w5942 = ( ~w5715 & w5934 ) | ( ~w5715 & w5941 ) | ( w5934 & w5941 ) ;
  assign w5943 = \pi066 ^ w5942 ;
  assign w5944 = \pi064 & ~w5716 ;
  assign w5945 = \pi031 ^ w5944 ;
  assign w5946 = ( ~\pi030 & \pi064 ) | ( ~\pi030 & w5943 ) | ( \pi064 & w5943 ) ;
  assign w5947 = ( \pi065 & ~w5945 ) | ( \pi065 & w5946 ) | ( ~w5945 & w5946 ) ;
  assign w5948 = w5943 | w5947 ;
  assign w5949 = \pi067 ^ w5930 ;
  assign w5950 = ( ~w5939 & w5948 ) | ( ~w5939 & w5949 ) | ( w5948 & w5949 ) ;
  assign w5951 = w5949 | w5950 ;
  assign w5952 = \pi068 ^ w5924 ;
  assign w5953 = ( ~w5931 & w5951 ) | ( ~w5931 & w5952 ) | ( w5951 & w5952 ) ;
  assign w5954 = w5952 | w5953 ;
  assign w5955 = \pi069 ^ w5917 ;
  assign w5956 = ( ~w5925 & w5954 ) | ( ~w5925 & w5955 ) | ( w5954 & w5955 ) ;
  assign w5957 = w5955 | w5956 ;
  assign w5958 = \pi070 ^ w5910 ;
  assign w5959 = ( ~w5918 & w5957 ) | ( ~w5918 & w5958 ) | ( w5957 & w5958 ) ;
  assign w5960 = w5958 | w5959 ;
  assign w5961 = \pi071 ^ w5903 ;
  assign w5962 = ( ~w5911 & w5960 ) | ( ~w5911 & w5961 ) | ( w5960 & w5961 ) ;
  assign w5963 = w5961 | w5962 ;
  assign w5964 = \pi072 ^ w5896 ;
  assign w5965 = ( ~w5904 & w5963 ) | ( ~w5904 & w5964 ) | ( w5963 & w5964 ) ;
  assign w5966 = w5964 | w5965 ;
  assign w5967 = \pi073 ^ w5889 ;
  assign w5968 = ( ~w5897 & w5966 ) | ( ~w5897 & w5967 ) | ( w5966 & w5967 ) ;
  assign w5969 = w5967 | w5968 ;
  assign w5970 = \pi074 ^ w5882 ;
  assign w5971 = ( ~w5890 & w5969 ) | ( ~w5890 & w5970 ) | ( w5969 & w5970 ) ;
  assign w5972 = w5970 | w5971 ;
  assign w5973 = \pi075 ^ w5875 ;
  assign w5974 = ( ~w5883 & w5972 ) | ( ~w5883 & w5973 ) | ( w5972 & w5973 ) ;
  assign w5975 = w5973 | w5974 ;
  assign w5976 = \pi076 ^ w5868 ;
  assign w5977 = ( ~w5876 & w5975 ) | ( ~w5876 & w5976 ) | ( w5975 & w5976 ) ;
  assign w5978 = w5976 | w5977 ;
  assign w5979 = \pi077 ^ w5861 ;
  assign w5980 = ( ~w5869 & w5978 ) | ( ~w5869 & w5979 ) | ( w5978 & w5979 ) ;
  assign w5981 = w5979 | w5980 ;
  assign w5982 = \pi078 ^ w5854 ;
  assign w5983 = ( ~w5862 & w5981 ) | ( ~w5862 & w5982 ) | ( w5981 & w5982 ) ;
  assign w5984 = w5982 | w5983 ;
  assign w5985 = \pi079 ^ w5847 ;
  assign w5986 = ( ~w5855 & w5984 ) | ( ~w5855 & w5985 ) | ( w5984 & w5985 ) ;
  assign w5987 = w5985 | w5986 ;
  assign w5988 = \pi080 ^ w5840 ;
  assign w5989 = ( ~w5848 & w5987 ) | ( ~w5848 & w5988 ) | ( w5987 & w5988 ) ;
  assign w5990 = w5988 | w5989 ;
  assign w5991 = \pi081 ^ w5833 ;
  assign w5992 = ( ~w5841 & w5990 ) | ( ~w5841 & w5991 ) | ( w5990 & w5991 ) ;
  assign w5993 = w5991 | w5992 ;
  assign w5994 = \pi082 ^ w5826 ;
  assign w5995 = ( ~w5834 & w5993 ) | ( ~w5834 & w5994 ) | ( w5993 & w5994 ) ;
  assign w5996 = w5994 | w5995 ;
  assign w5997 = \pi083 ^ w5819 ;
  assign w5998 = ( ~w5827 & w5996 ) | ( ~w5827 & w5997 ) | ( w5996 & w5997 ) ;
  assign w5999 = w5997 | w5998 ;
  assign w6000 = \pi084 ^ w5812 ;
  assign w6001 = ( ~w5820 & w5999 ) | ( ~w5820 & w6000 ) | ( w5999 & w6000 ) ;
  assign w6002 = w6000 | w6001 ;
  assign w6003 = \pi085 ^ w5805 ;
  assign w6004 = ( ~w5813 & w6002 ) | ( ~w5813 & w6003 ) | ( w6002 & w6003 ) ;
  assign w6005 = w6003 | w6004 ;
  assign w6006 = \pi086 ^ w5798 ;
  assign w6007 = ( ~w5806 & w6005 ) | ( ~w5806 & w6006 ) | ( w6005 & w6006 ) ;
  assign w6008 = w6006 | w6007 ;
  assign w6009 = \pi087 ^ w5791 ;
  assign w6010 = ( ~w5799 & w6008 ) | ( ~w5799 & w6009 ) | ( w6008 & w6009 ) ;
  assign w6011 = w6009 | w6010 ;
  assign w6012 = \pi088 ^ w5784 ;
  assign w6013 = ( ~w5792 & w6011 ) | ( ~w5792 & w6012 ) | ( w6011 & w6012 ) ;
  assign w6014 = w6012 | w6013 ;
  assign w6015 = \pi089 ^ w5777 ;
  assign w6016 = ( ~w5785 & w6014 ) | ( ~w5785 & w6015 ) | ( w6014 & w6015 ) ;
  assign w6017 = w6015 | w6016 ;
  assign w6018 = \pi090 ^ w5770 ;
  assign w6019 = ( ~w5778 & w6017 ) | ( ~w5778 & w6018 ) | ( w6017 & w6018 ) ;
  assign w6020 = w6018 | w6019 ;
  assign w6021 = \pi091 ^ w5763 ;
  assign w6022 = ( ~w5771 & w6020 ) | ( ~w5771 & w6021 ) | ( w6020 & w6021 ) ;
  assign w6023 = w6021 | w6022 ;
  assign w6024 = \pi092 ^ w5756 ;
  assign w6025 = ( ~w5764 & w6023 ) | ( ~w5764 & w6024 ) | ( w6023 & w6024 ) ;
  assign w6026 = w6024 | w6025 ;
  assign w6027 = \pi093 ^ w5749 ;
  assign w6028 = ( ~w5757 & w6026 ) | ( ~w5757 & w6027 ) | ( w6026 & w6027 ) ;
  assign w6029 = w6027 | w6028 ;
  assign w6030 = \pi094 ^ w5742 ;
  assign w6031 = ( ~w5750 & w6029 ) | ( ~w5750 & w6030 ) | ( w6029 & w6030 ) ;
  assign w6032 = w6030 | w6031 ;
  assign w6033 = \pi095 ^ w5735 ;
  assign w6034 = ( ~w5743 & w6032 ) | ( ~w5743 & w6033 ) | ( w6032 & w6033 ) ;
  assign w6035 = w6033 | w6034 ;
  assign w6036 = \pi096 ^ w5722 ;
  assign w6037 = ( ~w5736 & w6035 ) | ( ~w5736 & w6036 ) | ( w6035 & w6036 ) ;
  assign w6038 = w6036 | w6037 ;
  assign w6039 = \pi097 ^ w5728 ;
  assign w6040 = w5729 & ~w6039 ;
  assign w6041 = ( w6038 & w6039 ) | ( w6038 & ~w6040 ) | ( w6039 & ~w6040 ) ;
  assign w6042 = ~\pi097 & w5728 ;
  assign w6043 = w6041 & ~w6042 ;
  assign w6044 = \pi098 | \pi099 ;
  assign w6045 = w202 | w6044 ;
  assign w6046 = ( w161 & w201 ) | ( w161 & ~w202 ) | ( w201 & ~w202 ) ;
  assign w6047 = w6045 | w6046 ;
  assign w6048 = w6043 | w6047 ;
  assign w6049 = w5722 & w6048 ;
  assign w6050 = ~w5736 & w6035 ;
  assign w6051 = w6036 ^ w6050 ;
  assign w6052 = ~w6048 & w6051 ;
  assign w6053 = w6049 | w6052 ;
  assign w6054 = w5728 & w6048 ;
  assign w6055 = ~w5729 & w6038 ;
  assign w6056 = w6039 ^ w6055 ;
  assign w6057 = ~w6048 & w6056 ;
  assign w6058 = w6054 | w6057 ;
  assign w6059 = ~\pi097 & w6053 ;
  assign w6060 = w5735 & w6048 ;
  assign w6061 = ~w5743 & w6032 ;
  assign w6062 = w6033 ^ w6061 ;
  assign w6063 = ~w6048 & w6062 ;
  assign w6064 = w6060 | w6063 ;
  assign w6065 = ~\pi096 & w6064 ;
  assign w6066 = w5742 & w6048 ;
  assign w6067 = ~w5750 & w6029 ;
  assign w6068 = w6030 ^ w6067 ;
  assign w6069 = ~w6048 & w6068 ;
  assign w6070 = w6066 | w6069 ;
  assign w6071 = ~\pi095 & w6070 ;
  assign w6072 = w5749 & w6048 ;
  assign w6073 = ~w5757 & w6026 ;
  assign w6074 = w6027 ^ w6073 ;
  assign w6075 = ~w6048 & w6074 ;
  assign w6076 = w6072 | w6075 ;
  assign w6077 = ~\pi094 & w6076 ;
  assign w6078 = w5756 & w6048 ;
  assign w6079 = ~w5764 & w6023 ;
  assign w6080 = w6024 ^ w6079 ;
  assign w6081 = ~w6048 & w6080 ;
  assign w6082 = w6078 | w6081 ;
  assign w6083 = ~\pi093 & w6082 ;
  assign w6084 = w5763 & w6048 ;
  assign w6085 = ~w5771 & w6020 ;
  assign w6086 = w6021 ^ w6085 ;
  assign w6087 = ~w6048 & w6086 ;
  assign w6088 = w6084 | w6087 ;
  assign w6089 = ~\pi092 & w6088 ;
  assign w6090 = w5770 & w6048 ;
  assign w6091 = ~w5778 & w6017 ;
  assign w6092 = w6018 ^ w6091 ;
  assign w6093 = ~w6048 & w6092 ;
  assign w6094 = w6090 | w6093 ;
  assign w6095 = ~\pi091 & w6094 ;
  assign w6096 = w5777 & w6048 ;
  assign w6097 = ~w5785 & w6014 ;
  assign w6098 = w6015 ^ w6097 ;
  assign w6099 = ~w6048 & w6098 ;
  assign w6100 = w6096 | w6099 ;
  assign w6101 = ~\pi090 & w6100 ;
  assign w6102 = w5784 & w6048 ;
  assign w6103 = ~w5792 & w6011 ;
  assign w6104 = w6012 ^ w6103 ;
  assign w6105 = ~w6048 & w6104 ;
  assign w6106 = w6102 | w6105 ;
  assign w6107 = ~\pi089 & w6106 ;
  assign w6108 = w5791 & w6048 ;
  assign w6109 = ~w5799 & w6008 ;
  assign w6110 = w6009 ^ w6109 ;
  assign w6111 = ~w6048 & w6110 ;
  assign w6112 = w6108 | w6111 ;
  assign w6113 = ~\pi088 & w6112 ;
  assign w6114 = w5798 & w6048 ;
  assign w6115 = ~w5806 & w6005 ;
  assign w6116 = w6006 ^ w6115 ;
  assign w6117 = ~w6048 & w6116 ;
  assign w6118 = w6114 | w6117 ;
  assign w6119 = ~\pi087 & w6118 ;
  assign w6120 = w5805 & w6048 ;
  assign w6121 = ~w5813 & w6002 ;
  assign w6122 = w6003 ^ w6121 ;
  assign w6123 = ~w6048 & w6122 ;
  assign w6124 = w6120 | w6123 ;
  assign w6125 = ~\pi086 & w6124 ;
  assign w6126 = w5812 & w6048 ;
  assign w6127 = ~w5820 & w5999 ;
  assign w6128 = w6000 ^ w6127 ;
  assign w6129 = ~w6048 & w6128 ;
  assign w6130 = w6126 | w6129 ;
  assign w6131 = ~\pi085 & w6130 ;
  assign w6132 = w5819 & w6048 ;
  assign w6133 = ~w5827 & w5996 ;
  assign w6134 = w5997 ^ w6133 ;
  assign w6135 = ~w6048 & w6134 ;
  assign w6136 = w6132 | w6135 ;
  assign w6137 = ~\pi084 & w6136 ;
  assign w6138 = w5826 & w6048 ;
  assign w6139 = ~w5834 & w5993 ;
  assign w6140 = w5994 ^ w6139 ;
  assign w6141 = ~w6048 & w6140 ;
  assign w6142 = w6138 | w6141 ;
  assign w6143 = ~\pi083 & w6142 ;
  assign w6144 = w5833 & w6048 ;
  assign w6145 = ~w5841 & w5990 ;
  assign w6146 = w5991 ^ w6145 ;
  assign w6147 = ~w6048 & w6146 ;
  assign w6148 = w6144 | w6147 ;
  assign w6149 = ~\pi082 & w6148 ;
  assign w6150 = w5840 & w6048 ;
  assign w6151 = ~w5848 & w5987 ;
  assign w6152 = w5988 ^ w6151 ;
  assign w6153 = ~w6048 & w6152 ;
  assign w6154 = w6150 | w6153 ;
  assign w6155 = ~\pi081 & w6154 ;
  assign w6156 = w5847 & w6048 ;
  assign w6157 = ~w5855 & w5984 ;
  assign w6158 = w5985 ^ w6157 ;
  assign w6159 = ~w6048 & w6158 ;
  assign w6160 = w6156 | w6159 ;
  assign w6161 = ~\pi080 & w6160 ;
  assign w6162 = w5854 & w6048 ;
  assign w6163 = ~w5862 & w5981 ;
  assign w6164 = w5982 ^ w6163 ;
  assign w6165 = ~w6048 & w6164 ;
  assign w6166 = w6162 | w6165 ;
  assign w6167 = ~\pi079 & w6166 ;
  assign w6168 = w5861 & w6048 ;
  assign w6169 = ~w5869 & w5978 ;
  assign w6170 = w5979 ^ w6169 ;
  assign w6171 = ~w6048 & w6170 ;
  assign w6172 = w6168 | w6171 ;
  assign w6173 = ~\pi078 & w6172 ;
  assign w6174 = w5868 & w6048 ;
  assign w6175 = ~w5876 & w5975 ;
  assign w6176 = w5976 ^ w6175 ;
  assign w6177 = ~w6048 & w6176 ;
  assign w6178 = w6174 | w6177 ;
  assign w6179 = ~\pi077 & w6178 ;
  assign w6180 = w5875 & w6048 ;
  assign w6181 = ~w5883 & w5972 ;
  assign w6182 = w5973 ^ w6181 ;
  assign w6183 = ~w6048 & w6182 ;
  assign w6184 = w6180 | w6183 ;
  assign w6185 = ~\pi076 & w6184 ;
  assign w6186 = w5882 & w6048 ;
  assign w6187 = ~w5890 & w5969 ;
  assign w6188 = w5970 ^ w6187 ;
  assign w6189 = ~w6048 & w6188 ;
  assign w6190 = w6186 | w6189 ;
  assign w6191 = ~\pi075 & w6190 ;
  assign w6192 = w5889 & w6048 ;
  assign w6193 = ~w5897 & w5966 ;
  assign w6194 = w5967 ^ w6193 ;
  assign w6195 = ~w6048 & w6194 ;
  assign w6196 = w6192 | w6195 ;
  assign w6197 = ~\pi074 & w6196 ;
  assign w6198 = w5896 & w6048 ;
  assign w6199 = ~w5904 & w5963 ;
  assign w6200 = w5964 ^ w6199 ;
  assign w6201 = ~w6048 & w6200 ;
  assign w6202 = w6198 | w6201 ;
  assign w6203 = ~\pi073 & w6202 ;
  assign w6204 = w5903 & w6048 ;
  assign w6205 = ~w5911 & w5960 ;
  assign w6206 = w5961 ^ w6205 ;
  assign w6207 = ~w6048 & w6206 ;
  assign w6208 = w6204 | w6207 ;
  assign w6209 = ~\pi072 & w6208 ;
  assign w6210 = w5910 & w6048 ;
  assign w6211 = ~w5918 & w5957 ;
  assign w6212 = w5958 ^ w6211 ;
  assign w6213 = ~w6048 & w6212 ;
  assign w6214 = w6210 | w6213 ;
  assign w6215 = ~\pi071 & w6214 ;
  assign w6216 = w5917 & w6048 ;
  assign w6217 = ~w5925 & w5954 ;
  assign w6218 = w5955 ^ w6217 ;
  assign w6219 = ~w6048 & w6218 ;
  assign w6220 = w6216 | w6219 ;
  assign w6221 = ~\pi070 & w6220 ;
  assign w6222 = w5924 & w6048 ;
  assign w6223 = ~w5931 & w5951 ;
  assign w6224 = w5952 ^ w6223 ;
  assign w6225 = ~w6048 & w6224 ;
  assign w6226 = w6222 | w6225 ;
  assign w6227 = ~\pi069 & w6226 ;
  assign w6228 = w5930 & w6048 ;
  assign w6229 = ~w5939 & w5948 ;
  assign w6230 = w5949 ^ w6229 ;
  assign w6231 = ~w6048 & w6230 ;
  assign w6232 = w6228 | w6231 ;
  assign w6233 = ~\pi068 & w6232 ;
  assign w6234 = w5938 & w6048 ;
  assign w6235 = ~\pi030 & \pi064 ;
  assign w6236 = ( \pi065 & ~w5945 ) | ( \pi065 & w6235 ) | ( ~w5945 & w6235 ) ;
  assign w6237 = w5943 ^ w6236 ;
  assign w6238 = ( w6043 & w6047 ) | ( w6043 & w6237 ) | ( w6047 & w6237 ) ;
  assign w6239 = w6237 & ~w6238 ;
  assign w6240 = w6234 | w6239 ;
  assign w6241 = ~\pi067 & w6240 ;
  assign w6242 = \pi031 ^ \pi065 ;
  assign w6243 = \pi030 ^ w5716 ;
  assign w6244 = ( \pi064 & w6047 ) | ( \pi064 & w6243 ) | ( w6047 & w6243 ) ;
  assign w6245 = w6242 ^ w6244 ;
  assign w6246 = ~w6047 & w6245 ;
  assign w6247 = ~w6043 & w6246 ;
  assign w6248 = ( ~\pi064 & w5716 ) | ( ~\pi064 & w6048 ) | ( w5716 & w6048 ) ;
  assign w6249 = \pi031 ^ w6248 ;
  assign w6250 = w6048 & ~w6249 ;
  assign w6251 = w6247 | w6250 ;
  assign w6252 = ~\pi066 & w6251 ;
  assign w6253 = ( \pi064 & ~\pi098 ) | ( \pi064 & \pi099 ) | ( ~\pi098 & \pi099 ) ;
  assign w6254 = w278 | w288 ;
  assign w6255 = ( \pi099 & \pi100 ) | ( \pi099 & ~w278 ) | ( \pi100 & ~w278 ) ;
  assign w6256 = w6254 | w6255 ;
  assign w6257 = w6253 & ~w6256 ;
  assign w6258 = ~w275 & w6257 ;
  assign w6259 = ( \pi030 & w6043 ) | ( \pi030 & ~w6258 ) | ( w6043 & ~w6258 ) ;
  assign w6260 = \pi030 & w6259 ;
  assign w6261 = ( ~\pi030 & \pi064 ) | ( ~\pi030 & \pi098 ) | ( \pi064 & \pi098 ) ;
  assign w6262 = w161 | w202 ;
  assign w6263 = ( \pi098 & \pi099 ) | ( \pi098 & ~w161 ) | ( \pi099 & ~w161 ) ;
  assign w6264 = w6262 | w6263 ;
  assign w6265 = w6261 & ~w6264 ;
  assign w6266 = ~w201 & w6265 ;
  assign w6267 = ~w6043 & w6266 ;
  assign w6268 = w6260 | w6267 ;
  assign w6269 = ~\pi029 & \pi064 ;
  assign w6270 = \pi065 ^ w6268 ;
  assign w6271 = w6269 | w6270 ;
  assign w6272 = w6048 | w6247 ;
  assign w6273 = ( w5945 & w6247 ) | ( w5945 & w6272 ) | ( w6247 & w6272 ) ;
  assign w6274 = \pi066 ^ w6273 ;
  assign w6275 = ~\pi065 & w6268 ;
  assign w6276 = w6271 | w6275 ;
  assign w6277 = ( w6274 & ~w6275 ) | ( w6274 & w6276 ) | ( ~w6275 & w6276 ) ;
  assign w6278 = \pi067 ^ w6240 ;
  assign w6279 = ( ~w6252 & w6277 ) | ( ~w6252 & w6278 ) | ( w6277 & w6278 ) ;
  assign w6280 = w6278 | w6279 ;
  assign w6281 = \pi068 ^ w6232 ;
  assign w6282 = ( ~w6241 & w6280 ) | ( ~w6241 & w6281 ) | ( w6280 & w6281 ) ;
  assign w6283 = w6281 | w6282 ;
  assign w6284 = \pi069 ^ w6226 ;
  assign w6285 = ( ~w6233 & w6283 ) | ( ~w6233 & w6284 ) | ( w6283 & w6284 ) ;
  assign w6286 = w6284 | w6285 ;
  assign w6287 = \pi070 ^ w6220 ;
  assign w6288 = ( ~w6227 & w6286 ) | ( ~w6227 & w6287 ) | ( w6286 & w6287 ) ;
  assign w6289 = w6287 | w6288 ;
  assign w6290 = \pi071 ^ w6214 ;
  assign w6291 = ( ~w6221 & w6289 ) | ( ~w6221 & w6290 ) | ( w6289 & w6290 ) ;
  assign w6292 = w6290 | w6291 ;
  assign w6293 = \pi072 ^ w6208 ;
  assign w6294 = ( ~w6215 & w6292 ) | ( ~w6215 & w6293 ) | ( w6292 & w6293 ) ;
  assign w6295 = w6293 | w6294 ;
  assign w6296 = \pi073 ^ w6202 ;
  assign w6297 = ( ~w6209 & w6295 ) | ( ~w6209 & w6296 ) | ( w6295 & w6296 ) ;
  assign w6298 = w6296 | w6297 ;
  assign w6299 = \pi074 ^ w6196 ;
  assign w6300 = ( ~w6203 & w6298 ) | ( ~w6203 & w6299 ) | ( w6298 & w6299 ) ;
  assign w6301 = w6299 | w6300 ;
  assign w6302 = \pi075 ^ w6190 ;
  assign w6303 = ( ~w6197 & w6301 ) | ( ~w6197 & w6302 ) | ( w6301 & w6302 ) ;
  assign w6304 = w6302 | w6303 ;
  assign w6305 = \pi076 ^ w6184 ;
  assign w6306 = ( ~w6191 & w6304 ) | ( ~w6191 & w6305 ) | ( w6304 & w6305 ) ;
  assign w6307 = w6305 | w6306 ;
  assign w6308 = \pi077 ^ w6178 ;
  assign w6309 = ( ~w6185 & w6307 ) | ( ~w6185 & w6308 ) | ( w6307 & w6308 ) ;
  assign w6310 = w6308 | w6309 ;
  assign w6311 = \pi078 ^ w6172 ;
  assign w6312 = ( ~w6179 & w6310 ) | ( ~w6179 & w6311 ) | ( w6310 & w6311 ) ;
  assign w6313 = w6311 | w6312 ;
  assign w6314 = \pi079 ^ w6166 ;
  assign w6315 = ( ~w6173 & w6313 ) | ( ~w6173 & w6314 ) | ( w6313 & w6314 ) ;
  assign w6316 = w6314 | w6315 ;
  assign w6317 = \pi080 ^ w6160 ;
  assign w6318 = ( ~w6167 & w6316 ) | ( ~w6167 & w6317 ) | ( w6316 & w6317 ) ;
  assign w6319 = w6317 | w6318 ;
  assign w6320 = \pi081 ^ w6154 ;
  assign w6321 = ( ~w6161 & w6319 ) | ( ~w6161 & w6320 ) | ( w6319 & w6320 ) ;
  assign w6322 = w6320 | w6321 ;
  assign w6323 = \pi082 ^ w6148 ;
  assign w6324 = ( ~w6155 & w6322 ) | ( ~w6155 & w6323 ) | ( w6322 & w6323 ) ;
  assign w6325 = w6323 | w6324 ;
  assign w6326 = \pi083 ^ w6142 ;
  assign w6327 = ( ~w6149 & w6325 ) | ( ~w6149 & w6326 ) | ( w6325 & w6326 ) ;
  assign w6328 = w6326 | w6327 ;
  assign w6329 = \pi084 ^ w6136 ;
  assign w6330 = ( ~w6143 & w6328 ) | ( ~w6143 & w6329 ) | ( w6328 & w6329 ) ;
  assign w6331 = w6329 | w6330 ;
  assign w6332 = \pi085 ^ w6130 ;
  assign w6333 = ( ~w6137 & w6331 ) | ( ~w6137 & w6332 ) | ( w6331 & w6332 ) ;
  assign w6334 = w6332 | w6333 ;
  assign w6335 = \pi086 ^ w6124 ;
  assign w6336 = ( ~w6131 & w6334 ) | ( ~w6131 & w6335 ) | ( w6334 & w6335 ) ;
  assign w6337 = w6335 | w6336 ;
  assign w6338 = \pi087 ^ w6118 ;
  assign w6339 = ( ~w6125 & w6337 ) | ( ~w6125 & w6338 ) | ( w6337 & w6338 ) ;
  assign w6340 = w6338 | w6339 ;
  assign w6341 = \pi088 ^ w6112 ;
  assign w6342 = ( ~w6119 & w6340 ) | ( ~w6119 & w6341 ) | ( w6340 & w6341 ) ;
  assign w6343 = w6341 | w6342 ;
  assign w6344 = \pi089 ^ w6106 ;
  assign w6345 = ( ~w6113 & w6343 ) | ( ~w6113 & w6344 ) | ( w6343 & w6344 ) ;
  assign w6346 = w6344 | w6345 ;
  assign w6347 = \pi090 ^ w6100 ;
  assign w6348 = ( ~w6107 & w6346 ) | ( ~w6107 & w6347 ) | ( w6346 & w6347 ) ;
  assign w6349 = w6347 | w6348 ;
  assign w6350 = \pi091 ^ w6094 ;
  assign w6351 = ( ~w6101 & w6349 ) | ( ~w6101 & w6350 ) | ( w6349 & w6350 ) ;
  assign w6352 = w6350 | w6351 ;
  assign w6353 = \pi092 ^ w6088 ;
  assign w6354 = ( ~w6095 & w6352 ) | ( ~w6095 & w6353 ) | ( w6352 & w6353 ) ;
  assign w6355 = w6353 | w6354 ;
  assign w6356 = \pi093 ^ w6082 ;
  assign w6357 = ( ~w6089 & w6355 ) | ( ~w6089 & w6356 ) | ( w6355 & w6356 ) ;
  assign w6358 = w6356 | w6357 ;
  assign w6359 = \pi094 ^ w6076 ;
  assign w6360 = ( ~w6083 & w6358 ) | ( ~w6083 & w6359 ) | ( w6358 & w6359 ) ;
  assign w6361 = w6359 | w6360 ;
  assign w6362 = \pi095 ^ w6070 ;
  assign w6363 = ( ~w6077 & w6361 ) | ( ~w6077 & w6362 ) | ( w6361 & w6362 ) ;
  assign w6364 = w6362 | w6363 ;
  assign w6365 = \pi096 ^ w6064 ;
  assign w6366 = ( ~w6071 & w6364 ) | ( ~w6071 & w6365 ) | ( w6364 & w6365 ) ;
  assign w6367 = w6365 | w6366 ;
  assign w6368 = \pi097 ^ w6053 ;
  assign w6369 = ( ~w6065 & w6367 ) | ( ~w6065 & w6368 ) | ( w6367 & w6368 ) ;
  assign w6370 = w6368 | w6369 ;
  assign w6371 = \pi098 ^ w6058 ;
  assign w6372 = w6059 & ~w6371 ;
  assign w6373 = ( w6370 & w6371 ) | ( w6370 & ~w6372 ) | ( w6371 & ~w6372 ) ;
  assign w6374 = ~\pi098 & w6058 ;
  assign w6375 = w6373 & ~w6374 ;
  assign w6376 = \pi099 | \pi100 ;
  assign w6377 = w288 | w6376 ;
  assign w6378 = ( w275 & w278 ) | ( w275 & ~w288 ) | ( w278 & ~w288 ) ;
  assign w6379 = w6377 | w6378 ;
  assign w6380 = w6375 | w6379 ;
  assign w6381 = w6053 & w6380 ;
  assign w6382 = ~w6065 & w6367 ;
  assign w6383 = w6368 ^ w6382 ;
  assign w6384 = ~w6380 & w6383 ;
  assign w6385 = w6381 | w6384 ;
  assign w6386 = ~\pi098 & w6385 ;
  assign w6387 = w6064 & w6380 ;
  assign w6388 = ~w6071 & w6364 ;
  assign w6389 = w6365 ^ w6388 ;
  assign w6390 = ~w6380 & w6389 ;
  assign w6391 = w6387 | w6390 ;
  assign w6392 = ~\pi097 & w6391 ;
  assign w6393 = w6070 & w6380 ;
  assign w6394 = ~w6077 & w6361 ;
  assign w6395 = w6362 ^ w6394 ;
  assign w6396 = ~w6380 & w6395 ;
  assign w6397 = w6393 | w6396 ;
  assign w6398 = ~\pi096 & w6397 ;
  assign w6399 = w6076 & w6380 ;
  assign w6400 = ~w6083 & w6358 ;
  assign w6401 = w6359 ^ w6400 ;
  assign w6402 = ~w6380 & w6401 ;
  assign w6403 = w6399 | w6402 ;
  assign w6404 = ~\pi095 & w6403 ;
  assign w6405 = w6082 & w6380 ;
  assign w6406 = ~w6089 & w6355 ;
  assign w6407 = w6356 ^ w6406 ;
  assign w6408 = ~w6380 & w6407 ;
  assign w6409 = w6405 | w6408 ;
  assign w6410 = ~\pi094 & w6409 ;
  assign w6411 = w6088 & w6380 ;
  assign w6412 = ~w6095 & w6352 ;
  assign w6413 = w6353 ^ w6412 ;
  assign w6414 = ~w6380 & w6413 ;
  assign w6415 = w6411 | w6414 ;
  assign w6416 = ~\pi093 & w6415 ;
  assign w6417 = w6094 & w6380 ;
  assign w6418 = ~w6101 & w6349 ;
  assign w6419 = w6350 ^ w6418 ;
  assign w6420 = ~w6380 & w6419 ;
  assign w6421 = w6417 | w6420 ;
  assign w6422 = ~\pi092 & w6421 ;
  assign w6423 = w6100 & w6380 ;
  assign w6424 = ~w6107 & w6346 ;
  assign w6425 = w6347 ^ w6424 ;
  assign w6426 = ~w6380 & w6425 ;
  assign w6427 = w6423 | w6426 ;
  assign w6428 = ~\pi091 & w6427 ;
  assign w6429 = w6106 & w6380 ;
  assign w6430 = ~w6113 & w6343 ;
  assign w6431 = w6344 ^ w6430 ;
  assign w6432 = ~w6380 & w6431 ;
  assign w6433 = w6429 | w6432 ;
  assign w6434 = ~\pi090 & w6433 ;
  assign w6435 = w6112 & w6380 ;
  assign w6436 = ~w6119 & w6340 ;
  assign w6437 = w6341 ^ w6436 ;
  assign w6438 = ~w6380 & w6437 ;
  assign w6439 = w6435 | w6438 ;
  assign w6440 = ~\pi089 & w6439 ;
  assign w6441 = w6118 & w6380 ;
  assign w6442 = ~w6125 & w6337 ;
  assign w6443 = w6338 ^ w6442 ;
  assign w6444 = ~w6380 & w6443 ;
  assign w6445 = w6441 | w6444 ;
  assign w6446 = ~\pi088 & w6445 ;
  assign w6447 = w6124 & w6380 ;
  assign w6448 = ~w6131 & w6334 ;
  assign w6449 = w6335 ^ w6448 ;
  assign w6450 = ~w6380 & w6449 ;
  assign w6451 = w6447 | w6450 ;
  assign w6452 = ~\pi087 & w6451 ;
  assign w6453 = w6130 & w6380 ;
  assign w6454 = ~w6137 & w6331 ;
  assign w6455 = w6332 ^ w6454 ;
  assign w6456 = ~w6380 & w6455 ;
  assign w6457 = w6453 | w6456 ;
  assign w6458 = ~\pi086 & w6457 ;
  assign w6459 = w6136 & w6380 ;
  assign w6460 = ~w6143 & w6328 ;
  assign w6461 = w6329 ^ w6460 ;
  assign w6462 = ~w6380 & w6461 ;
  assign w6463 = w6459 | w6462 ;
  assign w6464 = ~\pi085 & w6463 ;
  assign w6465 = w6142 & w6380 ;
  assign w6466 = ~w6149 & w6325 ;
  assign w6467 = w6326 ^ w6466 ;
  assign w6468 = ~w6380 & w6467 ;
  assign w6469 = w6465 | w6468 ;
  assign w6470 = ~\pi084 & w6469 ;
  assign w6471 = w6148 & w6380 ;
  assign w6472 = ~w6155 & w6322 ;
  assign w6473 = w6323 ^ w6472 ;
  assign w6474 = ~w6380 & w6473 ;
  assign w6475 = w6471 | w6474 ;
  assign w6476 = ~\pi083 & w6475 ;
  assign w6477 = w6154 & w6380 ;
  assign w6478 = ~w6161 & w6319 ;
  assign w6479 = w6320 ^ w6478 ;
  assign w6480 = ~w6380 & w6479 ;
  assign w6481 = w6477 | w6480 ;
  assign w6482 = ~\pi082 & w6481 ;
  assign w6483 = w6160 & w6380 ;
  assign w6484 = ~w6167 & w6316 ;
  assign w6485 = w6317 ^ w6484 ;
  assign w6486 = ~w6380 & w6485 ;
  assign w6487 = w6483 | w6486 ;
  assign w6488 = ~\pi081 & w6487 ;
  assign w6489 = w6166 & w6380 ;
  assign w6490 = ~w6173 & w6313 ;
  assign w6491 = w6314 ^ w6490 ;
  assign w6492 = ~w6380 & w6491 ;
  assign w6493 = w6489 | w6492 ;
  assign w6494 = ~\pi080 & w6493 ;
  assign w6495 = w6172 & w6380 ;
  assign w6496 = ~w6179 & w6310 ;
  assign w6497 = w6311 ^ w6496 ;
  assign w6498 = ~w6380 & w6497 ;
  assign w6499 = w6495 | w6498 ;
  assign w6500 = ~\pi079 & w6499 ;
  assign w6501 = w6178 & w6380 ;
  assign w6502 = ~w6185 & w6307 ;
  assign w6503 = w6308 ^ w6502 ;
  assign w6504 = ~w6380 & w6503 ;
  assign w6505 = w6501 | w6504 ;
  assign w6506 = ~\pi078 & w6505 ;
  assign w6507 = w6184 & w6380 ;
  assign w6508 = ~w6191 & w6304 ;
  assign w6509 = w6305 ^ w6508 ;
  assign w6510 = ~w6380 & w6509 ;
  assign w6511 = w6507 | w6510 ;
  assign w6512 = ~\pi077 & w6511 ;
  assign w6513 = w6190 & w6380 ;
  assign w6514 = ~w6197 & w6301 ;
  assign w6515 = w6302 ^ w6514 ;
  assign w6516 = ~w6380 & w6515 ;
  assign w6517 = w6513 | w6516 ;
  assign w6518 = ~\pi076 & w6517 ;
  assign w6519 = w6196 & w6380 ;
  assign w6520 = ~w6203 & w6298 ;
  assign w6521 = w6299 ^ w6520 ;
  assign w6522 = ~w6380 & w6521 ;
  assign w6523 = w6519 | w6522 ;
  assign w6524 = ~\pi075 & w6523 ;
  assign w6525 = w6202 & w6380 ;
  assign w6526 = ~w6209 & w6295 ;
  assign w6527 = w6296 ^ w6526 ;
  assign w6528 = ~w6380 & w6527 ;
  assign w6529 = w6525 | w6528 ;
  assign w6530 = ~\pi074 & w6529 ;
  assign w6531 = w6208 & w6380 ;
  assign w6532 = ~w6215 & w6292 ;
  assign w6533 = w6293 ^ w6532 ;
  assign w6534 = ~w6380 & w6533 ;
  assign w6535 = w6531 | w6534 ;
  assign w6536 = ~\pi073 & w6535 ;
  assign w6537 = w6214 & w6380 ;
  assign w6538 = ~w6221 & w6289 ;
  assign w6539 = w6290 ^ w6538 ;
  assign w6540 = ~w6380 & w6539 ;
  assign w6541 = w6537 | w6540 ;
  assign w6542 = ~\pi072 & w6541 ;
  assign w6543 = w6220 & w6380 ;
  assign w6544 = ~w6227 & w6286 ;
  assign w6545 = w6287 ^ w6544 ;
  assign w6546 = ~w6380 & w6545 ;
  assign w6547 = w6543 | w6546 ;
  assign w6548 = ~\pi071 & w6547 ;
  assign w6549 = w6226 & w6380 ;
  assign w6550 = ~w6233 & w6283 ;
  assign w6551 = w6284 ^ w6550 ;
  assign w6552 = ~w6380 & w6551 ;
  assign w6553 = w6549 | w6552 ;
  assign w6554 = ~\pi070 & w6553 ;
  assign w6555 = w6232 & w6380 ;
  assign w6556 = ~w6241 & w6280 ;
  assign w6557 = w6281 ^ w6556 ;
  assign w6558 = ~w6380 & w6557 ;
  assign w6559 = w6555 | w6558 ;
  assign w6560 = ~\pi069 & w6559 ;
  assign w6561 = w6240 & w6380 ;
  assign w6562 = ~w6252 & w6277 ;
  assign w6563 = w6278 ^ w6562 ;
  assign w6564 = ~w6380 & w6563 ;
  assign w6565 = w6561 | w6564 ;
  assign w6566 = ~\pi068 & w6565 ;
  assign w6567 = w6251 & w6380 ;
  assign w6568 = ~w6268 & w6271 ;
  assign w6569 = ( \pi065 & w6271 ) | ( \pi065 & w6568 ) | ( w6271 & w6568 ) ;
  assign w6570 = w6274 ^ w6569 ;
  assign w6571 = ~w6380 & w6570 ;
  assign w6572 = w6567 | w6571 ;
  assign w6573 = ~\pi067 & w6572 ;
  assign w6574 = w6268 & w6380 ;
  assign w6575 = ( w6260 & w6267 ) | ( w6260 & ~w6379 ) | ( w6267 & ~w6379 ) ;
  assign w6576 = \pi065 ^ w6575 ;
  assign w6577 = ( w6269 & ~w6379 ) | ( w6269 & w6576 ) | ( ~w6379 & w6576 ) ;
  assign w6578 = ( w6269 & w6375 ) | ( w6269 & w6576 ) | ( w6375 & w6576 ) ;
  assign w6579 = w6577 & ~w6578 ;
  assign w6580 = w6574 | w6579 ;
  assign w6581 = ~\pi066 & w6580 ;
  assign w6582 = \pi064 & ~\pi099 ;
  assign w6583 = ~w202 & w6582 ;
  assign w6584 = ~w6046 & w6583 ;
  assign w6585 = ( \pi029 & w6375 ) | ( \pi029 & ~w6584 ) | ( w6375 & ~w6584 ) ;
  assign w6586 = \pi029 & w6585 ;
  assign w6587 = ( \pi099 & ~w278 ) | ( \pi099 & w6269 ) | ( ~w278 & w6269 ) ;
  assign w6588 = w275 | w288 ;
  assign w6589 = ( \pi099 & \pi100 ) | ( \pi099 & ~w288 ) | ( \pi100 & ~w288 ) ;
  assign w6590 = w6588 | w6589 ;
  assign w6591 = w6587 & ~w6590 ;
  assign w6592 = ~w6375 & w6591 ;
  assign w6593 = w6586 | w6592 ;
  assign w6594 = ~\pi028 & \pi064 ;
  assign w6595 = \pi065 ^ w6593 ;
  assign w6596 = w6594 | w6595 ;
  assign w6597 = \pi066 ^ w6580 ;
  assign w6598 = ~\pi065 & w6593 ;
  assign w6599 = w6596 | w6598 ;
  assign w6600 = ( w6597 & ~w6598 ) | ( w6597 & w6599 ) | ( ~w6598 & w6599 ) ;
  assign w6601 = \pi067 ^ w6572 ;
  assign w6602 = ( ~w6581 & w6600 ) | ( ~w6581 & w6601 ) | ( w6600 & w6601 ) ;
  assign w6603 = w6601 | w6602 ;
  assign w6604 = \pi068 ^ w6565 ;
  assign w6605 = ( ~w6573 & w6603 ) | ( ~w6573 & w6604 ) | ( w6603 & w6604 ) ;
  assign w6606 = w6604 | w6605 ;
  assign w6607 = \pi069 ^ w6559 ;
  assign w6608 = ( ~w6566 & w6606 ) | ( ~w6566 & w6607 ) | ( w6606 & w6607 ) ;
  assign w6609 = w6607 | w6608 ;
  assign w6610 = \pi070 ^ w6553 ;
  assign w6611 = ( ~w6560 & w6609 ) | ( ~w6560 & w6610 ) | ( w6609 & w6610 ) ;
  assign w6612 = w6610 | w6611 ;
  assign w6613 = \pi071 ^ w6547 ;
  assign w6614 = ( ~w6554 & w6612 ) | ( ~w6554 & w6613 ) | ( w6612 & w6613 ) ;
  assign w6615 = w6613 | w6614 ;
  assign w6616 = \pi072 ^ w6541 ;
  assign w6617 = ( ~w6548 & w6615 ) | ( ~w6548 & w6616 ) | ( w6615 & w6616 ) ;
  assign w6618 = w6616 | w6617 ;
  assign w6619 = \pi073 ^ w6535 ;
  assign w6620 = ( ~w6542 & w6618 ) | ( ~w6542 & w6619 ) | ( w6618 & w6619 ) ;
  assign w6621 = w6619 | w6620 ;
  assign w6622 = \pi074 ^ w6529 ;
  assign w6623 = ( ~w6536 & w6621 ) | ( ~w6536 & w6622 ) | ( w6621 & w6622 ) ;
  assign w6624 = w6622 | w6623 ;
  assign w6625 = \pi075 ^ w6523 ;
  assign w6626 = ( ~w6530 & w6624 ) | ( ~w6530 & w6625 ) | ( w6624 & w6625 ) ;
  assign w6627 = w6625 | w6626 ;
  assign w6628 = \pi076 ^ w6517 ;
  assign w6629 = ( ~w6524 & w6627 ) | ( ~w6524 & w6628 ) | ( w6627 & w6628 ) ;
  assign w6630 = w6628 | w6629 ;
  assign w6631 = \pi077 ^ w6511 ;
  assign w6632 = ( ~w6518 & w6630 ) | ( ~w6518 & w6631 ) | ( w6630 & w6631 ) ;
  assign w6633 = w6631 | w6632 ;
  assign w6634 = \pi078 ^ w6505 ;
  assign w6635 = ( ~w6512 & w6633 ) | ( ~w6512 & w6634 ) | ( w6633 & w6634 ) ;
  assign w6636 = w6634 | w6635 ;
  assign w6637 = \pi079 ^ w6499 ;
  assign w6638 = ( ~w6506 & w6636 ) | ( ~w6506 & w6637 ) | ( w6636 & w6637 ) ;
  assign w6639 = w6637 | w6638 ;
  assign w6640 = \pi080 ^ w6493 ;
  assign w6641 = ( ~w6500 & w6639 ) | ( ~w6500 & w6640 ) | ( w6639 & w6640 ) ;
  assign w6642 = w6640 | w6641 ;
  assign w6643 = \pi081 ^ w6487 ;
  assign w6644 = ( ~w6494 & w6642 ) | ( ~w6494 & w6643 ) | ( w6642 & w6643 ) ;
  assign w6645 = w6643 | w6644 ;
  assign w6646 = \pi082 ^ w6481 ;
  assign w6647 = ( ~w6488 & w6645 ) | ( ~w6488 & w6646 ) | ( w6645 & w6646 ) ;
  assign w6648 = w6646 | w6647 ;
  assign w6649 = \pi083 ^ w6475 ;
  assign w6650 = ( ~w6482 & w6648 ) | ( ~w6482 & w6649 ) | ( w6648 & w6649 ) ;
  assign w6651 = w6649 | w6650 ;
  assign w6652 = \pi084 ^ w6469 ;
  assign w6653 = ( ~w6476 & w6651 ) | ( ~w6476 & w6652 ) | ( w6651 & w6652 ) ;
  assign w6654 = w6652 | w6653 ;
  assign w6655 = \pi085 ^ w6463 ;
  assign w6656 = ( ~w6470 & w6654 ) | ( ~w6470 & w6655 ) | ( w6654 & w6655 ) ;
  assign w6657 = w6655 | w6656 ;
  assign w6658 = \pi086 ^ w6457 ;
  assign w6659 = ( ~w6464 & w6657 ) | ( ~w6464 & w6658 ) | ( w6657 & w6658 ) ;
  assign w6660 = w6658 | w6659 ;
  assign w6661 = \pi087 ^ w6451 ;
  assign w6662 = ( ~w6458 & w6660 ) | ( ~w6458 & w6661 ) | ( w6660 & w6661 ) ;
  assign w6663 = w6661 | w6662 ;
  assign w6664 = \pi088 ^ w6445 ;
  assign w6665 = ( ~w6452 & w6663 ) | ( ~w6452 & w6664 ) | ( w6663 & w6664 ) ;
  assign w6666 = w6664 | w6665 ;
  assign w6667 = \pi089 ^ w6439 ;
  assign w6668 = ( ~w6446 & w6666 ) | ( ~w6446 & w6667 ) | ( w6666 & w6667 ) ;
  assign w6669 = w6667 | w6668 ;
  assign w6670 = \pi090 ^ w6433 ;
  assign w6671 = ( ~w6440 & w6669 ) | ( ~w6440 & w6670 ) | ( w6669 & w6670 ) ;
  assign w6672 = w6670 | w6671 ;
  assign w6673 = \pi091 ^ w6427 ;
  assign w6674 = ( ~w6434 & w6672 ) | ( ~w6434 & w6673 ) | ( w6672 & w6673 ) ;
  assign w6675 = w6673 | w6674 ;
  assign w6676 = \pi092 ^ w6421 ;
  assign w6677 = ( ~w6428 & w6675 ) | ( ~w6428 & w6676 ) | ( w6675 & w6676 ) ;
  assign w6678 = w6676 | w6677 ;
  assign w6679 = \pi093 ^ w6415 ;
  assign w6680 = ( ~w6422 & w6678 ) | ( ~w6422 & w6679 ) | ( w6678 & w6679 ) ;
  assign w6681 = w6679 | w6680 ;
  assign w6682 = \pi094 ^ w6409 ;
  assign w6683 = ( ~w6416 & w6681 ) | ( ~w6416 & w6682 ) | ( w6681 & w6682 ) ;
  assign w6684 = w6682 | w6683 ;
  assign w6685 = \pi095 ^ w6403 ;
  assign w6686 = ( ~w6410 & w6684 ) | ( ~w6410 & w6685 ) | ( w6684 & w6685 ) ;
  assign w6687 = w6685 | w6686 ;
  assign w6688 = \pi096 ^ w6397 ;
  assign w6689 = ( ~w6404 & w6687 ) | ( ~w6404 & w6688 ) | ( w6687 & w6688 ) ;
  assign w6690 = w6688 | w6689 ;
  assign w6691 = \pi097 ^ w6391 ;
  assign w6692 = ( ~w6398 & w6690 ) | ( ~w6398 & w6691 ) | ( w6690 & w6691 ) ;
  assign w6693 = w6691 | w6692 ;
  assign w6694 = \pi098 ^ w6385 ;
  assign w6695 = ( ~w6392 & w6693 ) | ( ~w6392 & w6694 ) | ( w6693 & w6694 ) ;
  assign w6696 = w6694 | w6695 ;
  assign w6697 = w6058 & w6380 ;
  assign w6698 = ~w6059 & w6370 ;
  assign w6699 = w6371 ^ w6698 ;
  assign w6700 = ~w6380 & w6699 ;
  assign w6701 = w6697 | w6700 ;
  assign w6702 = ~\pi099 & w6701 ;
  assign w6703 = ( \pi099 & ~w6697 ) | ( \pi099 & w6700 ) | ( ~w6697 & w6700 ) ;
  assign w6704 = ~w6700 & w6703 ;
  assign w6705 = w6702 | w6704 ;
  assign w6706 = ( ~w6386 & w6696 ) | ( ~w6386 & w6705 ) | ( w6696 & w6705 ) ;
  assign w6707 = ( w368 & ~w6705 ) | ( w368 & w6706 ) | ( ~w6705 & w6706 ) ;
  assign w6708 = w6705 | w6707 ;
  assign w6709 = ~w6379 & w6701 ;
  assign w6710 = w6708 & ~w6709 ;
  assign w6711 = ~w6392 & w6693 ;
  assign w6712 = w6694 ^ w6711 ;
  assign w6713 = ~w6710 & w6712 ;
  assign w6714 = ( w6385 & w6708 ) | ( w6385 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6715 = ~w6709 & w6714 ;
  assign w6716 = w6713 | w6715 ;
  assign w6717 = ( ~w6386 & w6696 ) | ( ~w6386 & w6710 ) | ( w6696 & w6710 ) ;
  assign w6718 = w6705 ^ w6717 ;
  assign w6719 = ~w6710 & w6718 ;
  assign w6720 = ( w6379 & ~w6701 ) | ( w6379 & w6708 ) | ( ~w6701 & w6708 ) ;
  assign w6721 = w6701 & w6720 ;
  assign w6722 = w6719 | w6721 ;
  assign w6723 = ~\pi099 & w6716 ;
  assign w6724 = ~w6398 & w6690 ;
  assign w6725 = w6691 ^ w6724 ;
  assign w6726 = ~w6710 & w6725 ;
  assign w6727 = ( w6391 & w6708 ) | ( w6391 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6728 = ~w6709 & w6727 ;
  assign w6729 = w6726 | w6728 ;
  assign w6730 = ~\pi098 & w6729 ;
  assign w6731 = ~w6404 & w6687 ;
  assign w6732 = w6688 ^ w6731 ;
  assign w6733 = ~w6710 & w6732 ;
  assign w6734 = ( w6397 & w6708 ) | ( w6397 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6735 = ~w6709 & w6734 ;
  assign w6736 = w6733 | w6735 ;
  assign w6737 = ~\pi097 & w6736 ;
  assign w6738 = ~w6410 & w6684 ;
  assign w6739 = w6685 ^ w6738 ;
  assign w6740 = ~w6710 & w6739 ;
  assign w6741 = ( w6403 & w6708 ) | ( w6403 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6742 = ~w6709 & w6741 ;
  assign w6743 = w6740 | w6742 ;
  assign w6744 = ~\pi096 & w6743 ;
  assign w6745 = ~w6416 & w6681 ;
  assign w6746 = w6682 ^ w6745 ;
  assign w6747 = ~w6710 & w6746 ;
  assign w6748 = ( w6409 & w6708 ) | ( w6409 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6749 = ~w6709 & w6748 ;
  assign w6750 = w6747 | w6749 ;
  assign w6751 = ~\pi095 & w6750 ;
  assign w6752 = ~w6422 & w6678 ;
  assign w6753 = w6679 ^ w6752 ;
  assign w6754 = ~w6710 & w6753 ;
  assign w6755 = ( w6415 & w6708 ) | ( w6415 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6756 = ~w6709 & w6755 ;
  assign w6757 = w6754 | w6756 ;
  assign w6758 = ~\pi094 & w6757 ;
  assign w6759 = ~w6428 & w6675 ;
  assign w6760 = w6676 ^ w6759 ;
  assign w6761 = ~w6710 & w6760 ;
  assign w6762 = ( w6421 & w6708 ) | ( w6421 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6763 = ~w6709 & w6762 ;
  assign w6764 = w6761 | w6763 ;
  assign w6765 = ~\pi093 & w6764 ;
  assign w6766 = ~w6434 & w6672 ;
  assign w6767 = w6673 ^ w6766 ;
  assign w6768 = ~w6710 & w6767 ;
  assign w6769 = ( w6427 & w6708 ) | ( w6427 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6770 = ~w6709 & w6769 ;
  assign w6771 = w6768 | w6770 ;
  assign w6772 = ~\pi092 & w6771 ;
  assign w6773 = ~w6440 & w6669 ;
  assign w6774 = w6670 ^ w6773 ;
  assign w6775 = ~w6710 & w6774 ;
  assign w6776 = ( w6433 & w6708 ) | ( w6433 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6777 = ~w6709 & w6776 ;
  assign w6778 = w6775 | w6777 ;
  assign w6779 = ~\pi091 & w6778 ;
  assign w6780 = ~w6446 & w6666 ;
  assign w6781 = w6667 ^ w6780 ;
  assign w6782 = ~w6710 & w6781 ;
  assign w6783 = ( w6439 & w6708 ) | ( w6439 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6784 = ~w6709 & w6783 ;
  assign w6785 = w6782 | w6784 ;
  assign w6786 = ~\pi090 & w6785 ;
  assign w6787 = ~w6452 & w6663 ;
  assign w6788 = w6664 ^ w6787 ;
  assign w6789 = ~w6710 & w6788 ;
  assign w6790 = ( w6445 & w6708 ) | ( w6445 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6791 = ~w6709 & w6790 ;
  assign w6792 = w6789 | w6791 ;
  assign w6793 = ~\pi089 & w6792 ;
  assign w6794 = ~w6458 & w6660 ;
  assign w6795 = w6661 ^ w6794 ;
  assign w6796 = ~w6710 & w6795 ;
  assign w6797 = ( w6451 & w6708 ) | ( w6451 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6798 = ~w6709 & w6797 ;
  assign w6799 = w6796 | w6798 ;
  assign w6800 = ~\pi088 & w6799 ;
  assign w6801 = ~w6464 & w6657 ;
  assign w6802 = w6658 ^ w6801 ;
  assign w6803 = ~w6710 & w6802 ;
  assign w6804 = ( w6457 & w6708 ) | ( w6457 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6805 = ~w6709 & w6804 ;
  assign w6806 = w6803 | w6805 ;
  assign w6807 = ~\pi087 & w6806 ;
  assign w6808 = ~w6470 & w6654 ;
  assign w6809 = w6655 ^ w6808 ;
  assign w6810 = ~w6710 & w6809 ;
  assign w6811 = ( w6463 & w6708 ) | ( w6463 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6812 = ~w6709 & w6811 ;
  assign w6813 = w6810 | w6812 ;
  assign w6814 = ~\pi086 & w6813 ;
  assign w6815 = ~w6476 & w6651 ;
  assign w6816 = w6652 ^ w6815 ;
  assign w6817 = ~w6710 & w6816 ;
  assign w6818 = ( w6469 & w6708 ) | ( w6469 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6819 = ~w6709 & w6818 ;
  assign w6820 = w6817 | w6819 ;
  assign w6821 = ~\pi085 & w6820 ;
  assign w6822 = ~w6482 & w6648 ;
  assign w6823 = w6649 ^ w6822 ;
  assign w6824 = ~w6710 & w6823 ;
  assign w6825 = ( w6475 & w6708 ) | ( w6475 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6826 = ~w6709 & w6825 ;
  assign w6827 = w6824 | w6826 ;
  assign w6828 = ~\pi084 & w6827 ;
  assign w6829 = ~w6488 & w6645 ;
  assign w6830 = w6646 ^ w6829 ;
  assign w6831 = ~w6710 & w6830 ;
  assign w6832 = ( w6481 & w6708 ) | ( w6481 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6833 = ~w6709 & w6832 ;
  assign w6834 = w6831 | w6833 ;
  assign w6835 = ~\pi083 & w6834 ;
  assign w6836 = ~w6494 & w6642 ;
  assign w6837 = w6643 ^ w6836 ;
  assign w6838 = ~w6710 & w6837 ;
  assign w6839 = ( w6487 & w6708 ) | ( w6487 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6840 = ~w6709 & w6839 ;
  assign w6841 = w6838 | w6840 ;
  assign w6842 = ~\pi082 & w6841 ;
  assign w6843 = ~w6500 & w6639 ;
  assign w6844 = w6640 ^ w6843 ;
  assign w6845 = ~w6710 & w6844 ;
  assign w6846 = ( w6493 & w6708 ) | ( w6493 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6847 = ~w6709 & w6846 ;
  assign w6848 = w6845 | w6847 ;
  assign w6849 = ~\pi081 & w6848 ;
  assign w6850 = ~w6506 & w6636 ;
  assign w6851 = w6637 ^ w6850 ;
  assign w6852 = ~w6710 & w6851 ;
  assign w6853 = ( w6499 & w6708 ) | ( w6499 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6854 = ~w6709 & w6853 ;
  assign w6855 = w6852 | w6854 ;
  assign w6856 = ~\pi080 & w6855 ;
  assign w6857 = ~w6512 & w6633 ;
  assign w6858 = w6634 ^ w6857 ;
  assign w6859 = ~w6710 & w6858 ;
  assign w6860 = ( w6505 & w6708 ) | ( w6505 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6861 = ~w6709 & w6860 ;
  assign w6862 = w6859 | w6861 ;
  assign w6863 = ~\pi079 & w6862 ;
  assign w6864 = ~w6518 & w6630 ;
  assign w6865 = w6631 ^ w6864 ;
  assign w6866 = ~w6710 & w6865 ;
  assign w6867 = ( w6511 & w6708 ) | ( w6511 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6868 = ~w6709 & w6867 ;
  assign w6869 = w6866 | w6868 ;
  assign w6870 = ~\pi078 & w6869 ;
  assign w6871 = ~w6524 & w6627 ;
  assign w6872 = w6628 ^ w6871 ;
  assign w6873 = ~w6710 & w6872 ;
  assign w6874 = ( w6517 & w6708 ) | ( w6517 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6875 = ~w6709 & w6874 ;
  assign w6876 = w6873 | w6875 ;
  assign w6877 = ~\pi077 & w6876 ;
  assign w6878 = ~w6530 & w6624 ;
  assign w6879 = w6625 ^ w6878 ;
  assign w6880 = ~w6710 & w6879 ;
  assign w6881 = ( w6523 & w6708 ) | ( w6523 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6882 = ~w6709 & w6881 ;
  assign w6883 = w6880 | w6882 ;
  assign w6884 = ~\pi076 & w6883 ;
  assign w6885 = ~w6536 & w6621 ;
  assign w6886 = w6622 ^ w6885 ;
  assign w6887 = ~w6710 & w6886 ;
  assign w6888 = ( w6529 & w6708 ) | ( w6529 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6889 = ~w6709 & w6888 ;
  assign w6890 = w6887 | w6889 ;
  assign w6891 = ~\pi075 & w6890 ;
  assign w6892 = ~w6542 & w6618 ;
  assign w6893 = w6619 ^ w6892 ;
  assign w6894 = ~w6710 & w6893 ;
  assign w6895 = ( w6535 & w6708 ) | ( w6535 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6896 = ~w6709 & w6895 ;
  assign w6897 = w6894 | w6896 ;
  assign w6898 = ~\pi074 & w6897 ;
  assign w6899 = ~w6548 & w6615 ;
  assign w6900 = w6616 ^ w6899 ;
  assign w6901 = ~w6710 & w6900 ;
  assign w6902 = ( w6541 & w6708 ) | ( w6541 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6903 = ~w6709 & w6902 ;
  assign w6904 = w6901 | w6903 ;
  assign w6905 = ~\pi073 & w6904 ;
  assign w6906 = ~w6554 & w6612 ;
  assign w6907 = w6613 ^ w6906 ;
  assign w6908 = ~w6710 & w6907 ;
  assign w6909 = ( w6547 & w6708 ) | ( w6547 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6910 = ~w6709 & w6909 ;
  assign w6911 = w6908 | w6910 ;
  assign w6912 = ~\pi072 & w6911 ;
  assign w6913 = ~w6560 & w6609 ;
  assign w6914 = w6610 ^ w6913 ;
  assign w6915 = ~w6710 & w6914 ;
  assign w6916 = ( w6553 & w6708 ) | ( w6553 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6917 = ~w6709 & w6916 ;
  assign w6918 = w6915 | w6917 ;
  assign w6919 = ~\pi071 & w6918 ;
  assign w6920 = ~w6566 & w6606 ;
  assign w6921 = w6607 ^ w6920 ;
  assign w6922 = ~w6710 & w6921 ;
  assign w6923 = ( w6559 & w6708 ) | ( w6559 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6924 = ~w6709 & w6923 ;
  assign w6925 = w6922 | w6924 ;
  assign w6926 = ~\pi070 & w6925 ;
  assign w6927 = ~w6573 & w6603 ;
  assign w6928 = w6604 ^ w6927 ;
  assign w6929 = ~w6710 & w6928 ;
  assign w6930 = ( w6565 & w6708 ) | ( w6565 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6931 = ~w6709 & w6930 ;
  assign w6932 = w6929 | w6931 ;
  assign w6933 = ~\pi069 & w6932 ;
  assign w6934 = ~w6581 & w6600 ;
  assign w6935 = w6601 ^ w6934 ;
  assign w6936 = ~w6710 & w6935 ;
  assign w6937 = ( w6572 & w6708 ) | ( w6572 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6938 = ~w6709 & w6937 ;
  assign w6939 = w6936 | w6938 ;
  assign w6940 = ~\pi068 & w6939 ;
  assign w6941 = ( \pi065 & w6593 ) | ( \pi065 & ~w6710 ) | ( w6593 & ~w6710 ) ;
  assign w6942 = ( \pi065 & w6596 ) | ( \pi065 & ~w6941 ) | ( w6596 & ~w6941 ) ;
  assign w6943 = w6597 ^ w6942 ;
  assign w6944 = ~w6710 & w6943 ;
  assign w6945 = ( w6580 & w6708 ) | ( w6580 & w6709 ) | ( w6708 & w6709 ) ;
  assign w6946 = ~w6709 & w6945 ;
  assign w6947 = w6944 | w6946 ;
  assign w6948 = ~\pi067 & w6947 ;
  assign w6949 = w6593 ^ w6594 ;
  assign w6950 = \pi065 ^ w6949 ;
  assign w6951 = w6710 ^ w6950 ;
  assign w6952 = ( w6593 & w6950 ) | ( w6593 & w6951 ) | ( w6950 & w6951 ) ;
  assign w6953 = ~\pi066 & w6952 ;
  assign w6954 = w6593 ^ w6710 ;
  assign w6955 = ( w6593 & w6950 ) | ( w6593 & ~w6954 ) | ( w6950 & ~w6954 ) ;
  assign w6956 = \pi066 ^ w6955 ;
  assign w6957 = \pi064 & ~w6710 ;
  assign w6958 = \pi028 ^ w6957 ;
  assign w6959 = ( ~\pi027 & \pi064 ) | ( ~\pi027 & w6956 ) | ( \pi064 & w6956 ) ;
  assign w6960 = ( \pi065 & ~w6958 ) | ( \pi065 & w6959 ) | ( ~w6958 & w6959 ) ;
  assign w6961 = w6956 | w6960 ;
  assign w6962 = \pi067 ^ w6947 ;
  assign w6963 = ( ~w6953 & w6961 ) | ( ~w6953 & w6962 ) | ( w6961 & w6962 ) ;
  assign w6964 = w6962 | w6963 ;
  assign w6965 = \pi068 ^ w6939 ;
  assign w6966 = ( ~w6948 & w6964 ) | ( ~w6948 & w6965 ) | ( w6964 & w6965 ) ;
  assign w6967 = w6965 | w6966 ;
  assign w6968 = \pi069 ^ w6932 ;
  assign w6969 = ( ~w6940 & w6967 ) | ( ~w6940 & w6968 ) | ( w6967 & w6968 ) ;
  assign w6970 = w6968 | w6969 ;
  assign w6971 = \pi070 ^ w6925 ;
  assign w6972 = ( ~w6933 & w6970 ) | ( ~w6933 & w6971 ) | ( w6970 & w6971 ) ;
  assign w6973 = w6971 | w6972 ;
  assign w6974 = \pi071 ^ w6918 ;
  assign w6975 = ( ~w6926 & w6973 ) | ( ~w6926 & w6974 ) | ( w6973 & w6974 ) ;
  assign w6976 = w6974 | w6975 ;
  assign w6977 = \pi072 ^ w6911 ;
  assign w6978 = ( ~w6919 & w6976 ) | ( ~w6919 & w6977 ) | ( w6976 & w6977 ) ;
  assign w6979 = w6977 | w6978 ;
  assign w6980 = \pi073 ^ w6904 ;
  assign w6981 = ( ~w6912 & w6979 ) | ( ~w6912 & w6980 ) | ( w6979 & w6980 ) ;
  assign w6982 = w6980 | w6981 ;
  assign w6983 = \pi074 ^ w6897 ;
  assign w6984 = ( ~w6905 & w6982 ) | ( ~w6905 & w6983 ) | ( w6982 & w6983 ) ;
  assign w6985 = w6983 | w6984 ;
  assign w6986 = \pi075 ^ w6890 ;
  assign w6987 = ( ~w6898 & w6985 ) | ( ~w6898 & w6986 ) | ( w6985 & w6986 ) ;
  assign w6988 = w6986 | w6987 ;
  assign w6989 = \pi076 ^ w6883 ;
  assign w6990 = ( ~w6891 & w6988 ) | ( ~w6891 & w6989 ) | ( w6988 & w6989 ) ;
  assign w6991 = w6989 | w6990 ;
  assign w6992 = \pi077 ^ w6876 ;
  assign w6993 = ( ~w6884 & w6991 ) | ( ~w6884 & w6992 ) | ( w6991 & w6992 ) ;
  assign w6994 = w6992 | w6993 ;
  assign w6995 = \pi078 ^ w6869 ;
  assign w6996 = ( ~w6877 & w6994 ) | ( ~w6877 & w6995 ) | ( w6994 & w6995 ) ;
  assign w6997 = w6995 | w6996 ;
  assign w6998 = \pi079 ^ w6862 ;
  assign w6999 = ( ~w6870 & w6997 ) | ( ~w6870 & w6998 ) | ( w6997 & w6998 ) ;
  assign w7000 = w6998 | w6999 ;
  assign w7001 = \pi080 ^ w6855 ;
  assign w7002 = ( ~w6863 & w7000 ) | ( ~w6863 & w7001 ) | ( w7000 & w7001 ) ;
  assign w7003 = w7001 | w7002 ;
  assign w7004 = \pi081 ^ w6848 ;
  assign w7005 = ( ~w6856 & w7003 ) | ( ~w6856 & w7004 ) | ( w7003 & w7004 ) ;
  assign w7006 = w7004 | w7005 ;
  assign w7007 = \pi082 ^ w6841 ;
  assign w7008 = ( ~w6849 & w7006 ) | ( ~w6849 & w7007 ) | ( w7006 & w7007 ) ;
  assign w7009 = w7007 | w7008 ;
  assign w7010 = \pi083 ^ w6834 ;
  assign w7011 = ( ~w6842 & w7009 ) | ( ~w6842 & w7010 ) | ( w7009 & w7010 ) ;
  assign w7012 = w7010 | w7011 ;
  assign w7013 = \pi084 ^ w6827 ;
  assign w7014 = ( ~w6835 & w7012 ) | ( ~w6835 & w7013 ) | ( w7012 & w7013 ) ;
  assign w7015 = w7013 | w7014 ;
  assign w7016 = \pi085 ^ w6820 ;
  assign w7017 = ( ~w6828 & w7015 ) | ( ~w6828 & w7016 ) | ( w7015 & w7016 ) ;
  assign w7018 = w7016 | w7017 ;
  assign w7019 = \pi086 ^ w6813 ;
  assign w7020 = ( ~w6821 & w7018 ) | ( ~w6821 & w7019 ) | ( w7018 & w7019 ) ;
  assign w7021 = w7019 | w7020 ;
  assign w7022 = \pi087 ^ w6806 ;
  assign w7023 = ( ~w6814 & w7021 ) | ( ~w6814 & w7022 ) | ( w7021 & w7022 ) ;
  assign w7024 = w7022 | w7023 ;
  assign w7025 = \pi088 ^ w6799 ;
  assign w7026 = ( ~w6807 & w7024 ) | ( ~w6807 & w7025 ) | ( w7024 & w7025 ) ;
  assign w7027 = w7025 | w7026 ;
  assign w7028 = \pi089 ^ w6792 ;
  assign w7029 = ( ~w6800 & w7027 ) | ( ~w6800 & w7028 ) | ( w7027 & w7028 ) ;
  assign w7030 = w7028 | w7029 ;
  assign w7031 = \pi090 ^ w6785 ;
  assign w7032 = ( ~w6793 & w7030 ) | ( ~w6793 & w7031 ) | ( w7030 & w7031 ) ;
  assign w7033 = w7031 | w7032 ;
  assign w7034 = \pi091 ^ w6778 ;
  assign w7035 = ( ~w6786 & w7033 ) | ( ~w6786 & w7034 ) | ( w7033 & w7034 ) ;
  assign w7036 = w7034 | w7035 ;
  assign w7037 = \pi092 ^ w6771 ;
  assign w7038 = ( ~w6779 & w7036 ) | ( ~w6779 & w7037 ) | ( w7036 & w7037 ) ;
  assign w7039 = w7037 | w7038 ;
  assign w7040 = \pi093 ^ w6764 ;
  assign w7041 = ( ~w6772 & w7039 ) | ( ~w6772 & w7040 ) | ( w7039 & w7040 ) ;
  assign w7042 = w7040 | w7041 ;
  assign w7043 = \pi094 ^ w6757 ;
  assign w7044 = ( ~w6765 & w7042 ) | ( ~w6765 & w7043 ) | ( w7042 & w7043 ) ;
  assign w7045 = w7043 | w7044 ;
  assign w7046 = \pi095 ^ w6750 ;
  assign w7047 = ( ~w6758 & w7045 ) | ( ~w6758 & w7046 ) | ( w7045 & w7046 ) ;
  assign w7048 = w7046 | w7047 ;
  assign w7049 = \pi096 ^ w6743 ;
  assign w7050 = ( ~w6751 & w7048 ) | ( ~w6751 & w7049 ) | ( w7048 & w7049 ) ;
  assign w7051 = w7049 | w7050 ;
  assign w7052 = \pi097 ^ w6736 ;
  assign w7053 = ( ~w6744 & w7051 ) | ( ~w6744 & w7052 ) | ( w7051 & w7052 ) ;
  assign w7054 = w7052 | w7053 ;
  assign w7055 = \pi098 ^ w6729 ;
  assign w7056 = ( ~w6737 & w7054 ) | ( ~w6737 & w7055 ) | ( w7054 & w7055 ) ;
  assign w7057 = w7055 | w7056 ;
  assign w7058 = \pi099 ^ w6716 ;
  assign w7059 = ( ~w6730 & w7057 ) | ( ~w6730 & w7058 ) | ( w7057 & w7058 ) ;
  assign w7060 = w7058 | w7059 ;
  assign w7061 = \pi100 ^ w6722 ;
  assign w7062 = w6723 & ~w7061 ;
  assign w7063 = ( w7060 & w7061 ) | ( w7060 & ~w7062 ) | ( w7061 & ~w7062 ) ;
  assign w7064 = ~\pi100 & w6722 ;
  assign w7065 = w7063 & ~w7064 ;
  assign w7066 = w452 | w7065 ;
  assign w7067 = w6716 & w7066 ;
  assign w7068 = ~w6730 & w7057 ;
  assign w7069 = w7058 ^ w7068 ;
  assign w7070 = ~w7066 & w7069 ;
  assign w7071 = w7067 | w7070 ;
  assign w7072 = w6722 & w7066 ;
  assign w7073 = ~w6723 & w7060 ;
  assign w7074 = w7061 ^ w7073 ;
  assign w7075 = ~w7066 & w7074 ;
  assign w7076 = w7072 | w7075 ;
  assign w7077 = ~\pi100 & w7071 ;
  assign w7078 = w6729 & w7066 ;
  assign w7079 = ~w6737 & w7054 ;
  assign w7080 = w7055 ^ w7079 ;
  assign w7081 = ~w7066 & w7080 ;
  assign w7082 = w7078 | w7081 ;
  assign w7083 = ~\pi099 & w7082 ;
  assign w7084 = w6736 & w7066 ;
  assign w7085 = ~w6744 & w7051 ;
  assign w7086 = w7052 ^ w7085 ;
  assign w7087 = ~w7066 & w7086 ;
  assign w7088 = w7084 | w7087 ;
  assign w7089 = ~\pi098 & w7088 ;
  assign w7090 = w6743 & w7066 ;
  assign w7091 = ~w6751 & w7048 ;
  assign w7092 = w7049 ^ w7091 ;
  assign w7093 = ~w7066 & w7092 ;
  assign w7094 = w7090 | w7093 ;
  assign w7095 = ~\pi097 & w7094 ;
  assign w7096 = w6750 & w7066 ;
  assign w7097 = ~w6758 & w7045 ;
  assign w7098 = w7046 ^ w7097 ;
  assign w7099 = ~w7066 & w7098 ;
  assign w7100 = w7096 | w7099 ;
  assign w7101 = ~\pi096 & w7100 ;
  assign w7102 = w6757 & w7066 ;
  assign w7103 = ~w6765 & w7042 ;
  assign w7104 = w7043 ^ w7103 ;
  assign w7105 = ~w7066 & w7104 ;
  assign w7106 = w7102 | w7105 ;
  assign w7107 = ~\pi095 & w7106 ;
  assign w7108 = w6764 & w7066 ;
  assign w7109 = ~w6772 & w7039 ;
  assign w7110 = w7040 ^ w7109 ;
  assign w7111 = ~w7066 & w7110 ;
  assign w7112 = w7108 | w7111 ;
  assign w7113 = ~\pi094 & w7112 ;
  assign w7114 = w6771 & w7066 ;
  assign w7115 = ~w6779 & w7036 ;
  assign w7116 = w7037 ^ w7115 ;
  assign w7117 = ~w7066 & w7116 ;
  assign w7118 = w7114 | w7117 ;
  assign w7119 = ~\pi093 & w7118 ;
  assign w7120 = w6778 & w7066 ;
  assign w7121 = ~w6786 & w7033 ;
  assign w7122 = w7034 ^ w7121 ;
  assign w7123 = ~w7066 & w7122 ;
  assign w7124 = w7120 | w7123 ;
  assign w7125 = ~\pi092 & w7124 ;
  assign w7126 = w6785 & w7066 ;
  assign w7127 = ~w6793 & w7030 ;
  assign w7128 = w7031 ^ w7127 ;
  assign w7129 = ~w7066 & w7128 ;
  assign w7130 = w7126 | w7129 ;
  assign w7131 = ~\pi091 & w7130 ;
  assign w7132 = w6792 & w7066 ;
  assign w7133 = ~w6800 & w7027 ;
  assign w7134 = w7028 ^ w7133 ;
  assign w7135 = ~w7066 & w7134 ;
  assign w7136 = w7132 | w7135 ;
  assign w7137 = ~\pi090 & w7136 ;
  assign w7138 = w6799 & w7066 ;
  assign w7139 = ~w6807 & w7024 ;
  assign w7140 = w7025 ^ w7139 ;
  assign w7141 = ~w7066 & w7140 ;
  assign w7142 = w7138 | w7141 ;
  assign w7143 = ~\pi089 & w7142 ;
  assign w7144 = w6806 & w7066 ;
  assign w7145 = ~w6814 & w7021 ;
  assign w7146 = w7022 ^ w7145 ;
  assign w7147 = ~w7066 & w7146 ;
  assign w7148 = w7144 | w7147 ;
  assign w7149 = ~\pi088 & w7148 ;
  assign w7150 = w6813 & w7066 ;
  assign w7151 = ~w6821 & w7018 ;
  assign w7152 = w7019 ^ w7151 ;
  assign w7153 = ~w7066 & w7152 ;
  assign w7154 = w7150 | w7153 ;
  assign w7155 = ~\pi087 & w7154 ;
  assign w7156 = w6820 & w7066 ;
  assign w7157 = ~w6828 & w7015 ;
  assign w7158 = w7016 ^ w7157 ;
  assign w7159 = ~w7066 & w7158 ;
  assign w7160 = w7156 | w7159 ;
  assign w7161 = ~\pi086 & w7160 ;
  assign w7162 = w6827 & w7066 ;
  assign w7163 = ~w6835 & w7012 ;
  assign w7164 = w7013 ^ w7163 ;
  assign w7165 = ~w7066 & w7164 ;
  assign w7166 = w7162 | w7165 ;
  assign w7167 = ~\pi085 & w7166 ;
  assign w7168 = w6834 & w7066 ;
  assign w7169 = ~w6842 & w7009 ;
  assign w7170 = w7010 ^ w7169 ;
  assign w7171 = ~w7066 & w7170 ;
  assign w7172 = w7168 | w7171 ;
  assign w7173 = ~\pi084 & w7172 ;
  assign w7174 = w6841 & w7066 ;
  assign w7175 = ~w6849 & w7006 ;
  assign w7176 = w7007 ^ w7175 ;
  assign w7177 = ~w7066 & w7176 ;
  assign w7178 = w7174 | w7177 ;
  assign w7179 = ~\pi083 & w7178 ;
  assign w7180 = w6848 & w7066 ;
  assign w7181 = ~w6856 & w7003 ;
  assign w7182 = w7004 ^ w7181 ;
  assign w7183 = ~w7066 & w7182 ;
  assign w7184 = w7180 | w7183 ;
  assign w7185 = ~\pi082 & w7184 ;
  assign w7186 = w6855 & w7066 ;
  assign w7187 = ~w6863 & w7000 ;
  assign w7188 = w7001 ^ w7187 ;
  assign w7189 = ~w7066 & w7188 ;
  assign w7190 = w7186 | w7189 ;
  assign w7191 = ~\pi081 & w7190 ;
  assign w7192 = w6862 & w7066 ;
  assign w7193 = ~w6870 & w6997 ;
  assign w7194 = w6998 ^ w7193 ;
  assign w7195 = ~w7066 & w7194 ;
  assign w7196 = w7192 | w7195 ;
  assign w7197 = ~\pi080 & w7196 ;
  assign w7198 = w6869 & w7066 ;
  assign w7199 = ~w6877 & w6994 ;
  assign w7200 = w6995 ^ w7199 ;
  assign w7201 = ~w7066 & w7200 ;
  assign w7202 = w7198 | w7201 ;
  assign w7203 = ~\pi079 & w7202 ;
  assign w7204 = w6876 & w7066 ;
  assign w7205 = ~w6884 & w6991 ;
  assign w7206 = w6992 ^ w7205 ;
  assign w7207 = ~w7066 & w7206 ;
  assign w7208 = w7204 | w7207 ;
  assign w7209 = ~\pi078 & w7208 ;
  assign w7210 = w6883 & w7066 ;
  assign w7211 = ~w6891 & w6988 ;
  assign w7212 = w6989 ^ w7211 ;
  assign w7213 = ~w7066 & w7212 ;
  assign w7214 = w7210 | w7213 ;
  assign w7215 = ~\pi077 & w7214 ;
  assign w7216 = w6890 & w7066 ;
  assign w7217 = ~w6898 & w6985 ;
  assign w7218 = w6986 ^ w7217 ;
  assign w7219 = ~w7066 & w7218 ;
  assign w7220 = w7216 | w7219 ;
  assign w7221 = ~\pi076 & w7220 ;
  assign w7222 = w6897 & w7066 ;
  assign w7223 = ~w6905 & w6982 ;
  assign w7224 = w6983 ^ w7223 ;
  assign w7225 = ~w7066 & w7224 ;
  assign w7226 = w7222 | w7225 ;
  assign w7227 = ~\pi075 & w7226 ;
  assign w7228 = w6904 & w7066 ;
  assign w7229 = ~w6912 & w6979 ;
  assign w7230 = w6980 ^ w7229 ;
  assign w7231 = ~w7066 & w7230 ;
  assign w7232 = w7228 | w7231 ;
  assign w7233 = ~\pi074 & w7232 ;
  assign w7234 = w6911 & w7066 ;
  assign w7235 = ~w6919 & w6976 ;
  assign w7236 = w6977 ^ w7235 ;
  assign w7237 = ~w7066 & w7236 ;
  assign w7238 = w7234 | w7237 ;
  assign w7239 = ~\pi073 & w7238 ;
  assign w7240 = w6918 & w7066 ;
  assign w7241 = ~w6926 & w6973 ;
  assign w7242 = w6974 ^ w7241 ;
  assign w7243 = ~w7066 & w7242 ;
  assign w7244 = w7240 | w7243 ;
  assign w7245 = ~\pi072 & w7244 ;
  assign w7246 = w6925 & w7066 ;
  assign w7247 = ~w6933 & w6970 ;
  assign w7248 = w6971 ^ w7247 ;
  assign w7249 = ~w7066 & w7248 ;
  assign w7250 = w7246 | w7249 ;
  assign w7251 = ~\pi071 & w7250 ;
  assign w7252 = w6932 & w7066 ;
  assign w7253 = ~w6940 & w6967 ;
  assign w7254 = w6968 ^ w7253 ;
  assign w7255 = ~w7066 & w7254 ;
  assign w7256 = w7252 | w7255 ;
  assign w7257 = ~\pi070 & w7256 ;
  assign w7258 = w6939 & w7066 ;
  assign w7259 = ~w6948 & w6964 ;
  assign w7260 = w6965 ^ w7259 ;
  assign w7261 = ~w7066 & w7260 ;
  assign w7262 = w7258 | w7261 ;
  assign w7263 = ~\pi069 & w7262 ;
  assign w7264 = w6947 & w7066 ;
  assign w7265 = ~w6953 & w6961 ;
  assign w7266 = w6962 ^ w7265 ;
  assign w7267 = ~w7066 & w7266 ;
  assign w7268 = w7264 | w7267 ;
  assign w7269 = ~\pi068 & w7268 ;
  assign w7270 = w6952 & w7066 ;
  assign w7271 = ~\pi027 & \pi064 ;
  assign w7272 = ( \pi065 & ~w6958 ) | ( \pi065 & w7271 ) | ( ~w6958 & w7271 ) ;
  assign w7273 = w6956 ^ w7272 ;
  assign w7274 = ( w452 & w7065 ) | ( w452 & w7273 ) | ( w7065 & w7273 ) ;
  assign w7275 = w7273 & ~w7274 ;
  assign w7276 = w7270 | w7275 ;
  assign w7277 = ~\pi067 & w7276 ;
  assign w7278 = \pi028 ^ \pi065 ;
  assign w7279 = \pi027 ^ w6710 ;
  assign w7280 = ( \pi064 & w452 ) | ( \pi064 & w7279 ) | ( w452 & w7279 ) ;
  assign w7281 = w7278 ^ w7280 ;
  assign w7282 = ~w452 & w7281 ;
  assign w7283 = ~w7065 & w7282 ;
  assign w7284 = ( ~\pi064 & w6710 ) | ( ~\pi064 & w7066 ) | ( w6710 & w7066 ) ;
  assign w7285 = \pi028 ^ w7284 ;
  assign w7286 = w7066 & ~w7285 ;
  assign w7287 = w7283 | w7286 ;
  assign w7288 = ~\pi066 & w7287 ;
  assign w7289 = ( \pi064 & ~\pi101 ) | ( \pi064 & \pi102 ) | ( ~\pi101 & \pi102 ) ;
  assign w7290 = w158 | w168 ;
  assign w7291 = ( \pi102 & \pi103 ) | ( \pi102 & ~w158 ) | ( \pi103 & ~w158 ) ;
  assign w7292 = w7290 | w7291 ;
  assign w7293 = w7289 & ~w7292 ;
  assign w7294 = ~w155 & w7293 ;
  assign w7295 = ( \pi027 & w7065 ) | ( \pi027 & ~w7294 ) | ( w7065 & ~w7294 ) ;
  assign w7296 = \pi027 & w7295 ;
  assign w7297 = ( ~\pi027 & w278 ) | ( ~\pi027 & w288 ) | ( w278 & w288 ) ;
  assign w7298 = w275 | w7065 ;
  assign w7299 = ( ~\pi027 & \pi064 ) | ( ~\pi027 & w275 ) | ( \pi064 & w275 ) ;
  assign w7300 = ~w7298 & w7299 ;
  assign w7301 = ~w7297 & w7300 ;
  assign w7302 = ~\pi026 & \pi064 ;
  assign w7303 = w7066 | w7283 ;
  assign w7304 = ( w6958 & w7283 ) | ( w6958 & w7303 ) | ( w7283 & w7303 ) ;
  assign w7305 = \pi066 ^ w7304 ;
  assign w7306 = w7296 | w7301 ;
  assign w7307 = ( \pi065 & w7302 ) | ( \pi065 & ~w7306 ) | ( w7302 & ~w7306 ) ;
  assign w7308 = w7305 | w7307 ;
  assign w7309 = \pi067 ^ w7276 ;
  assign w7310 = ( ~w7288 & w7308 ) | ( ~w7288 & w7309 ) | ( w7308 & w7309 ) ;
  assign w7311 = w7309 | w7310 ;
  assign w7312 = \pi068 ^ w7268 ;
  assign w7313 = ( ~w7277 & w7311 ) | ( ~w7277 & w7312 ) | ( w7311 & w7312 ) ;
  assign w7314 = w7312 | w7313 ;
  assign w7315 = \pi069 ^ w7262 ;
  assign w7316 = ( ~w7269 & w7314 ) | ( ~w7269 & w7315 ) | ( w7314 & w7315 ) ;
  assign w7317 = w7315 | w7316 ;
  assign w7318 = \pi070 ^ w7256 ;
  assign w7319 = ( ~w7263 & w7317 ) | ( ~w7263 & w7318 ) | ( w7317 & w7318 ) ;
  assign w7320 = w7318 | w7319 ;
  assign w7321 = \pi071 ^ w7250 ;
  assign w7322 = ( ~w7257 & w7320 ) | ( ~w7257 & w7321 ) | ( w7320 & w7321 ) ;
  assign w7323 = w7321 | w7322 ;
  assign w7324 = \pi072 ^ w7244 ;
  assign w7325 = ( ~w7251 & w7323 ) | ( ~w7251 & w7324 ) | ( w7323 & w7324 ) ;
  assign w7326 = w7324 | w7325 ;
  assign w7327 = \pi073 ^ w7238 ;
  assign w7328 = ( ~w7245 & w7326 ) | ( ~w7245 & w7327 ) | ( w7326 & w7327 ) ;
  assign w7329 = w7327 | w7328 ;
  assign w7330 = \pi074 ^ w7232 ;
  assign w7331 = ( ~w7239 & w7329 ) | ( ~w7239 & w7330 ) | ( w7329 & w7330 ) ;
  assign w7332 = w7330 | w7331 ;
  assign w7333 = \pi075 ^ w7226 ;
  assign w7334 = ( ~w7233 & w7332 ) | ( ~w7233 & w7333 ) | ( w7332 & w7333 ) ;
  assign w7335 = w7333 | w7334 ;
  assign w7336 = \pi076 ^ w7220 ;
  assign w7337 = ( ~w7227 & w7335 ) | ( ~w7227 & w7336 ) | ( w7335 & w7336 ) ;
  assign w7338 = w7336 | w7337 ;
  assign w7339 = \pi077 ^ w7214 ;
  assign w7340 = ( ~w7221 & w7338 ) | ( ~w7221 & w7339 ) | ( w7338 & w7339 ) ;
  assign w7341 = w7339 | w7340 ;
  assign w7342 = \pi078 ^ w7208 ;
  assign w7343 = ( ~w7215 & w7341 ) | ( ~w7215 & w7342 ) | ( w7341 & w7342 ) ;
  assign w7344 = w7342 | w7343 ;
  assign w7345 = \pi079 ^ w7202 ;
  assign w7346 = ( ~w7209 & w7344 ) | ( ~w7209 & w7345 ) | ( w7344 & w7345 ) ;
  assign w7347 = w7345 | w7346 ;
  assign w7348 = \pi080 ^ w7196 ;
  assign w7349 = ( ~w7203 & w7347 ) | ( ~w7203 & w7348 ) | ( w7347 & w7348 ) ;
  assign w7350 = w7348 | w7349 ;
  assign w7351 = \pi081 ^ w7190 ;
  assign w7352 = ( ~w7197 & w7350 ) | ( ~w7197 & w7351 ) | ( w7350 & w7351 ) ;
  assign w7353 = w7351 | w7352 ;
  assign w7354 = \pi082 ^ w7184 ;
  assign w7355 = ( ~w7191 & w7353 ) | ( ~w7191 & w7354 ) | ( w7353 & w7354 ) ;
  assign w7356 = w7354 | w7355 ;
  assign w7357 = \pi083 ^ w7178 ;
  assign w7358 = ( ~w7185 & w7356 ) | ( ~w7185 & w7357 ) | ( w7356 & w7357 ) ;
  assign w7359 = w7357 | w7358 ;
  assign w7360 = \pi084 ^ w7172 ;
  assign w7361 = ( ~w7179 & w7359 ) | ( ~w7179 & w7360 ) | ( w7359 & w7360 ) ;
  assign w7362 = w7360 | w7361 ;
  assign w7363 = \pi085 ^ w7166 ;
  assign w7364 = ( ~w7173 & w7362 ) | ( ~w7173 & w7363 ) | ( w7362 & w7363 ) ;
  assign w7365 = w7363 | w7364 ;
  assign w7366 = \pi086 ^ w7160 ;
  assign w7367 = ( ~w7167 & w7365 ) | ( ~w7167 & w7366 ) | ( w7365 & w7366 ) ;
  assign w7368 = w7366 | w7367 ;
  assign w7369 = \pi087 ^ w7154 ;
  assign w7370 = ( ~w7161 & w7368 ) | ( ~w7161 & w7369 ) | ( w7368 & w7369 ) ;
  assign w7371 = w7369 | w7370 ;
  assign w7372 = \pi088 ^ w7148 ;
  assign w7373 = ( ~w7155 & w7371 ) | ( ~w7155 & w7372 ) | ( w7371 & w7372 ) ;
  assign w7374 = w7372 | w7373 ;
  assign w7375 = \pi089 ^ w7142 ;
  assign w7376 = ( ~w7149 & w7374 ) | ( ~w7149 & w7375 ) | ( w7374 & w7375 ) ;
  assign w7377 = w7375 | w7376 ;
  assign w7378 = \pi090 ^ w7136 ;
  assign w7379 = ( ~w7143 & w7377 ) | ( ~w7143 & w7378 ) | ( w7377 & w7378 ) ;
  assign w7380 = w7378 | w7379 ;
  assign w7381 = \pi091 ^ w7130 ;
  assign w7382 = ( ~w7137 & w7380 ) | ( ~w7137 & w7381 ) | ( w7380 & w7381 ) ;
  assign w7383 = w7381 | w7382 ;
  assign w7384 = \pi092 ^ w7124 ;
  assign w7385 = ( ~w7131 & w7383 ) | ( ~w7131 & w7384 ) | ( w7383 & w7384 ) ;
  assign w7386 = w7384 | w7385 ;
  assign w7387 = \pi093 ^ w7118 ;
  assign w7388 = ( ~w7125 & w7386 ) | ( ~w7125 & w7387 ) | ( w7386 & w7387 ) ;
  assign w7389 = w7387 | w7388 ;
  assign w7390 = \pi094 ^ w7112 ;
  assign w7391 = ( ~w7119 & w7389 ) | ( ~w7119 & w7390 ) | ( w7389 & w7390 ) ;
  assign w7392 = w7390 | w7391 ;
  assign w7393 = \pi095 ^ w7106 ;
  assign w7394 = ( ~w7113 & w7392 ) | ( ~w7113 & w7393 ) | ( w7392 & w7393 ) ;
  assign w7395 = w7393 | w7394 ;
  assign w7396 = \pi096 ^ w7100 ;
  assign w7397 = ( ~w7107 & w7395 ) | ( ~w7107 & w7396 ) | ( w7395 & w7396 ) ;
  assign w7398 = w7396 | w7397 ;
  assign w7399 = \pi097 ^ w7094 ;
  assign w7400 = ( ~w7101 & w7398 ) | ( ~w7101 & w7399 ) | ( w7398 & w7399 ) ;
  assign w7401 = w7399 | w7400 ;
  assign w7402 = \pi098 ^ w7088 ;
  assign w7403 = ( ~w7095 & w7401 ) | ( ~w7095 & w7402 ) | ( w7401 & w7402 ) ;
  assign w7404 = w7402 | w7403 ;
  assign w7405 = \pi099 ^ w7082 ;
  assign w7406 = ( ~w7089 & w7404 ) | ( ~w7089 & w7405 ) | ( w7404 & w7405 ) ;
  assign w7407 = w7405 | w7406 ;
  assign w7408 = \pi100 ^ w7071 ;
  assign w7409 = ( ~w7083 & w7407 ) | ( ~w7083 & w7408 ) | ( w7407 & w7408 ) ;
  assign w7410 = w7408 | w7409 ;
  assign w7411 = \pi101 ^ w7076 ;
  assign w7412 = w7077 & ~w7411 ;
  assign w7413 = ( w7410 & w7411 ) | ( w7410 & ~w7412 ) | ( w7411 & ~w7412 ) ;
  assign w7414 = ~\pi101 & w7076 ;
  assign w7415 = w7413 & ~w7414 ;
  assign w7416 = \pi102 | \pi103 ;
  assign w7417 = w168 | w7416 ;
  assign w7418 = ( w155 & w158 ) | ( w155 & ~w168 ) | ( w158 & ~w168 ) ;
  assign w7419 = w7417 | w7418 ;
  assign w7420 = w7415 | w7419 ;
  assign w7421 = w7071 & w7420 ;
  assign w7422 = ~w7083 & w7407 ;
  assign w7423 = w7408 ^ w7422 ;
  assign w7424 = ~w7420 & w7423 ;
  assign w7425 = w7421 | w7424 ;
  assign w7426 = ~\pi101 & w7425 ;
  assign w7427 = w7082 & w7420 ;
  assign w7428 = ~w7089 & w7404 ;
  assign w7429 = w7405 ^ w7428 ;
  assign w7430 = ~w7420 & w7429 ;
  assign w7431 = w7427 | w7430 ;
  assign w7432 = ~\pi100 & w7431 ;
  assign w7433 = w7088 & w7420 ;
  assign w7434 = ~w7095 & w7401 ;
  assign w7435 = w7402 ^ w7434 ;
  assign w7436 = ~w7420 & w7435 ;
  assign w7437 = w7433 | w7436 ;
  assign w7438 = ~\pi099 & w7437 ;
  assign w7439 = w7094 & w7420 ;
  assign w7440 = ~w7101 & w7398 ;
  assign w7441 = w7399 ^ w7440 ;
  assign w7442 = ~w7420 & w7441 ;
  assign w7443 = w7439 | w7442 ;
  assign w7444 = ~\pi098 & w7443 ;
  assign w7445 = w7100 & w7420 ;
  assign w7446 = ~w7107 & w7395 ;
  assign w7447 = w7396 ^ w7446 ;
  assign w7448 = ~w7420 & w7447 ;
  assign w7449 = w7445 | w7448 ;
  assign w7450 = ~\pi097 & w7449 ;
  assign w7451 = w7106 & w7420 ;
  assign w7452 = ~w7113 & w7392 ;
  assign w7453 = w7393 ^ w7452 ;
  assign w7454 = ~w7420 & w7453 ;
  assign w7455 = w7451 | w7454 ;
  assign w7456 = ~\pi096 & w7455 ;
  assign w7457 = w7112 & w7420 ;
  assign w7458 = ~w7119 & w7389 ;
  assign w7459 = w7390 ^ w7458 ;
  assign w7460 = ~w7420 & w7459 ;
  assign w7461 = w7457 | w7460 ;
  assign w7462 = ~\pi095 & w7461 ;
  assign w7463 = w7118 & w7420 ;
  assign w7464 = ~w7125 & w7386 ;
  assign w7465 = w7387 ^ w7464 ;
  assign w7466 = ~w7420 & w7465 ;
  assign w7467 = w7463 | w7466 ;
  assign w7468 = ~\pi094 & w7467 ;
  assign w7469 = w7124 & w7420 ;
  assign w7470 = ~w7131 & w7383 ;
  assign w7471 = w7384 ^ w7470 ;
  assign w7472 = ~w7420 & w7471 ;
  assign w7473 = w7469 | w7472 ;
  assign w7474 = ~\pi093 & w7473 ;
  assign w7475 = w7130 & w7420 ;
  assign w7476 = ~w7137 & w7380 ;
  assign w7477 = w7381 ^ w7476 ;
  assign w7478 = ~w7420 & w7477 ;
  assign w7479 = w7475 | w7478 ;
  assign w7480 = ~\pi092 & w7479 ;
  assign w7481 = w7136 & w7420 ;
  assign w7482 = ~w7143 & w7377 ;
  assign w7483 = w7378 ^ w7482 ;
  assign w7484 = ~w7420 & w7483 ;
  assign w7485 = w7481 | w7484 ;
  assign w7486 = ~\pi091 & w7485 ;
  assign w7487 = w7142 & w7420 ;
  assign w7488 = ~w7149 & w7374 ;
  assign w7489 = w7375 ^ w7488 ;
  assign w7490 = ~w7420 & w7489 ;
  assign w7491 = w7487 | w7490 ;
  assign w7492 = ~\pi090 & w7491 ;
  assign w7493 = w7148 & w7420 ;
  assign w7494 = ~w7155 & w7371 ;
  assign w7495 = w7372 ^ w7494 ;
  assign w7496 = ~w7420 & w7495 ;
  assign w7497 = w7493 | w7496 ;
  assign w7498 = ~\pi089 & w7497 ;
  assign w7499 = w7154 & w7420 ;
  assign w7500 = ~w7161 & w7368 ;
  assign w7501 = w7369 ^ w7500 ;
  assign w7502 = ~w7420 & w7501 ;
  assign w7503 = w7499 | w7502 ;
  assign w7504 = ~\pi088 & w7503 ;
  assign w7505 = w7160 & w7420 ;
  assign w7506 = ~w7167 & w7365 ;
  assign w7507 = w7366 ^ w7506 ;
  assign w7508 = ~w7420 & w7507 ;
  assign w7509 = w7505 | w7508 ;
  assign w7510 = ~\pi087 & w7509 ;
  assign w7511 = w7166 & w7420 ;
  assign w7512 = ~w7173 & w7362 ;
  assign w7513 = w7363 ^ w7512 ;
  assign w7514 = ~w7420 & w7513 ;
  assign w7515 = w7511 | w7514 ;
  assign w7516 = ~\pi086 & w7515 ;
  assign w7517 = w7172 & w7420 ;
  assign w7518 = ~w7179 & w7359 ;
  assign w7519 = w7360 ^ w7518 ;
  assign w7520 = ~w7420 & w7519 ;
  assign w7521 = w7517 | w7520 ;
  assign w7522 = ~\pi085 & w7521 ;
  assign w7523 = w7178 & w7420 ;
  assign w7524 = ~w7185 & w7356 ;
  assign w7525 = w7357 ^ w7524 ;
  assign w7526 = ~w7420 & w7525 ;
  assign w7527 = w7523 | w7526 ;
  assign w7528 = ~\pi084 & w7527 ;
  assign w7529 = w7184 & w7420 ;
  assign w7530 = ~w7191 & w7353 ;
  assign w7531 = w7354 ^ w7530 ;
  assign w7532 = ~w7420 & w7531 ;
  assign w7533 = w7529 | w7532 ;
  assign w7534 = ~\pi083 & w7533 ;
  assign w7535 = w7190 & w7420 ;
  assign w7536 = ~w7197 & w7350 ;
  assign w7537 = w7351 ^ w7536 ;
  assign w7538 = ~w7420 & w7537 ;
  assign w7539 = w7535 | w7538 ;
  assign w7540 = ~\pi082 & w7539 ;
  assign w7541 = w7196 & w7420 ;
  assign w7542 = ~w7203 & w7347 ;
  assign w7543 = w7348 ^ w7542 ;
  assign w7544 = ~w7420 & w7543 ;
  assign w7545 = w7541 | w7544 ;
  assign w7546 = ~\pi081 & w7545 ;
  assign w7547 = w7202 & w7420 ;
  assign w7548 = ~w7209 & w7344 ;
  assign w7549 = w7345 ^ w7548 ;
  assign w7550 = ~w7420 & w7549 ;
  assign w7551 = w7547 | w7550 ;
  assign w7552 = ~\pi080 & w7551 ;
  assign w7553 = w7208 & w7420 ;
  assign w7554 = ~w7215 & w7341 ;
  assign w7555 = w7342 ^ w7554 ;
  assign w7556 = ~w7420 & w7555 ;
  assign w7557 = w7553 | w7556 ;
  assign w7558 = ~\pi079 & w7557 ;
  assign w7559 = w7214 & w7420 ;
  assign w7560 = ~w7221 & w7338 ;
  assign w7561 = w7339 ^ w7560 ;
  assign w7562 = ~w7420 & w7561 ;
  assign w7563 = w7559 | w7562 ;
  assign w7564 = ~\pi078 & w7563 ;
  assign w7565 = w7220 & w7420 ;
  assign w7566 = ~w7227 & w7335 ;
  assign w7567 = w7336 ^ w7566 ;
  assign w7568 = ~w7420 & w7567 ;
  assign w7569 = w7565 | w7568 ;
  assign w7570 = ~\pi077 & w7569 ;
  assign w7571 = w7226 & w7420 ;
  assign w7572 = ~w7233 & w7332 ;
  assign w7573 = w7333 ^ w7572 ;
  assign w7574 = ~w7420 & w7573 ;
  assign w7575 = w7571 | w7574 ;
  assign w7576 = ~\pi076 & w7575 ;
  assign w7577 = w7232 & w7420 ;
  assign w7578 = ~w7239 & w7329 ;
  assign w7579 = w7330 ^ w7578 ;
  assign w7580 = ~w7420 & w7579 ;
  assign w7581 = w7577 | w7580 ;
  assign w7582 = ~\pi075 & w7581 ;
  assign w7583 = w7238 & w7420 ;
  assign w7584 = ~w7245 & w7326 ;
  assign w7585 = w7327 ^ w7584 ;
  assign w7586 = ~w7420 & w7585 ;
  assign w7587 = w7583 | w7586 ;
  assign w7588 = ~\pi074 & w7587 ;
  assign w7589 = w7244 & w7420 ;
  assign w7590 = ~w7251 & w7323 ;
  assign w7591 = w7324 ^ w7590 ;
  assign w7592 = ~w7420 & w7591 ;
  assign w7593 = w7589 | w7592 ;
  assign w7594 = ~\pi073 & w7593 ;
  assign w7595 = w7250 & w7420 ;
  assign w7596 = ~w7257 & w7320 ;
  assign w7597 = w7321 ^ w7596 ;
  assign w7598 = ~w7420 & w7597 ;
  assign w7599 = w7595 | w7598 ;
  assign w7600 = ~\pi072 & w7599 ;
  assign w7601 = w7256 & w7420 ;
  assign w7602 = ~w7263 & w7317 ;
  assign w7603 = w7318 ^ w7602 ;
  assign w7604 = ~w7420 & w7603 ;
  assign w7605 = w7601 | w7604 ;
  assign w7606 = ~\pi071 & w7605 ;
  assign w7607 = w7262 & w7420 ;
  assign w7608 = ~w7269 & w7314 ;
  assign w7609 = w7315 ^ w7608 ;
  assign w7610 = ~w7420 & w7609 ;
  assign w7611 = w7607 | w7610 ;
  assign w7612 = ~\pi070 & w7611 ;
  assign w7613 = w7268 & w7420 ;
  assign w7614 = ~w7277 & w7311 ;
  assign w7615 = w7312 ^ w7614 ;
  assign w7616 = ~w7420 & w7615 ;
  assign w7617 = w7613 | w7616 ;
  assign w7618 = ~\pi069 & w7617 ;
  assign w7619 = w7276 & w7420 ;
  assign w7620 = ~w7288 & w7308 ;
  assign w7621 = w7309 ^ w7620 ;
  assign w7622 = ~w7420 & w7621 ;
  assign w7623 = w7619 | w7622 ;
  assign w7624 = ~\pi068 & w7623 ;
  assign w7625 = w7287 & w7420 ;
  assign w7626 = w7305 ^ w7307 ;
  assign w7627 = ( w7415 & w7419 ) | ( w7415 & w7626 ) | ( w7419 & w7626 ) ;
  assign w7628 = w7626 & ~w7627 ;
  assign w7629 = w7625 | w7628 ;
  assign w7630 = ~\pi067 & w7629 ;
  assign w7631 = ( w7296 & w7301 ) | ( w7296 & ~w7419 ) | ( w7301 & ~w7419 ) ;
  assign w7632 = \pi065 ^ w7631 ;
  assign w7633 = ( w7302 & ~w7419 ) | ( w7302 & w7632 ) | ( ~w7419 & w7632 ) ;
  assign w7634 = ( w7302 & w7415 ) | ( w7302 & w7632 ) | ( w7415 & w7632 ) ;
  assign w7635 = w7633 & ~w7634 ;
  assign w7636 = w7306 & ~w7420 ;
  assign w7637 = ( w7306 & w7635 ) | ( w7306 & ~w7636 ) | ( w7635 & ~w7636 ) ;
  assign w7638 = ~\pi066 & w7637 ;
  assign w7639 = ( \pi064 & ~\pi102 ) | ( \pi064 & \pi103 ) | ( ~\pi102 & \pi103 ) ;
  assign w7640 = w287 | w449 ;
  assign w7641 = ( \pi103 & \pi104 ) | ( \pi103 & ~w287 ) | ( \pi104 & ~w287 ) ;
  assign w7642 = w7640 | w7641 ;
  assign w7643 = w7639 & ~w7642 ;
  assign w7644 = ~w448 & w7643 ;
  assign w7645 = ( \pi026 & w7415 ) | ( \pi026 & ~w7644 ) | ( w7415 & ~w7644 ) ;
  assign w7646 = \pi026 & w7645 ;
  assign w7647 = ( \pi102 & ~w158 ) | ( \pi102 & w7302 ) | ( ~w158 & w7302 ) ;
  assign w7648 = w155 | w168 ;
  assign w7649 = ( \pi102 & \pi103 ) | ( \pi102 & ~w168 ) | ( \pi103 & ~w168 ) ;
  assign w7650 = w7648 | w7649 ;
  assign w7651 = w7647 & ~w7650 ;
  assign w7652 = ~w7415 & w7651 ;
  assign w7653 = w7646 | w7652 ;
  assign w7654 = ~\pi025 & \pi064 ;
  assign w7655 = \pi065 ^ w7653 ;
  assign w7656 = w7654 | w7655 ;
  assign w7657 = \pi066 ^ w7637 ;
  assign w7658 = ~\pi065 & w7653 ;
  assign w7659 = w7656 | w7658 ;
  assign w7660 = ( w7657 & ~w7658 ) | ( w7657 & w7659 ) | ( ~w7658 & w7659 ) ;
  assign w7661 = \pi067 ^ w7629 ;
  assign w7662 = ( ~w7638 & w7660 ) | ( ~w7638 & w7661 ) | ( w7660 & w7661 ) ;
  assign w7663 = w7661 | w7662 ;
  assign w7664 = \pi068 ^ w7623 ;
  assign w7665 = ( ~w7630 & w7663 ) | ( ~w7630 & w7664 ) | ( w7663 & w7664 ) ;
  assign w7666 = w7664 | w7665 ;
  assign w7667 = \pi069 ^ w7617 ;
  assign w7668 = ( ~w7624 & w7666 ) | ( ~w7624 & w7667 ) | ( w7666 & w7667 ) ;
  assign w7669 = w7667 | w7668 ;
  assign w7670 = \pi070 ^ w7611 ;
  assign w7671 = ( ~w7618 & w7669 ) | ( ~w7618 & w7670 ) | ( w7669 & w7670 ) ;
  assign w7672 = w7670 | w7671 ;
  assign w7673 = \pi071 ^ w7605 ;
  assign w7674 = ( ~w7612 & w7672 ) | ( ~w7612 & w7673 ) | ( w7672 & w7673 ) ;
  assign w7675 = w7673 | w7674 ;
  assign w7676 = \pi072 ^ w7599 ;
  assign w7677 = ( ~w7606 & w7675 ) | ( ~w7606 & w7676 ) | ( w7675 & w7676 ) ;
  assign w7678 = w7676 | w7677 ;
  assign w7679 = \pi073 ^ w7593 ;
  assign w7680 = ( ~w7600 & w7678 ) | ( ~w7600 & w7679 ) | ( w7678 & w7679 ) ;
  assign w7681 = w7679 | w7680 ;
  assign w7682 = \pi074 ^ w7587 ;
  assign w7683 = ( ~w7594 & w7681 ) | ( ~w7594 & w7682 ) | ( w7681 & w7682 ) ;
  assign w7684 = w7682 | w7683 ;
  assign w7685 = \pi075 ^ w7581 ;
  assign w7686 = ( ~w7588 & w7684 ) | ( ~w7588 & w7685 ) | ( w7684 & w7685 ) ;
  assign w7687 = w7685 | w7686 ;
  assign w7688 = \pi076 ^ w7575 ;
  assign w7689 = ( ~w7582 & w7687 ) | ( ~w7582 & w7688 ) | ( w7687 & w7688 ) ;
  assign w7690 = w7688 | w7689 ;
  assign w7691 = \pi077 ^ w7569 ;
  assign w7692 = ( ~w7576 & w7690 ) | ( ~w7576 & w7691 ) | ( w7690 & w7691 ) ;
  assign w7693 = w7691 | w7692 ;
  assign w7694 = \pi078 ^ w7563 ;
  assign w7695 = ( ~w7570 & w7693 ) | ( ~w7570 & w7694 ) | ( w7693 & w7694 ) ;
  assign w7696 = w7694 | w7695 ;
  assign w7697 = \pi079 ^ w7557 ;
  assign w7698 = ( ~w7564 & w7696 ) | ( ~w7564 & w7697 ) | ( w7696 & w7697 ) ;
  assign w7699 = w7697 | w7698 ;
  assign w7700 = \pi080 ^ w7551 ;
  assign w7701 = ( ~w7558 & w7699 ) | ( ~w7558 & w7700 ) | ( w7699 & w7700 ) ;
  assign w7702 = w7700 | w7701 ;
  assign w7703 = \pi081 ^ w7545 ;
  assign w7704 = ( ~w7552 & w7702 ) | ( ~w7552 & w7703 ) | ( w7702 & w7703 ) ;
  assign w7705 = w7703 | w7704 ;
  assign w7706 = \pi082 ^ w7539 ;
  assign w7707 = ( ~w7546 & w7705 ) | ( ~w7546 & w7706 ) | ( w7705 & w7706 ) ;
  assign w7708 = w7706 | w7707 ;
  assign w7709 = \pi083 ^ w7533 ;
  assign w7710 = ( ~w7540 & w7708 ) | ( ~w7540 & w7709 ) | ( w7708 & w7709 ) ;
  assign w7711 = w7709 | w7710 ;
  assign w7712 = \pi084 ^ w7527 ;
  assign w7713 = ( ~w7534 & w7711 ) | ( ~w7534 & w7712 ) | ( w7711 & w7712 ) ;
  assign w7714 = w7712 | w7713 ;
  assign w7715 = \pi085 ^ w7521 ;
  assign w7716 = ( ~w7528 & w7714 ) | ( ~w7528 & w7715 ) | ( w7714 & w7715 ) ;
  assign w7717 = w7715 | w7716 ;
  assign w7718 = \pi086 ^ w7515 ;
  assign w7719 = ( ~w7522 & w7717 ) | ( ~w7522 & w7718 ) | ( w7717 & w7718 ) ;
  assign w7720 = w7718 | w7719 ;
  assign w7721 = \pi087 ^ w7509 ;
  assign w7722 = ( ~w7516 & w7720 ) | ( ~w7516 & w7721 ) | ( w7720 & w7721 ) ;
  assign w7723 = w7721 | w7722 ;
  assign w7724 = \pi088 ^ w7503 ;
  assign w7725 = ( ~w7510 & w7723 ) | ( ~w7510 & w7724 ) | ( w7723 & w7724 ) ;
  assign w7726 = w7724 | w7725 ;
  assign w7727 = \pi089 ^ w7497 ;
  assign w7728 = ( ~w7504 & w7726 ) | ( ~w7504 & w7727 ) | ( w7726 & w7727 ) ;
  assign w7729 = w7727 | w7728 ;
  assign w7730 = \pi090 ^ w7491 ;
  assign w7731 = ( ~w7498 & w7729 ) | ( ~w7498 & w7730 ) | ( w7729 & w7730 ) ;
  assign w7732 = w7730 | w7731 ;
  assign w7733 = \pi091 ^ w7485 ;
  assign w7734 = ( ~w7492 & w7732 ) | ( ~w7492 & w7733 ) | ( w7732 & w7733 ) ;
  assign w7735 = w7733 | w7734 ;
  assign w7736 = \pi092 ^ w7479 ;
  assign w7737 = ( ~w7486 & w7735 ) | ( ~w7486 & w7736 ) | ( w7735 & w7736 ) ;
  assign w7738 = w7736 | w7737 ;
  assign w7739 = \pi093 ^ w7473 ;
  assign w7740 = ( ~w7480 & w7738 ) | ( ~w7480 & w7739 ) | ( w7738 & w7739 ) ;
  assign w7741 = w7739 | w7740 ;
  assign w7742 = \pi094 ^ w7467 ;
  assign w7743 = ( ~w7474 & w7741 ) | ( ~w7474 & w7742 ) | ( w7741 & w7742 ) ;
  assign w7744 = w7742 | w7743 ;
  assign w7745 = \pi095 ^ w7461 ;
  assign w7746 = ( ~w7468 & w7744 ) | ( ~w7468 & w7745 ) | ( w7744 & w7745 ) ;
  assign w7747 = w7745 | w7746 ;
  assign w7748 = \pi096 ^ w7455 ;
  assign w7749 = ( ~w7462 & w7747 ) | ( ~w7462 & w7748 ) | ( w7747 & w7748 ) ;
  assign w7750 = w7748 | w7749 ;
  assign w7751 = \pi097 ^ w7449 ;
  assign w7752 = ( ~w7456 & w7750 ) | ( ~w7456 & w7751 ) | ( w7750 & w7751 ) ;
  assign w7753 = w7751 | w7752 ;
  assign w7754 = \pi098 ^ w7443 ;
  assign w7755 = ( ~w7450 & w7753 ) | ( ~w7450 & w7754 ) | ( w7753 & w7754 ) ;
  assign w7756 = w7754 | w7755 ;
  assign w7757 = \pi099 ^ w7437 ;
  assign w7758 = ( ~w7444 & w7756 ) | ( ~w7444 & w7757 ) | ( w7756 & w7757 ) ;
  assign w7759 = w7757 | w7758 ;
  assign w7760 = \pi100 ^ w7431 ;
  assign w7761 = ( ~w7438 & w7759 ) | ( ~w7438 & w7760 ) | ( w7759 & w7760 ) ;
  assign w7762 = w7760 | w7761 ;
  assign w7763 = \pi101 ^ w7425 ;
  assign w7764 = ( ~w7432 & w7762 ) | ( ~w7432 & w7763 ) | ( w7762 & w7763 ) ;
  assign w7765 = w7763 | w7764 ;
  assign w7766 = w7076 & w7420 ;
  assign w7767 = ~w7077 & w7410 ;
  assign w7768 = w7411 ^ w7767 ;
  assign w7769 = ~w7420 & w7768 ;
  assign w7770 = w7766 | w7769 ;
  assign w7771 = ~\pi102 & w7770 ;
  assign w7772 = ( \pi102 & ~w7766 ) | ( \pi102 & w7769 ) | ( ~w7766 & w7769 ) ;
  assign w7773 = ~w7769 & w7772 ;
  assign w7774 = \pi103 | \pi104 ;
  assign w7775 = w449 | w7774 ;
  assign w7776 = ( w287 & w448 ) | ( w287 & ~w449 ) | ( w448 & ~w449 ) ;
  assign w7777 = w7775 | w7776 ;
  assign w7778 = w7771 | w7773 ;
  assign w7779 = ( ~w7426 & w7765 ) | ( ~w7426 & w7778 ) | ( w7765 & w7778 ) ;
  assign w7780 = ( w7777 & ~w7778 ) | ( w7777 & w7779 ) | ( ~w7778 & w7779 ) ;
  assign w7781 = w7778 | w7780 ;
  assign w7782 = ~w7419 & w7770 ;
  assign w7783 = w7781 & ~w7782 ;
  assign w7784 = ~w7432 & w7762 ;
  assign w7785 = w7763 ^ w7784 ;
  assign w7786 = ~w7783 & w7785 ;
  assign w7787 = ( w7425 & w7781 ) | ( w7425 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7788 = ~w7782 & w7787 ;
  assign w7789 = w7786 | w7788 ;
  assign w7790 = ( ~w7426 & w7765 ) | ( ~w7426 & w7783 ) | ( w7765 & w7783 ) ;
  assign w7791 = w7778 ^ w7790 ;
  assign w7792 = ~w7783 & w7791 ;
  assign w7793 = ( w7419 & ~w7770 ) | ( w7419 & w7781 ) | ( ~w7770 & w7781 ) ;
  assign w7794 = w7770 & w7793 ;
  assign w7795 = w7792 | w7794 ;
  assign w7796 = ~\pi102 & w7789 ;
  assign w7797 = ~w7438 & w7759 ;
  assign w7798 = w7760 ^ w7797 ;
  assign w7799 = ~w7783 & w7798 ;
  assign w7800 = ( w7431 & w7781 ) | ( w7431 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7801 = ~w7782 & w7800 ;
  assign w7802 = w7799 | w7801 ;
  assign w7803 = ~\pi101 & w7802 ;
  assign w7804 = ~w7444 & w7756 ;
  assign w7805 = w7757 ^ w7804 ;
  assign w7806 = ~w7783 & w7805 ;
  assign w7807 = ( w7437 & w7781 ) | ( w7437 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7808 = ~w7782 & w7807 ;
  assign w7809 = w7806 | w7808 ;
  assign w7810 = ~\pi100 & w7809 ;
  assign w7811 = ~w7450 & w7753 ;
  assign w7812 = w7754 ^ w7811 ;
  assign w7813 = ~w7783 & w7812 ;
  assign w7814 = ( w7443 & w7781 ) | ( w7443 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7815 = ~w7782 & w7814 ;
  assign w7816 = w7813 | w7815 ;
  assign w7817 = ~\pi099 & w7816 ;
  assign w7818 = ~w7456 & w7750 ;
  assign w7819 = w7751 ^ w7818 ;
  assign w7820 = ~w7783 & w7819 ;
  assign w7821 = ( w7449 & w7781 ) | ( w7449 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7822 = ~w7782 & w7821 ;
  assign w7823 = w7820 | w7822 ;
  assign w7824 = ~\pi098 & w7823 ;
  assign w7825 = ~w7462 & w7747 ;
  assign w7826 = w7748 ^ w7825 ;
  assign w7827 = ~w7783 & w7826 ;
  assign w7828 = ( w7455 & w7781 ) | ( w7455 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7829 = ~w7782 & w7828 ;
  assign w7830 = w7827 | w7829 ;
  assign w7831 = ~\pi097 & w7830 ;
  assign w7832 = ~w7468 & w7744 ;
  assign w7833 = w7745 ^ w7832 ;
  assign w7834 = ~w7783 & w7833 ;
  assign w7835 = ( w7461 & w7781 ) | ( w7461 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7836 = ~w7782 & w7835 ;
  assign w7837 = w7834 | w7836 ;
  assign w7838 = ~\pi096 & w7837 ;
  assign w7839 = ~w7474 & w7741 ;
  assign w7840 = w7742 ^ w7839 ;
  assign w7841 = ~w7783 & w7840 ;
  assign w7842 = ( w7467 & w7781 ) | ( w7467 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7843 = ~w7782 & w7842 ;
  assign w7844 = w7841 | w7843 ;
  assign w7845 = ~\pi095 & w7844 ;
  assign w7846 = ~w7480 & w7738 ;
  assign w7847 = w7739 ^ w7846 ;
  assign w7848 = ~w7783 & w7847 ;
  assign w7849 = ( w7473 & w7781 ) | ( w7473 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7850 = ~w7782 & w7849 ;
  assign w7851 = w7848 | w7850 ;
  assign w7852 = ~\pi094 & w7851 ;
  assign w7853 = ~w7486 & w7735 ;
  assign w7854 = w7736 ^ w7853 ;
  assign w7855 = ~w7783 & w7854 ;
  assign w7856 = ( w7479 & w7781 ) | ( w7479 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7857 = ~w7782 & w7856 ;
  assign w7858 = w7855 | w7857 ;
  assign w7859 = ~\pi093 & w7858 ;
  assign w7860 = ~w7492 & w7732 ;
  assign w7861 = w7733 ^ w7860 ;
  assign w7862 = ~w7783 & w7861 ;
  assign w7863 = ( w7485 & w7781 ) | ( w7485 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7864 = ~w7782 & w7863 ;
  assign w7865 = w7862 | w7864 ;
  assign w7866 = ~\pi092 & w7865 ;
  assign w7867 = ~w7498 & w7729 ;
  assign w7868 = w7730 ^ w7867 ;
  assign w7869 = ~w7783 & w7868 ;
  assign w7870 = ( w7491 & w7781 ) | ( w7491 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7871 = ~w7782 & w7870 ;
  assign w7872 = w7869 | w7871 ;
  assign w7873 = ~\pi091 & w7872 ;
  assign w7874 = ~w7504 & w7726 ;
  assign w7875 = w7727 ^ w7874 ;
  assign w7876 = ~w7783 & w7875 ;
  assign w7877 = ( w7497 & w7781 ) | ( w7497 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7878 = ~w7782 & w7877 ;
  assign w7879 = w7876 | w7878 ;
  assign w7880 = ~\pi090 & w7879 ;
  assign w7881 = ~w7510 & w7723 ;
  assign w7882 = w7724 ^ w7881 ;
  assign w7883 = ~w7783 & w7882 ;
  assign w7884 = ( w7503 & w7781 ) | ( w7503 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7885 = ~w7782 & w7884 ;
  assign w7886 = w7883 | w7885 ;
  assign w7887 = ~\pi089 & w7886 ;
  assign w7888 = ~w7516 & w7720 ;
  assign w7889 = w7721 ^ w7888 ;
  assign w7890 = ~w7783 & w7889 ;
  assign w7891 = ( w7509 & w7781 ) | ( w7509 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7892 = ~w7782 & w7891 ;
  assign w7893 = w7890 | w7892 ;
  assign w7894 = ~\pi088 & w7893 ;
  assign w7895 = ~w7522 & w7717 ;
  assign w7896 = w7718 ^ w7895 ;
  assign w7897 = ~w7783 & w7896 ;
  assign w7898 = ( w7515 & w7781 ) | ( w7515 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7899 = ~w7782 & w7898 ;
  assign w7900 = w7897 | w7899 ;
  assign w7901 = ~\pi087 & w7900 ;
  assign w7902 = ~w7528 & w7714 ;
  assign w7903 = w7715 ^ w7902 ;
  assign w7904 = ~w7783 & w7903 ;
  assign w7905 = ( w7521 & w7781 ) | ( w7521 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7906 = ~w7782 & w7905 ;
  assign w7907 = w7904 | w7906 ;
  assign w7908 = ~\pi086 & w7907 ;
  assign w7909 = ~w7534 & w7711 ;
  assign w7910 = w7712 ^ w7909 ;
  assign w7911 = ~w7783 & w7910 ;
  assign w7912 = ( w7527 & w7781 ) | ( w7527 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7913 = ~w7782 & w7912 ;
  assign w7914 = w7911 | w7913 ;
  assign w7915 = ~\pi085 & w7914 ;
  assign w7916 = ~w7540 & w7708 ;
  assign w7917 = w7709 ^ w7916 ;
  assign w7918 = ~w7783 & w7917 ;
  assign w7919 = ( w7533 & w7781 ) | ( w7533 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7920 = ~w7782 & w7919 ;
  assign w7921 = w7918 | w7920 ;
  assign w7922 = ~\pi084 & w7921 ;
  assign w7923 = ~w7546 & w7705 ;
  assign w7924 = w7706 ^ w7923 ;
  assign w7925 = ~w7783 & w7924 ;
  assign w7926 = ( w7539 & w7781 ) | ( w7539 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7927 = ~w7782 & w7926 ;
  assign w7928 = w7925 | w7927 ;
  assign w7929 = ~\pi083 & w7928 ;
  assign w7930 = ~w7552 & w7702 ;
  assign w7931 = w7703 ^ w7930 ;
  assign w7932 = ~w7783 & w7931 ;
  assign w7933 = ( w7545 & w7781 ) | ( w7545 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7934 = ~w7782 & w7933 ;
  assign w7935 = w7932 | w7934 ;
  assign w7936 = ~\pi082 & w7935 ;
  assign w7937 = ~w7558 & w7699 ;
  assign w7938 = w7700 ^ w7937 ;
  assign w7939 = ~w7783 & w7938 ;
  assign w7940 = ( w7551 & w7781 ) | ( w7551 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7941 = ~w7782 & w7940 ;
  assign w7942 = w7939 | w7941 ;
  assign w7943 = ~\pi081 & w7942 ;
  assign w7944 = ~w7564 & w7696 ;
  assign w7945 = w7697 ^ w7944 ;
  assign w7946 = ~w7783 & w7945 ;
  assign w7947 = ( w7557 & w7781 ) | ( w7557 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7948 = ~w7782 & w7947 ;
  assign w7949 = w7946 | w7948 ;
  assign w7950 = ~\pi080 & w7949 ;
  assign w7951 = ~w7570 & w7693 ;
  assign w7952 = w7694 ^ w7951 ;
  assign w7953 = ~w7783 & w7952 ;
  assign w7954 = ( w7563 & w7781 ) | ( w7563 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7955 = ~w7782 & w7954 ;
  assign w7956 = w7953 | w7955 ;
  assign w7957 = ~\pi079 & w7956 ;
  assign w7958 = ~w7576 & w7690 ;
  assign w7959 = w7691 ^ w7958 ;
  assign w7960 = ~w7783 & w7959 ;
  assign w7961 = ( w7569 & w7781 ) | ( w7569 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7962 = ~w7782 & w7961 ;
  assign w7963 = w7960 | w7962 ;
  assign w7964 = ~\pi078 & w7963 ;
  assign w7965 = ~w7582 & w7687 ;
  assign w7966 = w7688 ^ w7965 ;
  assign w7967 = ~w7783 & w7966 ;
  assign w7968 = ( w7575 & w7781 ) | ( w7575 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7969 = ~w7782 & w7968 ;
  assign w7970 = w7967 | w7969 ;
  assign w7971 = ~\pi077 & w7970 ;
  assign w7972 = ~w7588 & w7684 ;
  assign w7973 = w7685 ^ w7972 ;
  assign w7974 = ~w7783 & w7973 ;
  assign w7975 = ( w7581 & w7781 ) | ( w7581 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7976 = ~w7782 & w7975 ;
  assign w7977 = w7974 | w7976 ;
  assign w7978 = ~\pi076 & w7977 ;
  assign w7979 = ~w7594 & w7681 ;
  assign w7980 = w7682 ^ w7979 ;
  assign w7981 = ~w7783 & w7980 ;
  assign w7982 = ( w7587 & w7781 ) | ( w7587 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7983 = ~w7782 & w7982 ;
  assign w7984 = w7981 | w7983 ;
  assign w7985 = ~\pi075 & w7984 ;
  assign w7986 = ~w7600 & w7678 ;
  assign w7987 = w7679 ^ w7986 ;
  assign w7988 = ~w7783 & w7987 ;
  assign w7989 = ( w7593 & w7781 ) | ( w7593 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7990 = ~w7782 & w7989 ;
  assign w7991 = w7988 | w7990 ;
  assign w7992 = ~\pi074 & w7991 ;
  assign w7993 = ~w7606 & w7675 ;
  assign w7994 = w7676 ^ w7993 ;
  assign w7995 = ~w7783 & w7994 ;
  assign w7996 = ( w7599 & w7781 ) | ( w7599 & w7782 ) | ( w7781 & w7782 ) ;
  assign w7997 = ~w7782 & w7996 ;
  assign w7998 = w7995 | w7997 ;
  assign w7999 = ~\pi073 & w7998 ;
  assign w8000 = ~w7612 & w7672 ;
  assign w8001 = w7673 ^ w8000 ;
  assign w8002 = ~w7783 & w8001 ;
  assign w8003 = ( w7605 & w7781 ) | ( w7605 & w7782 ) | ( w7781 & w7782 ) ;
  assign w8004 = ~w7782 & w8003 ;
  assign w8005 = w8002 | w8004 ;
  assign w8006 = ~\pi072 & w8005 ;
  assign w8007 = ~w7618 & w7669 ;
  assign w8008 = w7670 ^ w8007 ;
  assign w8009 = ~w7783 & w8008 ;
  assign w8010 = ( w7611 & w7781 ) | ( w7611 & w7782 ) | ( w7781 & w7782 ) ;
  assign w8011 = ~w7782 & w8010 ;
  assign w8012 = w8009 | w8011 ;
  assign w8013 = ~\pi071 & w8012 ;
  assign w8014 = ~w7624 & w7666 ;
  assign w8015 = w7667 ^ w8014 ;
  assign w8016 = ~w7783 & w8015 ;
  assign w8017 = ( w7617 & w7781 ) | ( w7617 & w7782 ) | ( w7781 & w7782 ) ;
  assign w8018 = ~w7782 & w8017 ;
  assign w8019 = w8016 | w8018 ;
  assign w8020 = ~\pi070 & w8019 ;
  assign w8021 = ~w7630 & w7663 ;
  assign w8022 = w7664 ^ w8021 ;
  assign w8023 = ~w7783 & w8022 ;
  assign w8024 = ( w7623 & w7781 ) | ( w7623 & w7782 ) | ( w7781 & w7782 ) ;
  assign w8025 = ~w7782 & w8024 ;
  assign w8026 = w8023 | w8025 ;
  assign w8027 = ~\pi069 & w8026 ;
  assign w8028 = ~w7638 & w7660 ;
  assign w8029 = w7661 ^ w8028 ;
  assign w8030 = ~w7783 & w8029 ;
  assign w8031 = ( w7629 & w7781 ) | ( w7629 & w7782 ) | ( w7781 & w7782 ) ;
  assign w8032 = ~w7782 & w8031 ;
  assign w8033 = w8030 | w8032 ;
  assign w8034 = ~\pi068 & w8033 ;
  assign w8035 = ( \pi065 & w7653 ) | ( \pi065 & ~w7783 ) | ( w7653 & ~w7783 ) ;
  assign w8036 = ( \pi065 & w7656 ) | ( \pi065 & ~w8035 ) | ( w7656 & ~w8035 ) ;
  assign w8037 = w7657 ^ w8036 ;
  assign w8038 = ~w7783 & w8037 ;
  assign w8039 = ( w7637 & w7781 ) | ( w7637 & w7782 ) | ( w7781 & w7782 ) ;
  assign w8040 = ~w7782 & w8039 ;
  assign w8041 = w8038 | w8040 ;
  assign w8042 = ~\pi067 & w8041 ;
  assign w8043 = w7653 ^ w7654 ;
  assign w8044 = \pi065 ^ w8043 ;
  assign w8045 = w7783 ^ w8044 ;
  assign w8046 = ( w7653 & w8044 ) | ( w7653 & w8045 ) | ( w8044 & w8045 ) ;
  assign w8047 = ~\pi066 & w8046 ;
  assign w8048 = w7653 ^ w7783 ;
  assign w8049 = ( w7653 & w8044 ) | ( w7653 & ~w8048 ) | ( w8044 & ~w8048 ) ;
  assign w8050 = \pi066 ^ w8049 ;
  assign w8051 = \pi064 & ~w7783 ;
  assign w8052 = \pi025 ^ w8051 ;
  assign w8053 = ( ~\pi024 & \pi064 ) | ( ~\pi024 & w8050 ) | ( \pi064 & w8050 ) ;
  assign w8054 = ( \pi065 & ~w8052 ) | ( \pi065 & w8053 ) | ( ~w8052 & w8053 ) ;
  assign w8055 = w8050 | w8054 ;
  assign w8056 = \pi067 ^ w8041 ;
  assign w8057 = ( ~w8047 & w8055 ) | ( ~w8047 & w8056 ) | ( w8055 & w8056 ) ;
  assign w8058 = w8056 | w8057 ;
  assign w8059 = \pi068 ^ w8033 ;
  assign w8060 = ( ~w8042 & w8058 ) | ( ~w8042 & w8059 ) | ( w8058 & w8059 ) ;
  assign w8061 = w8059 | w8060 ;
  assign w8062 = \pi069 ^ w8026 ;
  assign w8063 = ( ~w8034 & w8061 ) | ( ~w8034 & w8062 ) | ( w8061 & w8062 ) ;
  assign w8064 = w8062 | w8063 ;
  assign w8065 = \pi070 ^ w8019 ;
  assign w8066 = ( ~w8027 & w8064 ) | ( ~w8027 & w8065 ) | ( w8064 & w8065 ) ;
  assign w8067 = w8065 | w8066 ;
  assign w8068 = \pi071 ^ w8012 ;
  assign w8069 = ( ~w8020 & w8067 ) | ( ~w8020 & w8068 ) | ( w8067 & w8068 ) ;
  assign w8070 = w8068 | w8069 ;
  assign w8071 = \pi072 ^ w8005 ;
  assign w8072 = ( ~w8013 & w8070 ) | ( ~w8013 & w8071 ) | ( w8070 & w8071 ) ;
  assign w8073 = w8071 | w8072 ;
  assign w8074 = \pi073 ^ w7998 ;
  assign w8075 = ( ~w8006 & w8073 ) | ( ~w8006 & w8074 ) | ( w8073 & w8074 ) ;
  assign w8076 = w8074 | w8075 ;
  assign w8077 = \pi074 ^ w7991 ;
  assign w8078 = ( ~w7999 & w8076 ) | ( ~w7999 & w8077 ) | ( w8076 & w8077 ) ;
  assign w8079 = w8077 | w8078 ;
  assign w8080 = \pi075 ^ w7984 ;
  assign w8081 = ( ~w7992 & w8079 ) | ( ~w7992 & w8080 ) | ( w8079 & w8080 ) ;
  assign w8082 = w8080 | w8081 ;
  assign w8083 = \pi076 ^ w7977 ;
  assign w8084 = ( ~w7985 & w8082 ) | ( ~w7985 & w8083 ) | ( w8082 & w8083 ) ;
  assign w8085 = w8083 | w8084 ;
  assign w8086 = \pi077 ^ w7970 ;
  assign w8087 = ( ~w7978 & w8085 ) | ( ~w7978 & w8086 ) | ( w8085 & w8086 ) ;
  assign w8088 = w8086 | w8087 ;
  assign w8089 = \pi078 ^ w7963 ;
  assign w8090 = ( ~w7971 & w8088 ) | ( ~w7971 & w8089 ) | ( w8088 & w8089 ) ;
  assign w8091 = w8089 | w8090 ;
  assign w8092 = \pi079 ^ w7956 ;
  assign w8093 = ( ~w7964 & w8091 ) | ( ~w7964 & w8092 ) | ( w8091 & w8092 ) ;
  assign w8094 = w8092 | w8093 ;
  assign w8095 = \pi080 ^ w7949 ;
  assign w8096 = ( ~w7957 & w8094 ) | ( ~w7957 & w8095 ) | ( w8094 & w8095 ) ;
  assign w8097 = w8095 | w8096 ;
  assign w8098 = \pi081 ^ w7942 ;
  assign w8099 = ( ~w7950 & w8097 ) | ( ~w7950 & w8098 ) | ( w8097 & w8098 ) ;
  assign w8100 = w8098 | w8099 ;
  assign w8101 = \pi082 ^ w7935 ;
  assign w8102 = ( ~w7943 & w8100 ) | ( ~w7943 & w8101 ) | ( w8100 & w8101 ) ;
  assign w8103 = w8101 | w8102 ;
  assign w8104 = \pi083 ^ w7928 ;
  assign w8105 = ( ~w7936 & w8103 ) | ( ~w7936 & w8104 ) | ( w8103 & w8104 ) ;
  assign w8106 = w8104 | w8105 ;
  assign w8107 = \pi084 ^ w7921 ;
  assign w8108 = ( ~w7929 & w8106 ) | ( ~w7929 & w8107 ) | ( w8106 & w8107 ) ;
  assign w8109 = w8107 | w8108 ;
  assign w8110 = \pi085 ^ w7914 ;
  assign w8111 = ( ~w7922 & w8109 ) | ( ~w7922 & w8110 ) | ( w8109 & w8110 ) ;
  assign w8112 = w8110 | w8111 ;
  assign w8113 = \pi086 ^ w7907 ;
  assign w8114 = ( ~w7915 & w8112 ) | ( ~w7915 & w8113 ) | ( w8112 & w8113 ) ;
  assign w8115 = w8113 | w8114 ;
  assign w8116 = \pi087 ^ w7900 ;
  assign w8117 = ( ~w7908 & w8115 ) | ( ~w7908 & w8116 ) | ( w8115 & w8116 ) ;
  assign w8118 = w8116 | w8117 ;
  assign w8119 = \pi088 ^ w7893 ;
  assign w8120 = ( ~w7901 & w8118 ) | ( ~w7901 & w8119 ) | ( w8118 & w8119 ) ;
  assign w8121 = w8119 | w8120 ;
  assign w8122 = \pi089 ^ w7886 ;
  assign w8123 = ( ~w7894 & w8121 ) | ( ~w7894 & w8122 ) | ( w8121 & w8122 ) ;
  assign w8124 = w8122 | w8123 ;
  assign w8125 = \pi090 ^ w7879 ;
  assign w8126 = ( ~w7887 & w8124 ) | ( ~w7887 & w8125 ) | ( w8124 & w8125 ) ;
  assign w8127 = w8125 | w8126 ;
  assign w8128 = \pi091 ^ w7872 ;
  assign w8129 = ( ~w7880 & w8127 ) | ( ~w7880 & w8128 ) | ( w8127 & w8128 ) ;
  assign w8130 = w8128 | w8129 ;
  assign w8131 = \pi092 ^ w7865 ;
  assign w8132 = ( ~w7873 & w8130 ) | ( ~w7873 & w8131 ) | ( w8130 & w8131 ) ;
  assign w8133 = w8131 | w8132 ;
  assign w8134 = \pi093 ^ w7858 ;
  assign w8135 = ( ~w7866 & w8133 ) | ( ~w7866 & w8134 ) | ( w8133 & w8134 ) ;
  assign w8136 = w8134 | w8135 ;
  assign w8137 = \pi094 ^ w7851 ;
  assign w8138 = ( ~w7859 & w8136 ) | ( ~w7859 & w8137 ) | ( w8136 & w8137 ) ;
  assign w8139 = w8137 | w8138 ;
  assign w8140 = \pi095 ^ w7844 ;
  assign w8141 = ( ~w7852 & w8139 ) | ( ~w7852 & w8140 ) | ( w8139 & w8140 ) ;
  assign w8142 = w8140 | w8141 ;
  assign w8143 = \pi096 ^ w7837 ;
  assign w8144 = ( ~w7845 & w8142 ) | ( ~w7845 & w8143 ) | ( w8142 & w8143 ) ;
  assign w8145 = w8143 | w8144 ;
  assign w8146 = \pi097 ^ w7830 ;
  assign w8147 = ( ~w7838 & w8145 ) | ( ~w7838 & w8146 ) | ( w8145 & w8146 ) ;
  assign w8148 = w8146 | w8147 ;
  assign w8149 = \pi098 ^ w7823 ;
  assign w8150 = ( ~w7831 & w8148 ) | ( ~w7831 & w8149 ) | ( w8148 & w8149 ) ;
  assign w8151 = w8149 | w8150 ;
  assign w8152 = \pi099 ^ w7816 ;
  assign w8153 = ( ~w7824 & w8151 ) | ( ~w7824 & w8152 ) | ( w8151 & w8152 ) ;
  assign w8154 = w8152 | w8153 ;
  assign w8155 = \pi100 ^ w7809 ;
  assign w8156 = ( ~w7817 & w8154 ) | ( ~w7817 & w8155 ) | ( w8154 & w8155 ) ;
  assign w8157 = w8155 | w8156 ;
  assign w8158 = \pi101 ^ w7802 ;
  assign w8159 = ( ~w7810 & w8157 ) | ( ~w7810 & w8158 ) | ( w8157 & w8158 ) ;
  assign w8160 = w8158 | w8159 ;
  assign w8161 = \pi102 ^ w7789 ;
  assign w8162 = ( ~w7803 & w8160 ) | ( ~w7803 & w8161 ) | ( w8160 & w8161 ) ;
  assign w8163 = w8161 | w8162 ;
  assign w8164 = \pi103 ^ w7795 ;
  assign w8165 = w7796 & ~w8164 ;
  assign w8166 = ( w8163 & w8164 ) | ( w8163 & ~w8165 ) | ( w8164 & ~w8165 ) ;
  assign w8167 = ~\pi103 & w7795 ;
  assign w8168 = w8166 & ~w8167 ;
  assign w8169 = w201 | w202 ;
  assign w8170 = w8168 | w8169 ;
  assign w8171 = w7789 & w8170 ;
  assign w8172 = ~w7803 & w8160 ;
  assign w8173 = w8161 ^ w8172 ;
  assign w8174 = ~w8170 & w8173 ;
  assign w8175 = w8171 | w8174 ;
  assign w8176 = w7795 & w8170 ;
  assign w8177 = ~w7796 & w8163 ;
  assign w8178 = w8164 ^ w8177 ;
  assign w8179 = ~w8170 & w8178 ;
  assign w8180 = w8176 | w8179 ;
  assign w8181 = ~\pi103 & w8175 ;
  assign w8182 = w7802 & w8170 ;
  assign w8183 = ~w7810 & w8157 ;
  assign w8184 = w8158 ^ w8183 ;
  assign w8185 = ~w8170 & w8184 ;
  assign w8186 = w8182 | w8185 ;
  assign w8187 = ~\pi102 & w8186 ;
  assign w8188 = w7809 & w8170 ;
  assign w8189 = ~w7817 & w8154 ;
  assign w8190 = w8155 ^ w8189 ;
  assign w8191 = ~w8170 & w8190 ;
  assign w8192 = w8188 | w8191 ;
  assign w8193 = ~\pi101 & w8192 ;
  assign w8194 = w7816 & w8170 ;
  assign w8195 = ~w7824 & w8151 ;
  assign w8196 = w8152 ^ w8195 ;
  assign w8197 = ~w8170 & w8196 ;
  assign w8198 = w8194 | w8197 ;
  assign w8199 = ~\pi100 & w8198 ;
  assign w8200 = w7823 & w8170 ;
  assign w8201 = ~w7831 & w8148 ;
  assign w8202 = w8149 ^ w8201 ;
  assign w8203 = ~w8170 & w8202 ;
  assign w8204 = w8200 | w8203 ;
  assign w8205 = ~\pi099 & w8204 ;
  assign w8206 = w7830 & w8170 ;
  assign w8207 = ~w7838 & w8145 ;
  assign w8208 = w8146 ^ w8207 ;
  assign w8209 = ~w8170 & w8208 ;
  assign w8210 = w8206 | w8209 ;
  assign w8211 = ~\pi098 & w8210 ;
  assign w8212 = w7837 & w8170 ;
  assign w8213 = ~w7845 & w8142 ;
  assign w8214 = w8143 ^ w8213 ;
  assign w8215 = ~w8170 & w8214 ;
  assign w8216 = w8212 | w8215 ;
  assign w8217 = ~\pi097 & w8216 ;
  assign w8218 = w7844 & w8170 ;
  assign w8219 = ~w7852 & w8139 ;
  assign w8220 = w8140 ^ w8219 ;
  assign w8221 = ~w8170 & w8220 ;
  assign w8222 = w8218 | w8221 ;
  assign w8223 = ~\pi096 & w8222 ;
  assign w8224 = w7851 & w8170 ;
  assign w8225 = ~w7859 & w8136 ;
  assign w8226 = w8137 ^ w8225 ;
  assign w8227 = ~w8170 & w8226 ;
  assign w8228 = w8224 | w8227 ;
  assign w8229 = ~\pi095 & w8228 ;
  assign w8230 = w7858 & w8170 ;
  assign w8231 = ~w7866 & w8133 ;
  assign w8232 = w8134 ^ w8231 ;
  assign w8233 = ~w8170 & w8232 ;
  assign w8234 = w8230 | w8233 ;
  assign w8235 = ~\pi094 & w8234 ;
  assign w8236 = w7865 & w8170 ;
  assign w8237 = ~w7873 & w8130 ;
  assign w8238 = w8131 ^ w8237 ;
  assign w8239 = ~w8170 & w8238 ;
  assign w8240 = w8236 | w8239 ;
  assign w8241 = ~\pi093 & w8240 ;
  assign w8242 = w7872 & w8170 ;
  assign w8243 = ~w7880 & w8127 ;
  assign w8244 = w8128 ^ w8243 ;
  assign w8245 = ~w8170 & w8244 ;
  assign w8246 = w8242 | w8245 ;
  assign w8247 = ~\pi092 & w8246 ;
  assign w8248 = w7879 & w8170 ;
  assign w8249 = ~w7887 & w8124 ;
  assign w8250 = w8125 ^ w8249 ;
  assign w8251 = ~w8170 & w8250 ;
  assign w8252 = w8248 | w8251 ;
  assign w8253 = ~\pi091 & w8252 ;
  assign w8254 = w7886 & w8170 ;
  assign w8255 = ~w7894 & w8121 ;
  assign w8256 = w8122 ^ w8255 ;
  assign w8257 = ~w8170 & w8256 ;
  assign w8258 = w8254 | w8257 ;
  assign w8259 = ~\pi090 & w8258 ;
  assign w8260 = w7893 & w8170 ;
  assign w8261 = ~w7901 & w8118 ;
  assign w8262 = w8119 ^ w8261 ;
  assign w8263 = ~w8170 & w8262 ;
  assign w8264 = w8260 | w8263 ;
  assign w8265 = ~\pi089 & w8264 ;
  assign w8266 = w7900 & w8170 ;
  assign w8267 = ~w7908 & w8115 ;
  assign w8268 = w8116 ^ w8267 ;
  assign w8269 = ~w8170 & w8268 ;
  assign w8270 = w8266 | w8269 ;
  assign w8271 = ~\pi088 & w8270 ;
  assign w8272 = w7907 & w8170 ;
  assign w8273 = ~w7915 & w8112 ;
  assign w8274 = w8113 ^ w8273 ;
  assign w8275 = ~w8170 & w8274 ;
  assign w8276 = w8272 | w8275 ;
  assign w8277 = ~\pi087 & w8276 ;
  assign w8278 = w7914 & w8170 ;
  assign w8279 = ~w7922 & w8109 ;
  assign w8280 = w8110 ^ w8279 ;
  assign w8281 = ~w8170 & w8280 ;
  assign w8282 = w8278 | w8281 ;
  assign w8283 = ~\pi086 & w8282 ;
  assign w8284 = w7921 & w8170 ;
  assign w8285 = ~w7929 & w8106 ;
  assign w8286 = w8107 ^ w8285 ;
  assign w8287 = ~w8170 & w8286 ;
  assign w8288 = w8284 | w8287 ;
  assign w8289 = ~\pi085 & w8288 ;
  assign w8290 = w7928 & w8170 ;
  assign w8291 = ~w7936 & w8103 ;
  assign w8292 = w8104 ^ w8291 ;
  assign w8293 = ~w8170 & w8292 ;
  assign w8294 = w8290 | w8293 ;
  assign w8295 = ~\pi084 & w8294 ;
  assign w8296 = w7935 & w8170 ;
  assign w8297 = ~w7943 & w8100 ;
  assign w8298 = w8101 ^ w8297 ;
  assign w8299 = ~w8170 & w8298 ;
  assign w8300 = w8296 | w8299 ;
  assign w8301 = ~\pi083 & w8300 ;
  assign w8302 = w7942 & w8170 ;
  assign w8303 = ~w7950 & w8097 ;
  assign w8304 = w8098 ^ w8303 ;
  assign w8305 = ~w8170 & w8304 ;
  assign w8306 = w8302 | w8305 ;
  assign w8307 = ~\pi082 & w8306 ;
  assign w8308 = w7949 & w8170 ;
  assign w8309 = ~w7957 & w8094 ;
  assign w8310 = w8095 ^ w8309 ;
  assign w8311 = ~w8170 & w8310 ;
  assign w8312 = w8308 | w8311 ;
  assign w8313 = ~\pi081 & w8312 ;
  assign w8314 = w7956 & w8170 ;
  assign w8315 = ~w7964 & w8091 ;
  assign w8316 = w8092 ^ w8315 ;
  assign w8317 = ~w8170 & w8316 ;
  assign w8318 = w8314 | w8317 ;
  assign w8319 = ~\pi080 & w8318 ;
  assign w8320 = w7963 & w8170 ;
  assign w8321 = ~w7971 & w8088 ;
  assign w8322 = w8089 ^ w8321 ;
  assign w8323 = ~w8170 & w8322 ;
  assign w8324 = w8320 | w8323 ;
  assign w8325 = ~\pi079 & w8324 ;
  assign w8326 = w7970 & w8170 ;
  assign w8327 = ~w7978 & w8085 ;
  assign w8328 = w8086 ^ w8327 ;
  assign w8329 = ~w8170 & w8328 ;
  assign w8330 = w8326 | w8329 ;
  assign w8331 = ~\pi078 & w8330 ;
  assign w8332 = w7977 & w8170 ;
  assign w8333 = ~w7985 & w8082 ;
  assign w8334 = w8083 ^ w8333 ;
  assign w8335 = ~w8170 & w8334 ;
  assign w8336 = w8332 | w8335 ;
  assign w8337 = ~\pi077 & w8336 ;
  assign w8338 = w7984 & w8170 ;
  assign w8339 = ~w7992 & w8079 ;
  assign w8340 = w8080 ^ w8339 ;
  assign w8341 = ~w8170 & w8340 ;
  assign w8342 = w8338 | w8341 ;
  assign w8343 = ~\pi076 & w8342 ;
  assign w8344 = w7991 & w8170 ;
  assign w8345 = ~w7999 & w8076 ;
  assign w8346 = w8077 ^ w8345 ;
  assign w8347 = ~w8170 & w8346 ;
  assign w8348 = w8344 | w8347 ;
  assign w8349 = ~\pi075 & w8348 ;
  assign w8350 = w7998 & w8170 ;
  assign w8351 = ~w8006 & w8073 ;
  assign w8352 = w8074 ^ w8351 ;
  assign w8353 = ~w8170 & w8352 ;
  assign w8354 = w8350 | w8353 ;
  assign w8355 = ~\pi074 & w8354 ;
  assign w8356 = w8005 & w8170 ;
  assign w8357 = ~w8013 & w8070 ;
  assign w8358 = w8071 ^ w8357 ;
  assign w8359 = ~w8170 & w8358 ;
  assign w8360 = w8356 | w8359 ;
  assign w8361 = ~\pi073 & w8360 ;
  assign w8362 = w8012 & w8170 ;
  assign w8363 = ~w8020 & w8067 ;
  assign w8364 = w8068 ^ w8363 ;
  assign w8365 = ~w8170 & w8364 ;
  assign w8366 = w8362 | w8365 ;
  assign w8367 = ~\pi072 & w8366 ;
  assign w8368 = w8019 & w8170 ;
  assign w8369 = ~w8027 & w8064 ;
  assign w8370 = w8065 ^ w8369 ;
  assign w8371 = ~w8170 & w8370 ;
  assign w8372 = w8368 | w8371 ;
  assign w8373 = ~\pi071 & w8372 ;
  assign w8374 = w8026 & w8170 ;
  assign w8375 = ~w8034 & w8061 ;
  assign w8376 = w8062 ^ w8375 ;
  assign w8377 = ~w8170 & w8376 ;
  assign w8378 = w8374 | w8377 ;
  assign w8379 = ~\pi070 & w8378 ;
  assign w8380 = w8033 & w8170 ;
  assign w8381 = ~w8042 & w8058 ;
  assign w8382 = w8059 ^ w8381 ;
  assign w8383 = ~w8170 & w8382 ;
  assign w8384 = w8380 | w8383 ;
  assign w8385 = ~\pi069 & w8384 ;
  assign w8386 = w8041 & w8170 ;
  assign w8387 = ~w8047 & w8055 ;
  assign w8388 = w8056 ^ w8387 ;
  assign w8389 = ~w8170 & w8388 ;
  assign w8390 = w8386 | w8389 ;
  assign w8391 = ~\pi068 & w8390 ;
  assign w8392 = w8046 & w8170 ;
  assign w8393 = ~\pi024 & \pi064 ;
  assign w8394 = ( \pi065 & ~w8052 ) | ( \pi065 & w8393 ) | ( ~w8052 & w8393 ) ;
  assign w8395 = w8050 ^ w8394 ;
  assign w8396 = ( w8168 & w8169 ) | ( w8168 & w8395 ) | ( w8169 & w8395 ) ;
  assign w8397 = w8395 & ~w8396 ;
  assign w8398 = w8392 | w8397 ;
  assign w8399 = ~\pi067 & w8398 ;
  assign w8400 = \pi025 ^ \pi065 ;
  assign w8401 = \pi024 ^ w7783 ;
  assign w8402 = ( \pi064 & w8169 ) | ( \pi064 & w8401 ) | ( w8169 & w8401 ) ;
  assign w8403 = w8400 ^ w8402 ;
  assign w8404 = ~w8169 & w8403 ;
  assign w8405 = ~w8168 & w8404 ;
  assign w8406 = ( ~\pi064 & w7783 ) | ( ~\pi064 & w8170 ) | ( w7783 & w8170 ) ;
  assign w8407 = \pi025 ^ w8406 ;
  assign w8408 = w8170 & ~w8407 ;
  assign w8409 = w8405 | w8408 ;
  assign w8410 = ~\pi066 & w8409 ;
  assign w8411 = \pi064 & ~\pi104 ;
  assign w8412 = ~w449 & w8411 ;
  assign w8413 = ~w7776 & w8412 ;
  assign w8414 = ( \pi024 & w8168 ) | ( \pi024 & ~w8413 ) | ( w8168 & ~w8413 ) ;
  assign w8415 = \pi024 & w8414 ;
  assign w8416 = ( ~\pi024 & w158 ) | ( ~\pi024 & w168 ) | ( w158 & w168 ) ;
  assign w8417 = w155 | w8168 ;
  assign w8418 = ( ~\pi024 & \pi064 ) | ( ~\pi024 & w155 ) | ( \pi064 & w155 ) ;
  assign w8419 = ~w8417 & w8418 ;
  assign w8420 = ~w8416 & w8419 ;
  assign w8421 = w8415 | w8420 ;
  assign w8422 = ~\pi023 & \pi064 ;
  assign w8423 = w8170 | w8405 ;
  assign w8424 = ( w8052 & w8405 ) | ( w8052 & w8423 ) | ( w8405 & w8423 ) ;
  assign w8425 = \pi066 ^ w8424 ;
  assign w8426 = ( \pi065 & ~w8421 ) | ( \pi065 & w8422 ) | ( ~w8421 & w8422 ) ;
  assign w8427 = w8425 | w8426 ;
  assign w8428 = \pi067 ^ w8398 ;
  assign w8429 = ( ~w8410 & w8427 ) | ( ~w8410 & w8428 ) | ( w8427 & w8428 ) ;
  assign w8430 = w8428 | w8429 ;
  assign w8431 = \pi068 ^ w8390 ;
  assign w8432 = ( ~w8399 & w8430 ) | ( ~w8399 & w8431 ) | ( w8430 & w8431 ) ;
  assign w8433 = w8431 | w8432 ;
  assign w8434 = \pi069 ^ w8384 ;
  assign w8435 = ( ~w8391 & w8433 ) | ( ~w8391 & w8434 ) | ( w8433 & w8434 ) ;
  assign w8436 = w8434 | w8435 ;
  assign w8437 = \pi070 ^ w8378 ;
  assign w8438 = ( ~w8385 & w8436 ) | ( ~w8385 & w8437 ) | ( w8436 & w8437 ) ;
  assign w8439 = w8437 | w8438 ;
  assign w8440 = \pi071 ^ w8372 ;
  assign w8441 = ( ~w8379 & w8439 ) | ( ~w8379 & w8440 ) | ( w8439 & w8440 ) ;
  assign w8442 = w8440 | w8441 ;
  assign w8443 = \pi072 ^ w8366 ;
  assign w8444 = ( ~w8373 & w8442 ) | ( ~w8373 & w8443 ) | ( w8442 & w8443 ) ;
  assign w8445 = w8443 | w8444 ;
  assign w8446 = \pi073 ^ w8360 ;
  assign w8447 = ( ~w8367 & w8445 ) | ( ~w8367 & w8446 ) | ( w8445 & w8446 ) ;
  assign w8448 = w8446 | w8447 ;
  assign w8449 = \pi074 ^ w8354 ;
  assign w8450 = ( ~w8361 & w8448 ) | ( ~w8361 & w8449 ) | ( w8448 & w8449 ) ;
  assign w8451 = w8449 | w8450 ;
  assign w8452 = \pi075 ^ w8348 ;
  assign w8453 = ( ~w8355 & w8451 ) | ( ~w8355 & w8452 ) | ( w8451 & w8452 ) ;
  assign w8454 = w8452 | w8453 ;
  assign w8455 = \pi076 ^ w8342 ;
  assign w8456 = ( ~w8349 & w8454 ) | ( ~w8349 & w8455 ) | ( w8454 & w8455 ) ;
  assign w8457 = w8455 | w8456 ;
  assign w8458 = \pi077 ^ w8336 ;
  assign w8459 = ( ~w8343 & w8457 ) | ( ~w8343 & w8458 ) | ( w8457 & w8458 ) ;
  assign w8460 = w8458 | w8459 ;
  assign w8461 = \pi078 ^ w8330 ;
  assign w8462 = ( ~w8337 & w8460 ) | ( ~w8337 & w8461 ) | ( w8460 & w8461 ) ;
  assign w8463 = w8461 | w8462 ;
  assign w8464 = \pi079 ^ w8324 ;
  assign w8465 = ( ~w8331 & w8463 ) | ( ~w8331 & w8464 ) | ( w8463 & w8464 ) ;
  assign w8466 = w8464 | w8465 ;
  assign w8467 = \pi080 ^ w8318 ;
  assign w8468 = ( ~w8325 & w8466 ) | ( ~w8325 & w8467 ) | ( w8466 & w8467 ) ;
  assign w8469 = w8467 | w8468 ;
  assign w8470 = \pi081 ^ w8312 ;
  assign w8471 = ( ~w8319 & w8469 ) | ( ~w8319 & w8470 ) | ( w8469 & w8470 ) ;
  assign w8472 = w8470 | w8471 ;
  assign w8473 = \pi082 ^ w8306 ;
  assign w8474 = ( ~w8313 & w8472 ) | ( ~w8313 & w8473 ) | ( w8472 & w8473 ) ;
  assign w8475 = w8473 | w8474 ;
  assign w8476 = \pi083 ^ w8300 ;
  assign w8477 = ( ~w8307 & w8475 ) | ( ~w8307 & w8476 ) | ( w8475 & w8476 ) ;
  assign w8478 = w8476 | w8477 ;
  assign w8479 = \pi084 ^ w8294 ;
  assign w8480 = ( ~w8301 & w8478 ) | ( ~w8301 & w8479 ) | ( w8478 & w8479 ) ;
  assign w8481 = w8479 | w8480 ;
  assign w8482 = \pi085 ^ w8288 ;
  assign w8483 = ( ~w8295 & w8481 ) | ( ~w8295 & w8482 ) | ( w8481 & w8482 ) ;
  assign w8484 = w8482 | w8483 ;
  assign w8485 = \pi086 ^ w8282 ;
  assign w8486 = ( ~w8289 & w8484 ) | ( ~w8289 & w8485 ) | ( w8484 & w8485 ) ;
  assign w8487 = w8485 | w8486 ;
  assign w8488 = \pi087 ^ w8276 ;
  assign w8489 = ( ~w8283 & w8487 ) | ( ~w8283 & w8488 ) | ( w8487 & w8488 ) ;
  assign w8490 = w8488 | w8489 ;
  assign w8491 = \pi088 ^ w8270 ;
  assign w8492 = ( ~w8277 & w8490 ) | ( ~w8277 & w8491 ) | ( w8490 & w8491 ) ;
  assign w8493 = w8491 | w8492 ;
  assign w8494 = \pi089 ^ w8264 ;
  assign w8495 = ( ~w8271 & w8493 ) | ( ~w8271 & w8494 ) | ( w8493 & w8494 ) ;
  assign w8496 = w8494 | w8495 ;
  assign w8497 = \pi090 ^ w8258 ;
  assign w8498 = ( ~w8265 & w8496 ) | ( ~w8265 & w8497 ) | ( w8496 & w8497 ) ;
  assign w8499 = w8497 | w8498 ;
  assign w8500 = \pi091 ^ w8252 ;
  assign w8501 = ( ~w8259 & w8499 ) | ( ~w8259 & w8500 ) | ( w8499 & w8500 ) ;
  assign w8502 = w8500 | w8501 ;
  assign w8503 = \pi092 ^ w8246 ;
  assign w8504 = ( ~w8253 & w8502 ) | ( ~w8253 & w8503 ) | ( w8502 & w8503 ) ;
  assign w8505 = w8503 | w8504 ;
  assign w8506 = \pi093 ^ w8240 ;
  assign w8507 = ( ~w8247 & w8505 ) | ( ~w8247 & w8506 ) | ( w8505 & w8506 ) ;
  assign w8508 = w8506 | w8507 ;
  assign w8509 = \pi094 ^ w8234 ;
  assign w8510 = ( ~w8241 & w8508 ) | ( ~w8241 & w8509 ) | ( w8508 & w8509 ) ;
  assign w8511 = w8509 | w8510 ;
  assign w8512 = \pi095 ^ w8228 ;
  assign w8513 = ( ~w8235 & w8511 ) | ( ~w8235 & w8512 ) | ( w8511 & w8512 ) ;
  assign w8514 = w8512 | w8513 ;
  assign w8515 = \pi096 ^ w8222 ;
  assign w8516 = ( ~w8229 & w8514 ) | ( ~w8229 & w8515 ) | ( w8514 & w8515 ) ;
  assign w8517 = w8515 | w8516 ;
  assign w8518 = \pi097 ^ w8216 ;
  assign w8519 = ( ~w8223 & w8517 ) | ( ~w8223 & w8518 ) | ( w8517 & w8518 ) ;
  assign w8520 = w8518 | w8519 ;
  assign w8521 = \pi098 ^ w8210 ;
  assign w8522 = ( ~w8217 & w8520 ) | ( ~w8217 & w8521 ) | ( w8520 & w8521 ) ;
  assign w8523 = w8521 | w8522 ;
  assign w8524 = \pi099 ^ w8204 ;
  assign w8525 = ( ~w8211 & w8523 ) | ( ~w8211 & w8524 ) | ( w8523 & w8524 ) ;
  assign w8526 = w8524 | w8525 ;
  assign w8527 = \pi100 ^ w8198 ;
  assign w8528 = ( ~w8205 & w8526 ) | ( ~w8205 & w8527 ) | ( w8526 & w8527 ) ;
  assign w8529 = w8527 | w8528 ;
  assign w8530 = \pi101 ^ w8192 ;
  assign w8531 = ( ~w8199 & w8529 ) | ( ~w8199 & w8530 ) | ( w8529 & w8530 ) ;
  assign w8532 = w8530 | w8531 ;
  assign w8533 = \pi102 ^ w8186 ;
  assign w8534 = ( ~w8193 & w8532 ) | ( ~w8193 & w8533 ) | ( w8532 & w8533 ) ;
  assign w8535 = w8533 | w8534 ;
  assign w8536 = \pi103 ^ w8175 ;
  assign w8537 = ( ~w8187 & w8535 ) | ( ~w8187 & w8536 ) | ( w8535 & w8536 ) ;
  assign w8538 = w8536 | w8537 ;
  assign w8539 = \pi104 ^ w8180 ;
  assign w8540 = w8181 & ~w8539 ;
  assign w8541 = ( w8538 & w8539 ) | ( w8538 & ~w8540 ) | ( w8539 & ~w8540 ) ;
  assign w8542 = ~\pi104 & w8180 ;
  assign w8543 = w8541 & ~w8542 ;
  assign w8544 = w6588 | w8543 ;
  assign w8545 = w8175 & w8544 ;
  assign w8546 = ~w8187 & w8535 ;
  assign w8547 = w8536 ^ w8546 ;
  assign w8548 = ~w8544 & w8547 ;
  assign w8549 = w8545 | w8548 ;
  assign w8550 = ~\pi104 & w8549 ;
  assign w8551 = w8186 & w8544 ;
  assign w8552 = ~w8193 & w8532 ;
  assign w8553 = w8533 ^ w8552 ;
  assign w8554 = ~w8544 & w8553 ;
  assign w8555 = w8551 | w8554 ;
  assign w8556 = ~\pi103 & w8555 ;
  assign w8557 = w8192 & w8544 ;
  assign w8558 = ~w8199 & w8529 ;
  assign w8559 = w8530 ^ w8558 ;
  assign w8560 = ~w8544 & w8559 ;
  assign w8561 = w8557 | w8560 ;
  assign w8562 = ~\pi102 & w8561 ;
  assign w8563 = w8198 & w8544 ;
  assign w8564 = ~w8205 & w8526 ;
  assign w8565 = w8527 ^ w8564 ;
  assign w8566 = ~w8544 & w8565 ;
  assign w8567 = w8563 | w8566 ;
  assign w8568 = ~\pi101 & w8567 ;
  assign w8569 = w8204 & w8544 ;
  assign w8570 = ~w8211 & w8523 ;
  assign w8571 = w8524 ^ w8570 ;
  assign w8572 = ~w8544 & w8571 ;
  assign w8573 = w8569 | w8572 ;
  assign w8574 = ~\pi100 & w8573 ;
  assign w8575 = w8210 & w8544 ;
  assign w8576 = ~w8217 & w8520 ;
  assign w8577 = w8521 ^ w8576 ;
  assign w8578 = ~w8544 & w8577 ;
  assign w8579 = w8575 | w8578 ;
  assign w8580 = ~\pi099 & w8579 ;
  assign w8581 = w8216 & w8544 ;
  assign w8582 = ~w8223 & w8517 ;
  assign w8583 = w8518 ^ w8582 ;
  assign w8584 = ~w8544 & w8583 ;
  assign w8585 = w8581 | w8584 ;
  assign w8586 = ~\pi098 & w8585 ;
  assign w8587 = w8222 & w8544 ;
  assign w8588 = ~w8229 & w8514 ;
  assign w8589 = w8515 ^ w8588 ;
  assign w8590 = ~w8544 & w8589 ;
  assign w8591 = w8587 | w8590 ;
  assign w8592 = ~\pi097 & w8591 ;
  assign w8593 = w8228 & w8544 ;
  assign w8594 = ~w8235 & w8511 ;
  assign w8595 = w8512 ^ w8594 ;
  assign w8596 = ~w8544 & w8595 ;
  assign w8597 = w8593 | w8596 ;
  assign w8598 = ~\pi096 & w8597 ;
  assign w8599 = w8234 & w8544 ;
  assign w8600 = ~w8241 & w8508 ;
  assign w8601 = w8509 ^ w8600 ;
  assign w8602 = ~w8544 & w8601 ;
  assign w8603 = w8599 | w8602 ;
  assign w8604 = ~\pi095 & w8603 ;
  assign w8605 = w8240 & w8544 ;
  assign w8606 = ~w8247 & w8505 ;
  assign w8607 = w8506 ^ w8606 ;
  assign w8608 = ~w8544 & w8607 ;
  assign w8609 = w8605 | w8608 ;
  assign w8610 = ~\pi094 & w8609 ;
  assign w8611 = w8246 & w8544 ;
  assign w8612 = ~w8253 & w8502 ;
  assign w8613 = w8503 ^ w8612 ;
  assign w8614 = ~w8544 & w8613 ;
  assign w8615 = w8611 | w8614 ;
  assign w8616 = ~\pi093 & w8615 ;
  assign w8617 = w8252 & w8544 ;
  assign w8618 = ~w8259 & w8499 ;
  assign w8619 = w8500 ^ w8618 ;
  assign w8620 = ~w8544 & w8619 ;
  assign w8621 = w8617 | w8620 ;
  assign w8622 = ~\pi092 & w8621 ;
  assign w8623 = w8258 & w8544 ;
  assign w8624 = ~w8265 & w8496 ;
  assign w8625 = w8497 ^ w8624 ;
  assign w8626 = ~w8544 & w8625 ;
  assign w8627 = w8623 | w8626 ;
  assign w8628 = ~\pi091 & w8627 ;
  assign w8629 = w8264 & w8544 ;
  assign w8630 = ~w8271 & w8493 ;
  assign w8631 = w8494 ^ w8630 ;
  assign w8632 = ~w8544 & w8631 ;
  assign w8633 = w8629 | w8632 ;
  assign w8634 = ~\pi090 & w8633 ;
  assign w8635 = w8270 & w8544 ;
  assign w8636 = ~w8277 & w8490 ;
  assign w8637 = w8491 ^ w8636 ;
  assign w8638 = ~w8544 & w8637 ;
  assign w8639 = w8635 | w8638 ;
  assign w8640 = ~\pi089 & w8639 ;
  assign w8641 = w8276 & w8544 ;
  assign w8642 = ~w8283 & w8487 ;
  assign w8643 = w8488 ^ w8642 ;
  assign w8644 = ~w8544 & w8643 ;
  assign w8645 = w8641 | w8644 ;
  assign w8646 = ~\pi088 & w8645 ;
  assign w8647 = w8282 & w8544 ;
  assign w8648 = ~w8289 & w8484 ;
  assign w8649 = w8485 ^ w8648 ;
  assign w8650 = ~w8544 & w8649 ;
  assign w8651 = w8647 | w8650 ;
  assign w8652 = ~\pi087 & w8651 ;
  assign w8653 = w8288 & w8544 ;
  assign w8654 = ~w8295 & w8481 ;
  assign w8655 = w8482 ^ w8654 ;
  assign w8656 = ~w8544 & w8655 ;
  assign w8657 = w8653 | w8656 ;
  assign w8658 = ~\pi086 & w8657 ;
  assign w8659 = w8294 & w8544 ;
  assign w8660 = ~w8301 & w8478 ;
  assign w8661 = w8479 ^ w8660 ;
  assign w8662 = ~w8544 & w8661 ;
  assign w8663 = w8659 | w8662 ;
  assign w8664 = ~\pi085 & w8663 ;
  assign w8665 = w8300 & w8544 ;
  assign w8666 = ~w8307 & w8475 ;
  assign w8667 = w8476 ^ w8666 ;
  assign w8668 = ~w8544 & w8667 ;
  assign w8669 = w8665 | w8668 ;
  assign w8670 = ~\pi084 & w8669 ;
  assign w8671 = w8306 & w8544 ;
  assign w8672 = ~w8313 & w8472 ;
  assign w8673 = w8473 ^ w8672 ;
  assign w8674 = ~w8544 & w8673 ;
  assign w8675 = w8671 | w8674 ;
  assign w8676 = ~\pi083 & w8675 ;
  assign w8677 = w8312 & w8544 ;
  assign w8678 = ~w8319 & w8469 ;
  assign w8679 = w8470 ^ w8678 ;
  assign w8680 = ~w8544 & w8679 ;
  assign w8681 = w8677 | w8680 ;
  assign w8682 = ~\pi082 & w8681 ;
  assign w8683 = w8318 & w8544 ;
  assign w8684 = ~w8325 & w8466 ;
  assign w8685 = w8467 ^ w8684 ;
  assign w8686 = ~w8544 & w8685 ;
  assign w8687 = w8683 | w8686 ;
  assign w8688 = ~\pi081 & w8687 ;
  assign w8689 = w8324 & w8544 ;
  assign w8690 = ~w8331 & w8463 ;
  assign w8691 = w8464 ^ w8690 ;
  assign w8692 = ~w8544 & w8691 ;
  assign w8693 = w8689 | w8692 ;
  assign w8694 = ~\pi080 & w8693 ;
  assign w8695 = w8330 & w8544 ;
  assign w8696 = ~w8337 & w8460 ;
  assign w8697 = w8461 ^ w8696 ;
  assign w8698 = ~w8544 & w8697 ;
  assign w8699 = w8695 | w8698 ;
  assign w8700 = ~\pi079 & w8699 ;
  assign w8701 = w8336 & w8544 ;
  assign w8702 = ~w8343 & w8457 ;
  assign w8703 = w8458 ^ w8702 ;
  assign w8704 = ~w8544 & w8703 ;
  assign w8705 = w8701 | w8704 ;
  assign w8706 = ~\pi078 & w8705 ;
  assign w8707 = w8342 & w8544 ;
  assign w8708 = ~w8349 & w8454 ;
  assign w8709 = w8455 ^ w8708 ;
  assign w8710 = ~w8544 & w8709 ;
  assign w8711 = w8707 | w8710 ;
  assign w8712 = ~\pi077 & w8711 ;
  assign w8713 = w8348 & w8544 ;
  assign w8714 = ~w8355 & w8451 ;
  assign w8715 = w8452 ^ w8714 ;
  assign w8716 = ~w8544 & w8715 ;
  assign w8717 = w8713 | w8716 ;
  assign w8718 = ~\pi076 & w8717 ;
  assign w8719 = w8354 & w8544 ;
  assign w8720 = ~w8361 & w8448 ;
  assign w8721 = w8449 ^ w8720 ;
  assign w8722 = ~w8544 & w8721 ;
  assign w8723 = w8719 | w8722 ;
  assign w8724 = ~\pi075 & w8723 ;
  assign w8725 = w8360 & w8544 ;
  assign w8726 = ~w8367 & w8445 ;
  assign w8727 = w8446 ^ w8726 ;
  assign w8728 = ~w8544 & w8727 ;
  assign w8729 = w8725 | w8728 ;
  assign w8730 = ~\pi074 & w8729 ;
  assign w8731 = w8366 & w8544 ;
  assign w8732 = ~w8373 & w8442 ;
  assign w8733 = w8443 ^ w8732 ;
  assign w8734 = ~w8544 & w8733 ;
  assign w8735 = w8731 | w8734 ;
  assign w8736 = ~\pi073 & w8735 ;
  assign w8737 = w8372 & w8544 ;
  assign w8738 = ~w8379 & w8439 ;
  assign w8739 = w8440 ^ w8738 ;
  assign w8740 = ~w8544 & w8739 ;
  assign w8741 = w8737 | w8740 ;
  assign w8742 = ~\pi072 & w8741 ;
  assign w8743 = w8378 & w8544 ;
  assign w8744 = ~w8385 & w8436 ;
  assign w8745 = w8437 ^ w8744 ;
  assign w8746 = ~w8544 & w8745 ;
  assign w8747 = w8743 | w8746 ;
  assign w8748 = ~\pi071 & w8747 ;
  assign w8749 = w8384 & w8544 ;
  assign w8750 = ~w8391 & w8433 ;
  assign w8751 = w8434 ^ w8750 ;
  assign w8752 = ~w8544 & w8751 ;
  assign w8753 = w8749 | w8752 ;
  assign w8754 = ~\pi070 & w8753 ;
  assign w8755 = w8390 & w8544 ;
  assign w8756 = ~w8399 & w8430 ;
  assign w8757 = w8431 ^ w8756 ;
  assign w8758 = ~w8544 & w8757 ;
  assign w8759 = w8755 | w8758 ;
  assign w8760 = ~\pi069 & w8759 ;
  assign w8761 = w8398 & w8544 ;
  assign w8762 = ~w8410 & w8427 ;
  assign w8763 = w8428 ^ w8762 ;
  assign w8764 = ~w8544 & w8763 ;
  assign w8765 = w8761 | w8764 ;
  assign w8766 = ~\pi068 & w8765 ;
  assign w8767 = w8409 & w8544 ;
  assign w8768 = w8425 ^ w8426 ;
  assign w8769 = ( w6588 & w8543 ) | ( w6588 & w8768 ) | ( w8543 & w8768 ) ;
  assign w8770 = w8768 & ~w8769 ;
  assign w8771 = w8767 | w8770 ;
  assign w8772 = ~\pi067 & w8771 ;
  assign w8773 = ( ~w6588 & w8415 ) | ( ~w6588 & w8420 ) | ( w8415 & w8420 ) ;
  assign w8774 = \pi065 ^ w8773 ;
  assign w8775 = ( ~w6588 & w8422 ) | ( ~w6588 & w8774 ) | ( w8422 & w8774 ) ;
  assign w8776 = ( w8422 & w8543 ) | ( w8422 & w8774 ) | ( w8543 & w8774 ) ;
  assign w8777 = w8775 & ~w8776 ;
  assign w8778 = ( w8421 & w8544 ) | ( w8421 & w8777 ) | ( w8544 & w8777 ) ;
  assign w8779 = w8777 | w8778 ;
  assign w8780 = ~\pi066 & w8779 ;
  assign w8781 = ( \pi064 & ~\pi105 ) | ( \pi064 & \pi106 ) | ( ~\pi105 & \pi106 ) ;
  assign w8782 = w167 | w201 ;
  assign w8783 = ( \pi106 & \pi107 ) | ( \pi106 & ~w167 ) | ( \pi107 & ~w167 ) ;
  assign w8784 = w8782 | w8783 ;
  assign w8785 = w8781 & ~w8784 ;
  assign w8786 = ( \pi023 & w8543 ) | ( \pi023 & ~w8785 ) | ( w8543 & ~w8785 ) ;
  assign w8787 = \pi023 & w8786 ;
  assign w8788 = ~w449 & w8422 ;
  assign w8789 = ~w7776 & w8788 ;
  assign w8790 = ~w8543 & w8789 ;
  assign w8791 = w8787 | w8790 ;
  assign w8792 = ~\pi022 & \pi064 ;
  assign w8793 = \pi065 ^ w8791 ;
  assign w8794 = w8792 | w8793 ;
  assign w8795 = ~w8421 & w8544 ;
  assign w8796 = ( w8544 & w8777 ) | ( w8544 & ~w8795 ) | ( w8777 & ~w8795 ) ;
  assign w8797 = \pi066 ^ w8796 ;
  assign w8798 = ~\pi065 & w8791 ;
  assign w8799 = w8794 | w8798 ;
  assign w8800 = ( w8797 & ~w8798 ) | ( w8797 & w8799 ) | ( ~w8798 & w8799 ) ;
  assign w8801 = \pi067 ^ w8771 ;
  assign w8802 = ( ~w8780 & w8800 ) | ( ~w8780 & w8801 ) | ( w8800 & w8801 ) ;
  assign w8803 = w8801 | w8802 ;
  assign w8804 = \pi068 ^ w8765 ;
  assign w8805 = ( ~w8772 & w8803 ) | ( ~w8772 & w8804 ) | ( w8803 & w8804 ) ;
  assign w8806 = w8804 | w8805 ;
  assign w8807 = \pi069 ^ w8759 ;
  assign w8808 = ( ~w8766 & w8806 ) | ( ~w8766 & w8807 ) | ( w8806 & w8807 ) ;
  assign w8809 = w8807 | w8808 ;
  assign w8810 = \pi070 ^ w8753 ;
  assign w8811 = ( ~w8760 & w8809 ) | ( ~w8760 & w8810 ) | ( w8809 & w8810 ) ;
  assign w8812 = w8810 | w8811 ;
  assign w8813 = \pi071 ^ w8747 ;
  assign w8814 = ( ~w8754 & w8812 ) | ( ~w8754 & w8813 ) | ( w8812 & w8813 ) ;
  assign w8815 = w8813 | w8814 ;
  assign w8816 = \pi072 ^ w8741 ;
  assign w8817 = ( ~w8748 & w8815 ) | ( ~w8748 & w8816 ) | ( w8815 & w8816 ) ;
  assign w8818 = w8816 | w8817 ;
  assign w8819 = \pi073 ^ w8735 ;
  assign w8820 = ( ~w8742 & w8818 ) | ( ~w8742 & w8819 ) | ( w8818 & w8819 ) ;
  assign w8821 = w8819 | w8820 ;
  assign w8822 = \pi074 ^ w8729 ;
  assign w8823 = ( ~w8736 & w8821 ) | ( ~w8736 & w8822 ) | ( w8821 & w8822 ) ;
  assign w8824 = w8822 | w8823 ;
  assign w8825 = \pi075 ^ w8723 ;
  assign w8826 = ( ~w8730 & w8824 ) | ( ~w8730 & w8825 ) | ( w8824 & w8825 ) ;
  assign w8827 = w8825 | w8826 ;
  assign w8828 = \pi076 ^ w8717 ;
  assign w8829 = ( ~w8724 & w8827 ) | ( ~w8724 & w8828 ) | ( w8827 & w8828 ) ;
  assign w8830 = w8828 | w8829 ;
  assign w8831 = \pi077 ^ w8711 ;
  assign w8832 = ( ~w8718 & w8830 ) | ( ~w8718 & w8831 ) | ( w8830 & w8831 ) ;
  assign w8833 = w8831 | w8832 ;
  assign w8834 = \pi078 ^ w8705 ;
  assign w8835 = ( ~w8712 & w8833 ) | ( ~w8712 & w8834 ) | ( w8833 & w8834 ) ;
  assign w8836 = w8834 | w8835 ;
  assign w8837 = \pi079 ^ w8699 ;
  assign w8838 = ( ~w8706 & w8836 ) | ( ~w8706 & w8837 ) | ( w8836 & w8837 ) ;
  assign w8839 = w8837 | w8838 ;
  assign w8840 = \pi080 ^ w8693 ;
  assign w8841 = ( ~w8700 & w8839 ) | ( ~w8700 & w8840 ) | ( w8839 & w8840 ) ;
  assign w8842 = w8840 | w8841 ;
  assign w8843 = \pi081 ^ w8687 ;
  assign w8844 = ( ~w8694 & w8842 ) | ( ~w8694 & w8843 ) | ( w8842 & w8843 ) ;
  assign w8845 = w8843 | w8844 ;
  assign w8846 = \pi082 ^ w8681 ;
  assign w8847 = ( ~w8688 & w8845 ) | ( ~w8688 & w8846 ) | ( w8845 & w8846 ) ;
  assign w8848 = w8846 | w8847 ;
  assign w8849 = \pi083 ^ w8675 ;
  assign w8850 = ( ~w8682 & w8848 ) | ( ~w8682 & w8849 ) | ( w8848 & w8849 ) ;
  assign w8851 = w8849 | w8850 ;
  assign w8852 = \pi084 ^ w8669 ;
  assign w8853 = ( ~w8676 & w8851 ) | ( ~w8676 & w8852 ) | ( w8851 & w8852 ) ;
  assign w8854 = w8852 | w8853 ;
  assign w8855 = \pi085 ^ w8663 ;
  assign w8856 = ( ~w8670 & w8854 ) | ( ~w8670 & w8855 ) | ( w8854 & w8855 ) ;
  assign w8857 = w8855 | w8856 ;
  assign w8858 = \pi086 ^ w8657 ;
  assign w8859 = ( ~w8664 & w8857 ) | ( ~w8664 & w8858 ) | ( w8857 & w8858 ) ;
  assign w8860 = w8858 | w8859 ;
  assign w8861 = \pi087 ^ w8651 ;
  assign w8862 = ( ~w8658 & w8860 ) | ( ~w8658 & w8861 ) | ( w8860 & w8861 ) ;
  assign w8863 = w8861 | w8862 ;
  assign w8864 = \pi088 ^ w8645 ;
  assign w8865 = ( ~w8652 & w8863 ) | ( ~w8652 & w8864 ) | ( w8863 & w8864 ) ;
  assign w8866 = w8864 | w8865 ;
  assign w8867 = \pi089 ^ w8639 ;
  assign w8868 = ( ~w8646 & w8866 ) | ( ~w8646 & w8867 ) | ( w8866 & w8867 ) ;
  assign w8869 = w8867 | w8868 ;
  assign w8870 = \pi090 ^ w8633 ;
  assign w8871 = ( ~w8640 & w8869 ) | ( ~w8640 & w8870 ) | ( w8869 & w8870 ) ;
  assign w8872 = w8870 | w8871 ;
  assign w8873 = \pi091 ^ w8627 ;
  assign w8874 = ( ~w8634 & w8872 ) | ( ~w8634 & w8873 ) | ( w8872 & w8873 ) ;
  assign w8875 = w8873 | w8874 ;
  assign w8876 = \pi092 ^ w8621 ;
  assign w8877 = ( ~w8628 & w8875 ) | ( ~w8628 & w8876 ) | ( w8875 & w8876 ) ;
  assign w8878 = w8876 | w8877 ;
  assign w8879 = \pi093 ^ w8615 ;
  assign w8880 = ( ~w8622 & w8878 ) | ( ~w8622 & w8879 ) | ( w8878 & w8879 ) ;
  assign w8881 = w8879 | w8880 ;
  assign w8882 = \pi094 ^ w8609 ;
  assign w8883 = ( ~w8616 & w8881 ) | ( ~w8616 & w8882 ) | ( w8881 & w8882 ) ;
  assign w8884 = w8882 | w8883 ;
  assign w8885 = \pi095 ^ w8603 ;
  assign w8886 = ( ~w8610 & w8884 ) | ( ~w8610 & w8885 ) | ( w8884 & w8885 ) ;
  assign w8887 = w8885 | w8886 ;
  assign w8888 = \pi096 ^ w8597 ;
  assign w8889 = ( ~w8604 & w8887 ) | ( ~w8604 & w8888 ) | ( w8887 & w8888 ) ;
  assign w8890 = w8888 | w8889 ;
  assign w8891 = \pi097 ^ w8591 ;
  assign w8892 = ( ~w8598 & w8890 ) | ( ~w8598 & w8891 ) | ( w8890 & w8891 ) ;
  assign w8893 = w8891 | w8892 ;
  assign w8894 = \pi098 ^ w8585 ;
  assign w8895 = ( ~w8592 & w8893 ) | ( ~w8592 & w8894 ) | ( w8893 & w8894 ) ;
  assign w8896 = w8894 | w8895 ;
  assign w8897 = \pi099 ^ w8579 ;
  assign w8898 = ( ~w8586 & w8896 ) | ( ~w8586 & w8897 ) | ( w8896 & w8897 ) ;
  assign w8899 = w8897 | w8898 ;
  assign w8900 = \pi100 ^ w8573 ;
  assign w8901 = ( ~w8580 & w8899 ) | ( ~w8580 & w8900 ) | ( w8899 & w8900 ) ;
  assign w8902 = w8900 | w8901 ;
  assign w8903 = \pi101 ^ w8567 ;
  assign w8904 = ( ~w8574 & w8902 ) | ( ~w8574 & w8903 ) | ( w8902 & w8903 ) ;
  assign w8905 = w8903 | w8904 ;
  assign w8906 = \pi102 ^ w8561 ;
  assign w8907 = ( ~w8568 & w8905 ) | ( ~w8568 & w8906 ) | ( w8905 & w8906 ) ;
  assign w8908 = w8906 | w8907 ;
  assign w8909 = \pi103 ^ w8555 ;
  assign w8910 = ( ~w8562 & w8908 ) | ( ~w8562 & w8909 ) | ( w8908 & w8909 ) ;
  assign w8911 = w8909 | w8910 ;
  assign w8912 = \pi104 ^ w8549 ;
  assign w8913 = ( ~w8556 & w8911 ) | ( ~w8556 & w8912 ) | ( w8911 & w8912 ) ;
  assign w8914 = w8912 | w8913 ;
  assign w8915 = w8180 & w8544 ;
  assign w8916 = ~w8181 & w8538 ;
  assign w8917 = w8539 ^ w8916 ;
  assign w8918 = ~w8544 & w8917 ;
  assign w8919 = w8915 | w8918 ;
  assign w8920 = ~\pi105 & w8919 ;
  assign w8921 = ( \pi105 & ~w8915 ) | ( \pi105 & w8918 ) | ( ~w8915 & w8918 ) ;
  assign w8922 = ~w8918 & w8921 ;
  assign w8923 = ( ~\pi106 & \pi107 ) | ( ~\pi106 & w167 ) | ( \pi107 & w167 ) ;
  assign w8924 = \pi106 | w8923 ;
  assign w8925 = ( ~w8550 & w8914 ) | ( ~w8550 & w8920 ) | ( w8914 & w8920 ) ;
  assign w8926 = ( w8920 & w8924 ) | ( w8920 & ~w8925 ) | ( w8924 & ~w8925 ) ;
  assign w8927 = ( w201 & w8922 ) | ( w201 & ~w8925 ) | ( w8922 & ~w8925 ) ;
  assign w8928 = ( w8925 & ~w8926 ) | ( w8925 & w8927 ) | ( ~w8926 & w8927 ) ;
  assign w8929 = w8926 | w8928 ;
  assign w8930 = ~w6588 & w8919 ;
  assign w8931 = w8929 & ~w8930 ;
  assign w8932 = ~w8556 & w8911 ;
  assign w8933 = w8912 ^ w8932 ;
  assign w8934 = ~w8931 & w8933 ;
  assign w8935 = ( w8549 & w8929 ) | ( w8549 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8936 = ~w8930 & w8935 ;
  assign w8937 = w8934 | w8936 ;
  assign w8938 = w8920 | w8922 ;
  assign w8939 = ( ~w8550 & w8914 ) | ( ~w8550 & w8931 ) | ( w8914 & w8931 ) ;
  assign w8940 = w8938 ^ w8939 ;
  assign w8941 = ~w8931 & w8940 ;
  assign w8942 = ( w6588 & ~w8919 ) | ( w6588 & w8929 ) | ( ~w8919 & w8929 ) ;
  assign w8943 = w8919 & w8942 ;
  assign w8944 = w8941 | w8943 ;
  assign w8945 = ~\pi105 & w8937 ;
  assign w8946 = ~w8562 & w8908 ;
  assign w8947 = w8909 ^ w8946 ;
  assign w8948 = ~w8931 & w8947 ;
  assign w8949 = ( w8555 & w8929 ) | ( w8555 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8950 = ~w8930 & w8949 ;
  assign w8951 = w8948 | w8950 ;
  assign w8952 = ~\pi104 & w8951 ;
  assign w8953 = ~w8568 & w8905 ;
  assign w8954 = w8906 ^ w8953 ;
  assign w8955 = ~w8931 & w8954 ;
  assign w8956 = ( w8561 & w8929 ) | ( w8561 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8957 = ~w8930 & w8956 ;
  assign w8958 = w8955 | w8957 ;
  assign w8959 = ~\pi103 & w8958 ;
  assign w8960 = ~w8574 & w8902 ;
  assign w8961 = w8903 ^ w8960 ;
  assign w8962 = ~w8931 & w8961 ;
  assign w8963 = ( w8567 & w8929 ) | ( w8567 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8964 = ~w8930 & w8963 ;
  assign w8965 = w8962 | w8964 ;
  assign w8966 = ~\pi102 & w8965 ;
  assign w8967 = ~w8580 & w8899 ;
  assign w8968 = w8900 ^ w8967 ;
  assign w8969 = ~w8931 & w8968 ;
  assign w8970 = ( w8573 & w8929 ) | ( w8573 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8971 = ~w8930 & w8970 ;
  assign w8972 = w8969 | w8971 ;
  assign w8973 = ~\pi101 & w8972 ;
  assign w8974 = ~w8586 & w8896 ;
  assign w8975 = w8897 ^ w8974 ;
  assign w8976 = ~w8931 & w8975 ;
  assign w8977 = ( w8579 & w8929 ) | ( w8579 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8978 = ~w8930 & w8977 ;
  assign w8979 = w8976 | w8978 ;
  assign w8980 = ~\pi100 & w8979 ;
  assign w8981 = ~w8592 & w8893 ;
  assign w8982 = w8894 ^ w8981 ;
  assign w8983 = ~w8931 & w8982 ;
  assign w8984 = ( w8585 & w8929 ) | ( w8585 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8985 = ~w8930 & w8984 ;
  assign w8986 = w8983 | w8985 ;
  assign w8987 = ~\pi099 & w8986 ;
  assign w8988 = ~w8598 & w8890 ;
  assign w8989 = w8891 ^ w8988 ;
  assign w8990 = ~w8931 & w8989 ;
  assign w8991 = ( w8591 & w8929 ) | ( w8591 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8992 = ~w8930 & w8991 ;
  assign w8993 = w8990 | w8992 ;
  assign w8994 = ~\pi098 & w8993 ;
  assign w8995 = ~w8604 & w8887 ;
  assign w8996 = w8888 ^ w8995 ;
  assign w8997 = ~w8931 & w8996 ;
  assign w8998 = ( w8597 & w8929 ) | ( w8597 & w8930 ) | ( w8929 & w8930 ) ;
  assign w8999 = ~w8930 & w8998 ;
  assign w9000 = w8997 | w8999 ;
  assign w9001 = ~\pi097 & w9000 ;
  assign w9002 = ~w8610 & w8884 ;
  assign w9003 = w8885 ^ w9002 ;
  assign w9004 = ~w8931 & w9003 ;
  assign w9005 = ( w8603 & w8929 ) | ( w8603 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9006 = ~w8930 & w9005 ;
  assign w9007 = w9004 | w9006 ;
  assign w9008 = ~\pi096 & w9007 ;
  assign w9009 = ~w8616 & w8881 ;
  assign w9010 = w8882 ^ w9009 ;
  assign w9011 = ~w8931 & w9010 ;
  assign w9012 = ( w8609 & w8929 ) | ( w8609 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9013 = ~w8930 & w9012 ;
  assign w9014 = w9011 | w9013 ;
  assign w9015 = ~\pi095 & w9014 ;
  assign w9016 = ~w8622 & w8878 ;
  assign w9017 = w8879 ^ w9016 ;
  assign w9018 = ~w8931 & w9017 ;
  assign w9019 = ( w8615 & w8929 ) | ( w8615 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9020 = ~w8930 & w9019 ;
  assign w9021 = w9018 | w9020 ;
  assign w9022 = ~\pi094 & w9021 ;
  assign w9023 = ~w8628 & w8875 ;
  assign w9024 = w8876 ^ w9023 ;
  assign w9025 = ~w8931 & w9024 ;
  assign w9026 = ( w8621 & w8929 ) | ( w8621 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9027 = ~w8930 & w9026 ;
  assign w9028 = w9025 | w9027 ;
  assign w9029 = ~\pi093 & w9028 ;
  assign w9030 = ~w8634 & w8872 ;
  assign w9031 = w8873 ^ w9030 ;
  assign w9032 = ~w8931 & w9031 ;
  assign w9033 = ( w8627 & w8929 ) | ( w8627 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9034 = ~w8930 & w9033 ;
  assign w9035 = w9032 | w9034 ;
  assign w9036 = ~\pi092 & w9035 ;
  assign w9037 = ~w8640 & w8869 ;
  assign w9038 = w8870 ^ w9037 ;
  assign w9039 = ~w8931 & w9038 ;
  assign w9040 = ( w8633 & w8929 ) | ( w8633 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9041 = ~w8930 & w9040 ;
  assign w9042 = w9039 | w9041 ;
  assign w9043 = ~\pi091 & w9042 ;
  assign w9044 = ~w8646 & w8866 ;
  assign w9045 = w8867 ^ w9044 ;
  assign w9046 = ~w8931 & w9045 ;
  assign w9047 = ( w8639 & w8929 ) | ( w8639 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9048 = ~w8930 & w9047 ;
  assign w9049 = w9046 | w9048 ;
  assign w9050 = ~\pi090 & w9049 ;
  assign w9051 = ~w8652 & w8863 ;
  assign w9052 = w8864 ^ w9051 ;
  assign w9053 = ~w8931 & w9052 ;
  assign w9054 = ( w8645 & w8929 ) | ( w8645 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9055 = ~w8930 & w9054 ;
  assign w9056 = w9053 | w9055 ;
  assign w9057 = ~\pi089 & w9056 ;
  assign w9058 = ~w8658 & w8860 ;
  assign w9059 = w8861 ^ w9058 ;
  assign w9060 = ~w8931 & w9059 ;
  assign w9061 = ( w8651 & w8929 ) | ( w8651 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9062 = ~w8930 & w9061 ;
  assign w9063 = w9060 | w9062 ;
  assign w9064 = ~\pi088 & w9063 ;
  assign w9065 = ~w8664 & w8857 ;
  assign w9066 = w8858 ^ w9065 ;
  assign w9067 = ~w8931 & w9066 ;
  assign w9068 = ( w8657 & w8929 ) | ( w8657 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9069 = ~w8930 & w9068 ;
  assign w9070 = w9067 | w9069 ;
  assign w9071 = ~\pi087 & w9070 ;
  assign w9072 = ~w8670 & w8854 ;
  assign w9073 = w8855 ^ w9072 ;
  assign w9074 = ~w8931 & w9073 ;
  assign w9075 = ( w8663 & w8929 ) | ( w8663 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9076 = ~w8930 & w9075 ;
  assign w9077 = w9074 | w9076 ;
  assign w9078 = ~\pi086 & w9077 ;
  assign w9079 = ~w8676 & w8851 ;
  assign w9080 = w8852 ^ w9079 ;
  assign w9081 = ~w8931 & w9080 ;
  assign w9082 = ( w8669 & w8929 ) | ( w8669 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9083 = ~w8930 & w9082 ;
  assign w9084 = w9081 | w9083 ;
  assign w9085 = ~\pi085 & w9084 ;
  assign w9086 = ~w8682 & w8848 ;
  assign w9087 = w8849 ^ w9086 ;
  assign w9088 = ~w8931 & w9087 ;
  assign w9089 = ( w8675 & w8929 ) | ( w8675 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9090 = ~w8930 & w9089 ;
  assign w9091 = w9088 | w9090 ;
  assign w9092 = ~\pi084 & w9091 ;
  assign w9093 = ~w8688 & w8845 ;
  assign w9094 = w8846 ^ w9093 ;
  assign w9095 = ~w8931 & w9094 ;
  assign w9096 = ( w8681 & w8929 ) | ( w8681 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9097 = ~w8930 & w9096 ;
  assign w9098 = w9095 | w9097 ;
  assign w9099 = ~\pi083 & w9098 ;
  assign w9100 = ~w8694 & w8842 ;
  assign w9101 = w8843 ^ w9100 ;
  assign w9102 = ~w8931 & w9101 ;
  assign w9103 = ( w8687 & w8929 ) | ( w8687 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9104 = ~w8930 & w9103 ;
  assign w9105 = w9102 | w9104 ;
  assign w9106 = ~\pi082 & w9105 ;
  assign w9107 = ~w8700 & w8839 ;
  assign w9108 = w8840 ^ w9107 ;
  assign w9109 = ~w8931 & w9108 ;
  assign w9110 = ( w8693 & w8929 ) | ( w8693 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9111 = ~w8930 & w9110 ;
  assign w9112 = w9109 | w9111 ;
  assign w9113 = ~\pi081 & w9112 ;
  assign w9114 = ~w8706 & w8836 ;
  assign w9115 = w8837 ^ w9114 ;
  assign w9116 = ~w8931 & w9115 ;
  assign w9117 = ( w8699 & w8929 ) | ( w8699 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9118 = ~w8930 & w9117 ;
  assign w9119 = w9116 | w9118 ;
  assign w9120 = ~\pi080 & w9119 ;
  assign w9121 = ~w8712 & w8833 ;
  assign w9122 = w8834 ^ w9121 ;
  assign w9123 = ~w8931 & w9122 ;
  assign w9124 = ( w8705 & w8929 ) | ( w8705 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9125 = ~w8930 & w9124 ;
  assign w9126 = w9123 | w9125 ;
  assign w9127 = ~\pi079 & w9126 ;
  assign w9128 = ~w8718 & w8830 ;
  assign w9129 = w8831 ^ w9128 ;
  assign w9130 = ~w8931 & w9129 ;
  assign w9131 = ( w8711 & w8929 ) | ( w8711 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9132 = ~w8930 & w9131 ;
  assign w9133 = w9130 | w9132 ;
  assign w9134 = ~\pi078 & w9133 ;
  assign w9135 = ~w8724 & w8827 ;
  assign w9136 = w8828 ^ w9135 ;
  assign w9137 = ~w8931 & w9136 ;
  assign w9138 = ( w8717 & w8929 ) | ( w8717 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9139 = ~w8930 & w9138 ;
  assign w9140 = w9137 | w9139 ;
  assign w9141 = ~\pi077 & w9140 ;
  assign w9142 = ~w8730 & w8824 ;
  assign w9143 = w8825 ^ w9142 ;
  assign w9144 = ~w8931 & w9143 ;
  assign w9145 = ( w8723 & w8929 ) | ( w8723 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9146 = ~w8930 & w9145 ;
  assign w9147 = w9144 | w9146 ;
  assign w9148 = ~\pi076 & w9147 ;
  assign w9149 = ~w8736 & w8821 ;
  assign w9150 = w8822 ^ w9149 ;
  assign w9151 = ~w8931 & w9150 ;
  assign w9152 = ( w8729 & w8929 ) | ( w8729 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9153 = ~w8930 & w9152 ;
  assign w9154 = w9151 | w9153 ;
  assign w9155 = ~\pi075 & w9154 ;
  assign w9156 = ~w8742 & w8818 ;
  assign w9157 = w8819 ^ w9156 ;
  assign w9158 = ~w8931 & w9157 ;
  assign w9159 = ( w8735 & w8929 ) | ( w8735 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9160 = ~w8930 & w9159 ;
  assign w9161 = w9158 | w9160 ;
  assign w9162 = ~\pi074 & w9161 ;
  assign w9163 = ~w8748 & w8815 ;
  assign w9164 = w8816 ^ w9163 ;
  assign w9165 = ~w8931 & w9164 ;
  assign w9166 = ( w8741 & w8929 ) | ( w8741 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9167 = ~w8930 & w9166 ;
  assign w9168 = w9165 | w9167 ;
  assign w9169 = ~\pi073 & w9168 ;
  assign w9170 = ~w8754 & w8812 ;
  assign w9171 = w8813 ^ w9170 ;
  assign w9172 = ~w8931 & w9171 ;
  assign w9173 = ( w8747 & w8929 ) | ( w8747 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9174 = ~w8930 & w9173 ;
  assign w9175 = w9172 | w9174 ;
  assign w9176 = ~\pi072 & w9175 ;
  assign w9177 = ~w8760 & w8809 ;
  assign w9178 = w8810 ^ w9177 ;
  assign w9179 = ~w8931 & w9178 ;
  assign w9180 = ( w8753 & w8929 ) | ( w8753 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9181 = ~w8930 & w9180 ;
  assign w9182 = w9179 | w9181 ;
  assign w9183 = ~\pi071 & w9182 ;
  assign w9184 = ~w8766 & w8806 ;
  assign w9185 = w8807 ^ w9184 ;
  assign w9186 = ~w8931 & w9185 ;
  assign w9187 = ( w8759 & w8929 ) | ( w8759 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9188 = ~w8930 & w9187 ;
  assign w9189 = w9186 | w9188 ;
  assign w9190 = ~\pi070 & w9189 ;
  assign w9191 = ~w8772 & w8803 ;
  assign w9192 = w8804 ^ w9191 ;
  assign w9193 = ~w8931 & w9192 ;
  assign w9194 = ( w8765 & w8929 ) | ( w8765 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9195 = ~w8930 & w9194 ;
  assign w9196 = w9193 | w9195 ;
  assign w9197 = ~\pi069 & w9196 ;
  assign w9198 = ~w8780 & w8800 ;
  assign w9199 = w8801 ^ w9198 ;
  assign w9200 = ~w8931 & w9199 ;
  assign w9201 = ( w8771 & w8929 ) | ( w8771 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9202 = ~w8930 & w9201 ;
  assign w9203 = w9200 | w9202 ;
  assign w9204 = ~\pi068 & w9203 ;
  assign w9205 = ( \pi065 & w8791 ) | ( \pi065 & ~w8931 ) | ( w8791 & ~w8931 ) ;
  assign w9206 = ( \pi065 & w8794 ) | ( \pi065 & ~w9205 ) | ( w8794 & ~w9205 ) ;
  assign w9207 = w8797 ^ w9206 ;
  assign w9208 = ~w8931 & w9207 ;
  assign w9209 = ( w8779 & w8929 ) | ( w8779 & w8930 ) | ( w8929 & w8930 ) ;
  assign w9210 = ~w8930 & w9209 ;
  assign w9211 = w9208 | w9210 ;
  assign w9212 = ~\pi067 & w9211 ;
  assign w9213 = w8791 ^ w8792 ;
  assign w9214 = \pi065 ^ w9213 ;
  assign w9215 = w8931 ^ w9214 ;
  assign w9216 = ( w8791 & w9214 ) | ( w8791 & w9215 ) | ( w9214 & w9215 ) ;
  assign w9217 = ~\pi066 & w9216 ;
  assign w9218 = ~\pi021 & \pi064 ;
  assign w9219 = w8791 ^ w8931 ;
  assign w9220 = ( w8791 & w9214 ) | ( w8791 & ~w9219 ) | ( w9214 & ~w9219 ) ;
  assign w9221 = \pi066 ^ w9220 ;
  assign w9222 = \pi064 & ~w8931 ;
  assign w9223 = \pi022 ^ w9222 ;
  assign w9224 = ( ~\pi021 & \pi064 ) | ( ~\pi021 & w9221 ) | ( \pi064 & w9221 ) ;
  assign w9225 = ( \pi065 & ~w9223 ) | ( \pi065 & w9224 ) | ( ~w9223 & w9224 ) ;
  assign w9226 = w9221 | w9225 ;
  assign w9227 = \pi067 ^ w9211 ;
  assign w9228 = ( ~w9217 & w9226 ) | ( ~w9217 & w9227 ) | ( w9226 & w9227 ) ;
  assign w9229 = w9227 | w9228 ;
  assign w9230 = \pi068 ^ w9203 ;
  assign w9231 = ( ~w9212 & w9229 ) | ( ~w9212 & w9230 ) | ( w9229 & w9230 ) ;
  assign w9232 = w9230 | w9231 ;
  assign w9233 = \pi069 ^ w9196 ;
  assign w9234 = ( ~w9204 & w9232 ) | ( ~w9204 & w9233 ) | ( w9232 & w9233 ) ;
  assign w9235 = w9233 | w9234 ;
  assign w9236 = \pi070 ^ w9189 ;
  assign w9237 = ( ~w9197 & w9235 ) | ( ~w9197 & w9236 ) | ( w9235 & w9236 ) ;
  assign w9238 = w9236 | w9237 ;
  assign w9239 = \pi071 ^ w9182 ;
  assign w9240 = ( ~w9190 & w9238 ) | ( ~w9190 & w9239 ) | ( w9238 & w9239 ) ;
  assign w9241 = w9239 | w9240 ;
  assign w9242 = \pi072 ^ w9175 ;
  assign w9243 = ( ~w9183 & w9241 ) | ( ~w9183 & w9242 ) | ( w9241 & w9242 ) ;
  assign w9244 = w9242 | w9243 ;
  assign w9245 = \pi073 ^ w9168 ;
  assign w9246 = ( ~w9176 & w9244 ) | ( ~w9176 & w9245 ) | ( w9244 & w9245 ) ;
  assign w9247 = w9245 | w9246 ;
  assign w9248 = \pi074 ^ w9161 ;
  assign w9249 = ( ~w9169 & w9247 ) | ( ~w9169 & w9248 ) | ( w9247 & w9248 ) ;
  assign w9250 = w9248 | w9249 ;
  assign w9251 = \pi075 ^ w9154 ;
  assign w9252 = ( ~w9162 & w9250 ) | ( ~w9162 & w9251 ) | ( w9250 & w9251 ) ;
  assign w9253 = w9251 | w9252 ;
  assign w9254 = \pi076 ^ w9147 ;
  assign w9255 = ( ~w9155 & w9253 ) | ( ~w9155 & w9254 ) | ( w9253 & w9254 ) ;
  assign w9256 = w9254 | w9255 ;
  assign w9257 = \pi077 ^ w9140 ;
  assign w9258 = ( ~w9148 & w9256 ) | ( ~w9148 & w9257 ) | ( w9256 & w9257 ) ;
  assign w9259 = w9257 | w9258 ;
  assign w9260 = \pi078 ^ w9133 ;
  assign w9261 = ( ~w9141 & w9259 ) | ( ~w9141 & w9260 ) | ( w9259 & w9260 ) ;
  assign w9262 = w9260 | w9261 ;
  assign w9263 = \pi079 ^ w9126 ;
  assign w9264 = ( ~w9134 & w9262 ) | ( ~w9134 & w9263 ) | ( w9262 & w9263 ) ;
  assign w9265 = w9263 | w9264 ;
  assign w9266 = \pi080 ^ w9119 ;
  assign w9267 = ( ~w9127 & w9265 ) | ( ~w9127 & w9266 ) | ( w9265 & w9266 ) ;
  assign w9268 = w9266 | w9267 ;
  assign w9269 = \pi081 ^ w9112 ;
  assign w9270 = ( ~w9120 & w9268 ) | ( ~w9120 & w9269 ) | ( w9268 & w9269 ) ;
  assign w9271 = w9269 | w9270 ;
  assign w9272 = \pi082 ^ w9105 ;
  assign w9273 = ( ~w9113 & w9271 ) | ( ~w9113 & w9272 ) | ( w9271 & w9272 ) ;
  assign w9274 = w9272 | w9273 ;
  assign w9275 = \pi083 ^ w9098 ;
  assign w9276 = ( ~w9106 & w9274 ) | ( ~w9106 & w9275 ) | ( w9274 & w9275 ) ;
  assign w9277 = w9275 | w9276 ;
  assign w9278 = \pi084 ^ w9091 ;
  assign w9279 = ( ~w9099 & w9277 ) | ( ~w9099 & w9278 ) | ( w9277 & w9278 ) ;
  assign w9280 = w9278 | w9279 ;
  assign w9281 = \pi085 ^ w9084 ;
  assign w9282 = ( ~w9092 & w9280 ) | ( ~w9092 & w9281 ) | ( w9280 & w9281 ) ;
  assign w9283 = w9281 | w9282 ;
  assign w9284 = \pi086 ^ w9077 ;
  assign w9285 = ( ~w9085 & w9283 ) | ( ~w9085 & w9284 ) | ( w9283 & w9284 ) ;
  assign w9286 = w9284 | w9285 ;
  assign w9287 = \pi087 ^ w9070 ;
  assign w9288 = ( ~w9078 & w9286 ) | ( ~w9078 & w9287 ) | ( w9286 & w9287 ) ;
  assign w9289 = w9287 | w9288 ;
  assign w9290 = \pi088 ^ w9063 ;
  assign w9291 = ( ~w9071 & w9289 ) | ( ~w9071 & w9290 ) | ( w9289 & w9290 ) ;
  assign w9292 = w9290 | w9291 ;
  assign w9293 = \pi089 ^ w9056 ;
  assign w9294 = ( ~w9064 & w9292 ) | ( ~w9064 & w9293 ) | ( w9292 & w9293 ) ;
  assign w9295 = w9293 | w9294 ;
  assign w9296 = \pi090 ^ w9049 ;
  assign w9297 = ( ~w9057 & w9295 ) | ( ~w9057 & w9296 ) | ( w9295 & w9296 ) ;
  assign w9298 = w9296 | w9297 ;
  assign w9299 = \pi091 ^ w9042 ;
  assign w9300 = ( ~w9050 & w9298 ) | ( ~w9050 & w9299 ) | ( w9298 & w9299 ) ;
  assign w9301 = w9299 | w9300 ;
  assign w9302 = \pi092 ^ w9035 ;
  assign w9303 = ( ~w9043 & w9301 ) | ( ~w9043 & w9302 ) | ( w9301 & w9302 ) ;
  assign w9304 = w9302 | w9303 ;
  assign w9305 = \pi093 ^ w9028 ;
  assign w9306 = ( ~w9036 & w9304 ) | ( ~w9036 & w9305 ) | ( w9304 & w9305 ) ;
  assign w9307 = w9305 | w9306 ;
  assign w9308 = \pi094 ^ w9021 ;
  assign w9309 = ( ~w9029 & w9307 ) | ( ~w9029 & w9308 ) | ( w9307 & w9308 ) ;
  assign w9310 = w9308 | w9309 ;
  assign w9311 = \pi095 ^ w9014 ;
  assign w9312 = ( ~w9022 & w9310 ) | ( ~w9022 & w9311 ) | ( w9310 & w9311 ) ;
  assign w9313 = w9311 | w9312 ;
  assign w9314 = \pi096 ^ w9007 ;
  assign w9315 = ( ~w9015 & w9313 ) | ( ~w9015 & w9314 ) | ( w9313 & w9314 ) ;
  assign w9316 = w9314 | w9315 ;
  assign w9317 = \pi097 ^ w9000 ;
  assign w9318 = ( ~w9008 & w9316 ) | ( ~w9008 & w9317 ) | ( w9316 & w9317 ) ;
  assign w9319 = w9317 | w9318 ;
  assign w9320 = \pi098 ^ w8993 ;
  assign w9321 = ( ~w9001 & w9319 ) | ( ~w9001 & w9320 ) | ( w9319 & w9320 ) ;
  assign w9322 = w9320 | w9321 ;
  assign w9323 = \pi099 ^ w8986 ;
  assign w9324 = ( ~w8994 & w9322 ) | ( ~w8994 & w9323 ) | ( w9322 & w9323 ) ;
  assign w9325 = w9323 | w9324 ;
  assign w9326 = \pi100 ^ w8979 ;
  assign w9327 = ( ~w8987 & w9325 ) | ( ~w8987 & w9326 ) | ( w9325 & w9326 ) ;
  assign w9328 = w9326 | w9327 ;
  assign w9329 = \pi101 ^ w8972 ;
  assign w9330 = ( ~w8980 & w9328 ) | ( ~w8980 & w9329 ) | ( w9328 & w9329 ) ;
  assign w9331 = w9329 | w9330 ;
  assign w9332 = \pi102 ^ w8965 ;
  assign w9333 = ( ~w8973 & w9331 ) | ( ~w8973 & w9332 ) | ( w9331 & w9332 ) ;
  assign w9334 = w9332 | w9333 ;
  assign w9335 = \pi103 ^ w8958 ;
  assign w9336 = ( ~w8966 & w9334 ) | ( ~w8966 & w9335 ) | ( w9334 & w9335 ) ;
  assign w9337 = w9335 | w9336 ;
  assign w9338 = \pi104 ^ w8951 ;
  assign w9339 = ( ~w8959 & w9337 ) | ( ~w8959 & w9338 ) | ( w9337 & w9338 ) ;
  assign w9340 = w9338 | w9339 ;
  assign w9341 = \pi105 ^ w8937 ;
  assign w9342 = ( ~w8952 & w9340 ) | ( ~w8952 & w9341 ) | ( w9340 & w9341 ) ;
  assign w9343 = w9341 | w9342 ;
  assign w9344 = \pi106 ^ w8944 ;
  assign w9345 = w8945 & ~w9344 ;
  assign w9346 = ( w9343 & w9344 ) | ( w9343 & ~w9345 ) | ( w9344 & ~w9345 ) ;
  assign w9347 = ~\pi106 & w8944 ;
  assign w9348 = w9346 & ~w9347 ;
  assign w9349 = \pi108 | w284 ;
  assign w9350 = ( \pi107 & w275 ) | ( \pi107 & ~w284 ) | ( w275 & ~w284 ) ;
  assign w9351 = w9349 | w9350 ;
  assign w9352 = w9348 | w9351 ;
  assign w9353 = w8937 & w9352 ;
  assign w9354 = ~w8952 & w9340 ;
  assign w9355 = w9341 ^ w9354 ;
  assign w9356 = ~w9352 & w9355 ;
  assign w9357 = w9353 | w9356 ;
  assign w9358 = ~\pi106 & w9357 ;
  assign w9359 = w8951 & w9352 ;
  assign w9360 = ~w8959 & w9337 ;
  assign w9361 = w9338 ^ w9360 ;
  assign w9362 = ~w9352 & w9361 ;
  assign w9363 = w9359 | w9362 ;
  assign w9364 = ~\pi105 & w9363 ;
  assign w9365 = w8958 & w9352 ;
  assign w9366 = ~w8966 & w9334 ;
  assign w9367 = w9335 ^ w9366 ;
  assign w9368 = ~w9352 & w9367 ;
  assign w9369 = w9365 | w9368 ;
  assign w9370 = ~\pi104 & w9369 ;
  assign w9371 = w8965 & w9352 ;
  assign w9372 = ~w8973 & w9331 ;
  assign w9373 = w9332 ^ w9372 ;
  assign w9374 = ~w9352 & w9373 ;
  assign w9375 = w9371 | w9374 ;
  assign w9376 = ~\pi103 & w9375 ;
  assign w9377 = w8972 & w9352 ;
  assign w9378 = ~w8980 & w9328 ;
  assign w9379 = w9329 ^ w9378 ;
  assign w9380 = ~w9352 & w9379 ;
  assign w9381 = w9377 | w9380 ;
  assign w9382 = ~\pi102 & w9381 ;
  assign w9383 = w8979 & w9352 ;
  assign w9384 = ~w8987 & w9325 ;
  assign w9385 = w9326 ^ w9384 ;
  assign w9386 = ~w9352 & w9385 ;
  assign w9387 = w9383 | w9386 ;
  assign w9388 = ~\pi101 & w9387 ;
  assign w9389 = w8986 & w9352 ;
  assign w9390 = ~w8994 & w9322 ;
  assign w9391 = w9323 ^ w9390 ;
  assign w9392 = ~w9352 & w9391 ;
  assign w9393 = w9389 | w9392 ;
  assign w9394 = ~\pi100 & w9393 ;
  assign w9395 = w8993 & w9352 ;
  assign w9396 = ~w9001 & w9319 ;
  assign w9397 = w9320 ^ w9396 ;
  assign w9398 = ~w9352 & w9397 ;
  assign w9399 = w9395 | w9398 ;
  assign w9400 = ~\pi099 & w9399 ;
  assign w9401 = w9000 & w9352 ;
  assign w9402 = ~w9008 & w9316 ;
  assign w9403 = w9317 ^ w9402 ;
  assign w9404 = ~w9352 & w9403 ;
  assign w9405 = w9401 | w9404 ;
  assign w9406 = ~\pi098 & w9405 ;
  assign w9407 = w9007 & w9352 ;
  assign w9408 = ~w9015 & w9313 ;
  assign w9409 = w9314 ^ w9408 ;
  assign w9410 = ~w9352 & w9409 ;
  assign w9411 = w9407 | w9410 ;
  assign w9412 = ~\pi097 & w9411 ;
  assign w9413 = w9014 & w9352 ;
  assign w9414 = ~w9022 & w9310 ;
  assign w9415 = w9311 ^ w9414 ;
  assign w9416 = ~w9352 & w9415 ;
  assign w9417 = w9413 | w9416 ;
  assign w9418 = ~\pi096 & w9417 ;
  assign w9419 = w9021 & w9352 ;
  assign w9420 = ~w9029 & w9307 ;
  assign w9421 = w9308 ^ w9420 ;
  assign w9422 = ~w9352 & w9421 ;
  assign w9423 = w9419 | w9422 ;
  assign w9424 = ~\pi095 & w9423 ;
  assign w9425 = w9028 & w9352 ;
  assign w9426 = ~w9036 & w9304 ;
  assign w9427 = w9305 ^ w9426 ;
  assign w9428 = ~w9352 & w9427 ;
  assign w9429 = w9425 | w9428 ;
  assign w9430 = ~\pi094 & w9429 ;
  assign w9431 = w9035 & w9352 ;
  assign w9432 = ~w9043 & w9301 ;
  assign w9433 = w9302 ^ w9432 ;
  assign w9434 = ~w9352 & w9433 ;
  assign w9435 = w9431 | w9434 ;
  assign w9436 = ~\pi093 & w9435 ;
  assign w9437 = w9042 & w9352 ;
  assign w9438 = ~w9050 & w9298 ;
  assign w9439 = w9299 ^ w9438 ;
  assign w9440 = ~w9352 & w9439 ;
  assign w9441 = w9437 | w9440 ;
  assign w9442 = ~\pi092 & w9441 ;
  assign w9443 = w9049 & w9352 ;
  assign w9444 = ~w9057 & w9295 ;
  assign w9445 = w9296 ^ w9444 ;
  assign w9446 = ~w9352 & w9445 ;
  assign w9447 = w9443 | w9446 ;
  assign w9448 = ~\pi091 & w9447 ;
  assign w9449 = w9056 & w9352 ;
  assign w9450 = ~w9064 & w9292 ;
  assign w9451 = w9293 ^ w9450 ;
  assign w9452 = ~w9352 & w9451 ;
  assign w9453 = w9449 | w9452 ;
  assign w9454 = ~\pi090 & w9453 ;
  assign w9455 = w9063 & w9352 ;
  assign w9456 = ~w9071 & w9289 ;
  assign w9457 = w9290 ^ w9456 ;
  assign w9458 = ~w9352 & w9457 ;
  assign w9459 = w9455 | w9458 ;
  assign w9460 = ~\pi089 & w9459 ;
  assign w9461 = w9070 & w9352 ;
  assign w9462 = ~w9078 & w9286 ;
  assign w9463 = w9287 ^ w9462 ;
  assign w9464 = ~w9352 & w9463 ;
  assign w9465 = w9461 | w9464 ;
  assign w9466 = ~\pi088 & w9465 ;
  assign w9467 = w9077 & w9352 ;
  assign w9468 = ~w9085 & w9283 ;
  assign w9469 = w9284 ^ w9468 ;
  assign w9470 = ~w9352 & w9469 ;
  assign w9471 = w9467 | w9470 ;
  assign w9472 = ~\pi087 & w9471 ;
  assign w9473 = w9084 & w9352 ;
  assign w9474 = ~w9092 & w9280 ;
  assign w9475 = w9281 ^ w9474 ;
  assign w9476 = ~w9352 & w9475 ;
  assign w9477 = w9473 | w9476 ;
  assign w9478 = ~\pi086 & w9477 ;
  assign w9479 = w9091 & w9352 ;
  assign w9480 = ~w9099 & w9277 ;
  assign w9481 = w9278 ^ w9480 ;
  assign w9482 = ~w9352 & w9481 ;
  assign w9483 = w9479 | w9482 ;
  assign w9484 = ~\pi085 & w9483 ;
  assign w9485 = w9098 & w9352 ;
  assign w9486 = ~w9106 & w9274 ;
  assign w9487 = w9275 ^ w9486 ;
  assign w9488 = ~w9352 & w9487 ;
  assign w9489 = w9485 | w9488 ;
  assign w9490 = ~\pi084 & w9489 ;
  assign w9491 = w9105 & w9352 ;
  assign w9492 = ~w9113 & w9271 ;
  assign w9493 = w9272 ^ w9492 ;
  assign w9494 = ~w9352 & w9493 ;
  assign w9495 = w9491 | w9494 ;
  assign w9496 = ~\pi083 & w9495 ;
  assign w9497 = w9112 & w9352 ;
  assign w9498 = ~w9120 & w9268 ;
  assign w9499 = w9269 ^ w9498 ;
  assign w9500 = ~w9352 & w9499 ;
  assign w9501 = w9497 | w9500 ;
  assign w9502 = ~\pi082 & w9501 ;
  assign w9503 = w9119 & w9352 ;
  assign w9504 = ~w9127 & w9265 ;
  assign w9505 = w9266 ^ w9504 ;
  assign w9506 = ~w9352 & w9505 ;
  assign w9507 = w9503 | w9506 ;
  assign w9508 = ~\pi081 & w9507 ;
  assign w9509 = w9126 & w9352 ;
  assign w9510 = ~w9134 & w9262 ;
  assign w9511 = w9263 ^ w9510 ;
  assign w9512 = ~w9352 & w9511 ;
  assign w9513 = w9509 | w9512 ;
  assign w9514 = ~\pi080 & w9513 ;
  assign w9515 = w9133 & w9352 ;
  assign w9516 = ~w9141 & w9259 ;
  assign w9517 = w9260 ^ w9516 ;
  assign w9518 = ~w9352 & w9517 ;
  assign w9519 = w9515 | w9518 ;
  assign w9520 = ~\pi079 & w9519 ;
  assign w9521 = w9140 & w9352 ;
  assign w9522 = ~w9148 & w9256 ;
  assign w9523 = w9257 ^ w9522 ;
  assign w9524 = ~w9352 & w9523 ;
  assign w9525 = w9521 | w9524 ;
  assign w9526 = ~\pi078 & w9525 ;
  assign w9527 = w9147 & w9352 ;
  assign w9528 = ~w9155 & w9253 ;
  assign w9529 = w9254 ^ w9528 ;
  assign w9530 = ~w9352 & w9529 ;
  assign w9531 = w9527 | w9530 ;
  assign w9532 = ~\pi077 & w9531 ;
  assign w9533 = w9154 & w9352 ;
  assign w9534 = ~w9162 & w9250 ;
  assign w9535 = w9251 ^ w9534 ;
  assign w9536 = ~w9352 & w9535 ;
  assign w9537 = w9533 | w9536 ;
  assign w9538 = ~\pi076 & w9537 ;
  assign w9539 = w9161 & w9352 ;
  assign w9540 = ~w9169 & w9247 ;
  assign w9541 = w9248 ^ w9540 ;
  assign w9542 = ~w9352 & w9541 ;
  assign w9543 = w9539 | w9542 ;
  assign w9544 = ~\pi075 & w9543 ;
  assign w9545 = w9168 & w9352 ;
  assign w9546 = ~w9176 & w9244 ;
  assign w9547 = w9245 ^ w9546 ;
  assign w9548 = ~w9352 & w9547 ;
  assign w9549 = w9545 | w9548 ;
  assign w9550 = ~\pi074 & w9549 ;
  assign w9551 = w9175 & w9352 ;
  assign w9552 = ~w9183 & w9241 ;
  assign w9553 = w9242 ^ w9552 ;
  assign w9554 = ~w9352 & w9553 ;
  assign w9555 = w9551 | w9554 ;
  assign w9556 = ~\pi073 & w9555 ;
  assign w9557 = w9182 & w9352 ;
  assign w9558 = ~w9190 & w9238 ;
  assign w9559 = w9239 ^ w9558 ;
  assign w9560 = ~w9352 & w9559 ;
  assign w9561 = w9557 | w9560 ;
  assign w9562 = ~\pi072 & w9561 ;
  assign w9563 = w9189 & w9352 ;
  assign w9564 = ~w9197 & w9235 ;
  assign w9565 = w9236 ^ w9564 ;
  assign w9566 = ~w9352 & w9565 ;
  assign w9567 = w9563 | w9566 ;
  assign w9568 = ~\pi071 & w9567 ;
  assign w9569 = w9196 & w9352 ;
  assign w9570 = ~w9204 & w9232 ;
  assign w9571 = w9233 ^ w9570 ;
  assign w9572 = ~w9352 & w9571 ;
  assign w9573 = w9569 | w9572 ;
  assign w9574 = ~\pi070 & w9573 ;
  assign w9575 = w9203 & w9352 ;
  assign w9576 = ~w9212 & w9229 ;
  assign w9577 = w9230 ^ w9576 ;
  assign w9578 = ~w9352 & w9577 ;
  assign w9579 = w9575 | w9578 ;
  assign w9580 = ~\pi069 & w9579 ;
  assign w9581 = w9211 & w9352 ;
  assign w9582 = ~w9217 & w9226 ;
  assign w9583 = w9227 ^ w9582 ;
  assign w9584 = ~w9352 & w9583 ;
  assign w9585 = w9581 | w9584 ;
  assign w9586 = ~\pi068 & w9585 ;
  assign w9587 = w9216 & w9352 ;
  assign w9588 = ( \pi065 & w9218 ) | ( \pi065 & ~w9223 ) | ( w9218 & ~w9223 ) ;
  assign w9589 = w9221 ^ w9588 ;
  assign w9590 = ( w9348 & w9351 ) | ( w9348 & w9589 ) | ( w9351 & w9589 ) ;
  assign w9591 = w9589 & ~w9590 ;
  assign w9592 = w9587 | w9591 ;
  assign w9593 = ~\pi067 & w9592 ;
  assign w9594 = \pi022 ^ \pi065 ;
  assign w9595 = \pi021 ^ w8931 ;
  assign w9596 = ( \pi064 & w9351 ) | ( \pi064 & w9595 ) | ( w9351 & w9595 ) ;
  assign w9597 = w9594 ^ w9596 ;
  assign w9598 = ~w9351 & w9597 ;
  assign w9599 = ~w9348 & w9598 ;
  assign w9600 = ( ~\pi064 & w8931 ) | ( ~\pi064 & w9352 ) | ( w8931 & w9352 ) ;
  assign w9601 = \pi022 ^ w9600 ;
  assign w9602 = w9352 & ~w9601 ;
  assign w9603 = w9599 | w9602 ;
  assign w9604 = ~\pi066 & w9603 ;
  assign w9605 = ( \pi064 & w167 ) | ( \pi064 & w201 ) | ( w167 & w201 ) ;
  assign w9606 = \pi021 & \pi107 ;
  assign w9607 = ( \pi021 & w9605 ) | ( \pi021 & w9606 ) | ( w9605 & w9606 ) ;
  assign w9608 = ( \pi064 & w9348 ) | ( \pi064 & w9607 ) | ( w9348 & w9607 ) ;
  assign w9609 = ( \pi021 & ~\pi064 ) | ( \pi021 & w9608 ) | ( ~\pi064 & w9608 ) ;
  assign w9610 = ( \pi107 & ~w284 ) | ( \pi107 & w9218 ) | ( ~w284 & w9218 ) ;
  assign w9611 = w275 | w9348 ;
  assign w9612 = ( \pi107 & \pi108 ) | ( \pi107 & ~w275 ) | ( \pi108 & ~w275 ) ;
  assign w9613 = w9611 | w9612 ;
  assign w9614 = w9610 & ~w9613 ;
  assign w9615 = ~\pi020 & \pi064 ;
  assign w9616 = w9352 | w9599 ;
  assign w9617 = ( w9223 & w9599 ) | ( w9223 & w9616 ) | ( w9599 & w9616 ) ;
  assign w9618 = \pi066 ^ w9617 ;
  assign w9619 = w9609 | w9614 ;
  assign w9620 = ( \pi065 & w9615 ) | ( \pi065 & ~w9619 ) | ( w9615 & ~w9619 ) ;
  assign w9621 = w9618 | w9620 ;
  assign w9622 = \pi067 ^ w9592 ;
  assign w9623 = ( ~w9604 & w9621 ) | ( ~w9604 & w9622 ) | ( w9621 & w9622 ) ;
  assign w9624 = w9622 | w9623 ;
  assign w9625 = \pi068 ^ w9585 ;
  assign w9626 = ( ~w9593 & w9624 ) | ( ~w9593 & w9625 ) | ( w9624 & w9625 ) ;
  assign w9627 = w9625 | w9626 ;
  assign w9628 = \pi069 ^ w9579 ;
  assign w9629 = ( ~w9586 & w9627 ) | ( ~w9586 & w9628 ) | ( w9627 & w9628 ) ;
  assign w9630 = w9628 | w9629 ;
  assign w9631 = \pi070 ^ w9573 ;
  assign w9632 = ( ~w9580 & w9630 ) | ( ~w9580 & w9631 ) | ( w9630 & w9631 ) ;
  assign w9633 = w9631 | w9632 ;
  assign w9634 = \pi071 ^ w9567 ;
  assign w9635 = ( ~w9574 & w9633 ) | ( ~w9574 & w9634 ) | ( w9633 & w9634 ) ;
  assign w9636 = w9634 | w9635 ;
  assign w9637 = \pi072 ^ w9561 ;
  assign w9638 = ( ~w9568 & w9636 ) | ( ~w9568 & w9637 ) | ( w9636 & w9637 ) ;
  assign w9639 = w9637 | w9638 ;
  assign w9640 = \pi073 ^ w9555 ;
  assign w9641 = ( ~w9562 & w9639 ) | ( ~w9562 & w9640 ) | ( w9639 & w9640 ) ;
  assign w9642 = w9640 | w9641 ;
  assign w9643 = \pi074 ^ w9549 ;
  assign w9644 = ( ~w9556 & w9642 ) | ( ~w9556 & w9643 ) | ( w9642 & w9643 ) ;
  assign w9645 = w9643 | w9644 ;
  assign w9646 = \pi075 ^ w9543 ;
  assign w9647 = ( ~w9550 & w9645 ) | ( ~w9550 & w9646 ) | ( w9645 & w9646 ) ;
  assign w9648 = w9646 | w9647 ;
  assign w9649 = \pi076 ^ w9537 ;
  assign w9650 = ( ~w9544 & w9648 ) | ( ~w9544 & w9649 ) | ( w9648 & w9649 ) ;
  assign w9651 = w9649 | w9650 ;
  assign w9652 = \pi077 ^ w9531 ;
  assign w9653 = ( ~w9538 & w9651 ) | ( ~w9538 & w9652 ) | ( w9651 & w9652 ) ;
  assign w9654 = w9652 | w9653 ;
  assign w9655 = \pi078 ^ w9525 ;
  assign w9656 = ( ~w9532 & w9654 ) | ( ~w9532 & w9655 ) | ( w9654 & w9655 ) ;
  assign w9657 = w9655 | w9656 ;
  assign w9658 = \pi079 ^ w9519 ;
  assign w9659 = ( ~w9526 & w9657 ) | ( ~w9526 & w9658 ) | ( w9657 & w9658 ) ;
  assign w9660 = w9658 | w9659 ;
  assign w9661 = \pi080 ^ w9513 ;
  assign w9662 = ( ~w9520 & w9660 ) | ( ~w9520 & w9661 ) | ( w9660 & w9661 ) ;
  assign w9663 = w9661 | w9662 ;
  assign w9664 = \pi081 ^ w9507 ;
  assign w9665 = ( ~w9514 & w9663 ) | ( ~w9514 & w9664 ) | ( w9663 & w9664 ) ;
  assign w9666 = w9664 | w9665 ;
  assign w9667 = \pi082 ^ w9501 ;
  assign w9668 = ( ~w9508 & w9666 ) | ( ~w9508 & w9667 ) | ( w9666 & w9667 ) ;
  assign w9669 = w9667 | w9668 ;
  assign w9670 = \pi083 ^ w9495 ;
  assign w9671 = ( ~w9502 & w9669 ) | ( ~w9502 & w9670 ) | ( w9669 & w9670 ) ;
  assign w9672 = w9670 | w9671 ;
  assign w9673 = \pi084 ^ w9489 ;
  assign w9674 = ( ~w9496 & w9672 ) | ( ~w9496 & w9673 ) | ( w9672 & w9673 ) ;
  assign w9675 = w9673 | w9674 ;
  assign w9676 = \pi085 ^ w9483 ;
  assign w9677 = ( ~w9490 & w9675 ) | ( ~w9490 & w9676 ) | ( w9675 & w9676 ) ;
  assign w9678 = w9676 | w9677 ;
  assign w9679 = \pi086 ^ w9477 ;
  assign w9680 = ( ~w9484 & w9678 ) | ( ~w9484 & w9679 ) | ( w9678 & w9679 ) ;
  assign w9681 = w9679 | w9680 ;
  assign w9682 = \pi087 ^ w9471 ;
  assign w9683 = ( ~w9478 & w9681 ) | ( ~w9478 & w9682 ) | ( w9681 & w9682 ) ;
  assign w9684 = w9682 | w9683 ;
  assign w9685 = \pi088 ^ w9465 ;
  assign w9686 = ( ~w9472 & w9684 ) | ( ~w9472 & w9685 ) | ( w9684 & w9685 ) ;
  assign w9687 = w9685 | w9686 ;
  assign w9688 = \pi089 ^ w9459 ;
  assign w9689 = ( ~w9466 & w9687 ) | ( ~w9466 & w9688 ) | ( w9687 & w9688 ) ;
  assign w9690 = w9688 | w9689 ;
  assign w9691 = \pi090 ^ w9453 ;
  assign w9692 = ( ~w9460 & w9690 ) | ( ~w9460 & w9691 ) | ( w9690 & w9691 ) ;
  assign w9693 = w9691 | w9692 ;
  assign w9694 = \pi091 ^ w9447 ;
  assign w9695 = ( ~w9454 & w9693 ) | ( ~w9454 & w9694 ) | ( w9693 & w9694 ) ;
  assign w9696 = w9694 | w9695 ;
  assign w9697 = \pi092 ^ w9441 ;
  assign w9698 = ( ~w9448 & w9696 ) | ( ~w9448 & w9697 ) | ( w9696 & w9697 ) ;
  assign w9699 = w9697 | w9698 ;
  assign w9700 = \pi093 ^ w9435 ;
  assign w9701 = ( ~w9442 & w9699 ) | ( ~w9442 & w9700 ) | ( w9699 & w9700 ) ;
  assign w9702 = w9700 | w9701 ;
  assign w9703 = \pi094 ^ w9429 ;
  assign w9704 = ( ~w9436 & w9702 ) | ( ~w9436 & w9703 ) | ( w9702 & w9703 ) ;
  assign w9705 = w9703 | w9704 ;
  assign w9706 = \pi095 ^ w9423 ;
  assign w9707 = ( ~w9430 & w9705 ) | ( ~w9430 & w9706 ) | ( w9705 & w9706 ) ;
  assign w9708 = w9706 | w9707 ;
  assign w9709 = \pi096 ^ w9417 ;
  assign w9710 = ( ~w9424 & w9708 ) | ( ~w9424 & w9709 ) | ( w9708 & w9709 ) ;
  assign w9711 = w9709 | w9710 ;
  assign w9712 = \pi097 ^ w9411 ;
  assign w9713 = ( ~w9418 & w9711 ) | ( ~w9418 & w9712 ) | ( w9711 & w9712 ) ;
  assign w9714 = w9712 | w9713 ;
  assign w9715 = \pi098 ^ w9405 ;
  assign w9716 = ( ~w9412 & w9714 ) | ( ~w9412 & w9715 ) | ( w9714 & w9715 ) ;
  assign w9717 = w9715 | w9716 ;
  assign w9718 = \pi099 ^ w9399 ;
  assign w9719 = ( ~w9406 & w9717 ) | ( ~w9406 & w9718 ) | ( w9717 & w9718 ) ;
  assign w9720 = w9718 | w9719 ;
  assign w9721 = \pi100 ^ w9393 ;
  assign w9722 = ( ~w9400 & w9720 ) | ( ~w9400 & w9721 ) | ( w9720 & w9721 ) ;
  assign w9723 = w9721 | w9722 ;
  assign w9724 = \pi101 ^ w9387 ;
  assign w9725 = ( ~w9394 & w9723 ) | ( ~w9394 & w9724 ) | ( w9723 & w9724 ) ;
  assign w9726 = w9724 | w9725 ;
  assign w9727 = \pi102 ^ w9381 ;
  assign w9728 = ( ~w9388 & w9726 ) | ( ~w9388 & w9727 ) | ( w9726 & w9727 ) ;
  assign w9729 = w9727 | w9728 ;
  assign w9730 = \pi103 ^ w9375 ;
  assign w9731 = ( ~w9382 & w9729 ) | ( ~w9382 & w9730 ) | ( w9729 & w9730 ) ;
  assign w9732 = w9730 | w9731 ;
  assign w9733 = \pi104 ^ w9369 ;
  assign w9734 = ( ~w9376 & w9732 ) | ( ~w9376 & w9733 ) | ( w9732 & w9733 ) ;
  assign w9735 = w9733 | w9734 ;
  assign w9736 = \pi105 ^ w9363 ;
  assign w9737 = ( ~w9370 & w9735 ) | ( ~w9370 & w9736 ) | ( w9735 & w9736 ) ;
  assign w9738 = w9736 | w9737 ;
  assign w9739 = \pi106 ^ w9357 ;
  assign w9740 = ( ~w9364 & w9738 ) | ( ~w9364 & w9739 ) | ( w9738 & w9739 ) ;
  assign w9741 = w9739 | w9740 ;
  assign w9742 = w8944 & w9352 ;
  assign w9743 = ~w8945 & w9343 ;
  assign w9744 = w9344 ^ w9743 ;
  assign w9745 = ~w9352 & w9744 ;
  assign w9746 = w9742 | w9745 ;
  assign w9747 = ~\pi107 & w9746 ;
  assign w9748 = ( \pi107 & ~w9742 ) | ( \pi107 & w9745 ) | ( ~w9742 & w9745 ) ;
  assign w9749 = ~w9745 & w9748 ;
  assign w9750 = ( ~w9358 & w9741 ) | ( ~w9358 & w9747 ) | ( w9741 & w9747 ) ;
  assign w9751 = ( w168 & w9747 ) | ( w168 & ~w9750 ) | ( w9747 & ~w9750 ) ;
  assign w9752 = ( w155 & w9749 ) | ( w155 & ~w9750 ) | ( w9749 & ~w9750 ) ;
  assign w9753 = ( w9750 & ~w9751 ) | ( w9750 & w9752 ) | ( ~w9751 & w9752 ) ;
  assign w9754 = w9751 | w9753 ;
  assign w9755 = ~w9351 & w9746 ;
  assign w9756 = w9754 & ~w9755 ;
  assign w9757 = ~w9364 & w9738 ;
  assign w9758 = w9739 ^ w9757 ;
  assign w9759 = ~w9756 & w9758 ;
  assign w9760 = ( w9357 & w9754 ) | ( w9357 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9761 = ~w9755 & w9760 ;
  assign w9762 = w9759 | w9761 ;
  assign w9763 = ~\pi107 & w9762 ;
  assign w9764 = ~w9370 & w9735 ;
  assign w9765 = w9736 ^ w9764 ;
  assign w9766 = ~w9756 & w9765 ;
  assign w9767 = ( w9363 & w9754 ) | ( w9363 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9768 = ~w9755 & w9767 ;
  assign w9769 = w9766 | w9768 ;
  assign w9770 = ~\pi106 & w9769 ;
  assign w9771 = ~w9376 & w9732 ;
  assign w9772 = w9733 ^ w9771 ;
  assign w9773 = ~w9756 & w9772 ;
  assign w9774 = ( w9369 & w9754 ) | ( w9369 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9775 = ~w9755 & w9774 ;
  assign w9776 = w9773 | w9775 ;
  assign w9777 = ~\pi105 & w9776 ;
  assign w9778 = ~w9382 & w9729 ;
  assign w9779 = w9730 ^ w9778 ;
  assign w9780 = ~w9756 & w9779 ;
  assign w9781 = ( w9375 & w9754 ) | ( w9375 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9782 = ~w9755 & w9781 ;
  assign w9783 = w9780 | w9782 ;
  assign w9784 = ~\pi104 & w9783 ;
  assign w9785 = ~w9388 & w9726 ;
  assign w9786 = w9727 ^ w9785 ;
  assign w9787 = ~w9756 & w9786 ;
  assign w9788 = ( w9381 & w9754 ) | ( w9381 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9789 = ~w9755 & w9788 ;
  assign w9790 = w9787 | w9789 ;
  assign w9791 = ~\pi103 & w9790 ;
  assign w9792 = ~w9394 & w9723 ;
  assign w9793 = w9724 ^ w9792 ;
  assign w9794 = ~w9756 & w9793 ;
  assign w9795 = ( w9387 & w9754 ) | ( w9387 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9796 = ~w9755 & w9795 ;
  assign w9797 = w9794 | w9796 ;
  assign w9798 = ~\pi102 & w9797 ;
  assign w9799 = ~w9400 & w9720 ;
  assign w9800 = w9721 ^ w9799 ;
  assign w9801 = ~w9756 & w9800 ;
  assign w9802 = ( w9393 & w9754 ) | ( w9393 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9803 = ~w9755 & w9802 ;
  assign w9804 = w9801 | w9803 ;
  assign w9805 = ~\pi101 & w9804 ;
  assign w9806 = ~w9406 & w9717 ;
  assign w9807 = w9718 ^ w9806 ;
  assign w9808 = ~w9756 & w9807 ;
  assign w9809 = ( w9399 & w9754 ) | ( w9399 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9810 = ~w9755 & w9809 ;
  assign w9811 = w9808 | w9810 ;
  assign w9812 = ~\pi100 & w9811 ;
  assign w9813 = ~w9412 & w9714 ;
  assign w9814 = w9715 ^ w9813 ;
  assign w9815 = ~w9756 & w9814 ;
  assign w9816 = ( w9405 & w9754 ) | ( w9405 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9817 = ~w9755 & w9816 ;
  assign w9818 = w9815 | w9817 ;
  assign w9819 = ~\pi099 & w9818 ;
  assign w9820 = ~w9418 & w9711 ;
  assign w9821 = w9712 ^ w9820 ;
  assign w9822 = ~w9756 & w9821 ;
  assign w9823 = ( w9411 & w9754 ) | ( w9411 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9824 = ~w9755 & w9823 ;
  assign w9825 = w9822 | w9824 ;
  assign w9826 = ~\pi098 & w9825 ;
  assign w9827 = ~w9424 & w9708 ;
  assign w9828 = w9709 ^ w9827 ;
  assign w9829 = ~w9756 & w9828 ;
  assign w9830 = ( w9417 & w9754 ) | ( w9417 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9831 = ~w9755 & w9830 ;
  assign w9832 = w9829 | w9831 ;
  assign w9833 = ~\pi097 & w9832 ;
  assign w9834 = ~w9430 & w9705 ;
  assign w9835 = w9706 ^ w9834 ;
  assign w9836 = ~w9756 & w9835 ;
  assign w9837 = ( w9423 & w9754 ) | ( w9423 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9838 = ~w9755 & w9837 ;
  assign w9839 = w9836 | w9838 ;
  assign w9840 = ~\pi096 & w9839 ;
  assign w9841 = ~w9436 & w9702 ;
  assign w9842 = w9703 ^ w9841 ;
  assign w9843 = ~w9756 & w9842 ;
  assign w9844 = ( w9429 & w9754 ) | ( w9429 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9845 = ~w9755 & w9844 ;
  assign w9846 = w9843 | w9845 ;
  assign w9847 = ~\pi095 & w9846 ;
  assign w9848 = ~w9442 & w9699 ;
  assign w9849 = w9700 ^ w9848 ;
  assign w9850 = ~w9756 & w9849 ;
  assign w9851 = ( w9435 & w9754 ) | ( w9435 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9852 = ~w9755 & w9851 ;
  assign w9853 = w9850 | w9852 ;
  assign w9854 = ~\pi094 & w9853 ;
  assign w9855 = ~w9448 & w9696 ;
  assign w9856 = w9697 ^ w9855 ;
  assign w9857 = ~w9756 & w9856 ;
  assign w9858 = ( w9441 & w9754 ) | ( w9441 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9859 = ~w9755 & w9858 ;
  assign w9860 = w9857 | w9859 ;
  assign w9861 = ~\pi093 & w9860 ;
  assign w9862 = ~w9454 & w9693 ;
  assign w9863 = w9694 ^ w9862 ;
  assign w9864 = ~w9756 & w9863 ;
  assign w9865 = ( w9447 & w9754 ) | ( w9447 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9866 = ~w9755 & w9865 ;
  assign w9867 = w9864 | w9866 ;
  assign w9868 = ~\pi092 & w9867 ;
  assign w9869 = ~w9460 & w9690 ;
  assign w9870 = w9691 ^ w9869 ;
  assign w9871 = ~w9756 & w9870 ;
  assign w9872 = ( w9453 & w9754 ) | ( w9453 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9873 = ~w9755 & w9872 ;
  assign w9874 = w9871 | w9873 ;
  assign w9875 = ~\pi091 & w9874 ;
  assign w9876 = ~w9466 & w9687 ;
  assign w9877 = w9688 ^ w9876 ;
  assign w9878 = ~w9756 & w9877 ;
  assign w9879 = ( w9459 & w9754 ) | ( w9459 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9880 = ~w9755 & w9879 ;
  assign w9881 = w9878 | w9880 ;
  assign w9882 = ~\pi090 & w9881 ;
  assign w9883 = ~w9472 & w9684 ;
  assign w9884 = w9685 ^ w9883 ;
  assign w9885 = ~w9756 & w9884 ;
  assign w9886 = ( w9465 & w9754 ) | ( w9465 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9887 = ~w9755 & w9886 ;
  assign w9888 = w9885 | w9887 ;
  assign w9889 = ~\pi089 & w9888 ;
  assign w9890 = ~w9478 & w9681 ;
  assign w9891 = w9682 ^ w9890 ;
  assign w9892 = ~w9756 & w9891 ;
  assign w9893 = ( w9471 & w9754 ) | ( w9471 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9894 = ~w9755 & w9893 ;
  assign w9895 = w9892 | w9894 ;
  assign w9896 = ~\pi088 & w9895 ;
  assign w9897 = ~w9484 & w9678 ;
  assign w9898 = w9679 ^ w9897 ;
  assign w9899 = ~w9756 & w9898 ;
  assign w9900 = ( w9477 & w9754 ) | ( w9477 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9901 = ~w9755 & w9900 ;
  assign w9902 = w9899 | w9901 ;
  assign w9903 = ~\pi087 & w9902 ;
  assign w9904 = ~w9490 & w9675 ;
  assign w9905 = w9676 ^ w9904 ;
  assign w9906 = ~w9756 & w9905 ;
  assign w9907 = ( w9483 & w9754 ) | ( w9483 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9908 = ~w9755 & w9907 ;
  assign w9909 = w9906 | w9908 ;
  assign w9910 = ~\pi086 & w9909 ;
  assign w9911 = ~w9496 & w9672 ;
  assign w9912 = w9673 ^ w9911 ;
  assign w9913 = ~w9756 & w9912 ;
  assign w9914 = ( w9489 & w9754 ) | ( w9489 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9915 = ~w9755 & w9914 ;
  assign w9916 = w9913 | w9915 ;
  assign w9917 = ~\pi085 & w9916 ;
  assign w9918 = ~w9502 & w9669 ;
  assign w9919 = w9670 ^ w9918 ;
  assign w9920 = ~w9756 & w9919 ;
  assign w9921 = ( w9495 & w9754 ) | ( w9495 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9922 = ~w9755 & w9921 ;
  assign w9923 = w9920 | w9922 ;
  assign w9924 = ~\pi084 & w9923 ;
  assign w9925 = ~w9508 & w9666 ;
  assign w9926 = w9667 ^ w9925 ;
  assign w9927 = ~w9756 & w9926 ;
  assign w9928 = ( w9501 & w9754 ) | ( w9501 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9929 = ~w9755 & w9928 ;
  assign w9930 = w9927 | w9929 ;
  assign w9931 = ~\pi083 & w9930 ;
  assign w9932 = ~w9514 & w9663 ;
  assign w9933 = w9664 ^ w9932 ;
  assign w9934 = ~w9756 & w9933 ;
  assign w9935 = ( w9507 & w9754 ) | ( w9507 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9936 = ~w9755 & w9935 ;
  assign w9937 = w9934 | w9936 ;
  assign w9938 = ~\pi082 & w9937 ;
  assign w9939 = ~w9520 & w9660 ;
  assign w9940 = w9661 ^ w9939 ;
  assign w9941 = ~w9756 & w9940 ;
  assign w9942 = ( w9513 & w9754 ) | ( w9513 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9943 = ~w9755 & w9942 ;
  assign w9944 = w9941 | w9943 ;
  assign w9945 = ~\pi081 & w9944 ;
  assign w9946 = ~w9526 & w9657 ;
  assign w9947 = w9658 ^ w9946 ;
  assign w9948 = ~w9756 & w9947 ;
  assign w9949 = ( w9519 & w9754 ) | ( w9519 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9950 = ~w9755 & w9949 ;
  assign w9951 = w9948 | w9950 ;
  assign w9952 = ~\pi080 & w9951 ;
  assign w9953 = ~w9532 & w9654 ;
  assign w9954 = w9655 ^ w9953 ;
  assign w9955 = ~w9756 & w9954 ;
  assign w9956 = ( w9525 & w9754 ) | ( w9525 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9957 = ~w9755 & w9956 ;
  assign w9958 = w9955 | w9957 ;
  assign w9959 = ~\pi079 & w9958 ;
  assign w9960 = ~w9538 & w9651 ;
  assign w9961 = w9652 ^ w9960 ;
  assign w9962 = ~w9756 & w9961 ;
  assign w9963 = ( w9531 & w9754 ) | ( w9531 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9964 = ~w9755 & w9963 ;
  assign w9965 = w9962 | w9964 ;
  assign w9966 = ~\pi078 & w9965 ;
  assign w9967 = ~w9544 & w9648 ;
  assign w9968 = w9649 ^ w9967 ;
  assign w9969 = ~w9756 & w9968 ;
  assign w9970 = ( w9537 & w9754 ) | ( w9537 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9971 = ~w9755 & w9970 ;
  assign w9972 = w9969 | w9971 ;
  assign w9973 = ~\pi077 & w9972 ;
  assign w9974 = ~w9550 & w9645 ;
  assign w9975 = w9646 ^ w9974 ;
  assign w9976 = ~w9756 & w9975 ;
  assign w9977 = ( w9543 & w9754 ) | ( w9543 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9978 = ~w9755 & w9977 ;
  assign w9979 = w9976 | w9978 ;
  assign w9980 = ~\pi076 & w9979 ;
  assign w9981 = ~w9556 & w9642 ;
  assign w9982 = w9643 ^ w9981 ;
  assign w9983 = ~w9756 & w9982 ;
  assign w9984 = ( w9549 & w9754 ) | ( w9549 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9985 = ~w9755 & w9984 ;
  assign w9986 = w9983 | w9985 ;
  assign w9987 = ~\pi075 & w9986 ;
  assign w9988 = ~w9562 & w9639 ;
  assign w9989 = w9640 ^ w9988 ;
  assign w9990 = ~w9756 & w9989 ;
  assign w9991 = ( w9555 & w9754 ) | ( w9555 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9992 = ~w9755 & w9991 ;
  assign w9993 = w9990 | w9992 ;
  assign w9994 = ~\pi074 & w9993 ;
  assign w9995 = ~w9568 & w9636 ;
  assign w9996 = w9637 ^ w9995 ;
  assign w9997 = ~w9756 & w9996 ;
  assign w9998 = ( w9561 & w9754 ) | ( w9561 & w9755 ) | ( w9754 & w9755 ) ;
  assign w9999 = ~w9755 & w9998 ;
  assign w10000 = w9997 | w9999 ;
  assign w10001 = ~\pi073 & w10000 ;
  assign w10002 = ~w9574 & w9633 ;
  assign w10003 = w9634 ^ w10002 ;
  assign w10004 = ~w9756 & w10003 ;
  assign w10005 = ( w9567 & w9754 ) | ( w9567 & w9755 ) | ( w9754 & w9755 ) ;
  assign w10006 = ~w9755 & w10005 ;
  assign w10007 = w10004 | w10006 ;
  assign w10008 = ~\pi072 & w10007 ;
  assign w10009 = ~w9580 & w9630 ;
  assign w10010 = w9631 ^ w10009 ;
  assign w10011 = ~w9756 & w10010 ;
  assign w10012 = ( w9573 & w9754 ) | ( w9573 & w9755 ) | ( w9754 & w9755 ) ;
  assign w10013 = ~w9755 & w10012 ;
  assign w10014 = w10011 | w10013 ;
  assign w10015 = ~\pi071 & w10014 ;
  assign w10016 = ~w9586 & w9627 ;
  assign w10017 = w9628 ^ w10016 ;
  assign w10018 = ~w9756 & w10017 ;
  assign w10019 = ( w9579 & w9754 ) | ( w9579 & w9755 ) | ( w9754 & w9755 ) ;
  assign w10020 = ~w9755 & w10019 ;
  assign w10021 = w10018 | w10020 ;
  assign w10022 = ~\pi070 & w10021 ;
  assign w10023 = ~w9593 & w9624 ;
  assign w10024 = w9625 ^ w10023 ;
  assign w10025 = ~w9756 & w10024 ;
  assign w10026 = ( w9585 & w9754 ) | ( w9585 & w9755 ) | ( w9754 & w9755 ) ;
  assign w10027 = ~w9755 & w10026 ;
  assign w10028 = w10025 | w10027 ;
  assign w10029 = ~\pi069 & w10028 ;
  assign w10030 = ~w9604 & w9621 ;
  assign w10031 = w9622 ^ w10030 ;
  assign w10032 = ~w9756 & w10031 ;
  assign w10033 = ( w9592 & w9754 ) | ( w9592 & w9755 ) | ( w9754 & w9755 ) ;
  assign w10034 = ~w9755 & w10033 ;
  assign w10035 = w10032 | w10034 ;
  assign w10036 = ~\pi068 & w10035 ;
  assign w10037 = w9618 ^ w9620 ;
  assign w10038 = ~w9756 & w10037 ;
  assign w10039 = ( w9603 & w9754 ) | ( w9603 & w9755 ) | ( w9754 & w9755 ) ;
  assign w10040 = ~w9755 & w10039 ;
  assign w10041 = w10038 | w10040 ;
  assign w10042 = ~\pi067 & w10041 ;
  assign w10043 = w9615 ^ w9619 ;
  assign w10044 = \pi065 ^ w10043 ;
  assign w10045 = ~w9756 & w10044 ;
  assign w10046 = ( w9609 & w9614 ) | ( w9609 & ~w9755 ) | ( w9614 & ~w9755 ) ;
  assign w10047 = w9755 & w10046 ;
  assign w10048 = ( ~w9754 & w10046 ) | ( ~w9754 & w10047 ) | ( w10046 & w10047 ) ;
  assign w10049 = ( w10045 & w10046 ) | ( w10045 & ~w10048 ) | ( w10046 & ~w10048 ) ;
  assign w10050 = ~\pi066 & w10049 ;
  assign w10051 = w9754 | w9755 ;
  assign w10052 = ( w10045 & w10046 ) | ( w10045 & w10051 ) | ( w10046 & w10051 ) ;
  assign w10053 = ( ~w9755 & w10045 ) | ( ~w9755 & w10052 ) | ( w10045 & w10052 ) ;
  assign w10054 = \pi066 ^ w10053 ;
  assign w10055 = \pi064 & ~w9756 ;
  assign w10056 = \pi020 ^ w10055 ;
  assign w10057 = ( ~\pi019 & \pi064 ) | ( ~\pi019 & w10054 ) | ( \pi064 & w10054 ) ;
  assign w10058 = ( \pi065 & ~w10056 ) | ( \pi065 & w10057 ) | ( ~w10056 & w10057 ) ;
  assign w10059 = w10054 | w10058 ;
  assign w10060 = \pi067 ^ w10041 ;
  assign w10061 = ( ~w10050 & w10059 ) | ( ~w10050 & w10060 ) | ( w10059 & w10060 ) ;
  assign w10062 = w10060 | w10061 ;
  assign w10063 = \pi068 ^ w10035 ;
  assign w10064 = ( ~w10042 & w10062 ) | ( ~w10042 & w10063 ) | ( w10062 & w10063 ) ;
  assign w10065 = w10063 | w10064 ;
  assign w10066 = \pi069 ^ w10028 ;
  assign w10067 = ( ~w10036 & w10065 ) | ( ~w10036 & w10066 ) | ( w10065 & w10066 ) ;
  assign w10068 = w10066 | w10067 ;
  assign w10069 = \pi070 ^ w10021 ;
  assign w10070 = ( ~w10029 & w10068 ) | ( ~w10029 & w10069 ) | ( w10068 & w10069 ) ;
  assign w10071 = w10069 | w10070 ;
  assign w10072 = \pi071 ^ w10014 ;
  assign w10073 = ( ~w10022 & w10071 ) | ( ~w10022 & w10072 ) | ( w10071 & w10072 ) ;
  assign w10074 = w10072 | w10073 ;
  assign w10075 = \pi072 ^ w10007 ;
  assign w10076 = ( ~w10015 & w10074 ) | ( ~w10015 & w10075 ) | ( w10074 & w10075 ) ;
  assign w10077 = w10075 | w10076 ;
  assign w10078 = \pi073 ^ w10000 ;
  assign w10079 = ( ~w10008 & w10077 ) | ( ~w10008 & w10078 ) | ( w10077 & w10078 ) ;
  assign w10080 = w10078 | w10079 ;
  assign w10081 = \pi074 ^ w9993 ;
  assign w10082 = ( ~w10001 & w10080 ) | ( ~w10001 & w10081 ) | ( w10080 & w10081 ) ;
  assign w10083 = w10081 | w10082 ;
  assign w10084 = \pi075 ^ w9986 ;
  assign w10085 = ( ~w9994 & w10083 ) | ( ~w9994 & w10084 ) | ( w10083 & w10084 ) ;
  assign w10086 = w10084 | w10085 ;
  assign w10087 = \pi076 ^ w9979 ;
  assign w10088 = ( ~w9987 & w10086 ) | ( ~w9987 & w10087 ) | ( w10086 & w10087 ) ;
  assign w10089 = w10087 | w10088 ;
  assign w10090 = \pi077 ^ w9972 ;
  assign w10091 = ( ~w9980 & w10089 ) | ( ~w9980 & w10090 ) | ( w10089 & w10090 ) ;
  assign w10092 = w10090 | w10091 ;
  assign w10093 = \pi078 ^ w9965 ;
  assign w10094 = ( ~w9973 & w10092 ) | ( ~w9973 & w10093 ) | ( w10092 & w10093 ) ;
  assign w10095 = w10093 | w10094 ;
  assign w10096 = \pi079 ^ w9958 ;
  assign w10097 = ( ~w9966 & w10095 ) | ( ~w9966 & w10096 ) | ( w10095 & w10096 ) ;
  assign w10098 = w10096 | w10097 ;
  assign w10099 = \pi080 ^ w9951 ;
  assign w10100 = ( ~w9959 & w10098 ) | ( ~w9959 & w10099 ) | ( w10098 & w10099 ) ;
  assign w10101 = w10099 | w10100 ;
  assign w10102 = \pi081 ^ w9944 ;
  assign w10103 = ( ~w9952 & w10101 ) | ( ~w9952 & w10102 ) | ( w10101 & w10102 ) ;
  assign w10104 = w10102 | w10103 ;
  assign w10105 = \pi082 ^ w9937 ;
  assign w10106 = ( ~w9945 & w10104 ) | ( ~w9945 & w10105 ) | ( w10104 & w10105 ) ;
  assign w10107 = w10105 | w10106 ;
  assign w10108 = \pi083 ^ w9930 ;
  assign w10109 = ( ~w9938 & w10107 ) | ( ~w9938 & w10108 ) | ( w10107 & w10108 ) ;
  assign w10110 = w10108 | w10109 ;
  assign w10111 = \pi084 ^ w9923 ;
  assign w10112 = ( ~w9931 & w10110 ) | ( ~w9931 & w10111 ) | ( w10110 & w10111 ) ;
  assign w10113 = w10111 | w10112 ;
  assign w10114 = \pi085 ^ w9916 ;
  assign w10115 = ( ~w9924 & w10113 ) | ( ~w9924 & w10114 ) | ( w10113 & w10114 ) ;
  assign w10116 = w10114 | w10115 ;
  assign w10117 = \pi086 ^ w9909 ;
  assign w10118 = ( ~w9917 & w10116 ) | ( ~w9917 & w10117 ) | ( w10116 & w10117 ) ;
  assign w10119 = w10117 | w10118 ;
  assign w10120 = \pi087 ^ w9902 ;
  assign w10121 = ( ~w9910 & w10119 ) | ( ~w9910 & w10120 ) | ( w10119 & w10120 ) ;
  assign w10122 = w10120 | w10121 ;
  assign w10123 = \pi088 ^ w9895 ;
  assign w10124 = ( ~w9903 & w10122 ) | ( ~w9903 & w10123 ) | ( w10122 & w10123 ) ;
  assign w10125 = w10123 | w10124 ;
  assign w10126 = \pi089 ^ w9888 ;
  assign w10127 = ( ~w9896 & w10125 ) | ( ~w9896 & w10126 ) | ( w10125 & w10126 ) ;
  assign w10128 = w10126 | w10127 ;
  assign w10129 = \pi090 ^ w9881 ;
  assign w10130 = ( ~w9889 & w10128 ) | ( ~w9889 & w10129 ) | ( w10128 & w10129 ) ;
  assign w10131 = w10129 | w10130 ;
  assign w10132 = \pi091 ^ w9874 ;
  assign w10133 = ( ~w9882 & w10131 ) | ( ~w9882 & w10132 ) | ( w10131 & w10132 ) ;
  assign w10134 = w10132 | w10133 ;
  assign w10135 = \pi092 ^ w9867 ;
  assign w10136 = ( ~w9875 & w10134 ) | ( ~w9875 & w10135 ) | ( w10134 & w10135 ) ;
  assign w10137 = w10135 | w10136 ;
  assign w10138 = \pi093 ^ w9860 ;
  assign w10139 = ( ~w9868 & w10137 ) | ( ~w9868 & w10138 ) | ( w10137 & w10138 ) ;
  assign w10140 = w10138 | w10139 ;
  assign w10141 = \pi094 ^ w9853 ;
  assign w10142 = ( ~w9861 & w10140 ) | ( ~w9861 & w10141 ) | ( w10140 & w10141 ) ;
  assign w10143 = w10141 | w10142 ;
  assign w10144 = \pi095 ^ w9846 ;
  assign w10145 = ( ~w9854 & w10143 ) | ( ~w9854 & w10144 ) | ( w10143 & w10144 ) ;
  assign w10146 = w10144 | w10145 ;
  assign w10147 = \pi096 ^ w9839 ;
  assign w10148 = ( ~w9847 & w10146 ) | ( ~w9847 & w10147 ) | ( w10146 & w10147 ) ;
  assign w10149 = w10147 | w10148 ;
  assign w10150 = \pi097 ^ w9832 ;
  assign w10151 = ( ~w9840 & w10149 ) | ( ~w9840 & w10150 ) | ( w10149 & w10150 ) ;
  assign w10152 = w10150 | w10151 ;
  assign w10153 = \pi098 ^ w9825 ;
  assign w10154 = ( ~w9833 & w10152 ) | ( ~w9833 & w10153 ) | ( w10152 & w10153 ) ;
  assign w10155 = w10153 | w10154 ;
  assign w10156 = \pi099 ^ w9818 ;
  assign w10157 = ( ~w9826 & w10155 ) | ( ~w9826 & w10156 ) | ( w10155 & w10156 ) ;
  assign w10158 = w10156 | w10157 ;
  assign w10159 = \pi100 ^ w9811 ;
  assign w10160 = ( ~w9819 & w10158 ) | ( ~w9819 & w10159 ) | ( w10158 & w10159 ) ;
  assign w10161 = w10159 | w10160 ;
  assign w10162 = \pi101 ^ w9804 ;
  assign w10163 = ( ~w9812 & w10161 ) | ( ~w9812 & w10162 ) | ( w10161 & w10162 ) ;
  assign w10164 = w10162 | w10163 ;
  assign w10165 = \pi102 ^ w9797 ;
  assign w10166 = ( ~w9805 & w10164 ) | ( ~w9805 & w10165 ) | ( w10164 & w10165 ) ;
  assign w10167 = w10165 | w10166 ;
  assign w10168 = \pi103 ^ w9790 ;
  assign w10169 = ( ~w9798 & w10167 ) | ( ~w9798 & w10168 ) | ( w10167 & w10168 ) ;
  assign w10170 = w10168 | w10169 ;
  assign w10171 = \pi104 ^ w9783 ;
  assign w10172 = ( ~w9791 & w10170 ) | ( ~w9791 & w10171 ) | ( w10170 & w10171 ) ;
  assign w10173 = w10171 | w10172 ;
  assign w10174 = \pi105 ^ w9776 ;
  assign w10175 = ( ~w9784 & w10173 ) | ( ~w9784 & w10174 ) | ( w10173 & w10174 ) ;
  assign w10176 = w10174 | w10175 ;
  assign w10177 = \pi106 ^ w9769 ;
  assign w10178 = ( ~w9777 & w10176 ) | ( ~w9777 & w10177 ) | ( w10176 & w10177 ) ;
  assign w10179 = w10177 | w10178 ;
  assign w10180 = \pi107 ^ w9762 ;
  assign w10181 = ( ~w9770 & w10179 ) | ( ~w9770 & w10180 ) | ( w10179 & w10180 ) ;
  assign w10182 = w10180 | w10181 ;
  assign w10183 = w9747 | w9749 ;
  assign w10184 = ( ~w9358 & w9741 ) | ( ~w9358 & w9756 ) | ( w9741 & w9756 ) ;
  assign w10185 = w10183 ^ w10184 ;
  assign w10186 = ~w9756 & w10185 ;
  assign w10187 = ( w9351 & ~w9746 ) | ( w9351 & w9754 ) | ( ~w9746 & w9754 ) ;
  assign w10188 = w9746 & w10187 ;
  assign w10189 = w10186 | w10188 ;
  assign w10190 = ~\pi108 & w10189 ;
  assign w10191 = ( \pi108 & ~w10186 ) | ( \pi108 & w10188 ) | ( ~w10186 & w10188 ) ;
  assign w10192 = ~w10188 & w10191 ;
  assign w10193 = ( ~w9763 & w10182 ) | ( ~w9763 & w10190 ) | ( w10182 & w10190 ) ;
  assign w10194 = ( w449 & w10190 ) | ( w449 & ~w10193 ) | ( w10190 & ~w10193 ) ;
  assign w10195 = ( w448 & w10192 ) | ( w448 & ~w10193 ) | ( w10192 & ~w10193 ) ;
  assign w10196 = ( w10193 & ~w10194 ) | ( w10193 & w10195 ) | ( ~w10194 & w10195 ) ;
  assign w10197 = w10194 | w10196 ;
  assign w10198 = ( w155 & ~w168 ) | ( w155 & w10189 ) | ( ~w168 & w10189 ) ;
  assign w10199 = ~w155 & w10198 ;
  assign w10200 = w10197 & ~w10199 ;
  assign w10201 = ~w9770 & w10179 ;
  assign w10202 = w10180 ^ w10201 ;
  assign w10203 = ~w10200 & w10202 ;
  assign w10204 = ( w9762 & w10197 ) | ( w9762 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10205 = ~w10199 & w10204 ;
  assign w10206 = w10203 | w10205 ;
  assign w10207 = w10190 | w10192 ;
  assign w10208 = ( ~w9763 & w10182 ) | ( ~w9763 & w10200 ) | ( w10182 & w10200 ) ;
  assign w10209 = w10207 ^ w10208 ;
  assign w10210 = ~w10200 & w10209 ;
  assign w10211 = ( w10189 & w10197 ) | ( w10189 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10212 = ~w10199 & w10211 ;
  assign w10213 = w10210 | w10212 ;
  assign w10214 = ~\pi108 & w10206 ;
  assign w10215 = ~w9777 & w10176 ;
  assign w10216 = w10177 ^ w10215 ;
  assign w10217 = ~w10200 & w10216 ;
  assign w10218 = ( w9769 & w10197 ) | ( w9769 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10219 = ~w10199 & w10218 ;
  assign w10220 = w10217 | w10219 ;
  assign w10221 = ~\pi107 & w10220 ;
  assign w10222 = ~w9784 & w10173 ;
  assign w10223 = w10174 ^ w10222 ;
  assign w10224 = ~w10200 & w10223 ;
  assign w10225 = ( w9776 & w10197 ) | ( w9776 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10226 = ~w10199 & w10225 ;
  assign w10227 = w10224 | w10226 ;
  assign w10228 = ~\pi106 & w10227 ;
  assign w10229 = ~w9791 & w10170 ;
  assign w10230 = w10171 ^ w10229 ;
  assign w10231 = ~w10200 & w10230 ;
  assign w10232 = ( w9783 & w10197 ) | ( w9783 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10233 = ~w10199 & w10232 ;
  assign w10234 = w10231 | w10233 ;
  assign w10235 = ~\pi105 & w10234 ;
  assign w10236 = ~w9798 & w10167 ;
  assign w10237 = w10168 ^ w10236 ;
  assign w10238 = ~w10200 & w10237 ;
  assign w10239 = ( w9790 & w10197 ) | ( w9790 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10240 = ~w10199 & w10239 ;
  assign w10241 = w10238 | w10240 ;
  assign w10242 = ~\pi104 & w10241 ;
  assign w10243 = ~w9805 & w10164 ;
  assign w10244 = w10165 ^ w10243 ;
  assign w10245 = ~w10200 & w10244 ;
  assign w10246 = ( w9797 & w10197 ) | ( w9797 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10247 = ~w10199 & w10246 ;
  assign w10248 = w10245 | w10247 ;
  assign w10249 = ~\pi103 & w10248 ;
  assign w10250 = ~w9812 & w10161 ;
  assign w10251 = w10162 ^ w10250 ;
  assign w10252 = ~w10200 & w10251 ;
  assign w10253 = ( w9804 & w10197 ) | ( w9804 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10254 = ~w10199 & w10253 ;
  assign w10255 = w10252 | w10254 ;
  assign w10256 = ~\pi102 & w10255 ;
  assign w10257 = ~w9819 & w10158 ;
  assign w10258 = w10159 ^ w10257 ;
  assign w10259 = ~w10200 & w10258 ;
  assign w10260 = ( w9811 & w10197 ) | ( w9811 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10261 = ~w10199 & w10260 ;
  assign w10262 = w10259 | w10261 ;
  assign w10263 = ~\pi101 & w10262 ;
  assign w10264 = ~w9826 & w10155 ;
  assign w10265 = w10156 ^ w10264 ;
  assign w10266 = ~w10200 & w10265 ;
  assign w10267 = ( w9818 & w10197 ) | ( w9818 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10268 = ~w10199 & w10267 ;
  assign w10269 = w10266 | w10268 ;
  assign w10270 = ~\pi100 & w10269 ;
  assign w10271 = ~w9833 & w10152 ;
  assign w10272 = w10153 ^ w10271 ;
  assign w10273 = ~w10200 & w10272 ;
  assign w10274 = ( w9825 & w10197 ) | ( w9825 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10275 = ~w10199 & w10274 ;
  assign w10276 = w10273 | w10275 ;
  assign w10277 = ~\pi099 & w10276 ;
  assign w10278 = ~w9840 & w10149 ;
  assign w10279 = w10150 ^ w10278 ;
  assign w10280 = ~w10200 & w10279 ;
  assign w10281 = ( w9832 & w10197 ) | ( w9832 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10282 = ~w10199 & w10281 ;
  assign w10283 = w10280 | w10282 ;
  assign w10284 = ~\pi098 & w10283 ;
  assign w10285 = ~w9847 & w10146 ;
  assign w10286 = w10147 ^ w10285 ;
  assign w10287 = ~w10200 & w10286 ;
  assign w10288 = ( w9839 & w10197 ) | ( w9839 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10289 = ~w10199 & w10288 ;
  assign w10290 = w10287 | w10289 ;
  assign w10291 = ~\pi097 & w10290 ;
  assign w10292 = ~w9854 & w10143 ;
  assign w10293 = w10144 ^ w10292 ;
  assign w10294 = ~w10200 & w10293 ;
  assign w10295 = ( w9846 & w10197 ) | ( w9846 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10296 = ~w10199 & w10295 ;
  assign w10297 = w10294 | w10296 ;
  assign w10298 = ~\pi096 & w10297 ;
  assign w10299 = ~w9861 & w10140 ;
  assign w10300 = w10141 ^ w10299 ;
  assign w10301 = ~w10200 & w10300 ;
  assign w10302 = ( w9853 & w10197 ) | ( w9853 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10303 = ~w10199 & w10302 ;
  assign w10304 = w10301 | w10303 ;
  assign w10305 = ~\pi095 & w10304 ;
  assign w10306 = ~w9868 & w10137 ;
  assign w10307 = w10138 ^ w10306 ;
  assign w10308 = ~w10200 & w10307 ;
  assign w10309 = ( w9860 & w10197 ) | ( w9860 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10310 = ~w10199 & w10309 ;
  assign w10311 = w10308 | w10310 ;
  assign w10312 = ~\pi094 & w10311 ;
  assign w10313 = ~w9875 & w10134 ;
  assign w10314 = w10135 ^ w10313 ;
  assign w10315 = ~w10200 & w10314 ;
  assign w10316 = ( w9867 & w10197 ) | ( w9867 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10317 = ~w10199 & w10316 ;
  assign w10318 = w10315 | w10317 ;
  assign w10319 = ~\pi093 & w10318 ;
  assign w10320 = ~w9882 & w10131 ;
  assign w10321 = w10132 ^ w10320 ;
  assign w10322 = ~w10200 & w10321 ;
  assign w10323 = ( w9874 & w10197 ) | ( w9874 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10324 = ~w10199 & w10323 ;
  assign w10325 = w10322 | w10324 ;
  assign w10326 = ~\pi092 & w10325 ;
  assign w10327 = ~w9889 & w10128 ;
  assign w10328 = w10129 ^ w10327 ;
  assign w10329 = ~w10200 & w10328 ;
  assign w10330 = ( w9881 & w10197 ) | ( w9881 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10331 = ~w10199 & w10330 ;
  assign w10332 = w10329 | w10331 ;
  assign w10333 = ~\pi091 & w10332 ;
  assign w10334 = ~w9896 & w10125 ;
  assign w10335 = w10126 ^ w10334 ;
  assign w10336 = ~w10200 & w10335 ;
  assign w10337 = ( w9888 & w10197 ) | ( w9888 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10338 = ~w10199 & w10337 ;
  assign w10339 = w10336 | w10338 ;
  assign w10340 = ~\pi090 & w10339 ;
  assign w10341 = ~w9903 & w10122 ;
  assign w10342 = w10123 ^ w10341 ;
  assign w10343 = ~w10200 & w10342 ;
  assign w10344 = ( w9895 & w10197 ) | ( w9895 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10345 = ~w10199 & w10344 ;
  assign w10346 = w10343 | w10345 ;
  assign w10347 = ~\pi089 & w10346 ;
  assign w10348 = ~w9910 & w10119 ;
  assign w10349 = w10120 ^ w10348 ;
  assign w10350 = ~w10200 & w10349 ;
  assign w10351 = ( w9902 & w10197 ) | ( w9902 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10352 = ~w10199 & w10351 ;
  assign w10353 = w10350 | w10352 ;
  assign w10354 = ~\pi088 & w10353 ;
  assign w10355 = ~w9917 & w10116 ;
  assign w10356 = w10117 ^ w10355 ;
  assign w10357 = ~w10200 & w10356 ;
  assign w10358 = ( w9909 & w10197 ) | ( w9909 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10359 = ~w10199 & w10358 ;
  assign w10360 = w10357 | w10359 ;
  assign w10361 = ~\pi087 & w10360 ;
  assign w10362 = ~w9924 & w10113 ;
  assign w10363 = w10114 ^ w10362 ;
  assign w10364 = ~w10200 & w10363 ;
  assign w10365 = ( w9916 & w10197 ) | ( w9916 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10366 = ~w10199 & w10365 ;
  assign w10367 = w10364 | w10366 ;
  assign w10368 = ~\pi086 & w10367 ;
  assign w10369 = ~w9931 & w10110 ;
  assign w10370 = w10111 ^ w10369 ;
  assign w10371 = ~w10200 & w10370 ;
  assign w10372 = ( w9923 & w10197 ) | ( w9923 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10373 = ~w10199 & w10372 ;
  assign w10374 = w10371 | w10373 ;
  assign w10375 = ~\pi085 & w10374 ;
  assign w10376 = ~w9938 & w10107 ;
  assign w10377 = w10108 ^ w10376 ;
  assign w10378 = ~w10200 & w10377 ;
  assign w10379 = ( w9930 & w10197 ) | ( w9930 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10380 = ~w10199 & w10379 ;
  assign w10381 = w10378 | w10380 ;
  assign w10382 = ~\pi084 & w10381 ;
  assign w10383 = ~w9945 & w10104 ;
  assign w10384 = w10105 ^ w10383 ;
  assign w10385 = ~w10200 & w10384 ;
  assign w10386 = ( w9937 & w10197 ) | ( w9937 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10387 = ~w10199 & w10386 ;
  assign w10388 = w10385 | w10387 ;
  assign w10389 = ~\pi083 & w10388 ;
  assign w10390 = ~w9952 & w10101 ;
  assign w10391 = w10102 ^ w10390 ;
  assign w10392 = ~w10200 & w10391 ;
  assign w10393 = ( w9944 & w10197 ) | ( w9944 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10394 = ~w10199 & w10393 ;
  assign w10395 = w10392 | w10394 ;
  assign w10396 = ~\pi082 & w10395 ;
  assign w10397 = ~w9959 & w10098 ;
  assign w10398 = w10099 ^ w10397 ;
  assign w10399 = ~w10200 & w10398 ;
  assign w10400 = ( w9951 & w10197 ) | ( w9951 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10401 = ~w10199 & w10400 ;
  assign w10402 = w10399 | w10401 ;
  assign w10403 = ~\pi081 & w10402 ;
  assign w10404 = ~w9966 & w10095 ;
  assign w10405 = w10096 ^ w10404 ;
  assign w10406 = ~w10200 & w10405 ;
  assign w10407 = ( w9958 & w10197 ) | ( w9958 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10408 = ~w10199 & w10407 ;
  assign w10409 = w10406 | w10408 ;
  assign w10410 = ~\pi080 & w10409 ;
  assign w10411 = ~w9973 & w10092 ;
  assign w10412 = w10093 ^ w10411 ;
  assign w10413 = ~w10200 & w10412 ;
  assign w10414 = ( w9965 & w10197 ) | ( w9965 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10415 = ~w10199 & w10414 ;
  assign w10416 = w10413 | w10415 ;
  assign w10417 = ~\pi079 & w10416 ;
  assign w10418 = ~w9980 & w10089 ;
  assign w10419 = w10090 ^ w10418 ;
  assign w10420 = ~w10200 & w10419 ;
  assign w10421 = ( w9972 & w10197 ) | ( w9972 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10422 = ~w10199 & w10421 ;
  assign w10423 = w10420 | w10422 ;
  assign w10424 = ~\pi078 & w10423 ;
  assign w10425 = ~w9987 & w10086 ;
  assign w10426 = w10087 ^ w10425 ;
  assign w10427 = ~w10200 & w10426 ;
  assign w10428 = ( w9979 & w10197 ) | ( w9979 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10429 = ~w10199 & w10428 ;
  assign w10430 = w10427 | w10429 ;
  assign w10431 = ~\pi077 & w10430 ;
  assign w10432 = ~w9994 & w10083 ;
  assign w10433 = w10084 ^ w10432 ;
  assign w10434 = ~w10200 & w10433 ;
  assign w10435 = ( w9986 & w10197 ) | ( w9986 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10436 = ~w10199 & w10435 ;
  assign w10437 = w10434 | w10436 ;
  assign w10438 = ~\pi076 & w10437 ;
  assign w10439 = ~w10001 & w10080 ;
  assign w10440 = w10081 ^ w10439 ;
  assign w10441 = ~w10200 & w10440 ;
  assign w10442 = ( w9993 & w10197 ) | ( w9993 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10443 = ~w10199 & w10442 ;
  assign w10444 = w10441 | w10443 ;
  assign w10445 = ~\pi075 & w10444 ;
  assign w10446 = ~w10008 & w10077 ;
  assign w10447 = w10078 ^ w10446 ;
  assign w10448 = ~w10200 & w10447 ;
  assign w10449 = ( w10000 & w10197 ) | ( w10000 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10450 = ~w10199 & w10449 ;
  assign w10451 = w10448 | w10450 ;
  assign w10452 = ~\pi074 & w10451 ;
  assign w10453 = ~w10015 & w10074 ;
  assign w10454 = w10075 ^ w10453 ;
  assign w10455 = ~w10200 & w10454 ;
  assign w10456 = ( w10007 & w10197 ) | ( w10007 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10457 = ~w10199 & w10456 ;
  assign w10458 = w10455 | w10457 ;
  assign w10459 = ~\pi073 & w10458 ;
  assign w10460 = ~w10022 & w10071 ;
  assign w10461 = w10072 ^ w10460 ;
  assign w10462 = ~w10200 & w10461 ;
  assign w10463 = ( w10014 & w10197 ) | ( w10014 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10464 = ~w10199 & w10463 ;
  assign w10465 = w10462 | w10464 ;
  assign w10466 = ~\pi072 & w10465 ;
  assign w10467 = ~w10029 & w10068 ;
  assign w10468 = w10069 ^ w10467 ;
  assign w10469 = ~w10200 & w10468 ;
  assign w10470 = ( w10021 & w10197 ) | ( w10021 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10471 = ~w10199 & w10470 ;
  assign w10472 = w10469 | w10471 ;
  assign w10473 = ~\pi071 & w10472 ;
  assign w10474 = ~w10036 & w10065 ;
  assign w10475 = w10066 ^ w10474 ;
  assign w10476 = ~w10200 & w10475 ;
  assign w10477 = ( w10028 & w10197 ) | ( w10028 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10478 = ~w10199 & w10477 ;
  assign w10479 = w10476 | w10478 ;
  assign w10480 = ~\pi070 & w10479 ;
  assign w10481 = ~w10042 & w10062 ;
  assign w10482 = w10063 ^ w10481 ;
  assign w10483 = ~w10200 & w10482 ;
  assign w10484 = ( w10035 & w10197 ) | ( w10035 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10485 = ~w10199 & w10484 ;
  assign w10486 = w10483 | w10485 ;
  assign w10487 = ~\pi069 & w10486 ;
  assign w10488 = ~w10050 & w10059 ;
  assign w10489 = w10060 ^ w10488 ;
  assign w10490 = ~w10200 & w10489 ;
  assign w10491 = ( w10041 & w10197 ) | ( w10041 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10492 = ~w10199 & w10491 ;
  assign w10493 = w10490 | w10492 ;
  assign w10494 = ~\pi068 & w10493 ;
  assign w10495 = ~\pi019 & \pi064 ;
  assign w10496 = ( \pi065 & ~w10056 ) | ( \pi065 & w10495 ) | ( ~w10056 & w10495 ) ;
  assign w10497 = w10054 ^ w10496 ;
  assign w10498 = ~w10200 & w10497 ;
  assign w10499 = ( w10049 & w10197 ) | ( w10049 & w10199 ) | ( w10197 & w10199 ) ;
  assign w10500 = ~w10199 & w10499 ;
  assign w10501 = w10498 | w10500 ;
  assign w10502 = ~\pi067 & w10501 ;
  assign w10503 = \pi020 ^ \pi065 ;
  assign w10504 = \pi019 ^ w9756 ;
  assign w10505 = ( \pi064 & w10200 ) | ( \pi064 & w10504 ) | ( w10200 & w10504 ) ;
  assign w10506 = w10503 ^ w10505 ;
  assign w10507 = ~w10200 & w10506 ;
  assign w10508 = w10056 & w10200 ;
  assign w10509 = w10507 | w10508 ;
  assign w10510 = ~\pi066 & w10509 ;
  assign w10511 = \pi066 ^ w10509 ;
  assign w10512 = \pi064 & ~w10200 ;
  assign w10513 = \pi019 ^ w10512 ;
  assign w10514 = ( ~\pi018 & \pi064 ) | ( ~\pi018 & w10511 ) | ( \pi064 & w10511 ) ;
  assign w10515 = ( \pi065 & ~w10513 ) | ( \pi065 & w10514 ) | ( ~w10513 & w10514 ) ;
  assign w10516 = w10511 | w10515 ;
  assign w10517 = \pi067 ^ w10501 ;
  assign w10518 = ( ~w10510 & w10516 ) | ( ~w10510 & w10517 ) | ( w10516 & w10517 ) ;
  assign w10519 = w10517 | w10518 ;
  assign w10520 = \pi068 ^ w10493 ;
  assign w10521 = ( ~w10502 & w10519 ) | ( ~w10502 & w10520 ) | ( w10519 & w10520 ) ;
  assign w10522 = w10520 | w10521 ;
  assign w10523 = \pi069 ^ w10486 ;
  assign w10524 = ( ~w10494 & w10522 ) | ( ~w10494 & w10523 ) | ( w10522 & w10523 ) ;
  assign w10525 = w10523 | w10524 ;
  assign w10526 = \pi070 ^ w10479 ;
  assign w10527 = ( ~w10487 & w10525 ) | ( ~w10487 & w10526 ) | ( w10525 & w10526 ) ;
  assign w10528 = w10526 | w10527 ;
  assign w10529 = \pi071 ^ w10472 ;
  assign w10530 = ( ~w10480 & w10528 ) | ( ~w10480 & w10529 ) | ( w10528 & w10529 ) ;
  assign w10531 = w10529 | w10530 ;
  assign w10532 = \pi072 ^ w10465 ;
  assign w10533 = ( ~w10473 & w10531 ) | ( ~w10473 & w10532 ) | ( w10531 & w10532 ) ;
  assign w10534 = w10532 | w10533 ;
  assign w10535 = \pi073 ^ w10458 ;
  assign w10536 = ( ~w10466 & w10534 ) | ( ~w10466 & w10535 ) | ( w10534 & w10535 ) ;
  assign w10537 = w10535 | w10536 ;
  assign w10538 = \pi074 ^ w10451 ;
  assign w10539 = ( ~w10459 & w10537 ) | ( ~w10459 & w10538 ) | ( w10537 & w10538 ) ;
  assign w10540 = w10538 | w10539 ;
  assign w10541 = \pi075 ^ w10444 ;
  assign w10542 = ( ~w10452 & w10540 ) | ( ~w10452 & w10541 ) | ( w10540 & w10541 ) ;
  assign w10543 = w10541 | w10542 ;
  assign w10544 = \pi076 ^ w10437 ;
  assign w10545 = ( ~w10445 & w10543 ) | ( ~w10445 & w10544 ) | ( w10543 & w10544 ) ;
  assign w10546 = w10544 | w10545 ;
  assign w10547 = \pi077 ^ w10430 ;
  assign w10548 = ( ~w10438 & w10546 ) | ( ~w10438 & w10547 ) | ( w10546 & w10547 ) ;
  assign w10549 = w10547 | w10548 ;
  assign w10550 = \pi078 ^ w10423 ;
  assign w10551 = ( ~w10431 & w10549 ) | ( ~w10431 & w10550 ) | ( w10549 & w10550 ) ;
  assign w10552 = w10550 | w10551 ;
  assign w10553 = \pi079 ^ w10416 ;
  assign w10554 = ( ~w10424 & w10552 ) | ( ~w10424 & w10553 ) | ( w10552 & w10553 ) ;
  assign w10555 = w10553 | w10554 ;
  assign w10556 = \pi080 ^ w10409 ;
  assign w10557 = ( ~w10417 & w10555 ) | ( ~w10417 & w10556 ) | ( w10555 & w10556 ) ;
  assign w10558 = w10556 | w10557 ;
  assign w10559 = \pi081 ^ w10402 ;
  assign w10560 = ( ~w10410 & w10558 ) | ( ~w10410 & w10559 ) | ( w10558 & w10559 ) ;
  assign w10561 = w10559 | w10560 ;
  assign w10562 = \pi082 ^ w10395 ;
  assign w10563 = ( ~w10403 & w10561 ) | ( ~w10403 & w10562 ) | ( w10561 & w10562 ) ;
  assign w10564 = w10562 | w10563 ;
  assign w10565 = \pi083 ^ w10388 ;
  assign w10566 = ( ~w10396 & w10564 ) | ( ~w10396 & w10565 ) | ( w10564 & w10565 ) ;
  assign w10567 = w10565 | w10566 ;
  assign w10568 = \pi084 ^ w10381 ;
  assign w10569 = ( ~w10389 & w10567 ) | ( ~w10389 & w10568 ) | ( w10567 & w10568 ) ;
  assign w10570 = w10568 | w10569 ;
  assign w10571 = \pi085 ^ w10374 ;
  assign w10572 = ( ~w10382 & w10570 ) | ( ~w10382 & w10571 ) | ( w10570 & w10571 ) ;
  assign w10573 = w10571 | w10572 ;
  assign w10574 = \pi086 ^ w10367 ;
  assign w10575 = ( ~w10375 & w10573 ) | ( ~w10375 & w10574 ) | ( w10573 & w10574 ) ;
  assign w10576 = w10574 | w10575 ;
  assign w10577 = \pi087 ^ w10360 ;
  assign w10578 = ( ~w10368 & w10576 ) | ( ~w10368 & w10577 ) | ( w10576 & w10577 ) ;
  assign w10579 = w10577 | w10578 ;
  assign w10580 = \pi088 ^ w10353 ;
  assign w10581 = ( ~w10361 & w10579 ) | ( ~w10361 & w10580 ) | ( w10579 & w10580 ) ;
  assign w10582 = w10580 | w10581 ;
  assign w10583 = \pi089 ^ w10346 ;
  assign w10584 = ( ~w10354 & w10582 ) | ( ~w10354 & w10583 ) | ( w10582 & w10583 ) ;
  assign w10585 = w10583 | w10584 ;
  assign w10586 = \pi090 ^ w10339 ;
  assign w10587 = ( ~w10347 & w10585 ) | ( ~w10347 & w10586 ) | ( w10585 & w10586 ) ;
  assign w10588 = w10586 | w10587 ;
  assign w10589 = \pi091 ^ w10332 ;
  assign w10590 = ( ~w10340 & w10588 ) | ( ~w10340 & w10589 ) | ( w10588 & w10589 ) ;
  assign w10591 = w10589 | w10590 ;
  assign w10592 = \pi092 ^ w10325 ;
  assign w10593 = ( ~w10333 & w10591 ) | ( ~w10333 & w10592 ) | ( w10591 & w10592 ) ;
  assign w10594 = w10592 | w10593 ;
  assign w10595 = \pi093 ^ w10318 ;
  assign w10596 = ( ~w10326 & w10594 ) | ( ~w10326 & w10595 ) | ( w10594 & w10595 ) ;
  assign w10597 = w10595 | w10596 ;
  assign w10598 = \pi094 ^ w10311 ;
  assign w10599 = ( ~w10319 & w10597 ) | ( ~w10319 & w10598 ) | ( w10597 & w10598 ) ;
  assign w10600 = w10598 | w10599 ;
  assign w10601 = \pi095 ^ w10304 ;
  assign w10602 = ( ~w10312 & w10600 ) | ( ~w10312 & w10601 ) | ( w10600 & w10601 ) ;
  assign w10603 = w10601 | w10602 ;
  assign w10604 = \pi096 ^ w10297 ;
  assign w10605 = ( ~w10305 & w10603 ) | ( ~w10305 & w10604 ) | ( w10603 & w10604 ) ;
  assign w10606 = w10604 | w10605 ;
  assign w10607 = \pi097 ^ w10290 ;
  assign w10608 = ( ~w10298 & w10606 ) | ( ~w10298 & w10607 ) | ( w10606 & w10607 ) ;
  assign w10609 = w10607 | w10608 ;
  assign w10610 = \pi098 ^ w10283 ;
  assign w10611 = ( ~w10291 & w10609 ) | ( ~w10291 & w10610 ) | ( w10609 & w10610 ) ;
  assign w10612 = w10610 | w10611 ;
  assign w10613 = \pi099 ^ w10276 ;
  assign w10614 = ( ~w10284 & w10612 ) | ( ~w10284 & w10613 ) | ( w10612 & w10613 ) ;
  assign w10615 = w10613 | w10614 ;
  assign w10616 = \pi100 ^ w10269 ;
  assign w10617 = ( ~w10277 & w10615 ) | ( ~w10277 & w10616 ) | ( w10615 & w10616 ) ;
  assign w10618 = w10616 | w10617 ;
  assign w10619 = \pi101 ^ w10262 ;
  assign w10620 = ( ~w10270 & w10618 ) | ( ~w10270 & w10619 ) | ( w10618 & w10619 ) ;
  assign w10621 = w10619 | w10620 ;
  assign w10622 = \pi102 ^ w10255 ;
  assign w10623 = ( ~w10263 & w10621 ) | ( ~w10263 & w10622 ) | ( w10621 & w10622 ) ;
  assign w10624 = w10622 | w10623 ;
  assign w10625 = \pi103 ^ w10248 ;
  assign w10626 = ( ~w10256 & w10624 ) | ( ~w10256 & w10625 ) | ( w10624 & w10625 ) ;
  assign w10627 = w10625 | w10626 ;
  assign w10628 = \pi104 ^ w10241 ;
  assign w10629 = ( ~w10249 & w10627 ) | ( ~w10249 & w10628 ) | ( w10627 & w10628 ) ;
  assign w10630 = w10628 | w10629 ;
  assign w10631 = \pi105 ^ w10234 ;
  assign w10632 = ( ~w10242 & w10630 ) | ( ~w10242 & w10631 ) | ( w10630 & w10631 ) ;
  assign w10633 = w10631 | w10632 ;
  assign w10634 = \pi106 ^ w10227 ;
  assign w10635 = ( ~w10235 & w10633 ) | ( ~w10235 & w10634 ) | ( w10633 & w10634 ) ;
  assign w10636 = w10634 | w10635 ;
  assign w10637 = \pi107 ^ w10220 ;
  assign w10638 = ( ~w10228 & w10636 ) | ( ~w10228 & w10637 ) | ( w10636 & w10637 ) ;
  assign w10639 = w10637 | w10638 ;
  assign w10640 = \pi108 ^ w10206 ;
  assign w10641 = ( ~w10221 & w10639 ) | ( ~w10221 & w10640 ) | ( w10639 & w10640 ) ;
  assign w10642 = w10640 | w10641 ;
  assign w10643 = \pi109 ^ w10213 ;
  assign w10644 = w10214 & ~w10643 ;
  assign w10645 = ( w10642 & w10643 ) | ( w10642 & ~w10644 ) | ( w10643 & ~w10644 ) ;
  assign w10646 = ~\pi109 & w10213 ;
  assign w10647 = w10645 & ~w10646 ;
  assign w10648 = \pi111 | w164 ;
  assign w10649 = ( \pi110 & w155 ) | ( \pi110 & ~w164 ) | ( w155 & ~w164 ) ;
  assign w10650 = w10648 | w10649 ;
  assign w10651 = w10647 | w10650 ;
  assign w10652 = w10206 & w10651 ;
  assign w10653 = ~w10221 & w10639 ;
  assign w10654 = w10640 ^ w10653 ;
  assign w10655 = ~w10651 & w10654 ;
  assign w10656 = w10652 | w10655 ;
  assign w10657 = ~\pi109 & w10656 ;
  assign w10658 = w10220 & w10651 ;
  assign w10659 = ~w10228 & w10636 ;
  assign w10660 = w10637 ^ w10659 ;
  assign w10661 = ~w10651 & w10660 ;
  assign w10662 = w10658 | w10661 ;
  assign w10663 = ~\pi108 & w10662 ;
  assign w10664 = w10227 & w10651 ;
  assign w10665 = ~w10235 & w10633 ;
  assign w10666 = w10634 ^ w10665 ;
  assign w10667 = ~w10651 & w10666 ;
  assign w10668 = w10664 | w10667 ;
  assign w10669 = ~\pi107 & w10668 ;
  assign w10670 = w10234 & w10651 ;
  assign w10671 = ~w10242 & w10630 ;
  assign w10672 = w10631 ^ w10671 ;
  assign w10673 = ~w10651 & w10672 ;
  assign w10674 = w10670 | w10673 ;
  assign w10675 = ~\pi106 & w10674 ;
  assign w10676 = w10241 & w10651 ;
  assign w10677 = ~w10249 & w10627 ;
  assign w10678 = w10628 ^ w10677 ;
  assign w10679 = ~w10651 & w10678 ;
  assign w10680 = w10676 | w10679 ;
  assign w10681 = ~\pi105 & w10680 ;
  assign w10682 = w10248 & w10651 ;
  assign w10683 = ~w10256 & w10624 ;
  assign w10684 = w10625 ^ w10683 ;
  assign w10685 = ~w10651 & w10684 ;
  assign w10686 = w10682 | w10685 ;
  assign w10687 = ~\pi104 & w10686 ;
  assign w10688 = w10255 & w10651 ;
  assign w10689 = ~w10263 & w10621 ;
  assign w10690 = w10622 ^ w10689 ;
  assign w10691 = ~w10651 & w10690 ;
  assign w10692 = w10688 | w10691 ;
  assign w10693 = ~\pi103 & w10692 ;
  assign w10694 = w10262 & w10651 ;
  assign w10695 = ~w10270 & w10618 ;
  assign w10696 = w10619 ^ w10695 ;
  assign w10697 = ~w10651 & w10696 ;
  assign w10698 = w10694 | w10697 ;
  assign w10699 = ~\pi102 & w10698 ;
  assign w10700 = w10269 & w10651 ;
  assign w10701 = ~w10277 & w10615 ;
  assign w10702 = w10616 ^ w10701 ;
  assign w10703 = ~w10651 & w10702 ;
  assign w10704 = w10700 | w10703 ;
  assign w10705 = ~\pi101 & w10704 ;
  assign w10706 = w10276 & w10651 ;
  assign w10707 = ~w10284 & w10612 ;
  assign w10708 = w10613 ^ w10707 ;
  assign w10709 = ~w10651 & w10708 ;
  assign w10710 = w10706 | w10709 ;
  assign w10711 = ~\pi100 & w10710 ;
  assign w10712 = w10283 & w10651 ;
  assign w10713 = ~w10291 & w10609 ;
  assign w10714 = w10610 ^ w10713 ;
  assign w10715 = ~w10651 & w10714 ;
  assign w10716 = w10712 | w10715 ;
  assign w10717 = ~\pi099 & w10716 ;
  assign w10718 = w10290 & w10651 ;
  assign w10719 = ~w10298 & w10606 ;
  assign w10720 = w10607 ^ w10719 ;
  assign w10721 = ~w10651 & w10720 ;
  assign w10722 = w10718 | w10721 ;
  assign w10723 = ~\pi098 & w10722 ;
  assign w10724 = w10297 & w10651 ;
  assign w10725 = ~w10305 & w10603 ;
  assign w10726 = w10604 ^ w10725 ;
  assign w10727 = ~w10651 & w10726 ;
  assign w10728 = w10724 | w10727 ;
  assign w10729 = ~\pi097 & w10728 ;
  assign w10730 = w10304 & w10651 ;
  assign w10731 = ~w10312 & w10600 ;
  assign w10732 = w10601 ^ w10731 ;
  assign w10733 = ~w10651 & w10732 ;
  assign w10734 = w10730 | w10733 ;
  assign w10735 = ~\pi096 & w10734 ;
  assign w10736 = w10311 & w10651 ;
  assign w10737 = ~w10319 & w10597 ;
  assign w10738 = w10598 ^ w10737 ;
  assign w10739 = ~w10651 & w10738 ;
  assign w10740 = w10736 | w10739 ;
  assign w10741 = ~\pi095 & w10740 ;
  assign w10742 = w10318 & w10651 ;
  assign w10743 = ~w10326 & w10594 ;
  assign w10744 = w10595 ^ w10743 ;
  assign w10745 = ~w10651 & w10744 ;
  assign w10746 = w10742 | w10745 ;
  assign w10747 = ~\pi094 & w10746 ;
  assign w10748 = w10325 & w10651 ;
  assign w10749 = ~w10333 & w10591 ;
  assign w10750 = w10592 ^ w10749 ;
  assign w10751 = ~w10651 & w10750 ;
  assign w10752 = w10748 | w10751 ;
  assign w10753 = ~\pi093 & w10752 ;
  assign w10754 = w10332 & w10651 ;
  assign w10755 = ~w10340 & w10588 ;
  assign w10756 = w10589 ^ w10755 ;
  assign w10757 = ~w10651 & w10756 ;
  assign w10758 = w10754 | w10757 ;
  assign w10759 = ~\pi092 & w10758 ;
  assign w10760 = w10339 & w10651 ;
  assign w10761 = ~w10347 & w10585 ;
  assign w10762 = w10586 ^ w10761 ;
  assign w10763 = ~w10651 & w10762 ;
  assign w10764 = w10760 | w10763 ;
  assign w10765 = ~\pi091 & w10764 ;
  assign w10766 = w10346 & w10651 ;
  assign w10767 = ~w10354 & w10582 ;
  assign w10768 = w10583 ^ w10767 ;
  assign w10769 = ~w10651 & w10768 ;
  assign w10770 = w10766 | w10769 ;
  assign w10771 = ~\pi090 & w10770 ;
  assign w10772 = w10353 & w10651 ;
  assign w10773 = ~w10361 & w10579 ;
  assign w10774 = w10580 ^ w10773 ;
  assign w10775 = ~w10651 & w10774 ;
  assign w10776 = w10772 | w10775 ;
  assign w10777 = ~\pi089 & w10776 ;
  assign w10778 = w10360 & w10651 ;
  assign w10779 = ~w10368 & w10576 ;
  assign w10780 = w10577 ^ w10779 ;
  assign w10781 = ~w10651 & w10780 ;
  assign w10782 = w10778 | w10781 ;
  assign w10783 = ~\pi088 & w10782 ;
  assign w10784 = w10367 & w10651 ;
  assign w10785 = ~w10375 & w10573 ;
  assign w10786 = w10574 ^ w10785 ;
  assign w10787 = ~w10651 & w10786 ;
  assign w10788 = w10784 | w10787 ;
  assign w10789 = ~\pi087 & w10788 ;
  assign w10790 = w10374 & w10651 ;
  assign w10791 = ~w10382 & w10570 ;
  assign w10792 = w10571 ^ w10791 ;
  assign w10793 = ~w10651 & w10792 ;
  assign w10794 = w10790 | w10793 ;
  assign w10795 = ~\pi086 & w10794 ;
  assign w10796 = w10381 & w10651 ;
  assign w10797 = ~w10389 & w10567 ;
  assign w10798 = w10568 ^ w10797 ;
  assign w10799 = ~w10651 & w10798 ;
  assign w10800 = w10796 | w10799 ;
  assign w10801 = ~\pi085 & w10800 ;
  assign w10802 = w10388 & w10651 ;
  assign w10803 = ~w10396 & w10564 ;
  assign w10804 = w10565 ^ w10803 ;
  assign w10805 = ~w10651 & w10804 ;
  assign w10806 = w10802 | w10805 ;
  assign w10807 = ~\pi084 & w10806 ;
  assign w10808 = w10395 & w10651 ;
  assign w10809 = ~w10403 & w10561 ;
  assign w10810 = w10562 ^ w10809 ;
  assign w10811 = ~w10651 & w10810 ;
  assign w10812 = w10808 | w10811 ;
  assign w10813 = ~\pi083 & w10812 ;
  assign w10814 = w10402 & w10651 ;
  assign w10815 = ~w10410 & w10558 ;
  assign w10816 = w10559 ^ w10815 ;
  assign w10817 = ~w10651 & w10816 ;
  assign w10818 = w10814 | w10817 ;
  assign w10819 = ~\pi082 & w10818 ;
  assign w10820 = w10409 & w10651 ;
  assign w10821 = ~w10417 & w10555 ;
  assign w10822 = w10556 ^ w10821 ;
  assign w10823 = ~w10651 & w10822 ;
  assign w10824 = w10820 | w10823 ;
  assign w10825 = ~\pi081 & w10824 ;
  assign w10826 = w10416 & w10651 ;
  assign w10827 = ~w10424 & w10552 ;
  assign w10828 = w10553 ^ w10827 ;
  assign w10829 = ~w10651 & w10828 ;
  assign w10830 = w10826 | w10829 ;
  assign w10831 = ~\pi080 & w10830 ;
  assign w10832 = w10423 & w10651 ;
  assign w10833 = ~w10431 & w10549 ;
  assign w10834 = w10550 ^ w10833 ;
  assign w10835 = ~w10651 & w10834 ;
  assign w10836 = w10832 | w10835 ;
  assign w10837 = ~\pi079 & w10836 ;
  assign w10838 = w10430 & w10651 ;
  assign w10839 = ~w10438 & w10546 ;
  assign w10840 = w10547 ^ w10839 ;
  assign w10841 = ~w10651 & w10840 ;
  assign w10842 = w10838 | w10841 ;
  assign w10843 = ~\pi078 & w10842 ;
  assign w10844 = w10437 & w10651 ;
  assign w10845 = ~w10445 & w10543 ;
  assign w10846 = w10544 ^ w10845 ;
  assign w10847 = ~w10651 & w10846 ;
  assign w10848 = w10844 | w10847 ;
  assign w10849 = ~\pi077 & w10848 ;
  assign w10850 = w10444 & w10651 ;
  assign w10851 = ~w10452 & w10540 ;
  assign w10852 = w10541 ^ w10851 ;
  assign w10853 = ~w10651 & w10852 ;
  assign w10854 = w10850 | w10853 ;
  assign w10855 = ~\pi076 & w10854 ;
  assign w10856 = w10451 & w10651 ;
  assign w10857 = ~w10459 & w10537 ;
  assign w10858 = w10538 ^ w10857 ;
  assign w10859 = ~w10651 & w10858 ;
  assign w10860 = w10856 | w10859 ;
  assign w10861 = ~\pi075 & w10860 ;
  assign w10862 = w10458 & w10651 ;
  assign w10863 = ~w10466 & w10534 ;
  assign w10864 = w10535 ^ w10863 ;
  assign w10865 = ~w10651 & w10864 ;
  assign w10866 = w10862 | w10865 ;
  assign w10867 = ~\pi074 & w10866 ;
  assign w10868 = w10465 & w10651 ;
  assign w10869 = ~w10473 & w10531 ;
  assign w10870 = w10532 ^ w10869 ;
  assign w10871 = ~w10651 & w10870 ;
  assign w10872 = w10868 | w10871 ;
  assign w10873 = ~\pi073 & w10872 ;
  assign w10874 = w10472 & w10651 ;
  assign w10875 = ~w10480 & w10528 ;
  assign w10876 = w10529 ^ w10875 ;
  assign w10877 = ~w10651 & w10876 ;
  assign w10878 = w10874 | w10877 ;
  assign w10879 = ~\pi072 & w10878 ;
  assign w10880 = w10479 & w10651 ;
  assign w10881 = ~w10487 & w10525 ;
  assign w10882 = w10526 ^ w10881 ;
  assign w10883 = ~w10651 & w10882 ;
  assign w10884 = w10880 | w10883 ;
  assign w10885 = ~\pi071 & w10884 ;
  assign w10886 = w10486 & w10651 ;
  assign w10887 = ~w10494 & w10522 ;
  assign w10888 = w10523 ^ w10887 ;
  assign w10889 = ~w10651 & w10888 ;
  assign w10890 = w10886 | w10889 ;
  assign w10891 = ~\pi070 & w10890 ;
  assign w10892 = w10493 & w10651 ;
  assign w10893 = ~w10502 & w10519 ;
  assign w10894 = w10520 ^ w10893 ;
  assign w10895 = ~w10651 & w10894 ;
  assign w10896 = w10892 | w10895 ;
  assign w10897 = ~\pi069 & w10896 ;
  assign w10898 = w10501 & w10651 ;
  assign w10899 = ~w10510 & w10516 ;
  assign w10900 = w10517 ^ w10899 ;
  assign w10901 = ~w10651 & w10900 ;
  assign w10902 = w10898 | w10901 ;
  assign w10903 = ~\pi068 & w10902 ;
  assign w10904 = ~\pi018 & \pi064 ;
  assign w10905 = ( \pi065 & ~w10513 ) | ( \pi065 & w10904 ) | ( ~w10513 & w10904 ) ;
  assign w10906 = w10511 ^ w10905 ;
  assign w10907 = ( w10647 & w10650 ) | ( w10647 & w10906 ) | ( w10650 & w10906 ) ;
  assign w10908 = w10906 & ~w10907 ;
  assign w10909 = ( w10509 & w10651 ) | ( w10509 & w10908 ) | ( w10651 & w10908 ) ;
  assign w10910 = w10908 | w10909 ;
  assign w10911 = ~\pi067 & w10910 ;
  assign w10912 = \pi019 ^ \pi065 ;
  assign w10913 = \pi018 ^ w10200 ;
  assign w10914 = ( \pi064 & w10650 ) | ( \pi064 & w10913 ) | ( w10650 & w10913 ) ;
  assign w10915 = w10912 ^ w10914 ;
  assign w10916 = ~w10650 & w10915 ;
  assign w10917 = ~w10647 & w10916 ;
  assign w10918 = ( ~\pi064 & w10200 ) | ( ~\pi064 & w10651 ) | ( w10200 & w10651 ) ;
  assign w10919 = \pi019 ^ w10918 ;
  assign w10920 = w10651 & ~w10919 ;
  assign w10921 = w10917 | w10920 ;
  assign w10922 = ~\pi066 & w10921 ;
  assign w10923 = ( \pi064 & ~\pi110 ) | ( \pi064 & \pi111 ) | ( ~\pi110 & \pi111 ) ;
  assign w10924 = w267 | w448 ;
  assign w10925 = ( \pi111 & \pi112 ) | ( \pi111 & ~w267 ) | ( \pi112 & ~w267 ) ;
  assign w10926 = w10924 | w10925 ;
  assign w10927 = w10923 & ~w10926 ;
  assign w10928 = ( \pi018 & w10647 ) | ( \pi018 & ~w10927 ) | ( w10647 & ~w10927 ) ;
  assign w10929 = \pi018 & w10928 ;
  assign w10930 = ( ~\pi018 & \pi064 ) | ( ~\pi018 & \pi110 ) | ( \pi064 & \pi110 ) ;
  assign w10931 = w155 | w164 ;
  assign w10932 = ( \pi110 & \pi111 ) | ( \pi110 & ~w164 ) | ( \pi111 & ~w164 ) ;
  assign w10933 = w10931 | w10932 ;
  assign w10934 = w10930 & ~w10933 ;
  assign w10935 = ~w10647 & w10934 ;
  assign w10936 = w10929 | w10935 ;
  assign w10937 = ~\pi017 & \pi064 ;
  assign w10938 = \pi065 ^ w10936 ;
  assign w10939 = w10937 | w10938 ;
  assign w10940 = w10651 | w10917 ;
  assign w10941 = ( w10513 & w10917 ) | ( w10513 & w10940 ) | ( w10917 & w10940 ) ;
  assign w10942 = \pi066 ^ w10941 ;
  assign w10943 = ~\pi065 & w10936 ;
  assign w10944 = w10939 | w10943 ;
  assign w10945 = ( w10942 & ~w10943 ) | ( w10942 & w10944 ) | ( ~w10943 & w10944 ) ;
  assign w10946 = ~w10509 & w10651 ;
  assign w10947 = ( w10651 & w10908 ) | ( w10651 & ~w10946 ) | ( w10908 & ~w10946 ) ;
  assign w10948 = \pi067 ^ w10947 ;
  assign w10949 = ( ~w10922 & w10945 ) | ( ~w10922 & w10948 ) | ( w10945 & w10948 ) ;
  assign w10950 = w10948 | w10949 ;
  assign w10951 = \pi068 ^ w10902 ;
  assign w10952 = ( ~w10911 & w10950 ) | ( ~w10911 & w10951 ) | ( w10950 & w10951 ) ;
  assign w10953 = w10951 | w10952 ;
  assign w10954 = \pi069 ^ w10896 ;
  assign w10955 = ( ~w10903 & w10953 ) | ( ~w10903 & w10954 ) | ( w10953 & w10954 ) ;
  assign w10956 = w10954 | w10955 ;
  assign w10957 = \pi070 ^ w10890 ;
  assign w10958 = ( ~w10897 & w10956 ) | ( ~w10897 & w10957 ) | ( w10956 & w10957 ) ;
  assign w10959 = w10957 | w10958 ;
  assign w10960 = \pi071 ^ w10884 ;
  assign w10961 = ( ~w10891 & w10959 ) | ( ~w10891 & w10960 ) | ( w10959 & w10960 ) ;
  assign w10962 = w10960 | w10961 ;
  assign w10963 = \pi072 ^ w10878 ;
  assign w10964 = ( ~w10885 & w10962 ) | ( ~w10885 & w10963 ) | ( w10962 & w10963 ) ;
  assign w10965 = w10963 | w10964 ;
  assign w10966 = \pi073 ^ w10872 ;
  assign w10967 = ( ~w10879 & w10965 ) | ( ~w10879 & w10966 ) | ( w10965 & w10966 ) ;
  assign w10968 = w10966 | w10967 ;
  assign w10969 = \pi074 ^ w10866 ;
  assign w10970 = ( ~w10873 & w10968 ) | ( ~w10873 & w10969 ) | ( w10968 & w10969 ) ;
  assign w10971 = w10969 | w10970 ;
  assign w10972 = \pi075 ^ w10860 ;
  assign w10973 = ( ~w10867 & w10971 ) | ( ~w10867 & w10972 ) | ( w10971 & w10972 ) ;
  assign w10974 = w10972 | w10973 ;
  assign w10975 = \pi076 ^ w10854 ;
  assign w10976 = ( ~w10861 & w10974 ) | ( ~w10861 & w10975 ) | ( w10974 & w10975 ) ;
  assign w10977 = w10975 | w10976 ;
  assign w10978 = \pi077 ^ w10848 ;
  assign w10979 = ( ~w10855 & w10977 ) | ( ~w10855 & w10978 ) | ( w10977 & w10978 ) ;
  assign w10980 = w10978 | w10979 ;
  assign w10981 = \pi078 ^ w10842 ;
  assign w10982 = ( ~w10849 & w10980 ) | ( ~w10849 & w10981 ) | ( w10980 & w10981 ) ;
  assign w10983 = w10981 | w10982 ;
  assign w10984 = \pi079 ^ w10836 ;
  assign w10985 = ( ~w10843 & w10983 ) | ( ~w10843 & w10984 ) | ( w10983 & w10984 ) ;
  assign w10986 = w10984 | w10985 ;
  assign w10987 = \pi080 ^ w10830 ;
  assign w10988 = ( ~w10837 & w10986 ) | ( ~w10837 & w10987 ) | ( w10986 & w10987 ) ;
  assign w10989 = w10987 | w10988 ;
  assign w10990 = \pi081 ^ w10824 ;
  assign w10991 = ( ~w10831 & w10989 ) | ( ~w10831 & w10990 ) | ( w10989 & w10990 ) ;
  assign w10992 = w10990 | w10991 ;
  assign w10993 = \pi082 ^ w10818 ;
  assign w10994 = ( ~w10825 & w10992 ) | ( ~w10825 & w10993 ) | ( w10992 & w10993 ) ;
  assign w10995 = w10993 | w10994 ;
  assign w10996 = \pi083 ^ w10812 ;
  assign w10997 = ( ~w10819 & w10995 ) | ( ~w10819 & w10996 ) | ( w10995 & w10996 ) ;
  assign w10998 = w10996 | w10997 ;
  assign w10999 = \pi084 ^ w10806 ;
  assign w11000 = ( ~w10813 & w10998 ) | ( ~w10813 & w10999 ) | ( w10998 & w10999 ) ;
  assign w11001 = w10999 | w11000 ;
  assign w11002 = \pi085 ^ w10800 ;
  assign w11003 = ( ~w10807 & w11001 ) | ( ~w10807 & w11002 ) | ( w11001 & w11002 ) ;
  assign w11004 = w11002 | w11003 ;
  assign w11005 = \pi086 ^ w10794 ;
  assign w11006 = ( ~w10801 & w11004 ) | ( ~w10801 & w11005 ) | ( w11004 & w11005 ) ;
  assign w11007 = w11005 | w11006 ;
  assign w11008 = \pi087 ^ w10788 ;
  assign w11009 = ( ~w10795 & w11007 ) | ( ~w10795 & w11008 ) | ( w11007 & w11008 ) ;
  assign w11010 = w11008 | w11009 ;
  assign w11011 = \pi088 ^ w10782 ;
  assign w11012 = ( ~w10789 & w11010 ) | ( ~w10789 & w11011 ) | ( w11010 & w11011 ) ;
  assign w11013 = w11011 | w11012 ;
  assign w11014 = \pi089 ^ w10776 ;
  assign w11015 = ( ~w10783 & w11013 ) | ( ~w10783 & w11014 ) | ( w11013 & w11014 ) ;
  assign w11016 = w11014 | w11015 ;
  assign w11017 = \pi090 ^ w10770 ;
  assign w11018 = ( ~w10777 & w11016 ) | ( ~w10777 & w11017 ) | ( w11016 & w11017 ) ;
  assign w11019 = w11017 | w11018 ;
  assign w11020 = \pi091 ^ w10764 ;
  assign w11021 = ( ~w10771 & w11019 ) | ( ~w10771 & w11020 ) | ( w11019 & w11020 ) ;
  assign w11022 = w11020 | w11021 ;
  assign w11023 = \pi092 ^ w10758 ;
  assign w11024 = ( ~w10765 & w11022 ) | ( ~w10765 & w11023 ) | ( w11022 & w11023 ) ;
  assign w11025 = w11023 | w11024 ;
  assign w11026 = \pi093 ^ w10752 ;
  assign w11027 = ( ~w10759 & w11025 ) | ( ~w10759 & w11026 ) | ( w11025 & w11026 ) ;
  assign w11028 = w11026 | w11027 ;
  assign w11029 = \pi094 ^ w10746 ;
  assign w11030 = ( ~w10753 & w11028 ) | ( ~w10753 & w11029 ) | ( w11028 & w11029 ) ;
  assign w11031 = w11029 | w11030 ;
  assign w11032 = \pi095 ^ w10740 ;
  assign w11033 = ( ~w10747 & w11031 ) | ( ~w10747 & w11032 ) | ( w11031 & w11032 ) ;
  assign w11034 = w11032 | w11033 ;
  assign w11035 = \pi096 ^ w10734 ;
  assign w11036 = ( ~w10741 & w11034 ) | ( ~w10741 & w11035 ) | ( w11034 & w11035 ) ;
  assign w11037 = w11035 | w11036 ;
  assign w11038 = \pi097 ^ w10728 ;
  assign w11039 = ( ~w10735 & w11037 ) | ( ~w10735 & w11038 ) | ( w11037 & w11038 ) ;
  assign w11040 = w11038 | w11039 ;
  assign w11041 = \pi098 ^ w10722 ;
  assign w11042 = ( ~w10729 & w11040 ) | ( ~w10729 & w11041 ) | ( w11040 & w11041 ) ;
  assign w11043 = w11041 | w11042 ;
  assign w11044 = \pi099 ^ w10716 ;
  assign w11045 = ( ~w10723 & w11043 ) | ( ~w10723 & w11044 ) | ( w11043 & w11044 ) ;
  assign w11046 = w11044 | w11045 ;
  assign w11047 = \pi100 ^ w10710 ;
  assign w11048 = ( ~w10717 & w11046 ) | ( ~w10717 & w11047 ) | ( w11046 & w11047 ) ;
  assign w11049 = w11047 | w11048 ;
  assign w11050 = \pi101 ^ w10704 ;
  assign w11051 = ( ~w10711 & w11049 ) | ( ~w10711 & w11050 ) | ( w11049 & w11050 ) ;
  assign w11052 = w11050 | w11051 ;
  assign w11053 = \pi102 ^ w10698 ;
  assign w11054 = ( ~w10705 & w11052 ) | ( ~w10705 & w11053 ) | ( w11052 & w11053 ) ;
  assign w11055 = w11053 | w11054 ;
  assign w11056 = \pi103 ^ w10692 ;
  assign w11057 = ( ~w10699 & w11055 ) | ( ~w10699 & w11056 ) | ( w11055 & w11056 ) ;
  assign w11058 = w11056 | w11057 ;
  assign w11059 = \pi104 ^ w10686 ;
  assign w11060 = ( ~w10693 & w11058 ) | ( ~w10693 & w11059 ) | ( w11058 & w11059 ) ;
  assign w11061 = w11059 | w11060 ;
  assign w11062 = \pi105 ^ w10680 ;
  assign w11063 = ( ~w10687 & w11061 ) | ( ~w10687 & w11062 ) | ( w11061 & w11062 ) ;
  assign w11064 = w11062 | w11063 ;
  assign w11065 = \pi106 ^ w10674 ;
  assign w11066 = ( ~w10681 & w11064 ) | ( ~w10681 & w11065 ) | ( w11064 & w11065 ) ;
  assign w11067 = w11065 | w11066 ;
  assign w11068 = \pi107 ^ w10668 ;
  assign w11069 = ( ~w10675 & w11067 ) | ( ~w10675 & w11068 ) | ( w11067 & w11068 ) ;
  assign w11070 = w11068 | w11069 ;
  assign w11071 = \pi108 ^ w10662 ;
  assign w11072 = ( ~w10669 & w11070 ) | ( ~w10669 & w11071 ) | ( w11070 & w11071 ) ;
  assign w11073 = w11071 | w11072 ;
  assign w11074 = \pi109 ^ w10656 ;
  assign w11075 = ( ~w10663 & w11073 ) | ( ~w10663 & w11074 ) | ( w11073 & w11074 ) ;
  assign w11076 = w11074 | w11075 ;
  assign w11077 = w10213 & w10651 ;
  assign w11078 = ~w10214 & w10642 ;
  assign w11079 = w10643 ^ w11078 ;
  assign w11080 = ~w10651 & w11079 ;
  assign w11081 = w11077 | w11080 ;
  assign w11082 = ~\pi110 & w11081 ;
  assign w11083 = ( \pi110 & ~w11077 ) | ( \pi110 & w11080 ) | ( ~w11077 & w11080 ) ;
  assign w11084 = ~w11080 & w11083 ;
  assign w11085 = \pi112 | w267 ;
  assign w11086 = ( \pi111 & ~w267 ) | ( \pi111 & w448 ) | ( ~w267 & w448 ) ;
  assign w11087 = w11085 | w11086 ;
  assign w11088 = w11082 | w11084 ;
  assign w11089 = ( ~w10657 & w11076 ) | ( ~w10657 & w11088 ) | ( w11076 & w11088 ) ;
  assign w11090 = ( w11087 & ~w11088 ) | ( w11087 & w11089 ) | ( ~w11088 & w11089 ) ;
  assign w11091 = w11088 | w11090 ;
  assign w11092 = ~w10650 & w11081 ;
  assign w11093 = w11091 & ~w11092 ;
  assign w11094 = ~w10663 & w11073 ;
  assign w11095 = w11074 ^ w11094 ;
  assign w11096 = ~w11093 & w11095 ;
  assign w11097 = ( w10656 & w11091 ) | ( w10656 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11098 = ~w11092 & w11097 ;
  assign w11099 = w11096 | w11098 ;
  assign w11100 = ~\pi110 & w11099 ;
  assign w11101 = ~w10669 & w11070 ;
  assign w11102 = w11071 ^ w11101 ;
  assign w11103 = ~w11093 & w11102 ;
  assign w11104 = ( w10662 & w11091 ) | ( w10662 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11105 = ~w11092 & w11104 ;
  assign w11106 = w11103 | w11105 ;
  assign w11107 = ~\pi109 & w11106 ;
  assign w11108 = ~w10675 & w11067 ;
  assign w11109 = w11068 ^ w11108 ;
  assign w11110 = ~w11093 & w11109 ;
  assign w11111 = ( w10668 & w11091 ) | ( w10668 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11112 = ~w11092 & w11111 ;
  assign w11113 = w11110 | w11112 ;
  assign w11114 = ~\pi108 & w11113 ;
  assign w11115 = ~w10681 & w11064 ;
  assign w11116 = w11065 ^ w11115 ;
  assign w11117 = ~w11093 & w11116 ;
  assign w11118 = ( w10674 & w11091 ) | ( w10674 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11119 = ~w11092 & w11118 ;
  assign w11120 = w11117 | w11119 ;
  assign w11121 = ~\pi107 & w11120 ;
  assign w11122 = ~w10687 & w11061 ;
  assign w11123 = w11062 ^ w11122 ;
  assign w11124 = ~w11093 & w11123 ;
  assign w11125 = ( w10680 & w11091 ) | ( w10680 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11126 = ~w11092 & w11125 ;
  assign w11127 = w11124 | w11126 ;
  assign w11128 = ~\pi106 & w11127 ;
  assign w11129 = ~w10693 & w11058 ;
  assign w11130 = w11059 ^ w11129 ;
  assign w11131 = ~w11093 & w11130 ;
  assign w11132 = ( w10686 & w11091 ) | ( w10686 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11133 = ~w11092 & w11132 ;
  assign w11134 = w11131 | w11133 ;
  assign w11135 = ~\pi105 & w11134 ;
  assign w11136 = ~w10699 & w11055 ;
  assign w11137 = w11056 ^ w11136 ;
  assign w11138 = ~w11093 & w11137 ;
  assign w11139 = ( w10692 & w11091 ) | ( w10692 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11140 = ~w11092 & w11139 ;
  assign w11141 = w11138 | w11140 ;
  assign w11142 = ~\pi104 & w11141 ;
  assign w11143 = ~w10705 & w11052 ;
  assign w11144 = w11053 ^ w11143 ;
  assign w11145 = ~w11093 & w11144 ;
  assign w11146 = ( w10698 & w11091 ) | ( w10698 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11147 = ~w11092 & w11146 ;
  assign w11148 = w11145 | w11147 ;
  assign w11149 = ~\pi103 & w11148 ;
  assign w11150 = ~w10711 & w11049 ;
  assign w11151 = w11050 ^ w11150 ;
  assign w11152 = ~w11093 & w11151 ;
  assign w11153 = ( w10704 & w11091 ) | ( w10704 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11154 = ~w11092 & w11153 ;
  assign w11155 = w11152 | w11154 ;
  assign w11156 = ~\pi102 & w11155 ;
  assign w11157 = ~w10717 & w11046 ;
  assign w11158 = w11047 ^ w11157 ;
  assign w11159 = ~w11093 & w11158 ;
  assign w11160 = ( w10710 & w11091 ) | ( w10710 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11161 = ~w11092 & w11160 ;
  assign w11162 = w11159 | w11161 ;
  assign w11163 = ~\pi101 & w11162 ;
  assign w11164 = ~w10723 & w11043 ;
  assign w11165 = w11044 ^ w11164 ;
  assign w11166 = ~w11093 & w11165 ;
  assign w11167 = ( w10716 & w11091 ) | ( w10716 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11168 = ~w11092 & w11167 ;
  assign w11169 = w11166 | w11168 ;
  assign w11170 = ~\pi100 & w11169 ;
  assign w11171 = ~w10729 & w11040 ;
  assign w11172 = w11041 ^ w11171 ;
  assign w11173 = ~w11093 & w11172 ;
  assign w11174 = ( w10722 & w11091 ) | ( w10722 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11175 = ~w11092 & w11174 ;
  assign w11176 = w11173 | w11175 ;
  assign w11177 = ~\pi099 & w11176 ;
  assign w11178 = ~w10735 & w11037 ;
  assign w11179 = w11038 ^ w11178 ;
  assign w11180 = ~w11093 & w11179 ;
  assign w11181 = ( w10728 & w11091 ) | ( w10728 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11182 = ~w11092 & w11181 ;
  assign w11183 = w11180 | w11182 ;
  assign w11184 = ~\pi098 & w11183 ;
  assign w11185 = ~w10741 & w11034 ;
  assign w11186 = w11035 ^ w11185 ;
  assign w11187 = ~w11093 & w11186 ;
  assign w11188 = ( w10734 & w11091 ) | ( w10734 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11189 = ~w11092 & w11188 ;
  assign w11190 = w11187 | w11189 ;
  assign w11191 = ~\pi097 & w11190 ;
  assign w11192 = ~w10747 & w11031 ;
  assign w11193 = w11032 ^ w11192 ;
  assign w11194 = ~w11093 & w11193 ;
  assign w11195 = ( w10740 & w11091 ) | ( w10740 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11196 = ~w11092 & w11195 ;
  assign w11197 = w11194 | w11196 ;
  assign w11198 = ~\pi096 & w11197 ;
  assign w11199 = ~w10753 & w11028 ;
  assign w11200 = w11029 ^ w11199 ;
  assign w11201 = ~w11093 & w11200 ;
  assign w11202 = ( w10746 & w11091 ) | ( w10746 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11203 = ~w11092 & w11202 ;
  assign w11204 = w11201 | w11203 ;
  assign w11205 = ~\pi095 & w11204 ;
  assign w11206 = ~w10759 & w11025 ;
  assign w11207 = w11026 ^ w11206 ;
  assign w11208 = ~w11093 & w11207 ;
  assign w11209 = ( w10752 & w11091 ) | ( w10752 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11210 = ~w11092 & w11209 ;
  assign w11211 = w11208 | w11210 ;
  assign w11212 = ~\pi094 & w11211 ;
  assign w11213 = ~w10765 & w11022 ;
  assign w11214 = w11023 ^ w11213 ;
  assign w11215 = ~w11093 & w11214 ;
  assign w11216 = ( w10758 & w11091 ) | ( w10758 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11217 = ~w11092 & w11216 ;
  assign w11218 = w11215 | w11217 ;
  assign w11219 = ~\pi093 & w11218 ;
  assign w11220 = ~w10771 & w11019 ;
  assign w11221 = w11020 ^ w11220 ;
  assign w11222 = ~w11093 & w11221 ;
  assign w11223 = ( w10764 & w11091 ) | ( w10764 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11224 = ~w11092 & w11223 ;
  assign w11225 = w11222 | w11224 ;
  assign w11226 = ~\pi092 & w11225 ;
  assign w11227 = ~w10777 & w11016 ;
  assign w11228 = w11017 ^ w11227 ;
  assign w11229 = ~w11093 & w11228 ;
  assign w11230 = ( w10770 & w11091 ) | ( w10770 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11231 = ~w11092 & w11230 ;
  assign w11232 = w11229 | w11231 ;
  assign w11233 = ~\pi091 & w11232 ;
  assign w11234 = ~w10783 & w11013 ;
  assign w11235 = w11014 ^ w11234 ;
  assign w11236 = ~w11093 & w11235 ;
  assign w11237 = ( w10776 & w11091 ) | ( w10776 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11238 = ~w11092 & w11237 ;
  assign w11239 = w11236 | w11238 ;
  assign w11240 = ~\pi090 & w11239 ;
  assign w11241 = ~w10789 & w11010 ;
  assign w11242 = w11011 ^ w11241 ;
  assign w11243 = ~w11093 & w11242 ;
  assign w11244 = ( w10782 & w11091 ) | ( w10782 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11245 = ~w11092 & w11244 ;
  assign w11246 = w11243 | w11245 ;
  assign w11247 = ~\pi089 & w11246 ;
  assign w11248 = ~w10795 & w11007 ;
  assign w11249 = w11008 ^ w11248 ;
  assign w11250 = ~w11093 & w11249 ;
  assign w11251 = ( w10788 & w11091 ) | ( w10788 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11252 = ~w11092 & w11251 ;
  assign w11253 = w11250 | w11252 ;
  assign w11254 = ~\pi088 & w11253 ;
  assign w11255 = ~w10801 & w11004 ;
  assign w11256 = w11005 ^ w11255 ;
  assign w11257 = ~w11093 & w11256 ;
  assign w11258 = ( w10794 & w11091 ) | ( w10794 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11259 = ~w11092 & w11258 ;
  assign w11260 = w11257 | w11259 ;
  assign w11261 = ~\pi087 & w11260 ;
  assign w11262 = ~w10807 & w11001 ;
  assign w11263 = w11002 ^ w11262 ;
  assign w11264 = ~w11093 & w11263 ;
  assign w11265 = ( w10800 & w11091 ) | ( w10800 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11266 = ~w11092 & w11265 ;
  assign w11267 = w11264 | w11266 ;
  assign w11268 = ~\pi086 & w11267 ;
  assign w11269 = ~w10813 & w10998 ;
  assign w11270 = w10999 ^ w11269 ;
  assign w11271 = ~w11093 & w11270 ;
  assign w11272 = ( w10806 & w11091 ) | ( w10806 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11273 = ~w11092 & w11272 ;
  assign w11274 = w11271 | w11273 ;
  assign w11275 = ~\pi085 & w11274 ;
  assign w11276 = ~w10819 & w10995 ;
  assign w11277 = w10996 ^ w11276 ;
  assign w11278 = ~w11093 & w11277 ;
  assign w11279 = ( w10812 & w11091 ) | ( w10812 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11280 = ~w11092 & w11279 ;
  assign w11281 = w11278 | w11280 ;
  assign w11282 = ~\pi084 & w11281 ;
  assign w11283 = ~w10825 & w10992 ;
  assign w11284 = w10993 ^ w11283 ;
  assign w11285 = ~w11093 & w11284 ;
  assign w11286 = ( w10818 & w11091 ) | ( w10818 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11287 = ~w11092 & w11286 ;
  assign w11288 = w11285 | w11287 ;
  assign w11289 = ~\pi083 & w11288 ;
  assign w11290 = ~w10831 & w10989 ;
  assign w11291 = w10990 ^ w11290 ;
  assign w11292 = ~w11093 & w11291 ;
  assign w11293 = ( w10824 & w11091 ) | ( w10824 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11294 = ~w11092 & w11293 ;
  assign w11295 = w11292 | w11294 ;
  assign w11296 = ~\pi082 & w11295 ;
  assign w11297 = ~w10837 & w10986 ;
  assign w11298 = w10987 ^ w11297 ;
  assign w11299 = ~w11093 & w11298 ;
  assign w11300 = ( w10830 & w11091 ) | ( w10830 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11301 = ~w11092 & w11300 ;
  assign w11302 = w11299 | w11301 ;
  assign w11303 = ~\pi081 & w11302 ;
  assign w11304 = ~w10843 & w10983 ;
  assign w11305 = w10984 ^ w11304 ;
  assign w11306 = ~w11093 & w11305 ;
  assign w11307 = ( w10836 & w11091 ) | ( w10836 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11308 = ~w11092 & w11307 ;
  assign w11309 = w11306 | w11308 ;
  assign w11310 = ~\pi080 & w11309 ;
  assign w11311 = ~w10849 & w10980 ;
  assign w11312 = w10981 ^ w11311 ;
  assign w11313 = ~w11093 & w11312 ;
  assign w11314 = ( w10842 & w11091 ) | ( w10842 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11315 = ~w11092 & w11314 ;
  assign w11316 = w11313 | w11315 ;
  assign w11317 = ~\pi079 & w11316 ;
  assign w11318 = ~w10855 & w10977 ;
  assign w11319 = w10978 ^ w11318 ;
  assign w11320 = ~w11093 & w11319 ;
  assign w11321 = ( w10848 & w11091 ) | ( w10848 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11322 = ~w11092 & w11321 ;
  assign w11323 = w11320 | w11322 ;
  assign w11324 = ~\pi078 & w11323 ;
  assign w11325 = ~w10861 & w10974 ;
  assign w11326 = w10975 ^ w11325 ;
  assign w11327 = ~w11093 & w11326 ;
  assign w11328 = ( w10854 & w11091 ) | ( w10854 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11329 = ~w11092 & w11328 ;
  assign w11330 = w11327 | w11329 ;
  assign w11331 = ~\pi077 & w11330 ;
  assign w11332 = ~w10867 & w10971 ;
  assign w11333 = w10972 ^ w11332 ;
  assign w11334 = ~w11093 & w11333 ;
  assign w11335 = ( w10860 & w11091 ) | ( w10860 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11336 = ~w11092 & w11335 ;
  assign w11337 = w11334 | w11336 ;
  assign w11338 = ~\pi076 & w11337 ;
  assign w11339 = ~w10873 & w10968 ;
  assign w11340 = w10969 ^ w11339 ;
  assign w11341 = ~w11093 & w11340 ;
  assign w11342 = ( w10866 & w11091 ) | ( w10866 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11343 = ~w11092 & w11342 ;
  assign w11344 = w11341 | w11343 ;
  assign w11345 = ~\pi075 & w11344 ;
  assign w11346 = ~w10879 & w10965 ;
  assign w11347 = w10966 ^ w11346 ;
  assign w11348 = ~w11093 & w11347 ;
  assign w11349 = ( w10872 & w11091 ) | ( w10872 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11350 = ~w11092 & w11349 ;
  assign w11351 = w11348 | w11350 ;
  assign w11352 = ~\pi074 & w11351 ;
  assign w11353 = ~w10885 & w10962 ;
  assign w11354 = w10963 ^ w11353 ;
  assign w11355 = ~w11093 & w11354 ;
  assign w11356 = ( w10878 & w11091 ) | ( w10878 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11357 = ~w11092 & w11356 ;
  assign w11358 = w11355 | w11357 ;
  assign w11359 = ~\pi073 & w11358 ;
  assign w11360 = ~w10891 & w10959 ;
  assign w11361 = w10960 ^ w11360 ;
  assign w11362 = ~w11093 & w11361 ;
  assign w11363 = ( w10884 & w11091 ) | ( w10884 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11364 = ~w11092 & w11363 ;
  assign w11365 = w11362 | w11364 ;
  assign w11366 = ~\pi072 & w11365 ;
  assign w11367 = ~w10897 & w10956 ;
  assign w11368 = w10957 ^ w11367 ;
  assign w11369 = ~w11093 & w11368 ;
  assign w11370 = ( w10890 & w11091 ) | ( w10890 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11371 = ~w11092 & w11370 ;
  assign w11372 = w11369 | w11371 ;
  assign w11373 = ~\pi071 & w11372 ;
  assign w11374 = ~w10903 & w10953 ;
  assign w11375 = w10954 ^ w11374 ;
  assign w11376 = ~w11093 & w11375 ;
  assign w11377 = ( w10896 & w11091 ) | ( w10896 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11378 = ~w11092 & w11377 ;
  assign w11379 = w11376 | w11378 ;
  assign w11380 = ~\pi070 & w11379 ;
  assign w11381 = ~w10911 & w10950 ;
  assign w11382 = w10951 ^ w11381 ;
  assign w11383 = ~w11093 & w11382 ;
  assign w11384 = ( w10902 & w11091 ) | ( w10902 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11385 = ~w11092 & w11384 ;
  assign w11386 = w11383 | w11385 ;
  assign w11387 = ~\pi069 & w11386 ;
  assign w11388 = ~w10922 & w10945 ;
  assign w11389 = w10948 ^ w11388 ;
  assign w11390 = ~w11093 & w11389 ;
  assign w11391 = ( w10910 & w11091 ) | ( w10910 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11392 = ~w11092 & w11391 ;
  assign w11393 = w11390 | w11392 ;
  assign w11394 = ~\pi068 & w11393 ;
  assign w11395 = ( \pi065 & w10936 ) | ( \pi065 & ~w11093 ) | ( w10936 & ~w11093 ) ;
  assign w11396 = ( \pi065 & w10939 ) | ( \pi065 & ~w11395 ) | ( w10939 & ~w11395 ) ;
  assign w11397 = w10942 ^ w11396 ;
  assign w11398 = ~w11093 & w11397 ;
  assign w11399 = ( w10921 & w11091 ) | ( w10921 & w11092 ) | ( w11091 & w11092 ) ;
  assign w11400 = ~w11092 & w11399 ;
  assign w11401 = w11398 | w11400 ;
  assign w11402 = ~\pi067 & w11401 ;
  assign w11403 = w10936 ^ w10937 ;
  assign w11404 = \pi065 ^ w11403 ;
  assign w11405 = w11093 ^ w11404 ;
  assign w11406 = ( w10936 & w11404 ) | ( w10936 & w11405 ) | ( w11404 & w11405 ) ;
  assign w11407 = ~\pi066 & w11406 ;
  assign w11408 = w10936 ^ w11093 ;
  assign w11409 = ( w10936 & w11404 ) | ( w10936 & ~w11408 ) | ( w11404 & ~w11408 ) ;
  assign w11410 = \pi066 ^ w11409 ;
  assign w11411 = \pi064 & ~w11093 ;
  assign w11412 = \pi017 ^ w11411 ;
  assign w11413 = ( ~\pi016 & \pi064 ) | ( ~\pi016 & w11410 ) | ( \pi064 & w11410 ) ;
  assign w11414 = ( \pi065 & ~w11412 ) | ( \pi065 & w11413 ) | ( ~w11412 & w11413 ) ;
  assign w11415 = w11410 | w11414 ;
  assign w11416 = \pi067 ^ w11401 ;
  assign w11417 = ( ~w11407 & w11415 ) | ( ~w11407 & w11416 ) | ( w11415 & w11416 ) ;
  assign w11418 = w11416 | w11417 ;
  assign w11419 = \pi068 ^ w11393 ;
  assign w11420 = ( ~w11402 & w11418 ) | ( ~w11402 & w11419 ) | ( w11418 & w11419 ) ;
  assign w11421 = w11419 | w11420 ;
  assign w11422 = \pi069 ^ w11386 ;
  assign w11423 = ( ~w11394 & w11421 ) | ( ~w11394 & w11422 ) | ( w11421 & w11422 ) ;
  assign w11424 = w11422 | w11423 ;
  assign w11425 = \pi070 ^ w11379 ;
  assign w11426 = ( ~w11387 & w11424 ) | ( ~w11387 & w11425 ) | ( w11424 & w11425 ) ;
  assign w11427 = w11425 | w11426 ;
  assign w11428 = \pi071 ^ w11372 ;
  assign w11429 = ( ~w11380 & w11427 ) | ( ~w11380 & w11428 ) | ( w11427 & w11428 ) ;
  assign w11430 = w11428 | w11429 ;
  assign w11431 = \pi072 ^ w11365 ;
  assign w11432 = ( ~w11373 & w11430 ) | ( ~w11373 & w11431 ) | ( w11430 & w11431 ) ;
  assign w11433 = w11431 | w11432 ;
  assign w11434 = \pi073 ^ w11358 ;
  assign w11435 = ( ~w11366 & w11433 ) | ( ~w11366 & w11434 ) | ( w11433 & w11434 ) ;
  assign w11436 = w11434 | w11435 ;
  assign w11437 = \pi074 ^ w11351 ;
  assign w11438 = ( ~w11359 & w11436 ) | ( ~w11359 & w11437 ) | ( w11436 & w11437 ) ;
  assign w11439 = w11437 | w11438 ;
  assign w11440 = \pi075 ^ w11344 ;
  assign w11441 = ( ~w11352 & w11439 ) | ( ~w11352 & w11440 ) | ( w11439 & w11440 ) ;
  assign w11442 = w11440 | w11441 ;
  assign w11443 = \pi076 ^ w11337 ;
  assign w11444 = ( ~w11345 & w11442 ) | ( ~w11345 & w11443 ) | ( w11442 & w11443 ) ;
  assign w11445 = w11443 | w11444 ;
  assign w11446 = \pi077 ^ w11330 ;
  assign w11447 = ( ~w11338 & w11445 ) | ( ~w11338 & w11446 ) | ( w11445 & w11446 ) ;
  assign w11448 = w11446 | w11447 ;
  assign w11449 = \pi078 ^ w11323 ;
  assign w11450 = ( ~w11331 & w11448 ) | ( ~w11331 & w11449 ) | ( w11448 & w11449 ) ;
  assign w11451 = w11449 | w11450 ;
  assign w11452 = \pi079 ^ w11316 ;
  assign w11453 = ( ~w11324 & w11451 ) | ( ~w11324 & w11452 ) | ( w11451 & w11452 ) ;
  assign w11454 = w11452 | w11453 ;
  assign w11455 = \pi080 ^ w11309 ;
  assign w11456 = ( ~w11317 & w11454 ) | ( ~w11317 & w11455 ) | ( w11454 & w11455 ) ;
  assign w11457 = w11455 | w11456 ;
  assign w11458 = \pi081 ^ w11302 ;
  assign w11459 = ( ~w11310 & w11457 ) | ( ~w11310 & w11458 ) | ( w11457 & w11458 ) ;
  assign w11460 = w11458 | w11459 ;
  assign w11461 = \pi082 ^ w11295 ;
  assign w11462 = ( ~w11303 & w11460 ) | ( ~w11303 & w11461 ) | ( w11460 & w11461 ) ;
  assign w11463 = w11461 | w11462 ;
  assign w11464 = \pi083 ^ w11288 ;
  assign w11465 = ( ~w11296 & w11463 ) | ( ~w11296 & w11464 ) | ( w11463 & w11464 ) ;
  assign w11466 = w11464 | w11465 ;
  assign w11467 = \pi084 ^ w11281 ;
  assign w11468 = ( ~w11289 & w11466 ) | ( ~w11289 & w11467 ) | ( w11466 & w11467 ) ;
  assign w11469 = w11467 | w11468 ;
  assign w11470 = \pi085 ^ w11274 ;
  assign w11471 = ( ~w11282 & w11469 ) | ( ~w11282 & w11470 ) | ( w11469 & w11470 ) ;
  assign w11472 = w11470 | w11471 ;
  assign w11473 = \pi086 ^ w11267 ;
  assign w11474 = ( ~w11275 & w11472 ) | ( ~w11275 & w11473 ) | ( w11472 & w11473 ) ;
  assign w11475 = w11473 | w11474 ;
  assign w11476 = \pi087 ^ w11260 ;
  assign w11477 = ( ~w11268 & w11475 ) | ( ~w11268 & w11476 ) | ( w11475 & w11476 ) ;
  assign w11478 = w11476 | w11477 ;
  assign w11479 = \pi088 ^ w11253 ;
  assign w11480 = ( ~w11261 & w11478 ) | ( ~w11261 & w11479 ) | ( w11478 & w11479 ) ;
  assign w11481 = w11479 | w11480 ;
  assign w11482 = \pi089 ^ w11246 ;
  assign w11483 = ( ~w11254 & w11481 ) | ( ~w11254 & w11482 ) | ( w11481 & w11482 ) ;
  assign w11484 = w11482 | w11483 ;
  assign w11485 = \pi090 ^ w11239 ;
  assign w11486 = ( ~w11247 & w11484 ) | ( ~w11247 & w11485 ) | ( w11484 & w11485 ) ;
  assign w11487 = w11485 | w11486 ;
  assign w11488 = \pi091 ^ w11232 ;
  assign w11489 = ( ~w11240 & w11487 ) | ( ~w11240 & w11488 ) | ( w11487 & w11488 ) ;
  assign w11490 = w11488 | w11489 ;
  assign w11491 = \pi092 ^ w11225 ;
  assign w11492 = ( ~w11233 & w11490 ) | ( ~w11233 & w11491 ) | ( w11490 & w11491 ) ;
  assign w11493 = w11491 | w11492 ;
  assign w11494 = \pi093 ^ w11218 ;
  assign w11495 = ( ~w11226 & w11493 ) | ( ~w11226 & w11494 ) | ( w11493 & w11494 ) ;
  assign w11496 = w11494 | w11495 ;
  assign w11497 = \pi094 ^ w11211 ;
  assign w11498 = ( ~w11219 & w11496 ) | ( ~w11219 & w11497 ) | ( w11496 & w11497 ) ;
  assign w11499 = w11497 | w11498 ;
  assign w11500 = \pi095 ^ w11204 ;
  assign w11501 = ( ~w11212 & w11499 ) | ( ~w11212 & w11500 ) | ( w11499 & w11500 ) ;
  assign w11502 = w11500 | w11501 ;
  assign w11503 = \pi096 ^ w11197 ;
  assign w11504 = ( ~w11205 & w11502 ) | ( ~w11205 & w11503 ) | ( w11502 & w11503 ) ;
  assign w11505 = w11503 | w11504 ;
  assign w11506 = \pi097 ^ w11190 ;
  assign w11507 = ( ~w11198 & w11505 ) | ( ~w11198 & w11506 ) | ( w11505 & w11506 ) ;
  assign w11508 = w11506 | w11507 ;
  assign w11509 = \pi098 ^ w11183 ;
  assign w11510 = ( ~w11191 & w11508 ) | ( ~w11191 & w11509 ) | ( w11508 & w11509 ) ;
  assign w11511 = w11509 | w11510 ;
  assign w11512 = \pi099 ^ w11176 ;
  assign w11513 = ( ~w11184 & w11511 ) | ( ~w11184 & w11512 ) | ( w11511 & w11512 ) ;
  assign w11514 = w11512 | w11513 ;
  assign w11515 = \pi100 ^ w11169 ;
  assign w11516 = ( ~w11177 & w11514 ) | ( ~w11177 & w11515 ) | ( w11514 & w11515 ) ;
  assign w11517 = w11515 | w11516 ;
  assign w11518 = \pi101 ^ w11162 ;
  assign w11519 = ( ~w11170 & w11517 ) | ( ~w11170 & w11518 ) | ( w11517 & w11518 ) ;
  assign w11520 = w11518 | w11519 ;
  assign w11521 = \pi102 ^ w11155 ;
  assign w11522 = ( ~w11163 & w11520 ) | ( ~w11163 & w11521 ) | ( w11520 & w11521 ) ;
  assign w11523 = w11521 | w11522 ;
  assign w11524 = \pi103 ^ w11148 ;
  assign w11525 = ( ~w11156 & w11523 ) | ( ~w11156 & w11524 ) | ( w11523 & w11524 ) ;
  assign w11526 = w11524 | w11525 ;
  assign w11527 = \pi104 ^ w11141 ;
  assign w11528 = ( ~w11149 & w11526 ) | ( ~w11149 & w11527 ) | ( w11526 & w11527 ) ;
  assign w11529 = w11527 | w11528 ;
  assign w11530 = \pi105 ^ w11134 ;
  assign w11531 = ( ~w11142 & w11529 ) | ( ~w11142 & w11530 ) | ( w11529 & w11530 ) ;
  assign w11532 = w11530 | w11531 ;
  assign w11533 = \pi106 ^ w11127 ;
  assign w11534 = ( ~w11135 & w11532 ) | ( ~w11135 & w11533 ) | ( w11532 & w11533 ) ;
  assign w11535 = w11533 | w11534 ;
  assign w11536 = \pi107 ^ w11120 ;
  assign w11537 = ( ~w11128 & w11535 ) | ( ~w11128 & w11536 ) | ( w11535 & w11536 ) ;
  assign w11538 = w11536 | w11537 ;
  assign w11539 = \pi108 ^ w11113 ;
  assign w11540 = ( ~w11121 & w11538 ) | ( ~w11121 & w11539 ) | ( w11538 & w11539 ) ;
  assign w11541 = w11539 | w11540 ;
  assign w11542 = \pi109 ^ w11106 ;
  assign w11543 = ( ~w11114 & w11541 ) | ( ~w11114 & w11542 ) | ( w11541 & w11542 ) ;
  assign w11544 = w11542 | w11543 ;
  assign w11545 = \pi110 ^ w11099 ;
  assign w11546 = ( ~w11107 & w11544 ) | ( ~w11107 & w11545 ) | ( w11544 & w11545 ) ;
  assign w11547 = w11545 | w11546 ;
  assign w11548 = ( ~w10657 & w11076 ) | ( ~w10657 & w11093 ) | ( w11076 & w11093 ) ;
  assign w11549 = w11088 ^ w11548 ;
  assign w11550 = ~w11093 & w11549 ;
  assign w11551 = ( w10650 & ~w11081 ) | ( w10650 & w11091 ) | ( ~w11081 & w11091 ) ;
  assign w11552 = w11081 & w11551 ;
  assign w11553 = w11550 | w11552 ;
  assign w11554 = ~\pi111 & w11553 ;
  assign w11555 = ( \pi111 & ~w11550 ) | ( \pi111 & w11552 ) | ( ~w11550 & w11552 ) ;
  assign w11556 = ~w11552 & w11555 ;
  assign w11557 = w11554 | w11556 ;
  assign w11558 = ( ~w11100 & w11547 ) | ( ~w11100 & w11557 ) | ( w11547 & w11557 ) ;
  assign w11559 = ( w201 & ~w11557 ) | ( w201 & w11558 ) | ( ~w11557 & w11558 ) ;
  assign w11560 = w11557 | w11559 ;
  assign w11561 = ~w11087 & w11553 ;
  assign w11562 = w11560 & ~w11561 ;
  assign w11563 = ~w11107 & w11544 ;
  assign w11564 = w11545 ^ w11563 ;
  assign w11565 = ~w11562 & w11564 ;
  assign w11566 = ( w11099 & w11560 ) | ( w11099 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11567 = ~w11561 & w11566 ;
  assign w11568 = w11565 | w11567 ;
  assign w11569 = ( ~w11100 & w11547 ) | ( ~w11100 & w11562 ) | ( w11547 & w11562 ) ;
  assign w11570 = w11557 ^ w11569 ;
  assign w11571 = ~w11562 & w11570 ;
  assign w11572 = ( w11087 & ~w11553 ) | ( w11087 & w11560 ) | ( ~w11553 & w11560 ) ;
  assign w11573 = w11553 & w11572 ;
  assign w11574 = w11571 | w11573 ;
  assign w11575 = ~\pi111 & w11568 ;
  assign w11576 = ~w11114 & w11541 ;
  assign w11577 = w11542 ^ w11576 ;
  assign w11578 = ~w11562 & w11577 ;
  assign w11579 = ( w11106 & w11560 ) | ( w11106 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11580 = ~w11561 & w11579 ;
  assign w11581 = w11578 | w11580 ;
  assign w11582 = ~\pi110 & w11581 ;
  assign w11583 = ~w11121 & w11538 ;
  assign w11584 = w11539 ^ w11583 ;
  assign w11585 = ~w11562 & w11584 ;
  assign w11586 = ( w11113 & w11560 ) | ( w11113 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11587 = ~w11561 & w11586 ;
  assign w11588 = w11585 | w11587 ;
  assign w11589 = ~\pi109 & w11588 ;
  assign w11590 = ~w11128 & w11535 ;
  assign w11591 = w11536 ^ w11590 ;
  assign w11592 = ~w11562 & w11591 ;
  assign w11593 = ( w11120 & w11560 ) | ( w11120 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11594 = ~w11561 & w11593 ;
  assign w11595 = w11592 | w11594 ;
  assign w11596 = ~\pi108 & w11595 ;
  assign w11597 = ~w11135 & w11532 ;
  assign w11598 = w11533 ^ w11597 ;
  assign w11599 = ~w11562 & w11598 ;
  assign w11600 = ( w11127 & w11560 ) | ( w11127 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11601 = ~w11561 & w11600 ;
  assign w11602 = w11599 | w11601 ;
  assign w11603 = ~\pi107 & w11602 ;
  assign w11604 = ~w11142 & w11529 ;
  assign w11605 = w11530 ^ w11604 ;
  assign w11606 = ~w11562 & w11605 ;
  assign w11607 = ( w11134 & w11560 ) | ( w11134 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11608 = ~w11561 & w11607 ;
  assign w11609 = w11606 | w11608 ;
  assign w11610 = ~\pi106 & w11609 ;
  assign w11611 = ~w11149 & w11526 ;
  assign w11612 = w11527 ^ w11611 ;
  assign w11613 = ~w11562 & w11612 ;
  assign w11614 = ( w11141 & w11560 ) | ( w11141 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11615 = ~w11561 & w11614 ;
  assign w11616 = w11613 | w11615 ;
  assign w11617 = ~\pi105 & w11616 ;
  assign w11618 = ~w11156 & w11523 ;
  assign w11619 = w11524 ^ w11618 ;
  assign w11620 = ~w11562 & w11619 ;
  assign w11621 = ( w11148 & w11560 ) | ( w11148 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11622 = ~w11561 & w11621 ;
  assign w11623 = w11620 | w11622 ;
  assign w11624 = ~\pi104 & w11623 ;
  assign w11625 = ~w11163 & w11520 ;
  assign w11626 = w11521 ^ w11625 ;
  assign w11627 = ~w11562 & w11626 ;
  assign w11628 = ( w11155 & w11560 ) | ( w11155 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11629 = ~w11561 & w11628 ;
  assign w11630 = w11627 | w11629 ;
  assign w11631 = ~\pi103 & w11630 ;
  assign w11632 = ~w11170 & w11517 ;
  assign w11633 = w11518 ^ w11632 ;
  assign w11634 = ~w11562 & w11633 ;
  assign w11635 = ( w11162 & w11560 ) | ( w11162 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11636 = ~w11561 & w11635 ;
  assign w11637 = w11634 | w11636 ;
  assign w11638 = ~\pi102 & w11637 ;
  assign w11639 = ~w11177 & w11514 ;
  assign w11640 = w11515 ^ w11639 ;
  assign w11641 = ~w11562 & w11640 ;
  assign w11642 = ( w11169 & w11560 ) | ( w11169 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11643 = ~w11561 & w11642 ;
  assign w11644 = w11641 | w11643 ;
  assign w11645 = ~\pi101 & w11644 ;
  assign w11646 = ~w11184 & w11511 ;
  assign w11647 = w11512 ^ w11646 ;
  assign w11648 = ~w11562 & w11647 ;
  assign w11649 = ( w11176 & w11560 ) | ( w11176 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11650 = ~w11561 & w11649 ;
  assign w11651 = w11648 | w11650 ;
  assign w11652 = ~\pi100 & w11651 ;
  assign w11653 = ~w11191 & w11508 ;
  assign w11654 = w11509 ^ w11653 ;
  assign w11655 = ~w11562 & w11654 ;
  assign w11656 = ( w11183 & w11560 ) | ( w11183 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11657 = ~w11561 & w11656 ;
  assign w11658 = w11655 | w11657 ;
  assign w11659 = ~\pi099 & w11658 ;
  assign w11660 = ~w11198 & w11505 ;
  assign w11661 = w11506 ^ w11660 ;
  assign w11662 = ~w11562 & w11661 ;
  assign w11663 = ( w11190 & w11560 ) | ( w11190 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11664 = ~w11561 & w11663 ;
  assign w11665 = w11662 | w11664 ;
  assign w11666 = ~\pi098 & w11665 ;
  assign w11667 = ~w11205 & w11502 ;
  assign w11668 = w11503 ^ w11667 ;
  assign w11669 = ~w11562 & w11668 ;
  assign w11670 = ( w11197 & w11560 ) | ( w11197 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11671 = ~w11561 & w11670 ;
  assign w11672 = w11669 | w11671 ;
  assign w11673 = ~\pi097 & w11672 ;
  assign w11674 = ~w11212 & w11499 ;
  assign w11675 = w11500 ^ w11674 ;
  assign w11676 = ~w11562 & w11675 ;
  assign w11677 = ( w11204 & w11560 ) | ( w11204 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11678 = ~w11561 & w11677 ;
  assign w11679 = w11676 | w11678 ;
  assign w11680 = ~\pi096 & w11679 ;
  assign w11681 = ~w11219 & w11496 ;
  assign w11682 = w11497 ^ w11681 ;
  assign w11683 = ~w11562 & w11682 ;
  assign w11684 = ( w11211 & w11560 ) | ( w11211 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11685 = ~w11561 & w11684 ;
  assign w11686 = w11683 | w11685 ;
  assign w11687 = ~\pi095 & w11686 ;
  assign w11688 = ~w11226 & w11493 ;
  assign w11689 = w11494 ^ w11688 ;
  assign w11690 = ~w11562 & w11689 ;
  assign w11691 = ( w11218 & w11560 ) | ( w11218 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11692 = ~w11561 & w11691 ;
  assign w11693 = w11690 | w11692 ;
  assign w11694 = ~\pi094 & w11693 ;
  assign w11695 = ~w11233 & w11490 ;
  assign w11696 = w11491 ^ w11695 ;
  assign w11697 = ~w11562 & w11696 ;
  assign w11698 = ( w11225 & w11560 ) | ( w11225 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11699 = ~w11561 & w11698 ;
  assign w11700 = w11697 | w11699 ;
  assign w11701 = ~\pi093 & w11700 ;
  assign w11702 = ~w11240 & w11487 ;
  assign w11703 = w11488 ^ w11702 ;
  assign w11704 = ~w11562 & w11703 ;
  assign w11705 = ( w11232 & w11560 ) | ( w11232 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11706 = ~w11561 & w11705 ;
  assign w11707 = w11704 | w11706 ;
  assign w11708 = ~\pi092 & w11707 ;
  assign w11709 = ~w11247 & w11484 ;
  assign w11710 = w11485 ^ w11709 ;
  assign w11711 = ~w11562 & w11710 ;
  assign w11712 = ( w11239 & w11560 ) | ( w11239 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11713 = ~w11561 & w11712 ;
  assign w11714 = w11711 | w11713 ;
  assign w11715 = ~\pi091 & w11714 ;
  assign w11716 = ~w11254 & w11481 ;
  assign w11717 = w11482 ^ w11716 ;
  assign w11718 = ~w11562 & w11717 ;
  assign w11719 = ( w11246 & w11560 ) | ( w11246 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11720 = ~w11561 & w11719 ;
  assign w11721 = w11718 | w11720 ;
  assign w11722 = ~\pi090 & w11721 ;
  assign w11723 = ~w11261 & w11478 ;
  assign w11724 = w11479 ^ w11723 ;
  assign w11725 = ~w11562 & w11724 ;
  assign w11726 = ( w11253 & w11560 ) | ( w11253 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11727 = ~w11561 & w11726 ;
  assign w11728 = w11725 | w11727 ;
  assign w11729 = ~\pi089 & w11728 ;
  assign w11730 = ~w11268 & w11475 ;
  assign w11731 = w11476 ^ w11730 ;
  assign w11732 = ~w11562 & w11731 ;
  assign w11733 = ( w11260 & w11560 ) | ( w11260 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11734 = ~w11561 & w11733 ;
  assign w11735 = w11732 | w11734 ;
  assign w11736 = ~\pi088 & w11735 ;
  assign w11737 = ~w11275 & w11472 ;
  assign w11738 = w11473 ^ w11737 ;
  assign w11739 = ~w11562 & w11738 ;
  assign w11740 = ( w11267 & w11560 ) | ( w11267 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11741 = ~w11561 & w11740 ;
  assign w11742 = w11739 | w11741 ;
  assign w11743 = ~\pi087 & w11742 ;
  assign w11744 = ~w11282 & w11469 ;
  assign w11745 = w11470 ^ w11744 ;
  assign w11746 = ~w11562 & w11745 ;
  assign w11747 = ( w11274 & w11560 ) | ( w11274 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11748 = ~w11561 & w11747 ;
  assign w11749 = w11746 | w11748 ;
  assign w11750 = ~\pi086 & w11749 ;
  assign w11751 = ~w11289 & w11466 ;
  assign w11752 = w11467 ^ w11751 ;
  assign w11753 = ~w11562 & w11752 ;
  assign w11754 = ( w11281 & w11560 ) | ( w11281 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11755 = ~w11561 & w11754 ;
  assign w11756 = w11753 | w11755 ;
  assign w11757 = ~\pi085 & w11756 ;
  assign w11758 = ~w11296 & w11463 ;
  assign w11759 = w11464 ^ w11758 ;
  assign w11760 = ~w11562 & w11759 ;
  assign w11761 = ( w11288 & w11560 ) | ( w11288 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11762 = ~w11561 & w11761 ;
  assign w11763 = w11760 | w11762 ;
  assign w11764 = ~\pi084 & w11763 ;
  assign w11765 = ~w11303 & w11460 ;
  assign w11766 = w11461 ^ w11765 ;
  assign w11767 = ~w11562 & w11766 ;
  assign w11768 = ( w11295 & w11560 ) | ( w11295 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11769 = ~w11561 & w11768 ;
  assign w11770 = w11767 | w11769 ;
  assign w11771 = ~\pi083 & w11770 ;
  assign w11772 = ~w11310 & w11457 ;
  assign w11773 = w11458 ^ w11772 ;
  assign w11774 = ~w11562 & w11773 ;
  assign w11775 = ( w11302 & w11560 ) | ( w11302 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11776 = ~w11561 & w11775 ;
  assign w11777 = w11774 | w11776 ;
  assign w11778 = ~\pi082 & w11777 ;
  assign w11779 = ~w11317 & w11454 ;
  assign w11780 = w11455 ^ w11779 ;
  assign w11781 = ~w11562 & w11780 ;
  assign w11782 = ( w11309 & w11560 ) | ( w11309 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11783 = ~w11561 & w11782 ;
  assign w11784 = w11781 | w11783 ;
  assign w11785 = ~\pi081 & w11784 ;
  assign w11786 = ~w11324 & w11451 ;
  assign w11787 = w11452 ^ w11786 ;
  assign w11788 = ~w11562 & w11787 ;
  assign w11789 = ( w11316 & w11560 ) | ( w11316 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11790 = ~w11561 & w11789 ;
  assign w11791 = w11788 | w11790 ;
  assign w11792 = ~\pi080 & w11791 ;
  assign w11793 = ~w11331 & w11448 ;
  assign w11794 = w11449 ^ w11793 ;
  assign w11795 = ~w11562 & w11794 ;
  assign w11796 = ( w11323 & w11560 ) | ( w11323 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11797 = ~w11561 & w11796 ;
  assign w11798 = w11795 | w11797 ;
  assign w11799 = ~\pi079 & w11798 ;
  assign w11800 = ~w11338 & w11445 ;
  assign w11801 = w11446 ^ w11800 ;
  assign w11802 = ~w11562 & w11801 ;
  assign w11803 = ( w11330 & w11560 ) | ( w11330 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11804 = ~w11561 & w11803 ;
  assign w11805 = w11802 | w11804 ;
  assign w11806 = ~\pi078 & w11805 ;
  assign w11807 = ~w11345 & w11442 ;
  assign w11808 = w11443 ^ w11807 ;
  assign w11809 = ~w11562 & w11808 ;
  assign w11810 = ( w11337 & w11560 ) | ( w11337 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11811 = ~w11561 & w11810 ;
  assign w11812 = w11809 | w11811 ;
  assign w11813 = ~\pi077 & w11812 ;
  assign w11814 = ~w11352 & w11439 ;
  assign w11815 = w11440 ^ w11814 ;
  assign w11816 = ~w11562 & w11815 ;
  assign w11817 = ( w11344 & w11560 ) | ( w11344 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11818 = ~w11561 & w11817 ;
  assign w11819 = w11816 | w11818 ;
  assign w11820 = ~\pi076 & w11819 ;
  assign w11821 = ~w11359 & w11436 ;
  assign w11822 = w11437 ^ w11821 ;
  assign w11823 = ~w11562 & w11822 ;
  assign w11824 = ( w11351 & w11560 ) | ( w11351 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11825 = ~w11561 & w11824 ;
  assign w11826 = w11823 | w11825 ;
  assign w11827 = ~\pi075 & w11826 ;
  assign w11828 = ~w11366 & w11433 ;
  assign w11829 = w11434 ^ w11828 ;
  assign w11830 = ~w11562 & w11829 ;
  assign w11831 = ( w11358 & w11560 ) | ( w11358 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11832 = ~w11561 & w11831 ;
  assign w11833 = w11830 | w11832 ;
  assign w11834 = ~\pi074 & w11833 ;
  assign w11835 = ~w11373 & w11430 ;
  assign w11836 = w11431 ^ w11835 ;
  assign w11837 = ~w11562 & w11836 ;
  assign w11838 = ( w11365 & w11560 ) | ( w11365 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11839 = ~w11561 & w11838 ;
  assign w11840 = w11837 | w11839 ;
  assign w11841 = ~\pi073 & w11840 ;
  assign w11842 = ~w11380 & w11427 ;
  assign w11843 = w11428 ^ w11842 ;
  assign w11844 = ~w11562 & w11843 ;
  assign w11845 = ( w11372 & w11560 ) | ( w11372 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11846 = ~w11561 & w11845 ;
  assign w11847 = w11844 | w11846 ;
  assign w11848 = ~\pi072 & w11847 ;
  assign w11849 = ~w11387 & w11424 ;
  assign w11850 = w11425 ^ w11849 ;
  assign w11851 = ~w11562 & w11850 ;
  assign w11852 = ( w11379 & w11560 ) | ( w11379 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11853 = ~w11561 & w11852 ;
  assign w11854 = w11851 | w11853 ;
  assign w11855 = ~\pi071 & w11854 ;
  assign w11856 = ~w11394 & w11421 ;
  assign w11857 = w11422 ^ w11856 ;
  assign w11858 = ~w11562 & w11857 ;
  assign w11859 = ( w11386 & w11560 ) | ( w11386 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11860 = ~w11561 & w11859 ;
  assign w11861 = w11858 | w11860 ;
  assign w11862 = ~\pi070 & w11861 ;
  assign w11863 = ~w11402 & w11418 ;
  assign w11864 = w11419 ^ w11863 ;
  assign w11865 = ~w11562 & w11864 ;
  assign w11866 = ( w11393 & w11560 ) | ( w11393 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11867 = ~w11561 & w11866 ;
  assign w11868 = w11865 | w11867 ;
  assign w11869 = ~\pi069 & w11868 ;
  assign w11870 = ~w11407 & w11415 ;
  assign w11871 = w11416 ^ w11870 ;
  assign w11872 = ~w11562 & w11871 ;
  assign w11873 = ( w11401 & w11560 ) | ( w11401 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11874 = ~w11561 & w11873 ;
  assign w11875 = w11872 | w11874 ;
  assign w11876 = ~\pi068 & w11875 ;
  assign w11877 = ~\pi016 & \pi064 ;
  assign w11878 = ( \pi065 & ~w11412 ) | ( \pi065 & w11877 ) | ( ~w11412 & w11877 ) ;
  assign w11879 = w11410 ^ w11878 ;
  assign w11880 = ~w11562 & w11879 ;
  assign w11881 = ( w11406 & w11560 ) | ( w11406 & w11561 ) | ( w11560 & w11561 ) ;
  assign w11882 = ~w11561 & w11881 ;
  assign w11883 = w11880 | w11882 ;
  assign w11884 = ~\pi067 & w11883 ;
  assign w11885 = \pi017 ^ \pi065 ;
  assign w11886 = \pi016 ^ w11093 ;
  assign w11887 = ( \pi064 & w11562 ) | ( \pi064 & w11886 ) | ( w11562 & w11886 ) ;
  assign w11888 = w11885 ^ w11887 ;
  assign w11889 = ~w11562 & w11888 ;
  assign w11890 = w11412 & w11562 ;
  assign w11891 = w11889 | w11890 ;
  assign w11892 = ~\pi066 & w11891 ;
  assign w11893 = \pi066 ^ w11891 ;
  assign w11894 = \pi064 & ~w11562 ;
  assign w11895 = \pi016 ^ w11894 ;
  assign w11896 = ( ~\pi015 & \pi064 ) | ( ~\pi015 & w11893 ) | ( \pi064 & w11893 ) ;
  assign w11897 = ( \pi065 & ~w11895 ) | ( \pi065 & w11896 ) | ( ~w11895 & w11896 ) ;
  assign w11898 = w11893 | w11897 ;
  assign w11899 = \pi067 ^ w11883 ;
  assign w11900 = ( ~w11892 & w11898 ) | ( ~w11892 & w11899 ) | ( w11898 & w11899 ) ;
  assign w11901 = w11899 | w11900 ;
  assign w11902 = \pi068 ^ w11875 ;
  assign w11903 = ( ~w11884 & w11901 ) | ( ~w11884 & w11902 ) | ( w11901 & w11902 ) ;
  assign w11904 = w11902 | w11903 ;
  assign w11905 = \pi069 ^ w11868 ;
  assign w11906 = ( ~w11876 & w11904 ) | ( ~w11876 & w11905 ) | ( w11904 & w11905 ) ;
  assign w11907 = w11905 | w11906 ;
  assign w11908 = \pi070 ^ w11861 ;
  assign w11909 = ( ~w11869 & w11907 ) | ( ~w11869 & w11908 ) | ( w11907 & w11908 ) ;
  assign w11910 = w11908 | w11909 ;
  assign w11911 = \pi071 ^ w11854 ;
  assign w11912 = ( ~w11862 & w11910 ) | ( ~w11862 & w11911 ) | ( w11910 & w11911 ) ;
  assign w11913 = w11911 | w11912 ;
  assign w11914 = \pi072 ^ w11847 ;
  assign w11915 = ( ~w11855 & w11913 ) | ( ~w11855 & w11914 ) | ( w11913 & w11914 ) ;
  assign w11916 = w11914 | w11915 ;
  assign w11917 = \pi073 ^ w11840 ;
  assign w11918 = ( ~w11848 & w11916 ) | ( ~w11848 & w11917 ) | ( w11916 & w11917 ) ;
  assign w11919 = w11917 | w11918 ;
  assign w11920 = \pi074 ^ w11833 ;
  assign w11921 = ( ~w11841 & w11919 ) | ( ~w11841 & w11920 ) | ( w11919 & w11920 ) ;
  assign w11922 = w11920 | w11921 ;
  assign w11923 = \pi075 ^ w11826 ;
  assign w11924 = ( ~w11834 & w11922 ) | ( ~w11834 & w11923 ) | ( w11922 & w11923 ) ;
  assign w11925 = w11923 | w11924 ;
  assign w11926 = \pi076 ^ w11819 ;
  assign w11927 = ( ~w11827 & w11925 ) | ( ~w11827 & w11926 ) | ( w11925 & w11926 ) ;
  assign w11928 = w11926 | w11927 ;
  assign w11929 = \pi077 ^ w11812 ;
  assign w11930 = ( ~w11820 & w11928 ) | ( ~w11820 & w11929 ) | ( w11928 & w11929 ) ;
  assign w11931 = w11929 | w11930 ;
  assign w11932 = \pi078 ^ w11805 ;
  assign w11933 = ( ~w11813 & w11931 ) | ( ~w11813 & w11932 ) | ( w11931 & w11932 ) ;
  assign w11934 = w11932 | w11933 ;
  assign w11935 = \pi079 ^ w11798 ;
  assign w11936 = ( ~w11806 & w11934 ) | ( ~w11806 & w11935 ) | ( w11934 & w11935 ) ;
  assign w11937 = w11935 | w11936 ;
  assign w11938 = \pi080 ^ w11791 ;
  assign w11939 = ( ~w11799 & w11937 ) | ( ~w11799 & w11938 ) | ( w11937 & w11938 ) ;
  assign w11940 = w11938 | w11939 ;
  assign w11941 = \pi081 ^ w11784 ;
  assign w11942 = ( ~w11792 & w11940 ) | ( ~w11792 & w11941 ) | ( w11940 & w11941 ) ;
  assign w11943 = w11941 | w11942 ;
  assign w11944 = \pi082 ^ w11777 ;
  assign w11945 = ( ~w11785 & w11943 ) | ( ~w11785 & w11944 ) | ( w11943 & w11944 ) ;
  assign w11946 = w11944 | w11945 ;
  assign w11947 = \pi083 ^ w11770 ;
  assign w11948 = ( ~w11778 & w11946 ) | ( ~w11778 & w11947 ) | ( w11946 & w11947 ) ;
  assign w11949 = w11947 | w11948 ;
  assign w11950 = \pi084 ^ w11763 ;
  assign w11951 = ( ~w11771 & w11949 ) | ( ~w11771 & w11950 ) | ( w11949 & w11950 ) ;
  assign w11952 = w11950 | w11951 ;
  assign w11953 = \pi085 ^ w11756 ;
  assign w11954 = ( ~w11764 & w11952 ) | ( ~w11764 & w11953 ) | ( w11952 & w11953 ) ;
  assign w11955 = w11953 | w11954 ;
  assign w11956 = \pi086 ^ w11749 ;
  assign w11957 = ( ~w11757 & w11955 ) | ( ~w11757 & w11956 ) | ( w11955 & w11956 ) ;
  assign w11958 = w11956 | w11957 ;
  assign w11959 = \pi087 ^ w11742 ;
  assign w11960 = ( ~w11750 & w11958 ) | ( ~w11750 & w11959 ) | ( w11958 & w11959 ) ;
  assign w11961 = w11959 | w11960 ;
  assign w11962 = \pi088 ^ w11735 ;
  assign w11963 = ( ~w11743 & w11961 ) | ( ~w11743 & w11962 ) | ( w11961 & w11962 ) ;
  assign w11964 = w11962 | w11963 ;
  assign w11965 = \pi089 ^ w11728 ;
  assign w11966 = ( ~w11736 & w11964 ) | ( ~w11736 & w11965 ) | ( w11964 & w11965 ) ;
  assign w11967 = w11965 | w11966 ;
  assign w11968 = \pi090 ^ w11721 ;
  assign w11969 = ( ~w11729 & w11967 ) | ( ~w11729 & w11968 ) | ( w11967 & w11968 ) ;
  assign w11970 = w11968 | w11969 ;
  assign w11971 = \pi091 ^ w11714 ;
  assign w11972 = ( ~w11722 & w11970 ) | ( ~w11722 & w11971 ) | ( w11970 & w11971 ) ;
  assign w11973 = w11971 | w11972 ;
  assign w11974 = \pi092 ^ w11707 ;
  assign w11975 = ( ~w11715 & w11973 ) | ( ~w11715 & w11974 ) | ( w11973 & w11974 ) ;
  assign w11976 = w11974 | w11975 ;
  assign w11977 = \pi093 ^ w11700 ;
  assign w11978 = ( ~w11708 & w11976 ) | ( ~w11708 & w11977 ) | ( w11976 & w11977 ) ;
  assign w11979 = w11977 | w11978 ;
  assign w11980 = \pi094 ^ w11693 ;
  assign w11981 = ( ~w11701 & w11979 ) | ( ~w11701 & w11980 ) | ( w11979 & w11980 ) ;
  assign w11982 = w11980 | w11981 ;
  assign w11983 = \pi095 ^ w11686 ;
  assign w11984 = ( ~w11694 & w11982 ) | ( ~w11694 & w11983 ) | ( w11982 & w11983 ) ;
  assign w11985 = w11983 | w11984 ;
  assign w11986 = \pi096 ^ w11679 ;
  assign w11987 = ( ~w11687 & w11985 ) | ( ~w11687 & w11986 ) | ( w11985 & w11986 ) ;
  assign w11988 = w11986 | w11987 ;
  assign w11989 = \pi097 ^ w11672 ;
  assign w11990 = ( ~w11680 & w11988 ) | ( ~w11680 & w11989 ) | ( w11988 & w11989 ) ;
  assign w11991 = w11989 | w11990 ;
  assign w11992 = \pi098 ^ w11665 ;
  assign w11993 = ( ~w11673 & w11991 ) | ( ~w11673 & w11992 ) | ( w11991 & w11992 ) ;
  assign w11994 = w11992 | w11993 ;
  assign w11995 = \pi099 ^ w11658 ;
  assign w11996 = ( ~w11666 & w11994 ) | ( ~w11666 & w11995 ) | ( w11994 & w11995 ) ;
  assign w11997 = w11995 | w11996 ;
  assign w11998 = \pi100 ^ w11651 ;
  assign w11999 = ( ~w11659 & w11997 ) | ( ~w11659 & w11998 ) | ( w11997 & w11998 ) ;
  assign w12000 = w11998 | w11999 ;
  assign w12001 = \pi101 ^ w11644 ;
  assign w12002 = ( ~w11652 & w12000 ) | ( ~w11652 & w12001 ) | ( w12000 & w12001 ) ;
  assign w12003 = w12001 | w12002 ;
  assign w12004 = \pi102 ^ w11637 ;
  assign w12005 = ( ~w11645 & w12003 ) | ( ~w11645 & w12004 ) | ( w12003 & w12004 ) ;
  assign w12006 = w12004 | w12005 ;
  assign w12007 = \pi103 ^ w11630 ;
  assign w12008 = ( ~w11638 & w12006 ) | ( ~w11638 & w12007 ) | ( w12006 & w12007 ) ;
  assign w12009 = w12007 | w12008 ;
  assign w12010 = \pi104 ^ w11623 ;
  assign w12011 = ( ~w11631 & w12009 ) | ( ~w11631 & w12010 ) | ( w12009 & w12010 ) ;
  assign w12012 = w12010 | w12011 ;
  assign w12013 = \pi105 ^ w11616 ;
  assign w12014 = ( ~w11624 & w12012 ) | ( ~w11624 & w12013 ) | ( w12012 & w12013 ) ;
  assign w12015 = w12013 | w12014 ;
  assign w12016 = \pi106 ^ w11609 ;
  assign w12017 = ( ~w11617 & w12015 ) | ( ~w11617 & w12016 ) | ( w12015 & w12016 ) ;
  assign w12018 = w12016 | w12017 ;
  assign w12019 = \pi107 ^ w11602 ;
  assign w12020 = ( ~w11610 & w12018 ) | ( ~w11610 & w12019 ) | ( w12018 & w12019 ) ;
  assign w12021 = w12019 | w12020 ;
  assign w12022 = \pi108 ^ w11595 ;
  assign w12023 = ( ~w11603 & w12021 ) | ( ~w11603 & w12022 ) | ( w12021 & w12022 ) ;
  assign w12024 = w12022 | w12023 ;
  assign w12025 = \pi109 ^ w11588 ;
  assign w12026 = ( ~w11596 & w12024 ) | ( ~w11596 & w12025 ) | ( w12024 & w12025 ) ;
  assign w12027 = w12025 | w12026 ;
  assign w12028 = \pi110 ^ w11581 ;
  assign w12029 = ( ~w11589 & w12027 ) | ( ~w11589 & w12028 ) | ( w12027 & w12028 ) ;
  assign w12030 = w12028 | w12029 ;
  assign w12031 = \pi111 ^ w11568 ;
  assign w12032 = ( ~w11582 & w12030 ) | ( ~w11582 & w12031 ) | ( w12030 & w12031 ) ;
  assign w12033 = w12031 | w12032 ;
  assign w12034 = \pi112 ^ w11574 ;
  assign w12035 = w11575 & ~w12034 ;
  assign w12036 = ( w12033 & w12034 ) | ( w12033 & ~w12035 ) | ( w12034 & ~w12035 ) ;
  assign w12037 = ~\pi112 & w11574 ;
  assign w12038 = w12036 & ~w12037 ;
  assign w12039 = w275 | w12038 ;
  assign w12040 = w11568 & w12039 ;
  assign w12041 = ~w11582 & w12030 ;
  assign w12042 = w12031 ^ w12041 ;
  assign w12043 = ~w12039 & w12042 ;
  assign w12044 = w12040 | w12043 ;
  assign w12045 = ~\pi112 & w12044 ;
  assign w12046 = w11581 & w12039 ;
  assign w12047 = ~w11589 & w12027 ;
  assign w12048 = w12028 ^ w12047 ;
  assign w12049 = ~w12039 & w12048 ;
  assign w12050 = w12046 | w12049 ;
  assign w12051 = ~\pi111 & w12050 ;
  assign w12052 = w11588 & w12039 ;
  assign w12053 = ~w11596 & w12024 ;
  assign w12054 = w12025 ^ w12053 ;
  assign w12055 = ~w12039 & w12054 ;
  assign w12056 = w12052 | w12055 ;
  assign w12057 = ~\pi110 & w12056 ;
  assign w12058 = w11595 & w12039 ;
  assign w12059 = ~w11603 & w12021 ;
  assign w12060 = w12022 ^ w12059 ;
  assign w12061 = ~w12039 & w12060 ;
  assign w12062 = w12058 | w12061 ;
  assign w12063 = ~\pi109 & w12062 ;
  assign w12064 = w11602 & w12039 ;
  assign w12065 = ~w11610 & w12018 ;
  assign w12066 = w12019 ^ w12065 ;
  assign w12067 = ~w12039 & w12066 ;
  assign w12068 = w12064 | w12067 ;
  assign w12069 = ~\pi108 & w12068 ;
  assign w12070 = w11609 & w12039 ;
  assign w12071 = ~w11617 & w12015 ;
  assign w12072 = w12016 ^ w12071 ;
  assign w12073 = ~w12039 & w12072 ;
  assign w12074 = w12070 | w12073 ;
  assign w12075 = ~\pi107 & w12074 ;
  assign w12076 = w11616 & w12039 ;
  assign w12077 = ~w11624 & w12012 ;
  assign w12078 = w12013 ^ w12077 ;
  assign w12079 = ~w12039 & w12078 ;
  assign w12080 = w12076 | w12079 ;
  assign w12081 = ~\pi106 & w12080 ;
  assign w12082 = w11623 & w12039 ;
  assign w12083 = ~w11631 & w12009 ;
  assign w12084 = w12010 ^ w12083 ;
  assign w12085 = ~w12039 & w12084 ;
  assign w12086 = w12082 | w12085 ;
  assign w12087 = ~\pi105 & w12086 ;
  assign w12088 = w11630 & w12039 ;
  assign w12089 = ~w11638 & w12006 ;
  assign w12090 = w12007 ^ w12089 ;
  assign w12091 = ~w12039 & w12090 ;
  assign w12092 = w12088 | w12091 ;
  assign w12093 = ~\pi104 & w12092 ;
  assign w12094 = w11637 & w12039 ;
  assign w12095 = ~w11645 & w12003 ;
  assign w12096 = w12004 ^ w12095 ;
  assign w12097 = ~w12039 & w12096 ;
  assign w12098 = w12094 | w12097 ;
  assign w12099 = ~\pi103 & w12098 ;
  assign w12100 = w11644 & w12039 ;
  assign w12101 = ~w11652 & w12000 ;
  assign w12102 = w12001 ^ w12101 ;
  assign w12103 = ~w12039 & w12102 ;
  assign w12104 = w12100 | w12103 ;
  assign w12105 = ~\pi102 & w12104 ;
  assign w12106 = w11651 & w12039 ;
  assign w12107 = ~w11659 & w11997 ;
  assign w12108 = w11998 ^ w12107 ;
  assign w12109 = ~w12039 & w12108 ;
  assign w12110 = w12106 | w12109 ;
  assign w12111 = ~\pi101 & w12110 ;
  assign w12112 = w11658 & w12039 ;
  assign w12113 = ~w11666 & w11994 ;
  assign w12114 = w11995 ^ w12113 ;
  assign w12115 = ~w12039 & w12114 ;
  assign w12116 = w12112 | w12115 ;
  assign w12117 = ~\pi100 & w12116 ;
  assign w12118 = w11665 & w12039 ;
  assign w12119 = ~w11673 & w11991 ;
  assign w12120 = w11992 ^ w12119 ;
  assign w12121 = ~w12039 & w12120 ;
  assign w12122 = w12118 | w12121 ;
  assign w12123 = ~\pi099 & w12122 ;
  assign w12124 = w11672 & w12039 ;
  assign w12125 = ~w11680 & w11988 ;
  assign w12126 = w11989 ^ w12125 ;
  assign w12127 = ~w12039 & w12126 ;
  assign w12128 = w12124 | w12127 ;
  assign w12129 = ~\pi098 & w12128 ;
  assign w12130 = w11679 & w12039 ;
  assign w12131 = ~w11687 & w11985 ;
  assign w12132 = w11986 ^ w12131 ;
  assign w12133 = ~w12039 & w12132 ;
  assign w12134 = w12130 | w12133 ;
  assign w12135 = ~\pi097 & w12134 ;
  assign w12136 = w11686 & w12039 ;
  assign w12137 = ~w11694 & w11982 ;
  assign w12138 = w11983 ^ w12137 ;
  assign w12139 = ~w12039 & w12138 ;
  assign w12140 = w12136 | w12139 ;
  assign w12141 = ~\pi096 & w12140 ;
  assign w12142 = w11693 & w12039 ;
  assign w12143 = ~w11701 & w11979 ;
  assign w12144 = w11980 ^ w12143 ;
  assign w12145 = ~w12039 & w12144 ;
  assign w12146 = w12142 | w12145 ;
  assign w12147 = ~\pi095 & w12146 ;
  assign w12148 = w11700 & w12039 ;
  assign w12149 = ~w11708 & w11976 ;
  assign w12150 = w11977 ^ w12149 ;
  assign w12151 = ~w12039 & w12150 ;
  assign w12152 = w12148 | w12151 ;
  assign w12153 = ~\pi094 & w12152 ;
  assign w12154 = w11707 & w12039 ;
  assign w12155 = ~w11715 & w11973 ;
  assign w12156 = w11974 ^ w12155 ;
  assign w12157 = ~w12039 & w12156 ;
  assign w12158 = w12154 | w12157 ;
  assign w12159 = ~\pi093 & w12158 ;
  assign w12160 = w11714 & w12039 ;
  assign w12161 = ~w11722 & w11970 ;
  assign w12162 = w11971 ^ w12161 ;
  assign w12163 = ~w12039 & w12162 ;
  assign w12164 = w12160 | w12163 ;
  assign w12165 = ~\pi092 & w12164 ;
  assign w12166 = w11721 & w12039 ;
  assign w12167 = ~w11729 & w11967 ;
  assign w12168 = w11968 ^ w12167 ;
  assign w12169 = ~w12039 & w12168 ;
  assign w12170 = w12166 | w12169 ;
  assign w12171 = ~\pi091 & w12170 ;
  assign w12172 = w11728 & w12039 ;
  assign w12173 = ~w11736 & w11964 ;
  assign w12174 = w11965 ^ w12173 ;
  assign w12175 = ~w12039 & w12174 ;
  assign w12176 = w12172 | w12175 ;
  assign w12177 = ~\pi090 & w12176 ;
  assign w12178 = w11735 & w12039 ;
  assign w12179 = ~w11743 & w11961 ;
  assign w12180 = w11962 ^ w12179 ;
  assign w12181 = ~w12039 & w12180 ;
  assign w12182 = w12178 | w12181 ;
  assign w12183 = ~\pi089 & w12182 ;
  assign w12184 = w11742 & w12039 ;
  assign w12185 = ~w11750 & w11958 ;
  assign w12186 = w11959 ^ w12185 ;
  assign w12187 = ~w12039 & w12186 ;
  assign w12188 = w12184 | w12187 ;
  assign w12189 = ~\pi088 & w12188 ;
  assign w12190 = w11749 & w12039 ;
  assign w12191 = ~w11757 & w11955 ;
  assign w12192 = w11956 ^ w12191 ;
  assign w12193 = ~w12039 & w12192 ;
  assign w12194 = w12190 | w12193 ;
  assign w12195 = ~\pi087 & w12194 ;
  assign w12196 = w11756 & w12039 ;
  assign w12197 = ~w11764 & w11952 ;
  assign w12198 = w11953 ^ w12197 ;
  assign w12199 = ~w12039 & w12198 ;
  assign w12200 = w12196 | w12199 ;
  assign w12201 = ~\pi086 & w12200 ;
  assign w12202 = w11763 & w12039 ;
  assign w12203 = ~w11771 & w11949 ;
  assign w12204 = w11950 ^ w12203 ;
  assign w12205 = ~w12039 & w12204 ;
  assign w12206 = w12202 | w12205 ;
  assign w12207 = ~\pi085 & w12206 ;
  assign w12208 = w11770 & w12039 ;
  assign w12209 = ~w11778 & w11946 ;
  assign w12210 = w11947 ^ w12209 ;
  assign w12211 = ~w12039 & w12210 ;
  assign w12212 = w12208 | w12211 ;
  assign w12213 = ~\pi084 & w12212 ;
  assign w12214 = w11777 & w12039 ;
  assign w12215 = ~w11785 & w11943 ;
  assign w12216 = w11944 ^ w12215 ;
  assign w12217 = ~w12039 & w12216 ;
  assign w12218 = w12214 | w12217 ;
  assign w12219 = ~\pi083 & w12218 ;
  assign w12220 = w11784 & w12039 ;
  assign w12221 = ~w11792 & w11940 ;
  assign w12222 = w11941 ^ w12221 ;
  assign w12223 = ~w12039 & w12222 ;
  assign w12224 = w12220 | w12223 ;
  assign w12225 = ~\pi082 & w12224 ;
  assign w12226 = w11791 & w12039 ;
  assign w12227 = ~w11799 & w11937 ;
  assign w12228 = w11938 ^ w12227 ;
  assign w12229 = ~w12039 & w12228 ;
  assign w12230 = w12226 | w12229 ;
  assign w12231 = ~\pi081 & w12230 ;
  assign w12232 = w11798 & w12039 ;
  assign w12233 = ~w11806 & w11934 ;
  assign w12234 = w11935 ^ w12233 ;
  assign w12235 = ~w12039 & w12234 ;
  assign w12236 = w12232 | w12235 ;
  assign w12237 = ~\pi080 & w12236 ;
  assign w12238 = w11805 & w12039 ;
  assign w12239 = ~w11813 & w11931 ;
  assign w12240 = w11932 ^ w12239 ;
  assign w12241 = ~w12039 & w12240 ;
  assign w12242 = w12238 | w12241 ;
  assign w12243 = ~\pi079 & w12242 ;
  assign w12244 = w11812 & w12039 ;
  assign w12245 = ~w11820 & w11928 ;
  assign w12246 = w11929 ^ w12245 ;
  assign w12247 = ~w12039 & w12246 ;
  assign w12248 = w12244 | w12247 ;
  assign w12249 = ~\pi078 & w12248 ;
  assign w12250 = w11819 & w12039 ;
  assign w12251 = ~w11827 & w11925 ;
  assign w12252 = w11926 ^ w12251 ;
  assign w12253 = ~w12039 & w12252 ;
  assign w12254 = w12250 | w12253 ;
  assign w12255 = ~\pi077 & w12254 ;
  assign w12256 = w11826 & w12039 ;
  assign w12257 = ~w11834 & w11922 ;
  assign w12258 = w11923 ^ w12257 ;
  assign w12259 = ~w12039 & w12258 ;
  assign w12260 = w12256 | w12259 ;
  assign w12261 = ~\pi076 & w12260 ;
  assign w12262 = w11833 & w12039 ;
  assign w12263 = ~w11841 & w11919 ;
  assign w12264 = w11920 ^ w12263 ;
  assign w12265 = ~w12039 & w12264 ;
  assign w12266 = w12262 | w12265 ;
  assign w12267 = ~\pi075 & w12266 ;
  assign w12268 = w11840 & w12039 ;
  assign w12269 = ~w11848 & w11916 ;
  assign w12270 = w11917 ^ w12269 ;
  assign w12271 = ~w12039 & w12270 ;
  assign w12272 = w12268 | w12271 ;
  assign w12273 = ~\pi074 & w12272 ;
  assign w12274 = w11847 & w12039 ;
  assign w12275 = ~w11855 & w11913 ;
  assign w12276 = w11914 ^ w12275 ;
  assign w12277 = ~w12039 & w12276 ;
  assign w12278 = w12274 | w12277 ;
  assign w12279 = ~\pi073 & w12278 ;
  assign w12280 = w11854 & w12039 ;
  assign w12281 = ~w11862 & w11910 ;
  assign w12282 = w11911 ^ w12281 ;
  assign w12283 = ~w12039 & w12282 ;
  assign w12284 = w12280 | w12283 ;
  assign w12285 = ~\pi072 & w12284 ;
  assign w12286 = w11861 & w12039 ;
  assign w12287 = ~w11869 & w11907 ;
  assign w12288 = w11908 ^ w12287 ;
  assign w12289 = ~w12039 & w12288 ;
  assign w12290 = w12286 | w12289 ;
  assign w12291 = ~\pi071 & w12290 ;
  assign w12292 = w11868 & w12039 ;
  assign w12293 = ~w11876 & w11904 ;
  assign w12294 = w11905 ^ w12293 ;
  assign w12295 = ~w12039 & w12294 ;
  assign w12296 = w12292 | w12295 ;
  assign w12297 = ~\pi070 & w12296 ;
  assign w12298 = w11875 & w12039 ;
  assign w12299 = ~w11884 & w11901 ;
  assign w12300 = w11902 ^ w12299 ;
  assign w12301 = ~w12039 & w12300 ;
  assign w12302 = w12298 | w12301 ;
  assign w12303 = ~\pi069 & w12302 ;
  assign w12304 = w11883 & w12039 ;
  assign w12305 = ~w11892 & w11898 ;
  assign w12306 = w11899 ^ w12305 ;
  assign w12307 = ~w12039 & w12306 ;
  assign w12308 = w12304 | w12307 ;
  assign w12309 = ~\pi068 & w12308 ;
  assign w12310 = ~\pi015 & \pi064 ;
  assign w12311 = ( \pi065 & ~w11895 ) | ( \pi065 & w12310 ) | ( ~w11895 & w12310 ) ;
  assign w12312 = w11893 ^ w12311 ;
  assign w12313 = ( w275 & w12038 ) | ( w275 & w12312 ) | ( w12038 & w12312 ) ;
  assign w12314 = w12312 & ~w12313 ;
  assign w12315 = ( w11891 & w12039 ) | ( w11891 & w12314 ) | ( w12039 & w12314 ) ;
  assign w12316 = w12314 | w12315 ;
  assign w12317 = ~\pi067 & w12316 ;
  assign w12318 = \pi016 ^ \pi065 ;
  assign w12319 = \pi015 ^ w11562 ;
  assign w12320 = ( \pi064 & w275 ) | ( \pi064 & w12319 ) | ( w275 & w12319 ) ;
  assign w12321 = w12318 ^ w12320 ;
  assign w12322 = ~w275 & w12321 ;
  assign w12323 = ~w12038 & w12322 ;
  assign w12324 = ( ~\pi064 & w11562 ) | ( ~\pi064 & w12039 ) | ( w11562 & w12039 ) ;
  assign w12325 = \pi016 ^ w12324 ;
  assign w12326 = w12039 & ~w12325 ;
  assign w12327 = w12323 | w12326 ;
  assign w12328 = ~\pi066 & w12327 ;
  assign w12329 = ( \pi064 & ~\pi113 ) | ( \pi064 & \pi114 ) | ( ~\pi113 & \pi114 ) ;
  assign w12330 = w153 | w199 ;
  assign w12331 = ( \pi114 & \pi115 ) | ( \pi114 & ~w153 ) | ( \pi115 & ~w153 ) ;
  assign w12332 = w12330 | w12331 ;
  assign w12333 = w12329 & ~w12332 ;
  assign w12334 = ( \pi015 & w12038 ) | ( \pi015 & ~w12333 ) | ( w12038 & ~w12333 ) ;
  assign w12335 = \pi015 & w12334 ;
  assign w12336 = ~w448 & w12310 ;
  assign w12337 = ( w267 & ~w448 ) | ( w267 & w12038 ) | ( ~w448 & w12038 ) ;
  assign w12338 = w12336 & ~w12337 ;
  assign w12339 = ~\pi014 & \pi064 ;
  assign w12340 = w12039 | w12323 ;
  assign w12341 = ( w11895 & w12323 ) | ( w11895 & w12340 ) | ( w12323 & w12340 ) ;
  assign w12342 = \pi066 ^ w12341 ;
  assign w12343 = w12335 | w12338 ;
  assign w12344 = ( \pi065 & w12339 ) | ( \pi065 & ~w12343 ) | ( w12339 & ~w12343 ) ;
  assign w12345 = w12342 | w12344 ;
  assign w12346 = ~w11891 & w12039 ;
  assign w12347 = ( w12039 & w12314 ) | ( w12039 & ~w12346 ) | ( w12314 & ~w12346 ) ;
  assign w12348 = \pi067 ^ w12347 ;
  assign w12349 = ( ~w12328 & w12345 ) | ( ~w12328 & w12348 ) | ( w12345 & w12348 ) ;
  assign w12350 = w12348 | w12349 ;
  assign w12351 = \pi068 ^ w12308 ;
  assign w12352 = ( ~w12317 & w12350 ) | ( ~w12317 & w12351 ) | ( w12350 & w12351 ) ;
  assign w12353 = w12351 | w12352 ;
  assign w12354 = \pi069 ^ w12302 ;
  assign w12355 = ( ~w12309 & w12353 ) | ( ~w12309 & w12354 ) | ( w12353 & w12354 ) ;
  assign w12356 = w12354 | w12355 ;
  assign w12357 = \pi070 ^ w12296 ;
  assign w12358 = ( ~w12303 & w12356 ) | ( ~w12303 & w12357 ) | ( w12356 & w12357 ) ;
  assign w12359 = w12357 | w12358 ;
  assign w12360 = \pi071 ^ w12290 ;
  assign w12361 = ( ~w12297 & w12359 ) | ( ~w12297 & w12360 ) | ( w12359 & w12360 ) ;
  assign w12362 = w12360 | w12361 ;
  assign w12363 = \pi072 ^ w12284 ;
  assign w12364 = ( ~w12291 & w12362 ) | ( ~w12291 & w12363 ) | ( w12362 & w12363 ) ;
  assign w12365 = w12363 | w12364 ;
  assign w12366 = \pi073 ^ w12278 ;
  assign w12367 = ( ~w12285 & w12365 ) | ( ~w12285 & w12366 ) | ( w12365 & w12366 ) ;
  assign w12368 = w12366 | w12367 ;
  assign w12369 = \pi074 ^ w12272 ;
  assign w12370 = ( ~w12279 & w12368 ) | ( ~w12279 & w12369 ) | ( w12368 & w12369 ) ;
  assign w12371 = w12369 | w12370 ;
  assign w12372 = \pi075 ^ w12266 ;
  assign w12373 = ( ~w12273 & w12371 ) | ( ~w12273 & w12372 ) | ( w12371 & w12372 ) ;
  assign w12374 = w12372 | w12373 ;
  assign w12375 = \pi076 ^ w12260 ;
  assign w12376 = ( ~w12267 & w12374 ) | ( ~w12267 & w12375 ) | ( w12374 & w12375 ) ;
  assign w12377 = w12375 | w12376 ;
  assign w12378 = \pi077 ^ w12254 ;
  assign w12379 = ( ~w12261 & w12377 ) | ( ~w12261 & w12378 ) | ( w12377 & w12378 ) ;
  assign w12380 = w12378 | w12379 ;
  assign w12381 = \pi078 ^ w12248 ;
  assign w12382 = ( ~w12255 & w12380 ) | ( ~w12255 & w12381 ) | ( w12380 & w12381 ) ;
  assign w12383 = w12381 | w12382 ;
  assign w12384 = \pi079 ^ w12242 ;
  assign w12385 = ( ~w12249 & w12383 ) | ( ~w12249 & w12384 ) | ( w12383 & w12384 ) ;
  assign w12386 = w12384 | w12385 ;
  assign w12387 = \pi080 ^ w12236 ;
  assign w12388 = ( ~w12243 & w12386 ) | ( ~w12243 & w12387 ) | ( w12386 & w12387 ) ;
  assign w12389 = w12387 | w12388 ;
  assign w12390 = \pi081 ^ w12230 ;
  assign w12391 = ( ~w12237 & w12389 ) | ( ~w12237 & w12390 ) | ( w12389 & w12390 ) ;
  assign w12392 = w12390 | w12391 ;
  assign w12393 = \pi082 ^ w12224 ;
  assign w12394 = ( ~w12231 & w12392 ) | ( ~w12231 & w12393 ) | ( w12392 & w12393 ) ;
  assign w12395 = w12393 | w12394 ;
  assign w12396 = \pi083 ^ w12218 ;
  assign w12397 = ( ~w12225 & w12395 ) | ( ~w12225 & w12396 ) | ( w12395 & w12396 ) ;
  assign w12398 = w12396 | w12397 ;
  assign w12399 = \pi084 ^ w12212 ;
  assign w12400 = ( ~w12219 & w12398 ) | ( ~w12219 & w12399 ) | ( w12398 & w12399 ) ;
  assign w12401 = w12399 | w12400 ;
  assign w12402 = \pi085 ^ w12206 ;
  assign w12403 = ( ~w12213 & w12401 ) | ( ~w12213 & w12402 ) | ( w12401 & w12402 ) ;
  assign w12404 = w12402 | w12403 ;
  assign w12405 = \pi086 ^ w12200 ;
  assign w12406 = ( ~w12207 & w12404 ) | ( ~w12207 & w12405 ) | ( w12404 & w12405 ) ;
  assign w12407 = w12405 | w12406 ;
  assign w12408 = \pi087 ^ w12194 ;
  assign w12409 = ( ~w12201 & w12407 ) | ( ~w12201 & w12408 ) | ( w12407 & w12408 ) ;
  assign w12410 = w12408 | w12409 ;
  assign w12411 = \pi088 ^ w12188 ;
  assign w12412 = ( ~w12195 & w12410 ) | ( ~w12195 & w12411 ) | ( w12410 & w12411 ) ;
  assign w12413 = w12411 | w12412 ;
  assign w12414 = \pi089 ^ w12182 ;
  assign w12415 = ( ~w12189 & w12413 ) | ( ~w12189 & w12414 ) | ( w12413 & w12414 ) ;
  assign w12416 = w12414 | w12415 ;
  assign w12417 = \pi090 ^ w12176 ;
  assign w12418 = ( ~w12183 & w12416 ) | ( ~w12183 & w12417 ) | ( w12416 & w12417 ) ;
  assign w12419 = w12417 | w12418 ;
  assign w12420 = \pi091 ^ w12170 ;
  assign w12421 = ( ~w12177 & w12419 ) | ( ~w12177 & w12420 ) | ( w12419 & w12420 ) ;
  assign w12422 = w12420 | w12421 ;
  assign w12423 = \pi092 ^ w12164 ;
  assign w12424 = ( ~w12171 & w12422 ) | ( ~w12171 & w12423 ) | ( w12422 & w12423 ) ;
  assign w12425 = w12423 | w12424 ;
  assign w12426 = \pi093 ^ w12158 ;
  assign w12427 = ( ~w12165 & w12425 ) | ( ~w12165 & w12426 ) | ( w12425 & w12426 ) ;
  assign w12428 = w12426 | w12427 ;
  assign w12429 = \pi094 ^ w12152 ;
  assign w12430 = ( ~w12159 & w12428 ) | ( ~w12159 & w12429 ) | ( w12428 & w12429 ) ;
  assign w12431 = w12429 | w12430 ;
  assign w12432 = \pi095 ^ w12146 ;
  assign w12433 = ( ~w12153 & w12431 ) | ( ~w12153 & w12432 ) | ( w12431 & w12432 ) ;
  assign w12434 = w12432 | w12433 ;
  assign w12435 = \pi096 ^ w12140 ;
  assign w12436 = ( ~w12147 & w12434 ) | ( ~w12147 & w12435 ) | ( w12434 & w12435 ) ;
  assign w12437 = w12435 | w12436 ;
  assign w12438 = \pi097 ^ w12134 ;
  assign w12439 = ( ~w12141 & w12437 ) | ( ~w12141 & w12438 ) | ( w12437 & w12438 ) ;
  assign w12440 = w12438 | w12439 ;
  assign w12441 = \pi098 ^ w12128 ;
  assign w12442 = ( ~w12135 & w12440 ) | ( ~w12135 & w12441 ) | ( w12440 & w12441 ) ;
  assign w12443 = w12441 | w12442 ;
  assign w12444 = \pi099 ^ w12122 ;
  assign w12445 = ( ~w12129 & w12443 ) | ( ~w12129 & w12444 ) | ( w12443 & w12444 ) ;
  assign w12446 = w12444 | w12445 ;
  assign w12447 = \pi100 ^ w12116 ;
  assign w12448 = ( ~w12123 & w12446 ) | ( ~w12123 & w12447 ) | ( w12446 & w12447 ) ;
  assign w12449 = w12447 | w12448 ;
  assign w12450 = \pi101 ^ w12110 ;
  assign w12451 = ( ~w12117 & w12449 ) | ( ~w12117 & w12450 ) | ( w12449 & w12450 ) ;
  assign w12452 = w12450 | w12451 ;
  assign w12453 = \pi102 ^ w12104 ;
  assign w12454 = ( ~w12111 & w12452 ) | ( ~w12111 & w12453 ) | ( w12452 & w12453 ) ;
  assign w12455 = w12453 | w12454 ;
  assign w12456 = \pi103 ^ w12098 ;
  assign w12457 = ( ~w12105 & w12455 ) | ( ~w12105 & w12456 ) | ( w12455 & w12456 ) ;
  assign w12458 = w12456 | w12457 ;
  assign w12459 = \pi104 ^ w12092 ;
  assign w12460 = ( ~w12099 & w12458 ) | ( ~w12099 & w12459 ) | ( w12458 & w12459 ) ;
  assign w12461 = w12459 | w12460 ;
  assign w12462 = \pi105 ^ w12086 ;
  assign w12463 = ( ~w12093 & w12461 ) | ( ~w12093 & w12462 ) | ( w12461 & w12462 ) ;
  assign w12464 = w12462 | w12463 ;
  assign w12465 = \pi106 ^ w12080 ;
  assign w12466 = ( ~w12087 & w12464 ) | ( ~w12087 & w12465 ) | ( w12464 & w12465 ) ;
  assign w12467 = w12465 | w12466 ;
  assign w12468 = \pi107 ^ w12074 ;
  assign w12469 = ( ~w12081 & w12467 ) | ( ~w12081 & w12468 ) | ( w12467 & w12468 ) ;
  assign w12470 = w12468 | w12469 ;
  assign w12471 = \pi108 ^ w12068 ;
  assign w12472 = ( ~w12075 & w12470 ) | ( ~w12075 & w12471 ) | ( w12470 & w12471 ) ;
  assign w12473 = w12471 | w12472 ;
  assign w12474 = \pi109 ^ w12062 ;
  assign w12475 = ( ~w12069 & w12473 ) | ( ~w12069 & w12474 ) | ( w12473 & w12474 ) ;
  assign w12476 = w12474 | w12475 ;
  assign w12477 = \pi110 ^ w12056 ;
  assign w12478 = ( ~w12063 & w12476 ) | ( ~w12063 & w12477 ) | ( w12476 & w12477 ) ;
  assign w12479 = w12477 | w12478 ;
  assign w12480 = \pi111 ^ w12050 ;
  assign w12481 = ( ~w12057 & w12479 ) | ( ~w12057 & w12480 ) | ( w12479 & w12480 ) ;
  assign w12482 = w12480 | w12481 ;
  assign w12483 = \pi112 ^ w12044 ;
  assign w12484 = ( ~w12051 & w12482 ) | ( ~w12051 & w12483 ) | ( w12482 & w12483 ) ;
  assign w12485 = w12483 | w12484 ;
  assign w12486 = w11574 & w12039 ;
  assign w12487 = ~w11575 & w12033 ;
  assign w12488 = w12034 ^ w12487 ;
  assign w12489 = ~w12039 & w12488 ;
  assign w12490 = w12486 | w12489 ;
  assign w12491 = ~\pi113 & w12490 ;
  assign w12492 = ( \pi113 & ~w12486 ) | ( \pi113 & w12489 ) | ( ~w12486 & w12489 ) ;
  assign w12493 = ~w12489 & w12492 ;
  assign w12494 = \pi115 | w153 ;
  assign w12495 = ( \pi114 & ~w153 ) | ( \pi114 & w199 ) | ( ~w153 & w199 ) ;
  assign w12496 = w12494 | w12495 ;
  assign w12497 = w12491 | w12493 ;
  assign w12498 = ( ~w12045 & w12485 ) | ( ~w12045 & w12497 ) | ( w12485 & w12497 ) ;
  assign w12499 = ( w12496 & ~w12497 ) | ( w12496 & w12498 ) | ( ~w12497 & w12498 ) ;
  assign w12500 = w12497 | w12499 ;
  assign w12501 = ~w275 & w12490 ;
  assign w12502 = w12500 & ~w12501 ;
  assign w12503 = ~w12051 & w12482 ;
  assign w12504 = w12483 ^ w12503 ;
  assign w12505 = ~w12502 & w12504 ;
  assign w12506 = ( w12044 & w12500 ) | ( w12044 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12507 = ~w12501 & w12506 ;
  assign w12508 = w12505 | w12507 ;
  assign w12509 = ~\pi113 & w12508 ;
  assign w12510 = ~w12057 & w12479 ;
  assign w12511 = w12480 ^ w12510 ;
  assign w12512 = ~w12502 & w12511 ;
  assign w12513 = ( w12050 & w12500 ) | ( w12050 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12514 = ~w12501 & w12513 ;
  assign w12515 = w12512 | w12514 ;
  assign w12516 = ~\pi112 & w12515 ;
  assign w12517 = ~w12063 & w12476 ;
  assign w12518 = w12477 ^ w12517 ;
  assign w12519 = ~w12502 & w12518 ;
  assign w12520 = ( w12056 & w12500 ) | ( w12056 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12521 = ~w12501 & w12520 ;
  assign w12522 = w12519 | w12521 ;
  assign w12523 = ~\pi111 & w12522 ;
  assign w12524 = ~w12069 & w12473 ;
  assign w12525 = w12474 ^ w12524 ;
  assign w12526 = ~w12502 & w12525 ;
  assign w12527 = ( w12062 & w12500 ) | ( w12062 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12528 = ~w12501 & w12527 ;
  assign w12529 = w12526 | w12528 ;
  assign w12530 = ~\pi110 & w12529 ;
  assign w12531 = ~w12075 & w12470 ;
  assign w12532 = w12471 ^ w12531 ;
  assign w12533 = ~w12502 & w12532 ;
  assign w12534 = ( w12068 & w12500 ) | ( w12068 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12535 = ~w12501 & w12534 ;
  assign w12536 = w12533 | w12535 ;
  assign w12537 = ~\pi109 & w12536 ;
  assign w12538 = ~w12081 & w12467 ;
  assign w12539 = w12468 ^ w12538 ;
  assign w12540 = ~w12502 & w12539 ;
  assign w12541 = ( w12074 & w12500 ) | ( w12074 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12542 = ~w12501 & w12541 ;
  assign w12543 = w12540 | w12542 ;
  assign w12544 = ~\pi108 & w12543 ;
  assign w12545 = ~w12087 & w12464 ;
  assign w12546 = w12465 ^ w12545 ;
  assign w12547 = ~w12502 & w12546 ;
  assign w12548 = ( w12080 & w12500 ) | ( w12080 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12549 = ~w12501 & w12548 ;
  assign w12550 = w12547 | w12549 ;
  assign w12551 = ~\pi107 & w12550 ;
  assign w12552 = ~w12093 & w12461 ;
  assign w12553 = w12462 ^ w12552 ;
  assign w12554 = ~w12502 & w12553 ;
  assign w12555 = ( w12086 & w12500 ) | ( w12086 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12556 = ~w12501 & w12555 ;
  assign w12557 = w12554 | w12556 ;
  assign w12558 = ~\pi106 & w12557 ;
  assign w12559 = ~w12099 & w12458 ;
  assign w12560 = w12459 ^ w12559 ;
  assign w12561 = ~w12502 & w12560 ;
  assign w12562 = ( w12092 & w12500 ) | ( w12092 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12563 = ~w12501 & w12562 ;
  assign w12564 = w12561 | w12563 ;
  assign w12565 = ~\pi105 & w12564 ;
  assign w12566 = ~w12105 & w12455 ;
  assign w12567 = w12456 ^ w12566 ;
  assign w12568 = ~w12502 & w12567 ;
  assign w12569 = ( w12098 & w12500 ) | ( w12098 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12570 = ~w12501 & w12569 ;
  assign w12571 = w12568 | w12570 ;
  assign w12572 = ~\pi104 & w12571 ;
  assign w12573 = ~w12111 & w12452 ;
  assign w12574 = w12453 ^ w12573 ;
  assign w12575 = ~w12502 & w12574 ;
  assign w12576 = ( w12104 & w12500 ) | ( w12104 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12577 = ~w12501 & w12576 ;
  assign w12578 = w12575 | w12577 ;
  assign w12579 = ~\pi103 & w12578 ;
  assign w12580 = ~w12117 & w12449 ;
  assign w12581 = w12450 ^ w12580 ;
  assign w12582 = ~w12502 & w12581 ;
  assign w12583 = ( w12110 & w12500 ) | ( w12110 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12584 = ~w12501 & w12583 ;
  assign w12585 = w12582 | w12584 ;
  assign w12586 = ~\pi102 & w12585 ;
  assign w12587 = ~w12123 & w12446 ;
  assign w12588 = w12447 ^ w12587 ;
  assign w12589 = ~w12502 & w12588 ;
  assign w12590 = ( w12116 & w12500 ) | ( w12116 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12591 = ~w12501 & w12590 ;
  assign w12592 = w12589 | w12591 ;
  assign w12593 = ~\pi101 & w12592 ;
  assign w12594 = ~w12129 & w12443 ;
  assign w12595 = w12444 ^ w12594 ;
  assign w12596 = ~w12502 & w12595 ;
  assign w12597 = ( w12122 & w12500 ) | ( w12122 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12598 = ~w12501 & w12597 ;
  assign w12599 = w12596 | w12598 ;
  assign w12600 = ~\pi100 & w12599 ;
  assign w12601 = ~w12135 & w12440 ;
  assign w12602 = w12441 ^ w12601 ;
  assign w12603 = ~w12502 & w12602 ;
  assign w12604 = ( w12128 & w12500 ) | ( w12128 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12605 = ~w12501 & w12604 ;
  assign w12606 = w12603 | w12605 ;
  assign w12607 = ~\pi099 & w12606 ;
  assign w12608 = ~w12141 & w12437 ;
  assign w12609 = w12438 ^ w12608 ;
  assign w12610 = ~w12502 & w12609 ;
  assign w12611 = ( w12134 & w12500 ) | ( w12134 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12612 = ~w12501 & w12611 ;
  assign w12613 = w12610 | w12612 ;
  assign w12614 = ~\pi098 & w12613 ;
  assign w12615 = ~w12147 & w12434 ;
  assign w12616 = w12435 ^ w12615 ;
  assign w12617 = ~w12502 & w12616 ;
  assign w12618 = ( w12140 & w12500 ) | ( w12140 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12619 = ~w12501 & w12618 ;
  assign w12620 = w12617 | w12619 ;
  assign w12621 = ~\pi097 & w12620 ;
  assign w12622 = ~w12153 & w12431 ;
  assign w12623 = w12432 ^ w12622 ;
  assign w12624 = ~w12502 & w12623 ;
  assign w12625 = ( w12146 & w12500 ) | ( w12146 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12626 = ~w12501 & w12625 ;
  assign w12627 = w12624 | w12626 ;
  assign w12628 = ~\pi096 & w12627 ;
  assign w12629 = ~w12159 & w12428 ;
  assign w12630 = w12429 ^ w12629 ;
  assign w12631 = ~w12502 & w12630 ;
  assign w12632 = ( w12152 & w12500 ) | ( w12152 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12633 = ~w12501 & w12632 ;
  assign w12634 = w12631 | w12633 ;
  assign w12635 = ~\pi095 & w12634 ;
  assign w12636 = ~w12165 & w12425 ;
  assign w12637 = w12426 ^ w12636 ;
  assign w12638 = ~w12502 & w12637 ;
  assign w12639 = ( w12158 & w12500 ) | ( w12158 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12640 = ~w12501 & w12639 ;
  assign w12641 = w12638 | w12640 ;
  assign w12642 = ~\pi094 & w12641 ;
  assign w12643 = ~w12171 & w12422 ;
  assign w12644 = w12423 ^ w12643 ;
  assign w12645 = ~w12502 & w12644 ;
  assign w12646 = ( w12164 & w12500 ) | ( w12164 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12647 = ~w12501 & w12646 ;
  assign w12648 = w12645 | w12647 ;
  assign w12649 = ~\pi093 & w12648 ;
  assign w12650 = ~w12177 & w12419 ;
  assign w12651 = w12420 ^ w12650 ;
  assign w12652 = ~w12502 & w12651 ;
  assign w12653 = ( w12170 & w12500 ) | ( w12170 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12654 = ~w12501 & w12653 ;
  assign w12655 = w12652 | w12654 ;
  assign w12656 = ~\pi092 & w12655 ;
  assign w12657 = ~w12183 & w12416 ;
  assign w12658 = w12417 ^ w12657 ;
  assign w12659 = ~w12502 & w12658 ;
  assign w12660 = ( w12176 & w12500 ) | ( w12176 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12661 = ~w12501 & w12660 ;
  assign w12662 = w12659 | w12661 ;
  assign w12663 = ~\pi091 & w12662 ;
  assign w12664 = ~w12189 & w12413 ;
  assign w12665 = w12414 ^ w12664 ;
  assign w12666 = ~w12502 & w12665 ;
  assign w12667 = ( w12182 & w12500 ) | ( w12182 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12668 = ~w12501 & w12667 ;
  assign w12669 = w12666 | w12668 ;
  assign w12670 = ~\pi090 & w12669 ;
  assign w12671 = ~w12195 & w12410 ;
  assign w12672 = w12411 ^ w12671 ;
  assign w12673 = ~w12502 & w12672 ;
  assign w12674 = ( w12188 & w12500 ) | ( w12188 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12675 = ~w12501 & w12674 ;
  assign w12676 = w12673 | w12675 ;
  assign w12677 = ~\pi089 & w12676 ;
  assign w12678 = ~w12201 & w12407 ;
  assign w12679 = w12408 ^ w12678 ;
  assign w12680 = ~w12502 & w12679 ;
  assign w12681 = ( w12194 & w12500 ) | ( w12194 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12682 = ~w12501 & w12681 ;
  assign w12683 = w12680 | w12682 ;
  assign w12684 = ~\pi088 & w12683 ;
  assign w12685 = ~w12207 & w12404 ;
  assign w12686 = w12405 ^ w12685 ;
  assign w12687 = ~w12502 & w12686 ;
  assign w12688 = ( w12200 & w12500 ) | ( w12200 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12689 = ~w12501 & w12688 ;
  assign w12690 = w12687 | w12689 ;
  assign w12691 = ~\pi087 & w12690 ;
  assign w12692 = ~w12213 & w12401 ;
  assign w12693 = w12402 ^ w12692 ;
  assign w12694 = ~w12502 & w12693 ;
  assign w12695 = ( w12206 & w12500 ) | ( w12206 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12696 = ~w12501 & w12695 ;
  assign w12697 = w12694 | w12696 ;
  assign w12698 = ~\pi086 & w12697 ;
  assign w12699 = ~w12219 & w12398 ;
  assign w12700 = w12399 ^ w12699 ;
  assign w12701 = ~w12502 & w12700 ;
  assign w12702 = ( w12212 & w12500 ) | ( w12212 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12703 = ~w12501 & w12702 ;
  assign w12704 = w12701 | w12703 ;
  assign w12705 = ~\pi085 & w12704 ;
  assign w12706 = ~w12225 & w12395 ;
  assign w12707 = w12396 ^ w12706 ;
  assign w12708 = ~w12502 & w12707 ;
  assign w12709 = ( w12218 & w12500 ) | ( w12218 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12710 = ~w12501 & w12709 ;
  assign w12711 = w12708 | w12710 ;
  assign w12712 = ~\pi084 & w12711 ;
  assign w12713 = ~w12231 & w12392 ;
  assign w12714 = w12393 ^ w12713 ;
  assign w12715 = ~w12502 & w12714 ;
  assign w12716 = ( w12224 & w12500 ) | ( w12224 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12717 = ~w12501 & w12716 ;
  assign w12718 = w12715 | w12717 ;
  assign w12719 = ~\pi083 & w12718 ;
  assign w12720 = ~w12237 & w12389 ;
  assign w12721 = w12390 ^ w12720 ;
  assign w12722 = ~w12502 & w12721 ;
  assign w12723 = ( w12230 & w12500 ) | ( w12230 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12724 = ~w12501 & w12723 ;
  assign w12725 = w12722 | w12724 ;
  assign w12726 = ~\pi082 & w12725 ;
  assign w12727 = ~w12243 & w12386 ;
  assign w12728 = w12387 ^ w12727 ;
  assign w12729 = ~w12502 & w12728 ;
  assign w12730 = ( w12236 & w12500 ) | ( w12236 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12731 = ~w12501 & w12730 ;
  assign w12732 = w12729 | w12731 ;
  assign w12733 = ~\pi081 & w12732 ;
  assign w12734 = ~w12249 & w12383 ;
  assign w12735 = w12384 ^ w12734 ;
  assign w12736 = ~w12502 & w12735 ;
  assign w12737 = ( w12242 & w12500 ) | ( w12242 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12738 = ~w12501 & w12737 ;
  assign w12739 = w12736 | w12738 ;
  assign w12740 = ~\pi080 & w12739 ;
  assign w12741 = ~w12255 & w12380 ;
  assign w12742 = w12381 ^ w12741 ;
  assign w12743 = ~w12502 & w12742 ;
  assign w12744 = ( w12248 & w12500 ) | ( w12248 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12745 = ~w12501 & w12744 ;
  assign w12746 = w12743 | w12745 ;
  assign w12747 = ~\pi079 & w12746 ;
  assign w12748 = ~w12261 & w12377 ;
  assign w12749 = w12378 ^ w12748 ;
  assign w12750 = ~w12502 & w12749 ;
  assign w12751 = ( w12254 & w12500 ) | ( w12254 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12752 = ~w12501 & w12751 ;
  assign w12753 = w12750 | w12752 ;
  assign w12754 = ~\pi078 & w12753 ;
  assign w12755 = ~w12267 & w12374 ;
  assign w12756 = w12375 ^ w12755 ;
  assign w12757 = ~w12502 & w12756 ;
  assign w12758 = ( w12260 & w12500 ) | ( w12260 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12759 = ~w12501 & w12758 ;
  assign w12760 = w12757 | w12759 ;
  assign w12761 = ~\pi077 & w12760 ;
  assign w12762 = ~w12273 & w12371 ;
  assign w12763 = w12372 ^ w12762 ;
  assign w12764 = ~w12502 & w12763 ;
  assign w12765 = ( w12266 & w12500 ) | ( w12266 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12766 = ~w12501 & w12765 ;
  assign w12767 = w12764 | w12766 ;
  assign w12768 = ~\pi076 & w12767 ;
  assign w12769 = ~w12279 & w12368 ;
  assign w12770 = w12369 ^ w12769 ;
  assign w12771 = ~w12502 & w12770 ;
  assign w12772 = ( w12272 & w12500 ) | ( w12272 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12773 = ~w12501 & w12772 ;
  assign w12774 = w12771 | w12773 ;
  assign w12775 = ~\pi075 & w12774 ;
  assign w12776 = ~w12285 & w12365 ;
  assign w12777 = w12366 ^ w12776 ;
  assign w12778 = ~w12502 & w12777 ;
  assign w12779 = ( w12278 & w12500 ) | ( w12278 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12780 = ~w12501 & w12779 ;
  assign w12781 = w12778 | w12780 ;
  assign w12782 = ~\pi074 & w12781 ;
  assign w12783 = ~w12291 & w12362 ;
  assign w12784 = w12363 ^ w12783 ;
  assign w12785 = ~w12502 & w12784 ;
  assign w12786 = ( w12284 & w12500 ) | ( w12284 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12787 = ~w12501 & w12786 ;
  assign w12788 = w12785 | w12787 ;
  assign w12789 = ~\pi073 & w12788 ;
  assign w12790 = ~w12297 & w12359 ;
  assign w12791 = w12360 ^ w12790 ;
  assign w12792 = ~w12502 & w12791 ;
  assign w12793 = ( w12290 & w12500 ) | ( w12290 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12794 = ~w12501 & w12793 ;
  assign w12795 = w12792 | w12794 ;
  assign w12796 = ~\pi072 & w12795 ;
  assign w12797 = ~w12303 & w12356 ;
  assign w12798 = w12357 ^ w12797 ;
  assign w12799 = ~w12502 & w12798 ;
  assign w12800 = ( w12296 & w12500 ) | ( w12296 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12801 = ~w12501 & w12800 ;
  assign w12802 = w12799 | w12801 ;
  assign w12803 = ~\pi071 & w12802 ;
  assign w12804 = ~w12309 & w12353 ;
  assign w12805 = w12354 ^ w12804 ;
  assign w12806 = ~w12502 & w12805 ;
  assign w12807 = ( w12302 & w12500 ) | ( w12302 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12808 = ~w12501 & w12807 ;
  assign w12809 = w12806 | w12808 ;
  assign w12810 = ~\pi070 & w12809 ;
  assign w12811 = ~w12317 & w12350 ;
  assign w12812 = w12351 ^ w12811 ;
  assign w12813 = ~w12502 & w12812 ;
  assign w12814 = ( w12308 & w12500 ) | ( w12308 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12815 = ~w12501 & w12814 ;
  assign w12816 = w12813 | w12815 ;
  assign w12817 = ~\pi069 & w12816 ;
  assign w12818 = ~w12328 & w12345 ;
  assign w12819 = w12348 ^ w12818 ;
  assign w12820 = ~w12502 & w12819 ;
  assign w12821 = ( w12316 & w12500 ) | ( w12316 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12822 = ~w12501 & w12821 ;
  assign w12823 = w12820 | w12822 ;
  assign w12824 = ~\pi068 & w12823 ;
  assign w12825 = w12342 ^ w12344 ;
  assign w12826 = ~w12502 & w12825 ;
  assign w12827 = ( w12327 & w12500 ) | ( w12327 & w12501 ) | ( w12500 & w12501 ) ;
  assign w12828 = ~w12501 & w12827 ;
  assign w12829 = w12826 | w12828 ;
  assign w12830 = ~\pi067 & w12829 ;
  assign w12831 = w12339 ^ w12343 ;
  assign w12832 = \pi065 ^ w12831 ;
  assign w12833 = w12502 ^ w12832 ;
  assign w12834 = ( w12343 & w12832 ) | ( w12343 & w12833 ) | ( w12832 & w12833 ) ;
  assign w12835 = ~\pi066 & w12834 ;
  assign w12836 = w12343 ^ w12502 ;
  assign w12837 = ( w12343 & w12832 ) | ( w12343 & ~w12836 ) | ( w12832 & ~w12836 ) ;
  assign w12838 = \pi066 ^ w12837 ;
  assign w12839 = \pi064 & ~w12502 ;
  assign w12840 = \pi014 ^ w12839 ;
  assign w12841 = ( ~\pi013 & \pi064 ) | ( ~\pi013 & w12838 ) | ( \pi064 & w12838 ) ;
  assign w12842 = ( \pi065 & ~w12840 ) | ( \pi065 & w12841 ) | ( ~w12840 & w12841 ) ;
  assign w12843 = w12838 | w12842 ;
  assign w12844 = \pi067 ^ w12829 ;
  assign w12845 = ( ~w12835 & w12843 ) | ( ~w12835 & w12844 ) | ( w12843 & w12844 ) ;
  assign w12846 = w12844 | w12845 ;
  assign w12847 = \pi068 ^ w12823 ;
  assign w12848 = ( ~w12830 & w12846 ) | ( ~w12830 & w12847 ) | ( w12846 & w12847 ) ;
  assign w12849 = w12847 | w12848 ;
  assign w12850 = \pi069 ^ w12816 ;
  assign w12851 = ( ~w12824 & w12849 ) | ( ~w12824 & w12850 ) | ( w12849 & w12850 ) ;
  assign w12852 = w12850 | w12851 ;
  assign w12853 = \pi070 ^ w12809 ;
  assign w12854 = ( ~w12817 & w12852 ) | ( ~w12817 & w12853 ) | ( w12852 & w12853 ) ;
  assign w12855 = w12853 | w12854 ;
  assign w12856 = \pi071 ^ w12802 ;
  assign w12857 = ( ~w12810 & w12855 ) | ( ~w12810 & w12856 ) | ( w12855 & w12856 ) ;
  assign w12858 = w12856 | w12857 ;
  assign w12859 = \pi072 ^ w12795 ;
  assign w12860 = ( ~w12803 & w12858 ) | ( ~w12803 & w12859 ) | ( w12858 & w12859 ) ;
  assign w12861 = w12859 | w12860 ;
  assign w12862 = \pi073 ^ w12788 ;
  assign w12863 = ( ~w12796 & w12861 ) | ( ~w12796 & w12862 ) | ( w12861 & w12862 ) ;
  assign w12864 = w12862 | w12863 ;
  assign w12865 = \pi074 ^ w12781 ;
  assign w12866 = ( ~w12789 & w12864 ) | ( ~w12789 & w12865 ) | ( w12864 & w12865 ) ;
  assign w12867 = w12865 | w12866 ;
  assign w12868 = \pi075 ^ w12774 ;
  assign w12869 = ( ~w12782 & w12867 ) | ( ~w12782 & w12868 ) | ( w12867 & w12868 ) ;
  assign w12870 = w12868 | w12869 ;
  assign w12871 = \pi076 ^ w12767 ;
  assign w12872 = ( ~w12775 & w12870 ) | ( ~w12775 & w12871 ) | ( w12870 & w12871 ) ;
  assign w12873 = w12871 | w12872 ;
  assign w12874 = \pi077 ^ w12760 ;
  assign w12875 = ( ~w12768 & w12873 ) | ( ~w12768 & w12874 ) | ( w12873 & w12874 ) ;
  assign w12876 = w12874 | w12875 ;
  assign w12877 = \pi078 ^ w12753 ;
  assign w12878 = ( ~w12761 & w12876 ) | ( ~w12761 & w12877 ) | ( w12876 & w12877 ) ;
  assign w12879 = w12877 | w12878 ;
  assign w12880 = \pi079 ^ w12746 ;
  assign w12881 = ( ~w12754 & w12879 ) | ( ~w12754 & w12880 ) | ( w12879 & w12880 ) ;
  assign w12882 = w12880 | w12881 ;
  assign w12883 = \pi080 ^ w12739 ;
  assign w12884 = ( ~w12747 & w12882 ) | ( ~w12747 & w12883 ) | ( w12882 & w12883 ) ;
  assign w12885 = w12883 | w12884 ;
  assign w12886 = \pi081 ^ w12732 ;
  assign w12887 = ( ~w12740 & w12885 ) | ( ~w12740 & w12886 ) | ( w12885 & w12886 ) ;
  assign w12888 = w12886 | w12887 ;
  assign w12889 = \pi082 ^ w12725 ;
  assign w12890 = ( ~w12733 & w12888 ) | ( ~w12733 & w12889 ) | ( w12888 & w12889 ) ;
  assign w12891 = w12889 | w12890 ;
  assign w12892 = \pi083 ^ w12718 ;
  assign w12893 = ( ~w12726 & w12891 ) | ( ~w12726 & w12892 ) | ( w12891 & w12892 ) ;
  assign w12894 = w12892 | w12893 ;
  assign w12895 = \pi084 ^ w12711 ;
  assign w12896 = ( ~w12719 & w12894 ) | ( ~w12719 & w12895 ) | ( w12894 & w12895 ) ;
  assign w12897 = w12895 | w12896 ;
  assign w12898 = \pi085 ^ w12704 ;
  assign w12899 = ( ~w12712 & w12897 ) | ( ~w12712 & w12898 ) | ( w12897 & w12898 ) ;
  assign w12900 = w12898 | w12899 ;
  assign w12901 = \pi086 ^ w12697 ;
  assign w12902 = ( ~w12705 & w12900 ) | ( ~w12705 & w12901 ) | ( w12900 & w12901 ) ;
  assign w12903 = w12901 | w12902 ;
  assign w12904 = \pi087 ^ w12690 ;
  assign w12905 = ( ~w12698 & w12903 ) | ( ~w12698 & w12904 ) | ( w12903 & w12904 ) ;
  assign w12906 = w12904 | w12905 ;
  assign w12907 = \pi088 ^ w12683 ;
  assign w12908 = ( ~w12691 & w12906 ) | ( ~w12691 & w12907 ) | ( w12906 & w12907 ) ;
  assign w12909 = w12907 | w12908 ;
  assign w12910 = \pi089 ^ w12676 ;
  assign w12911 = ( ~w12684 & w12909 ) | ( ~w12684 & w12910 ) | ( w12909 & w12910 ) ;
  assign w12912 = w12910 | w12911 ;
  assign w12913 = \pi090 ^ w12669 ;
  assign w12914 = ( ~w12677 & w12912 ) | ( ~w12677 & w12913 ) | ( w12912 & w12913 ) ;
  assign w12915 = w12913 | w12914 ;
  assign w12916 = \pi091 ^ w12662 ;
  assign w12917 = ( ~w12670 & w12915 ) | ( ~w12670 & w12916 ) | ( w12915 & w12916 ) ;
  assign w12918 = w12916 | w12917 ;
  assign w12919 = \pi092 ^ w12655 ;
  assign w12920 = ( ~w12663 & w12918 ) | ( ~w12663 & w12919 ) | ( w12918 & w12919 ) ;
  assign w12921 = w12919 | w12920 ;
  assign w12922 = \pi093 ^ w12648 ;
  assign w12923 = ( ~w12656 & w12921 ) | ( ~w12656 & w12922 ) | ( w12921 & w12922 ) ;
  assign w12924 = w12922 | w12923 ;
  assign w12925 = \pi094 ^ w12641 ;
  assign w12926 = ( ~w12649 & w12924 ) | ( ~w12649 & w12925 ) | ( w12924 & w12925 ) ;
  assign w12927 = w12925 | w12926 ;
  assign w12928 = \pi095 ^ w12634 ;
  assign w12929 = ( ~w12642 & w12927 ) | ( ~w12642 & w12928 ) | ( w12927 & w12928 ) ;
  assign w12930 = w12928 | w12929 ;
  assign w12931 = \pi096 ^ w12627 ;
  assign w12932 = ( ~w12635 & w12930 ) | ( ~w12635 & w12931 ) | ( w12930 & w12931 ) ;
  assign w12933 = w12931 | w12932 ;
  assign w12934 = \pi097 ^ w12620 ;
  assign w12935 = ( ~w12628 & w12933 ) | ( ~w12628 & w12934 ) | ( w12933 & w12934 ) ;
  assign w12936 = w12934 | w12935 ;
  assign w12937 = \pi098 ^ w12613 ;
  assign w12938 = ( ~w12621 & w12936 ) | ( ~w12621 & w12937 ) | ( w12936 & w12937 ) ;
  assign w12939 = w12937 | w12938 ;
  assign w12940 = \pi099 ^ w12606 ;
  assign w12941 = ( ~w12614 & w12939 ) | ( ~w12614 & w12940 ) | ( w12939 & w12940 ) ;
  assign w12942 = w12940 | w12941 ;
  assign w12943 = \pi100 ^ w12599 ;
  assign w12944 = ( ~w12607 & w12942 ) | ( ~w12607 & w12943 ) | ( w12942 & w12943 ) ;
  assign w12945 = w12943 | w12944 ;
  assign w12946 = \pi101 ^ w12592 ;
  assign w12947 = ( ~w12600 & w12945 ) | ( ~w12600 & w12946 ) | ( w12945 & w12946 ) ;
  assign w12948 = w12946 | w12947 ;
  assign w12949 = \pi102 ^ w12585 ;
  assign w12950 = ( ~w12593 & w12948 ) | ( ~w12593 & w12949 ) | ( w12948 & w12949 ) ;
  assign w12951 = w12949 | w12950 ;
  assign w12952 = \pi103 ^ w12578 ;
  assign w12953 = ( ~w12586 & w12951 ) | ( ~w12586 & w12952 ) | ( w12951 & w12952 ) ;
  assign w12954 = w12952 | w12953 ;
  assign w12955 = \pi104 ^ w12571 ;
  assign w12956 = ( ~w12579 & w12954 ) | ( ~w12579 & w12955 ) | ( w12954 & w12955 ) ;
  assign w12957 = w12955 | w12956 ;
  assign w12958 = \pi105 ^ w12564 ;
  assign w12959 = ( ~w12572 & w12957 ) | ( ~w12572 & w12958 ) | ( w12957 & w12958 ) ;
  assign w12960 = w12958 | w12959 ;
  assign w12961 = \pi106 ^ w12557 ;
  assign w12962 = ( ~w12565 & w12960 ) | ( ~w12565 & w12961 ) | ( w12960 & w12961 ) ;
  assign w12963 = w12961 | w12962 ;
  assign w12964 = \pi107 ^ w12550 ;
  assign w12965 = ( ~w12558 & w12963 ) | ( ~w12558 & w12964 ) | ( w12963 & w12964 ) ;
  assign w12966 = w12964 | w12965 ;
  assign w12967 = \pi108 ^ w12543 ;
  assign w12968 = ( ~w12551 & w12966 ) | ( ~w12551 & w12967 ) | ( w12966 & w12967 ) ;
  assign w12969 = w12967 | w12968 ;
  assign w12970 = \pi109 ^ w12536 ;
  assign w12971 = ( ~w12544 & w12969 ) | ( ~w12544 & w12970 ) | ( w12969 & w12970 ) ;
  assign w12972 = w12970 | w12971 ;
  assign w12973 = \pi110 ^ w12529 ;
  assign w12974 = ( ~w12537 & w12972 ) | ( ~w12537 & w12973 ) | ( w12972 & w12973 ) ;
  assign w12975 = w12973 | w12974 ;
  assign w12976 = \pi111 ^ w12522 ;
  assign w12977 = ( ~w12530 & w12975 ) | ( ~w12530 & w12976 ) | ( w12975 & w12976 ) ;
  assign w12978 = w12976 | w12977 ;
  assign w12979 = \pi112 ^ w12515 ;
  assign w12980 = ( ~w12523 & w12978 ) | ( ~w12523 & w12979 ) | ( w12978 & w12979 ) ;
  assign w12981 = w12979 | w12980 ;
  assign w12982 = \pi113 ^ w12508 ;
  assign w12983 = ( ~w12516 & w12981 ) | ( ~w12516 & w12982 ) | ( w12981 & w12982 ) ;
  assign w12984 = w12982 | w12983 ;
  assign w12985 = ( ~w12045 & w12485 ) | ( ~w12045 & w12502 ) | ( w12485 & w12502 ) ;
  assign w12986 = w12497 ^ w12985 ;
  assign w12987 = ~w12502 & w12986 ;
  assign w12988 = ( w275 & ~w12490 ) | ( w275 & w12500 ) | ( ~w12490 & w12500 ) ;
  assign w12989 = w12490 & w12988 ;
  assign w12990 = w12987 | w12989 ;
  assign w12991 = ~\pi114 & w12990 ;
  assign w12992 = ( \pi114 & ~w12987 ) | ( \pi114 & w12989 ) | ( ~w12987 & w12989 ) ;
  assign w12993 = ~w12989 & w12992 ;
  assign w12994 = \pi116 | w264 ;
  assign w12995 = ( \pi115 & ~w264 ) | ( \pi115 & w273 ) | ( ~w264 & w273 ) ;
  assign w12996 = w12994 | w12995 ;
  assign w12997 = w12991 | w12993 ;
  assign w12998 = ( ~w12509 & w12984 ) | ( ~w12509 & w12997 ) | ( w12984 & w12997 ) ;
  assign w12999 = ( w12996 & ~w12997 ) | ( w12996 & w12998 ) | ( ~w12997 & w12998 ) ;
  assign w13000 = w12997 | w12999 ;
  assign w13001 = ~w12496 & w12990 ;
  assign w13002 = w13000 & ~w13001 ;
  assign w13003 = ~w12516 & w12981 ;
  assign w13004 = w12982 ^ w13003 ;
  assign w13005 = ~w13002 & w13004 ;
  assign w13006 = ( w12508 & w13000 ) | ( w12508 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13007 = ~w13001 & w13006 ;
  assign w13008 = w13005 | w13007 ;
  assign w13009 = ( ~w12509 & w12984 ) | ( ~w12509 & w13002 ) | ( w12984 & w13002 ) ;
  assign w13010 = w12997 ^ w13009 ;
  assign w13011 = ~w13002 & w13010 ;
  assign w13012 = ( w12496 & ~w12990 ) | ( w12496 & w13000 ) | ( ~w12990 & w13000 ) ;
  assign w13013 = w12990 & w13012 ;
  assign w13014 = w13011 | w13013 ;
  assign w13015 = ~\pi114 & w13008 ;
  assign w13016 = ~w12523 & w12978 ;
  assign w13017 = w12979 ^ w13016 ;
  assign w13018 = ~w13002 & w13017 ;
  assign w13019 = ( w12515 & w13000 ) | ( w12515 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13020 = ~w13001 & w13019 ;
  assign w13021 = w13018 | w13020 ;
  assign w13022 = ~\pi113 & w13021 ;
  assign w13023 = ~w12530 & w12975 ;
  assign w13024 = w12976 ^ w13023 ;
  assign w13025 = ~w13002 & w13024 ;
  assign w13026 = ( w12522 & w13000 ) | ( w12522 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13027 = ~w13001 & w13026 ;
  assign w13028 = w13025 | w13027 ;
  assign w13029 = ~\pi112 & w13028 ;
  assign w13030 = ~w12537 & w12972 ;
  assign w13031 = w12973 ^ w13030 ;
  assign w13032 = ~w13002 & w13031 ;
  assign w13033 = ( w12529 & w13000 ) | ( w12529 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13034 = ~w13001 & w13033 ;
  assign w13035 = w13032 | w13034 ;
  assign w13036 = ~\pi111 & w13035 ;
  assign w13037 = ~w12544 & w12969 ;
  assign w13038 = w12970 ^ w13037 ;
  assign w13039 = ~w13002 & w13038 ;
  assign w13040 = ( w12536 & w13000 ) | ( w12536 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13041 = ~w13001 & w13040 ;
  assign w13042 = w13039 | w13041 ;
  assign w13043 = ~\pi110 & w13042 ;
  assign w13044 = ~w12551 & w12966 ;
  assign w13045 = w12967 ^ w13044 ;
  assign w13046 = ~w13002 & w13045 ;
  assign w13047 = ( w12543 & w13000 ) | ( w12543 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13048 = ~w13001 & w13047 ;
  assign w13049 = w13046 | w13048 ;
  assign w13050 = ~\pi109 & w13049 ;
  assign w13051 = ~w12558 & w12963 ;
  assign w13052 = w12964 ^ w13051 ;
  assign w13053 = ~w13002 & w13052 ;
  assign w13054 = ( w12550 & w13000 ) | ( w12550 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13055 = ~w13001 & w13054 ;
  assign w13056 = w13053 | w13055 ;
  assign w13057 = ~\pi108 & w13056 ;
  assign w13058 = ~w12565 & w12960 ;
  assign w13059 = w12961 ^ w13058 ;
  assign w13060 = ~w13002 & w13059 ;
  assign w13061 = ( w12557 & w13000 ) | ( w12557 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13062 = ~w13001 & w13061 ;
  assign w13063 = w13060 | w13062 ;
  assign w13064 = ~\pi107 & w13063 ;
  assign w13065 = ~w12572 & w12957 ;
  assign w13066 = w12958 ^ w13065 ;
  assign w13067 = ~w13002 & w13066 ;
  assign w13068 = ( w12564 & w13000 ) | ( w12564 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13069 = ~w13001 & w13068 ;
  assign w13070 = w13067 | w13069 ;
  assign w13071 = ~\pi106 & w13070 ;
  assign w13072 = ~w12579 & w12954 ;
  assign w13073 = w12955 ^ w13072 ;
  assign w13074 = ~w13002 & w13073 ;
  assign w13075 = ( w12571 & w13000 ) | ( w12571 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13076 = ~w13001 & w13075 ;
  assign w13077 = w13074 | w13076 ;
  assign w13078 = ~\pi105 & w13077 ;
  assign w13079 = ~w12586 & w12951 ;
  assign w13080 = w12952 ^ w13079 ;
  assign w13081 = ~w13002 & w13080 ;
  assign w13082 = ( w12578 & w13000 ) | ( w12578 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13083 = ~w13001 & w13082 ;
  assign w13084 = w13081 | w13083 ;
  assign w13085 = ~\pi104 & w13084 ;
  assign w13086 = ~w12593 & w12948 ;
  assign w13087 = w12949 ^ w13086 ;
  assign w13088 = ~w13002 & w13087 ;
  assign w13089 = ( w12585 & w13000 ) | ( w12585 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13090 = ~w13001 & w13089 ;
  assign w13091 = w13088 | w13090 ;
  assign w13092 = ~\pi103 & w13091 ;
  assign w13093 = ~w12600 & w12945 ;
  assign w13094 = w12946 ^ w13093 ;
  assign w13095 = ~w13002 & w13094 ;
  assign w13096 = ( w12592 & w13000 ) | ( w12592 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13097 = ~w13001 & w13096 ;
  assign w13098 = w13095 | w13097 ;
  assign w13099 = ~\pi102 & w13098 ;
  assign w13100 = ~w12607 & w12942 ;
  assign w13101 = w12943 ^ w13100 ;
  assign w13102 = ~w13002 & w13101 ;
  assign w13103 = ( w12599 & w13000 ) | ( w12599 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13104 = ~w13001 & w13103 ;
  assign w13105 = w13102 | w13104 ;
  assign w13106 = ~\pi101 & w13105 ;
  assign w13107 = ~w12614 & w12939 ;
  assign w13108 = w12940 ^ w13107 ;
  assign w13109 = ~w13002 & w13108 ;
  assign w13110 = ( w12606 & w13000 ) | ( w12606 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13111 = ~w13001 & w13110 ;
  assign w13112 = w13109 | w13111 ;
  assign w13113 = ~\pi100 & w13112 ;
  assign w13114 = ~w12621 & w12936 ;
  assign w13115 = w12937 ^ w13114 ;
  assign w13116 = ~w13002 & w13115 ;
  assign w13117 = ( w12613 & w13000 ) | ( w12613 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13118 = ~w13001 & w13117 ;
  assign w13119 = w13116 | w13118 ;
  assign w13120 = ~\pi099 & w13119 ;
  assign w13121 = ~w12628 & w12933 ;
  assign w13122 = w12934 ^ w13121 ;
  assign w13123 = ~w13002 & w13122 ;
  assign w13124 = ( w12620 & w13000 ) | ( w12620 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13125 = ~w13001 & w13124 ;
  assign w13126 = w13123 | w13125 ;
  assign w13127 = ~\pi098 & w13126 ;
  assign w13128 = ~w12635 & w12930 ;
  assign w13129 = w12931 ^ w13128 ;
  assign w13130 = ~w13002 & w13129 ;
  assign w13131 = ( w12627 & w13000 ) | ( w12627 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13132 = ~w13001 & w13131 ;
  assign w13133 = w13130 | w13132 ;
  assign w13134 = ~\pi097 & w13133 ;
  assign w13135 = ~w12642 & w12927 ;
  assign w13136 = w12928 ^ w13135 ;
  assign w13137 = ~w13002 & w13136 ;
  assign w13138 = ( w12634 & w13000 ) | ( w12634 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13139 = ~w13001 & w13138 ;
  assign w13140 = w13137 | w13139 ;
  assign w13141 = ~\pi096 & w13140 ;
  assign w13142 = ~w12649 & w12924 ;
  assign w13143 = w12925 ^ w13142 ;
  assign w13144 = ~w13002 & w13143 ;
  assign w13145 = ( w12641 & w13000 ) | ( w12641 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13146 = ~w13001 & w13145 ;
  assign w13147 = w13144 | w13146 ;
  assign w13148 = ~\pi095 & w13147 ;
  assign w13149 = ~w12656 & w12921 ;
  assign w13150 = w12922 ^ w13149 ;
  assign w13151 = ~w13002 & w13150 ;
  assign w13152 = ( w12648 & w13000 ) | ( w12648 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13153 = ~w13001 & w13152 ;
  assign w13154 = w13151 | w13153 ;
  assign w13155 = ~\pi094 & w13154 ;
  assign w13156 = ~w12663 & w12918 ;
  assign w13157 = w12919 ^ w13156 ;
  assign w13158 = ~w13002 & w13157 ;
  assign w13159 = ( w12655 & w13000 ) | ( w12655 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13160 = ~w13001 & w13159 ;
  assign w13161 = w13158 | w13160 ;
  assign w13162 = ~\pi093 & w13161 ;
  assign w13163 = ~w12670 & w12915 ;
  assign w13164 = w12916 ^ w13163 ;
  assign w13165 = ~w13002 & w13164 ;
  assign w13166 = ( w12662 & w13000 ) | ( w12662 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13167 = ~w13001 & w13166 ;
  assign w13168 = w13165 | w13167 ;
  assign w13169 = ~\pi092 & w13168 ;
  assign w13170 = ~w12677 & w12912 ;
  assign w13171 = w12913 ^ w13170 ;
  assign w13172 = ~w13002 & w13171 ;
  assign w13173 = ( w12669 & w13000 ) | ( w12669 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13174 = ~w13001 & w13173 ;
  assign w13175 = w13172 | w13174 ;
  assign w13176 = ~\pi091 & w13175 ;
  assign w13177 = ~w12684 & w12909 ;
  assign w13178 = w12910 ^ w13177 ;
  assign w13179 = ~w13002 & w13178 ;
  assign w13180 = ( w12676 & w13000 ) | ( w12676 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13181 = ~w13001 & w13180 ;
  assign w13182 = w13179 | w13181 ;
  assign w13183 = ~\pi090 & w13182 ;
  assign w13184 = ~w12691 & w12906 ;
  assign w13185 = w12907 ^ w13184 ;
  assign w13186 = ~w13002 & w13185 ;
  assign w13187 = ( w12683 & w13000 ) | ( w12683 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13188 = ~w13001 & w13187 ;
  assign w13189 = w13186 | w13188 ;
  assign w13190 = ~\pi089 & w13189 ;
  assign w13191 = ~w12698 & w12903 ;
  assign w13192 = w12904 ^ w13191 ;
  assign w13193 = ~w13002 & w13192 ;
  assign w13194 = ( w12690 & w13000 ) | ( w12690 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13195 = ~w13001 & w13194 ;
  assign w13196 = w13193 | w13195 ;
  assign w13197 = ~\pi088 & w13196 ;
  assign w13198 = ~w12705 & w12900 ;
  assign w13199 = w12901 ^ w13198 ;
  assign w13200 = ~w13002 & w13199 ;
  assign w13201 = ( w12697 & w13000 ) | ( w12697 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13202 = ~w13001 & w13201 ;
  assign w13203 = w13200 | w13202 ;
  assign w13204 = ~\pi087 & w13203 ;
  assign w13205 = ~w12712 & w12897 ;
  assign w13206 = w12898 ^ w13205 ;
  assign w13207 = ~w13002 & w13206 ;
  assign w13208 = ( w12704 & w13000 ) | ( w12704 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13209 = ~w13001 & w13208 ;
  assign w13210 = w13207 | w13209 ;
  assign w13211 = ~\pi086 & w13210 ;
  assign w13212 = ~w12719 & w12894 ;
  assign w13213 = w12895 ^ w13212 ;
  assign w13214 = ~w13002 & w13213 ;
  assign w13215 = ( w12711 & w13000 ) | ( w12711 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13216 = ~w13001 & w13215 ;
  assign w13217 = w13214 | w13216 ;
  assign w13218 = ~\pi085 & w13217 ;
  assign w13219 = ~w12726 & w12891 ;
  assign w13220 = w12892 ^ w13219 ;
  assign w13221 = ~w13002 & w13220 ;
  assign w13222 = ( w12718 & w13000 ) | ( w12718 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13223 = ~w13001 & w13222 ;
  assign w13224 = w13221 | w13223 ;
  assign w13225 = ~\pi084 & w13224 ;
  assign w13226 = ~w12733 & w12888 ;
  assign w13227 = w12889 ^ w13226 ;
  assign w13228 = ~w13002 & w13227 ;
  assign w13229 = ( w12725 & w13000 ) | ( w12725 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13230 = ~w13001 & w13229 ;
  assign w13231 = w13228 | w13230 ;
  assign w13232 = ~\pi083 & w13231 ;
  assign w13233 = ~w12740 & w12885 ;
  assign w13234 = w12886 ^ w13233 ;
  assign w13235 = ~w13002 & w13234 ;
  assign w13236 = ( w12732 & w13000 ) | ( w12732 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13237 = ~w13001 & w13236 ;
  assign w13238 = w13235 | w13237 ;
  assign w13239 = ~\pi082 & w13238 ;
  assign w13240 = ~w12747 & w12882 ;
  assign w13241 = w12883 ^ w13240 ;
  assign w13242 = ~w13002 & w13241 ;
  assign w13243 = ( w12739 & w13000 ) | ( w12739 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13244 = ~w13001 & w13243 ;
  assign w13245 = w13242 | w13244 ;
  assign w13246 = ~\pi081 & w13245 ;
  assign w13247 = ~w12754 & w12879 ;
  assign w13248 = w12880 ^ w13247 ;
  assign w13249 = ~w13002 & w13248 ;
  assign w13250 = ( w12746 & w13000 ) | ( w12746 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13251 = ~w13001 & w13250 ;
  assign w13252 = w13249 | w13251 ;
  assign w13253 = ~\pi080 & w13252 ;
  assign w13254 = ~w12761 & w12876 ;
  assign w13255 = w12877 ^ w13254 ;
  assign w13256 = ~w13002 & w13255 ;
  assign w13257 = ( w12753 & w13000 ) | ( w12753 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13258 = ~w13001 & w13257 ;
  assign w13259 = w13256 | w13258 ;
  assign w13260 = ~\pi079 & w13259 ;
  assign w13261 = ~w12768 & w12873 ;
  assign w13262 = w12874 ^ w13261 ;
  assign w13263 = ~w13002 & w13262 ;
  assign w13264 = ( w12760 & w13000 ) | ( w12760 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13265 = ~w13001 & w13264 ;
  assign w13266 = w13263 | w13265 ;
  assign w13267 = ~\pi078 & w13266 ;
  assign w13268 = ~w12775 & w12870 ;
  assign w13269 = w12871 ^ w13268 ;
  assign w13270 = ~w13002 & w13269 ;
  assign w13271 = ( w12767 & w13000 ) | ( w12767 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13272 = ~w13001 & w13271 ;
  assign w13273 = w13270 | w13272 ;
  assign w13274 = ~\pi077 & w13273 ;
  assign w13275 = ~w12782 & w12867 ;
  assign w13276 = w12868 ^ w13275 ;
  assign w13277 = ~w13002 & w13276 ;
  assign w13278 = ( w12774 & w13000 ) | ( w12774 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13279 = ~w13001 & w13278 ;
  assign w13280 = w13277 | w13279 ;
  assign w13281 = ~\pi076 & w13280 ;
  assign w13282 = ~w12789 & w12864 ;
  assign w13283 = w12865 ^ w13282 ;
  assign w13284 = ~w13002 & w13283 ;
  assign w13285 = ( w12781 & w13000 ) | ( w12781 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13286 = ~w13001 & w13285 ;
  assign w13287 = w13284 | w13286 ;
  assign w13288 = ~\pi075 & w13287 ;
  assign w13289 = ~w12796 & w12861 ;
  assign w13290 = w12862 ^ w13289 ;
  assign w13291 = ~w13002 & w13290 ;
  assign w13292 = ( w12788 & w13000 ) | ( w12788 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13293 = ~w13001 & w13292 ;
  assign w13294 = w13291 | w13293 ;
  assign w13295 = ~\pi074 & w13294 ;
  assign w13296 = ~w12803 & w12858 ;
  assign w13297 = w12859 ^ w13296 ;
  assign w13298 = ~w13002 & w13297 ;
  assign w13299 = ( w12795 & w13000 ) | ( w12795 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13300 = ~w13001 & w13299 ;
  assign w13301 = w13298 | w13300 ;
  assign w13302 = ~\pi073 & w13301 ;
  assign w13303 = ~w12810 & w12855 ;
  assign w13304 = w12856 ^ w13303 ;
  assign w13305 = ~w13002 & w13304 ;
  assign w13306 = ( w12802 & w13000 ) | ( w12802 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13307 = ~w13001 & w13306 ;
  assign w13308 = w13305 | w13307 ;
  assign w13309 = ~\pi072 & w13308 ;
  assign w13310 = ~w12817 & w12852 ;
  assign w13311 = w12853 ^ w13310 ;
  assign w13312 = ~w13002 & w13311 ;
  assign w13313 = ( w12809 & w13000 ) | ( w12809 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13314 = ~w13001 & w13313 ;
  assign w13315 = w13312 | w13314 ;
  assign w13316 = ~\pi071 & w13315 ;
  assign w13317 = ~w12824 & w12849 ;
  assign w13318 = w12850 ^ w13317 ;
  assign w13319 = ~w13002 & w13318 ;
  assign w13320 = ( w12816 & w13000 ) | ( w12816 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13321 = ~w13001 & w13320 ;
  assign w13322 = w13319 | w13321 ;
  assign w13323 = ~\pi070 & w13322 ;
  assign w13324 = ~w12830 & w12846 ;
  assign w13325 = w12847 ^ w13324 ;
  assign w13326 = ~w13002 & w13325 ;
  assign w13327 = ( w12823 & w13000 ) | ( w12823 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13328 = ~w13001 & w13327 ;
  assign w13329 = w13326 | w13328 ;
  assign w13330 = ~\pi069 & w13329 ;
  assign w13331 = ~w12835 & w12843 ;
  assign w13332 = w12844 ^ w13331 ;
  assign w13333 = ~w13002 & w13332 ;
  assign w13334 = ( w12829 & w13000 ) | ( w12829 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13335 = ~w13001 & w13334 ;
  assign w13336 = w13333 | w13335 ;
  assign w13337 = ~\pi068 & w13336 ;
  assign w13338 = ~\pi013 & \pi064 ;
  assign w13339 = ( \pi065 & ~w12840 ) | ( \pi065 & w13338 ) | ( ~w12840 & w13338 ) ;
  assign w13340 = w12838 ^ w13339 ;
  assign w13341 = ~w13002 & w13340 ;
  assign w13342 = ( w12834 & w13000 ) | ( w12834 & w13001 ) | ( w13000 & w13001 ) ;
  assign w13343 = ~w13001 & w13342 ;
  assign w13344 = w13341 | w13343 ;
  assign w13345 = ~\pi067 & w13344 ;
  assign w13346 = \pi014 ^ \pi065 ;
  assign w13347 = \pi013 ^ w12502 ;
  assign w13348 = ( \pi064 & w13002 ) | ( \pi064 & w13347 ) | ( w13002 & w13347 ) ;
  assign w13349 = w13346 ^ w13348 ;
  assign w13350 = ~w13002 & w13349 ;
  assign w13351 = w12840 & w13002 ;
  assign w13352 = w13350 | w13351 ;
  assign w13353 = ~\pi066 & w13352 ;
  assign w13354 = \pi066 ^ w13352 ;
  assign w13355 = \pi064 & ~w13002 ;
  assign w13356 = \pi013 ^ w13355 ;
  assign w13357 = ( ~\pi012 & \pi064 ) | ( ~\pi012 & w13354 ) | ( \pi064 & w13354 ) ;
  assign w13358 = ( \pi065 & ~w13356 ) | ( \pi065 & w13357 ) | ( ~w13356 & w13357 ) ;
  assign w13359 = w13354 | w13358 ;
  assign w13360 = \pi067 ^ w13344 ;
  assign w13361 = ( ~w13353 & w13359 ) | ( ~w13353 & w13360 ) | ( w13359 & w13360 ) ;
  assign w13362 = w13360 | w13361 ;
  assign w13363 = \pi068 ^ w13336 ;
  assign w13364 = ( ~w13345 & w13362 ) | ( ~w13345 & w13363 ) | ( w13362 & w13363 ) ;
  assign w13365 = w13363 | w13364 ;
  assign w13366 = \pi069 ^ w13329 ;
  assign w13367 = ( ~w13337 & w13365 ) | ( ~w13337 & w13366 ) | ( w13365 & w13366 ) ;
  assign w13368 = w13366 | w13367 ;
  assign w13369 = \pi070 ^ w13322 ;
  assign w13370 = ( ~w13330 & w13368 ) | ( ~w13330 & w13369 ) | ( w13368 & w13369 ) ;
  assign w13371 = w13369 | w13370 ;
  assign w13372 = \pi071 ^ w13315 ;
  assign w13373 = ( ~w13323 & w13371 ) | ( ~w13323 & w13372 ) | ( w13371 & w13372 ) ;
  assign w13374 = w13372 | w13373 ;
  assign w13375 = \pi072 ^ w13308 ;
  assign w13376 = ( ~w13316 & w13374 ) | ( ~w13316 & w13375 ) | ( w13374 & w13375 ) ;
  assign w13377 = w13375 | w13376 ;
  assign w13378 = \pi073 ^ w13301 ;
  assign w13379 = ( ~w13309 & w13377 ) | ( ~w13309 & w13378 ) | ( w13377 & w13378 ) ;
  assign w13380 = w13378 | w13379 ;
  assign w13381 = \pi074 ^ w13294 ;
  assign w13382 = ( ~w13302 & w13380 ) | ( ~w13302 & w13381 ) | ( w13380 & w13381 ) ;
  assign w13383 = w13381 | w13382 ;
  assign w13384 = \pi075 ^ w13287 ;
  assign w13385 = ( ~w13295 & w13383 ) | ( ~w13295 & w13384 ) | ( w13383 & w13384 ) ;
  assign w13386 = w13384 | w13385 ;
  assign w13387 = \pi076 ^ w13280 ;
  assign w13388 = ( ~w13288 & w13386 ) | ( ~w13288 & w13387 ) | ( w13386 & w13387 ) ;
  assign w13389 = w13387 | w13388 ;
  assign w13390 = \pi077 ^ w13273 ;
  assign w13391 = ( ~w13281 & w13389 ) | ( ~w13281 & w13390 ) | ( w13389 & w13390 ) ;
  assign w13392 = w13390 | w13391 ;
  assign w13393 = \pi078 ^ w13266 ;
  assign w13394 = ( ~w13274 & w13392 ) | ( ~w13274 & w13393 ) | ( w13392 & w13393 ) ;
  assign w13395 = w13393 | w13394 ;
  assign w13396 = \pi079 ^ w13259 ;
  assign w13397 = ( ~w13267 & w13395 ) | ( ~w13267 & w13396 ) | ( w13395 & w13396 ) ;
  assign w13398 = w13396 | w13397 ;
  assign w13399 = \pi080 ^ w13252 ;
  assign w13400 = ( ~w13260 & w13398 ) | ( ~w13260 & w13399 ) | ( w13398 & w13399 ) ;
  assign w13401 = w13399 | w13400 ;
  assign w13402 = \pi081 ^ w13245 ;
  assign w13403 = ( ~w13253 & w13401 ) | ( ~w13253 & w13402 ) | ( w13401 & w13402 ) ;
  assign w13404 = w13402 | w13403 ;
  assign w13405 = \pi082 ^ w13238 ;
  assign w13406 = ( ~w13246 & w13404 ) | ( ~w13246 & w13405 ) | ( w13404 & w13405 ) ;
  assign w13407 = w13405 | w13406 ;
  assign w13408 = \pi083 ^ w13231 ;
  assign w13409 = ( ~w13239 & w13407 ) | ( ~w13239 & w13408 ) | ( w13407 & w13408 ) ;
  assign w13410 = w13408 | w13409 ;
  assign w13411 = \pi084 ^ w13224 ;
  assign w13412 = ( ~w13232 & w13410 ) | ( ~w13232 & w13411 ) | ( w13410 & w13411 ) ;
  assign w13413 = w13411 | w13412 ;
  assign w13414 = \pi085 ^ w13217 ;
  assign w13415 = ( ~w13225 & w13413 ) | ( ~w13225 & w13414 ) | ( w13413 & w13414 ) ;
  assign w13416 = w13414 | w13415 ;
  assign w13417 = \pi086 ^ w13210 ;
  assign w13418 = ( ~w13218 & w13416 ) | ( ~w13218 & w13417 ) | ( w13416 & w13417 ) ;
  assign w13419 = w13417 | w13418 ;
  assign w13420 = \pi087 ^ w13203 ;
  assign w13421 = ( ~w13211 & w13419 ) | ( ~w13211 & w13420 ) | ( w13419 & w13420 ) ;
  assign w13422 = w13420 | w13421 ;
  assign w13423 = \pi088 ^ w13196 ;
  assign w13424 = ( ~w13204 & w13422 ) | ( ~w13204 & w13423 ) | ( w13422 & w13423 ) ;
  assign w13425 = w13423 | w13424 ;
  assign w13426 = \pi089 ^ w13189 ;
  assign w13427 = ( ~w13197 & w13425 ) | ( ~w13197 & w13426 ) | ( w13425 & w13426 ) ;
  assign w13428 = w13426 | w13427 ;
  assign w13429 = \pi090 ^ w13182 ;
  assign w13430 = ( ~w13190 & w13428 ) | ( ~w13190 & w13429 ) | ( w13428 & w13429 ) ;
  assign w13431 = w13429 | w13430 ;
  assign w13432 = \pi091 ^ w13175 ;
  assign w13433 = ( ~w13183 & w13431 ) | ( ~w13183 & w13432 ) | ( w13431 & w13432 ) ;
  assign w13434 = w13432 | w13433 ;
  assign w13435 = \pi092 ^ w13168 ;
  assign w13436 = ( ~w13176 & w13434 ) | ( ~w13176 & w13435 ) | ( w13434 & w13435 ) ;
  assign w13437 = w13435 | w13436 ;
  assign w13438 = \pi093 ^ w13161 ;
  assign w13439 = ( ~w13169 & w13437 ) | ( ~w13169 & w13438 ) | ( w13437 & w13438 ) ;
  assign w13440 = w13438 | w13439 ;
  assign w13441 = \pi094 ^ w13154 ;
  assign w13442 = ( ~w13162 & w13440 ) | ( ~w13162 & w13441 ) | ( w13440 & w13441 ) ;
  assign w13443 = w13441 | w13442 ;
  assign w13444 = \pi095 ^ w13147 ;
  assign w13445 = ( ~w13155 & w13443 ) | ( ~w13155 & w13444 ) | ( w13443 & w13444 ) ;
  assign w13446 = w13444 | w13445 ;
  assign w13447 = \pi096 ^ w13140 ;
  assign w13448 = ( ~w13148 & w13446 ) | ( ~w13148 & w13447 ) | ( w13446 & w13447 ) ;
  assign w13449 = w13447 | w13448 ;
  assign w13450 = \pi097 ^ w13133 ;
  assign w13451 = ( ~w13141 & w13449 ) | ( ~w13141 & w13450 ) | ( w13449 & w13450 ) ;
  assign w13452 = w13450 | w13451 ;
  assign w13453 = \pi098 ^ w13126 ;
  assign w13454 = ( ~w13134 & w13452 ) | ( ~w13134 & w13453 ) | ( w13452 & w13453 ) ;
  assign w13455 = w13453 | w13454 ;
  assign w13456 = \pi099 ^ w13119 ;
  assign w13457 = ( ~w13127 & w13455 ) | ( ~w13127 & w13456 ) | ( w13455 & w13456 ) ;
  assign w13458 = w13456 | w13457 ;
  assign w13459 = \pi100 ^ w13112 ;
  assign w13460 = ( ~w13120 & w13458 ) | ( ~w13120 & w13459 ) | ( w13458 & w13459 ) ;
  assign w13461 = w13459 | w13460 ;
  assign w13462 = \pi101 ^ w13105 ;
  assign w13463 = ( ~w13113 & w13461 ) | ( ~w13113 & w13462 ) | ( w13461 & w13462 ) ;
  assign w13464 = w13462 | w13463 ;
  assign w13465 = \pi102 ^ w13098 ;
  assign w13466 = ( ~w13106 & w13464 ) | ( ~w13106 & w13465 ) | ( w13464 & w13465 ) ;
  assign w13467 = w13465 | w13466 ;
  assign w13468 = \pi103 ^ w13091 ;
  assign w13469 = ( ~w13099 & w13467 ) | ( ~w13099 & w13468 ) | ( w13467 & w13468 ) ;
  assign w13470 = w13468 | w13469 ;
  assign w13471 = \pi104 ^ w13084 ;
  assign w13472 = ( ~w13092 & w13470 ) | ( ~w13092 & w13471 ) | ( w13470 & w13471 ) ;
  assign w13473 = w13471 | w13472 ;
  assign w13474 = \pi105 ^ w13077 ;
  assign w13475 = ( ~w13085 & w13473 ) | ( ~w13085 & w13474 ) | ( w13473 & w13474 ) ;
  assign w13476 = w13474 | w13475 ;
  assign w13477 = \pi106 ^ w13070 ;
  assign w13478 = ( ~w13078 & w13476 ) | ( ~w13078 & w13477 ) | ( w13476 & w13477 ) ;
  assign w13479 = w13477 | w13478 ;
  assign w13480 = \pi107 ^ w13063 ;
  assign w13481 = ( ~w13071 & w13479 ) | ( ~w13071 & w13480 ) | ( w13479 & w13480 ) ;
  assign w13482 = w13480 | w13481 ;
  assign w13483 = \pi108 ^ w13056 ;
  assign w13484 = ( ~w13064 & w13482 ) | ( ~w13064 & w13483 ) | ( w13482 & w13483 ) ;
  assign w13485 = w13483 | w13484 ;
  assign w13486 = \pi109 ^ w13049 ;
  assign w13487 = ( ~w13057 & w13485 ) | ( ~w13057 & w13486 ) | ( w13485 & w13486 ) ;
  assign w13488 = w13486 | w13487 ;
  assign w13489 = \pi110 ^ w13042 ;
  assign w13490 = ( ~w13050 & w13488 ) | ( ~w13050 & w13489 ) | ( w13488 & w13489 ) ;
  assign w13491 = w13489 | w13490 ;
  assign w13492 = \pi111 ^ w13035 ;
  assign w13493 = ( ~w13043 & w13491 ) | ( ~w13043 & w13492 ) | ( w13491 & w13492 ) ;
  assign w13494 = w13492 | w13493 ;
  assign w13495 = \pi112 ^ w13028 ;
  assign w13496 = ( ~w13036 & w13494 ) | ( ~w13036 & w13495 ) | ( w13494 & w13495 ) ;
  assign w13497 = w13495 | w13496 ;
  assign w13498 = \pi113 ^ w13021 ;
  assign w13499 = ( ~w13029 & w13497 ) | ( ~w13029 & w13498 ) | ( w13497 & w13498 ) ;
  assign w13500 = w13498 | w13499 ;
  assign w13501 = \pi114 ^ w13008 ;
  assign w13502 = ( ~w13022 & w13500 ) | ( ~w13022 & w13501 ) | ( w13500 & w13501 ) ;
  assign w13503 = w13501 | w13502 ;
  assign w13504 = \pi115 ^ w13014 ;
  assign w13505 = w13015 & ~w13504 ;
  assign w13506 = ( w13503 & w13504 ) | ( w13503 & ~w13505 ) | ( w13504 & ~w13505 ) ;
  assign w13507 = ~\pi115 & w13014 ;
  assign w13508 = w13506 & ~w13507 ;
  assign w13509 = w155 | w13508 ;
  assign w13510 = w13008 & w13509 ;
  assign w13511 = ~w13022 & w13500 ;
  assign w13512 = w13501 ^ w13511 ;
  assign w13513 = ~w13509 & w13512 ;
  assign w13514 = w13510 | w13513 ;
  assign w13515 = ~\pi115 & w13514 ;
  assign w13516 = w13021 & w13509 ;
  assign w13517 = ~w13029 & w13497 ;
  assign w13518 = w13498 ^ w13517 ;
  assign w13519 = ~w13509 & w13518 ;
  assign w13520 = w13516 | w13519 ;
  assign w13521 = ~\pi114 & w13520 ;
  assign w13522 = w13028 & w13509 ;
  assign w13523 = ~w13036 & w13494 ;
  assign w13524 = w13495 ^ w13523 ;
  assign w13525 = ~w13509 & w13524 ;
  assign w13526 = w13522 | w13525 ;
  assign w13527 = ~\pi113 & w13526 ;
  assign w13528 = w13035 & w13509 ;
  assign w13529 = ~w13043 & w13491 ;
  assign w13530 = w13492 ^ w13529 ;
  assign w13531 = ~w13509 & w13530 ;
  assign w13532 = w13528 | w13531 ;
  assign w13533 = ~\pi112 & w13532 ;
  assign w13534 = w13042 & w13509 ;
  assign w13535 = ~w13050 & w13488 ;
  assign w13536 = w13489 ^ w13535 ;
  assign w13537 = ~w13509 & w13536 ;
  assign w13538 = w13534 | w13537 ;
  assign w13539 = ~\pi111 & w13538 ;
  assign w13540 = w13049 & w13509 ;
  assign w13541 = ~w13057 & w13485 ;
  assign w13542 = w13486 ^ w13541 ;
  assign w13543 = ~w13509 & w13542 ;
  assign w13544 = w13540 | w13543 ;
  assign w13545 = ~\pi110 & w13544 ;
  assign w13546 = w13056 & w13509 ;
  assign w13547 = ~w13064 & w13482 ;
  assign w13548 = w13483 ^ w13547 ;
  assign w13549 = ~w13509 & w13548 ;
  assign w13550 = w13546 | w13549 ;
  assign w13551 = ~\pi109 & w13550 ;
  assign w13552 = w13063 & w13509 ;
  assign w13553 = ~w13071 & w13479 ;
  assign w13554 = w13480 ^ w13553 ;
  assign w13555 = ~w13509 & w13554 ;
  assign w13556 = w13552 | w13555 ;
  assign w13557 = ~\pi108 & w13556 ;
  assign w13558 = w13070 & w13509 ;
  assign w13559 = ~w13078 & w13476 ;
  assign w13560 = w13477 ^ w13559 ;
  assign w13561 = ~w13509 & w13560 ;
  assign w13562 = w13558 | w13561 ;
  assign w13563 = ~\pi107 & w13562 ;
  assign w13564 = w13077 & w13509 ;
  assign w13565 = ~w13085 & w13473 ;
  assign w13566 = w13474 ^ w13565 ;
  assign w13567 = ~w13509 & w13566 ;
  assign w13568 = w13564 | w13567 ;
  assign w13569 = ~\pi106 & w13568 ;
  assign w13570 = w13084 & w13509 ;
  assign w13571 = ~w13092 & w13470 ;
  assign w13572 = w13471 ^ w13571 ;
  assign w13573 = ~w13509 & w13572 ;
  assign w13574 = w13570 | w13573 ;
  assign w13575 = ~\pi105 & w13574 ;
  assign w13576 = w13091 & w13509 ;
  assign w13577 = ~w13099 & w13467 ;
  assign w13578 = w13468 ^ w13577 ;
  assign w13579 = ~w13509 & w13578 ;
  assign w13580 = w13576 | w13579 ;
  assign w13581 = ~\pi104 & w13580 ;
  assign w13582 = w13098 & w13509 ;
  assign w13583 = ~w13106 & w13464 ;
  assign w13584 = w13465 ^ w13583 ;
  assign w13585 = ~w13509 & w13584 ;
  assign w13586 = w13582 | w13585 ;
  assign w13587 = ~\pi103 & w13586 ;
  assign w13588 = w13105 & w13509 ;
  assign w13589 = ~w13113 & w13461 ;
  assign w13590 = w13462 ^ w13589 ;
  assign w13591 = ~w13509 & w13590 ;
  assign w13592 = w13588 | w13591 ;
  assign w13593 = ~\pi102 & w13592 ;
  assign w13594 = w13112 & w13509 ;
  assign w13595 = ~w13120 & w13458 ;
  assign w13596 = w13459 ^ w13595 ;
  assign w13597 = ~w13509 & w13596 ;
  assign w13598 = w13594 | w13597 ;
  assign w13599 = ~\pi101 & w13598 ;
  assign w13600 = w13119 & w13509 ;
  assign w13601 = ~w13127 & w13455 ;
  assign w13602 = w13456 ^ w13601 ;
  assign w13603 = ~w13509 & w13602 ;
  assign w13604 = w13600 | w13603 ;
  assign w13605 = ~\pi100 & w13604 ;
  assign w13606 = w13126 & w13509 ;
  assign w13607 = ~w13134 & w13452 ;
  assign w13608 = w13453 ^ w13607 ;
  assign w13609 = ~w13509 & w13608 ;
  assign w13610 = w13606 | w13609 ;
  assign w13611 = ~\pi099 & w13610 ;
  assign w13612 = w13133 & w13509 ;
  assign w13613 = ~w13141 & w13449 ;
  assign w13614 = w13450 ^ w13613 ;
  assign w13615 = ~w13509 & w13614 ;
  assign w13616 = w13612 | w13615 ;
  assign w13617 = ~\pi098 & w13616 ;
  assign w13618 = w13140 & w13509 ;
  assign w13619 = ~w13148 & w13446 ;
  assign w13620 = w13447 ^ w13619 ;
  assign w13621 = ~w13509 & w13620 ;
  assign w13622 = w13618 | w13621 ;
  assign w13623 = ~\pi097 & w13622 ;
  assign w13624 = w13147 & w13509 ;
  assign w13625 = ~w13155 & w13443 ;
  assign w13626 = w13444 ^ w13625 ;
  assign w13627 = ~w13509 & w13626 ;
  assign w13628 = w13624 | w13627 ;
  assign w13629 = ~\pi096 & w13628 ;
  assign w13630 = w13154 & w13509 ;
  assign w13631 = ~w13162 & w13440 ;
  assign w13632 = w13441 ^ w13631 ;
  assign w13633 = ~w13509 & w13632 ;
  assign w13634 = w13630 | w13633 ;
  assign w13635 = ~\pi095 & w13634 ;
  assign w13636 = w13161 & w13509 ;
  assign w13637 = ~w13169 & w13437 ;
  assign w13638 = w13438 ^ w13637 ;
  assign w13639 = ~w13509 & w13638 ;
  assign w13640 = w13636 | w13639 ;
  assign w13641 = ~\pi094 & w13640 ;
  assign w13642 = w13168 & w13509 ;
  assign w13643 = ~w13176 & w13434 ;
  assign w13644 = w13435 ^ w13643 ;
  assign w13645 = ~w13509 & w13644 ;
  assign w13646 = w13642 | w13645 ;
  assign w13647 = ~\pi093 & w13646 ;
  assign w13648 = w13175 & w13509 ;
  assign w13649 = ~w13183 & w13431 ;
  assign w13650 = w13432 ^ w13649 ;
  assign w13651 = ~w13509 & w13650 ;
  assign w13652 = w13648 | w13651 ;
  assign w13653 = ~\pi092 & w13652 ;
  assign w13654 = w13182 & w13509 ;
  assign w13655 = ~w13190 & w13428 ;
  assign w13656 = w13429 ^ w13655 ;
  assign w13657 = ~w13509 & w13656 ;
  assign w13658 = w13654 | w13657 ;
  assign w13659 = ~\pi091 & w13658 ;
  assign w13660 = w13189 & w13509 ;
  assign w13661 = ~w13197 & w13425 ;
  assign w13662 = w13426 ^ w13661 ;
  assign w13663 = ~w13509 & w13662 ;
  assign w13664 = w13660 | w13663 ;
  assign w13665 = ~\pi090 & w13664 ;
  assign w13666 = w13196 & w13509 ;
  assign w13667 = ~w13204 & w13422 ;
  assign w13668 = w13423 ^ w13667 ;
  assign w13669 = ~w13509 & w13668 ;
  assign w13670 = w13666 | w13669 ;
  assign w13671 = ~\pi089 & w13670 ;
  assign w13672 = w13203 & w13509 ;
  assign w13673 = ~w13211 & w13419 ;
  assign w13674 = w13420 ^ w13673 ;
  assign w13675 = ~w13509 & w13674 ;
  assign w13676 = w13672 | w13675 ;
  assign w13677 = ~\pi088 & w13676 ;
  assign w13678 = w13210 & w13509 ;
  assign w13679 = ~w13218 & w13416 ;
  assign w13680 = w13417 ^ w13679 ;
  assign w13681 = ~w13509 & w13680 ;
  assign w13682 = w13678 | w13681 ;
  assign w13683 = ~\pi087 & w13682 ;
  assign w13684 = w13217 & w13509 ;
  assign w13685 = ~w13225 & w13413 ;
  assign w13686 = w13414 ^ w13685 ;
  assign w13687 = ~w13509 & w13686 ;
  assign w13688 = w13684 | w13687 ;
  assign w13689 = ~\pi086 & w13688 ;
  assign w13690 = w13224 & w13509 ;
  assign w13691 = ~w13232 & w13410 ;
  assign w13692 = w13411 ^ w13691 ;
  assign w13693 = ~w13509 & w13692 ;
  assign w13694 = w13690 | w13693 ;
  assign w13695 = ~\pi085 & w13694 ;
  assign w13696 = w13231 & w13509 ;
  assign w13697 = ~w13239 & w13407 ;
  assign w13698 = w13408 ^ w13697 ;
  assign w13699 = ~w13509 & w13698 ;
  assign w13700 = w13696 | w13699 ;
  assign w13701 = ~\pi084 & w13700 ;
  assign w13702 = w13238 & w13509 ;
  assign w13703 = ~w13246 & w13404 ;
  assign w13704 = w13405 ^ w13703 ;
  assign w13705 = ~w13509 & w13704 ;
  assign w13706 = w13702 | w13705 ;
  assign w13707 = ~\pi083 & w13706 ;
  assign w13708 = w13245 & w13509 ;
  assign w13709 = ~w13253 & w13401 ;
  assign w13710 = w13402 ^ w13709 ;
  assign w13711 = ~w13509 & w13710 ;
  assign w13712 = w13708 | w13711 ;
  assign w13713 = ~\pi082 & w13712 ;
  assign w13714 = w13252 & w13509 ;
  assign w13715 = ~w13260 & w13398 ;
  assign w13716 = w13399 ^ w13715 ;
  assign w13717 = ~w13509 & w13716 ;
  assign w13718 = w13714 | w13717 ;
  assign w13719 = ~\pi081 & w13718 ;
  assign w13720 = w13259 & w13509 ;
  assign w13721 = ~w13267 & w13395 ;
  assign w13722 = w13396 ^ w13721 ;
  assign w13723 = ~w13509 & w13722 ;
  assign w13724 = w13720 | w13723 ;
  assign w13725 = ~\pi080 & w13724 ;
  assign w13726 = w13266 & w13509 ;
  assign w13727 = ~w13274 & w13392 ;
  assign w13728 = w13393 ^ w13727 ;
  assign w13729 = ~w13509 & w13728 ;
  assign w13730 = w13726 | w13729 ;
  assign w13731 = ~\pi079 & w13730 ;
  assign w13732 = w13273 & w13509 ;
  assign w13733 = ~w13281 & w13389 ;
  assign w13734 = w13390 ^ w13733 ;
  assign w13735 = ~w13509 & w13734 ;
  assign w13736 = w13732 | w13735 ;
  assign w13737 = ~\pi078 & w13736 ;
  assign w13738 = w13280 & w13509 ;
  assign w13739 = ~w13288 & w13386 ;
  assign w13740 = w13387 ^ w13739 ;
  assign w13741 = ~w13509 & w13740 ;
  assign w13742 = w13738 | w13741 ;
  assign w13743 = ~\pi077 & w13742 ;
  assign w13744 = w13287 & w13509 ;
  assign w13745 = ~w13295 & w13383 ;
  assign w13746 = w13384 ^ w13745 ;
  assign w13747 = ~w13509 & w13746 ;
  assign w13748 = w13744 | w13747 ;
  assign w13749 = ~\pi076 & w13748 ;
  assign w13750 = w13294 & w13509 ;
  assign w13751 = ~w13302 & w13380 ;
  assign w13752 = w13381 ^ w13751 ;
  assign w13753 = ~w13509 & w13752 ;
  assign w13754 = w13750 | w13753 ;
  assign w13755 = ~\pi075 & w13754 ;
  assign w13756 = w13301 & w13509 ;
  assign w13757 = ~w13309 & w13377 ;
  assign w13758 = w13378 ^ w13757 ;
  assign w13759 = ~w13509 & w13758 ;
  assign w13760 = w13756 | w13759 ;
  assign w13761 = ~\pi074 & w13760 ;
  assign w13762 = w13308 & w13509 ;
  assign w13763 = ~w13316 & w13374 ;
  assign w13764 = w13375 ^ w13763 ;
  assign w13765 = ~w13509 & w13764 ;
  assign w13766 = w13762 | w13765 ;
  assign w13767 = ~\pi073 & w13766 ;
  assign w13768 = w13315 & w13509 ;
  assign w13769 = ~w13323 & w13371 ;
  assign w13770 = w13372 ^ w13769 ;
  assign w13771 = ~w13509 & w13770 ;
  assign w13772 = w13768 | w13771 ;
  assign w13773 = ~\pi072 & w13772 ;
  assign w13774 = w13322 & w13509 ;
  assign w13775 = ~w13330 & w13368 ;
  assign w13776 = w13369 ^ w13775 ;
  assign w13777 = ~w13509 & w13776 ;
  assign w13778 = w13774 | w13777 ;
  assign w13779 = ~\pi071 & w13778 ;
  assign w13780 = w13329 & w13509 ;
  assign w13781 = ~w13337 & w13365 ;
  assign w13782 = w13366 ^ w13781 ;
  assign w13783 = ~w13509 & w13782 ;
  assign w13784 = w13780 | w13783 ;
  assign w13785 = ~\pi070 & w13784 ;
  assign w13786 = w13336 & w13509 ;
  assign w13787 = ~w13345 & w13362 ;
  assign w13788 = w13363 ^ w13787 ;
  assign w13789 = ~w13509 & w13788 ;
  assign w13790 = w13786 | w13789 ;
  assign w13791 = ~\pi069 & w13790 ;
  assign w13792 = w13344 & w13509 ;
  assign w13793 = ~w13353 & w13359 ;
  assign w13794 = w13360 ^ w13793 ;
  assign w13795 = ~w13509 & w13794 ;
  assign w13796 = w13792 | w13795 ;
  assign w13797 = ~\pi068 & w13796 ;
  assign w13798 = ~\pi012 & \pi064 ;
  assign w13799 = ( \pi065 & ~w13356 ) | ( \pi065 & w13798 ) | ( ~w13356 & w13798 ) ;
  assign w13800 = w13354 ^ w13799 ;
  assign w13801 = ( w155 & w13508 ) | ( w155 & w13800 ) | ( w13508 & w13800 ) ;
  assign w13802 = w13800 & ~w13801 ;
  assign w13803 = ( w13352 & w13509 ) | ( w13352 & w13802 ) | ( w13509 & w13802 ) ;
  assign w13804 = w13802 | w13803 ;
  assign w13805 = ~\pi067 & w13804 ;
  assign w13806 = \pi013 ^ \pi065 ;
  assign w13807 = \pi012 ^ w13002 ;
  assign w13808 = ( \pi064 & w155 ) | ( \pi064 & w13807 ) | ( w155 & w13807 ) ;
  assign w13809 = w13806 ^ w13808 ;
  assign w13810 = ~w155 & w13809 ;
  assign w13811 = ~w13508 & w13810 ;
  assign w13812 = ( ~\pi064 & w13002 ) | ( ~\pi064 & w13509 ) | ( w13002 & w13509 ) ;
  assign w13813 = \pi013 ^ w13812 ;
  assign w13814 = w13509 & ~w13813 ;
  assign w13815 = w13811 | w13814 ;
  assign w13816 = ~\pi066 & w13815 ;
  assign w13817 = ( \pi064 & w264 ) | ( \pi064 & w273 ) | ( w264 & w273 ) ;
  assign w13818 = \pi012 & \pi116 ;
  assign w13819 = ( \pi012 & w13817 ) | ( \pi012 & w13818 ) | ( w13817 & w13818 ) ;
  assign w13820 = ( \pi064 & w13508 ) | ( \pi064 & w13819 ) | ( w13508 & w13819 ) ;
  assign w13821 = ( \pi012 & ~\pi064 ) | ( \pi012 & w13820 ) | ( ~\pi064 & w13820 ) ;
  assign w13822 = ~w199 & w13798 ;
  assign w13823 = ( w153 & ~w199 ) | ( w153 & w13508 ) | ( ~w199 & w13508 ) ;
  assign w13824 = w13822 & ~w13823 ;
  assign w13825 = ~\pi011 & \pi064 ;
  assign w13826 = w13509 | w13811 ;
  assign w13827 = ( w13356 & w13811 ) | ( w13356 & w13826 ) | ( w13811 & w13826 ) ;
  assign w13828 = \pi066 ^ w13827 ;
  assign w13829 = w13821 | w13824 ;
  assign w13830 = ( \pi065 & w13825 ) | ( \pi065 & ~w13829 ) | ( w13825 & ~w13829 ) ;
  assign w13831 = w13828 | w13830 ;
  assign w13832 = ~w13352 & w13509 ;
  assign w13833 = ( w13509 & w13802 ) | ( w13509 & ~w13832 ) | ( w13802 & ~w13832 ) ;
  assign w13834 = \pi067 ^ w13833 ;
  assign w13835 = ( ~w13816 & w13831 ) | ( ~w13816 & w13834 ) | ( w13831 & w13834 ) ;
  assign w13836 = w13834 | w13835 ;
  assign w13837 = \pi068 ^ w13796 ;
  assign w13838 = ( ~w13805 & w13836 ) | ( ~w13805 & w13837 ) | ( w13836 & w13837 ) ;
  assign w13839 = w13837 | w13838 ;
  assign w13840 = \pi069 ^ w13790 ;
  assign w13841 = ( ~w13797 & w13839 ) | ( ~w13797 & w13840 ) | ( w13839 & w13840 ) ;
  assign w13842 = w13840 | w13841 ;
  assign w13843 = \pi070 ^ w13784 ;
  assign w13844 = ( ~w13791 & w13842 ) | ( ~w13791 & w13843 ) | ( w13842 & w13843 ) ;
  assign w13845 = w13843 | w13844 ;
  assign w13846 = \pi071 ^ w13778 ;
  assign w13847 = ( ~w13785 & w13845 ) | ( ~w13785 & w13846 ) | ( w13845 & w13846 ) ;
  assign w13848 = w13846 | w13847 ;
  assign w13849 = \pi072 ^ w13772 ;
  assign w13850 = ( ~w13779 & w13848 ) | ( ~w13779 & w13849 ) | ( w13848 & w13849 ) ;
  assign w13851 = w13849 | w13850 ;
  assign w13852 = \pi073 ^ w13766 ;
  assign w13853 = ( ~w13773 & w13851 ) | ( ~w13773 & w13852 ) | ( w13851 & w13852 ) ;
  assign w13854 = w13852 | w13853 ;
  assign w13855 = \pi074 ^ w13760 ;
  assign w13856 = ( ~w13767 & w13854 ) | ( ~w13767 & w13855 ) | ( w13854 & w13855 ) ;
  assign w13857 = w13855 | w13856 ;
  assign w13858 = \pi075 ^ w13754 ;
  assign w13859 = ( ~w13761 & w13857 ) | ( ~w13761 & w13858 ) | ( w13857 & w13858 ) ;
  assign w13860 = w13858 | w13859 ;
  assign w13861 = \pi076 ^ w13748 ;
  assign w13862 = ( ~w13755 & w13860 ) | ( ~w13755 & w13861 ) | ( w13860 & w13861 ) ;
  assign w13863 = w13861 | w13862 ;
  assign w13864 = \pi077 ^ w13742 ;
  assign w13865 = ( ~w13749 & w13863 ) | ( ~w13749 & w13864 ) | ( w13863 & w13864 ) ;
  assign w13866 = w13864 | w13865 ;
  assign w13867 = \pi078 ^ w13736 ;
  assign w13868 = ( ~w13743 & w13866 ) | ( ~w13743 & w13867 ) | ( w13866 & w13867 ) ;
  assign w13869 = w13867 | w13868 ;
  assign w13870 = \pi079 ^ w13730 ;
  assign w13871 = ( ~w13737 & w13869 ) | ( ~w13737 & w13870 ) | ( w13869 & w13870 ) ;
  assign w13872 = w13870 | w13871 ;
  assign w13873 = \pi080 ^ w13724 ;
  assign w13874 = ( ~w13731 & w13872 ) | ( ~w13731 & w13873 ) | ( w13872 & w13873 ) ;
  assign w13875 = w13873 | w13874 ;
  assign w13876 = \pi081 ^ w13718 ;
  assign w13877 = ( ~w13725 & w13875 ) | ( ~w13725 & w13876 ) | ( w13875 & w13876 ) ;
  assign w13878 = w13876 | w13877 ;
  assign w13879 = \pi082 ^ w13712 ;
  assign w13880 = ( ~w13719 & w13878 ) | ( ~w13719 & w13879 ) | ( w13878 & w13879 ) ;
  assign w13881 = w13879 | w13880 ;
  assign w13882 = \pi083 ^ w13706 ;
  assign w13883 = ( ~w13713 & w13881 ) | ( ~w13713 & w13882 ) | ( w13881 & w13882 ) ;
  assign w13884 = w13882 | w13883 ;
  assign w13885 = \pi084 ^ w13700 ;
  assign w13886 = ( ~w13707 & w13884 ) | ( ~w13707 & w13885 ) | ( w13884 & w13885 ) ;
  assign w13887 = w13885 | w13886 ;
  assign w13888 = \pi085 ^ w13694 ;
  assign w13889 = ( ~w13701 & w13887 ) | ( ~w13701 & w13888 ) | ( w13887 & w13888 ) ;
  assign w13890 = w13888 | w13889 ;
  assign w13891 = \pi086 ^ w13688 ;
  assign w13892 = ( ~w13695 & w13890 ) | ( ~w13695 & w13891 ) | ( w13890 & w13891 ) ;
  assign w13893 = w13891 | w13892 ;
  assign w13894 = \pi087 ^ w13682 ;
  assign w13895 = ( ~w13689 & w13893 ) | ( ~w13689 & w13894 ) | ( w13893 & w13894 ) ;
  assign w13896 = w13894 | w13895 ;
  assign w13897 = \pi088 ^ w13676 ;
  assign w13898 = ( ~w13683 & w13896 ) | ( ~w13683 & w13897 ) | ( w13896 & w13897 ) ;
  assign w13899 = w13897 | w13898 ;
  assign w13900 = \pi089 ^ w13670 ;
  assign w13901 = ( ~w13677 & w13899 ) | ( ~w13677 & w13900 ) | ( w13899 & w13900 ) ;
  assign w13902 = w13900 | w13901 ;
  assign w13903 = \pi090 ^ w13664 ;
  assign w13904 = ( ~w13671 & w13902 ) | ( ~w13671 & w13903 ) | ( w13902 & w13903 ) ;
  assign w13905 = w13903 | w13904 ;
  assign w13906 = \pi091 ^ w13658 ;
  assign w13907 = ( ~w13665 & w13905 ) | ( ~w13665 & w13906 ) | ( w13905 & w13906 ) ;
  assign w13908 = w13906 | w13907 ;
  assign w13909 = \pi092 ^ w13652 ;
  assign w13910 = ( ~w13659 & w13908 ) | ( ~w13659 & w13909 ) | ( w13908 & w13909 ) ;
  assign w13911 = w13909 | w13910 ;
  assign w13912 = \pi093 ^ w13646 ;
  assign w13913 = ( ~w13653 & w13911 ) | ( ~w13653 & w13912 ) | ( w13911 & w13912 ) ;
  assign w13914 = w13912 | w13913 ;
  assign w13915 = \pi094 ^ w13640 ;
  assign w13916 = ( ~w13647 & w13914 ) | ( ~w13647 & w13915 ) | ( w13914 & w13915 ) ;
  assign w13917 = w13915 | w13916 ;
  assign w13918 = \pi095 ^ w13634 ;
  assign w13919 = ( ~w13641 & w13917 ) | ( ~w13641 & w13918 ) | ( w13917 & w13918 ) ;
  assign w13920 = w13918 | w13919 ;
  assign w13921 = \pi096 ^ w13628 ;
  assign w13922 = ( ~w13635 & w13920 ) | ( ~w13635 & w13921 ) | ( w13920 & w13921 ) ;
  assign w13923 = w13921 | w13922 ;
  assign w13924 = \pi097 ^ w13622 ;
  assign w13925 = ( ~w13629 & w13923 ) | ( ~w13629 & w13924 ) | ( w13923 & w13924 ) ;
  assign w13926 = w13924 | w13925 ;
  assign w13927 = \pi098 ^ w13616 ;
  assign w13928 = ( ~w13623 & w13926 ) | ( ~w13623 & w13927 ) | ( w13926 & w13927 ) ;
  assign w13929 = w13927 | w13928 ;
  assign w13930 = \pi099 ^ w13610 ;
  assign w13931 = ( ~w13617 & w13929 ) | ( ~w13617 & w13930 ) | ( w13929 & w13930 ) ;
  assign w13932 = w13930 | w13931 ;
  assign w13933 = \pi100 ^ w13604 ;
  assign w13934 = ( ~w13611 & w13932 ) | ( ~w13611 & w13933 ) | ( w13932 & w13933 ) ;
  assign w13935 = w13933 | w13934 ;
  assign w13936 = \pi101 ^ w13598 ;
  assign w13937 = ( ~w13605 & w13935 ) | ( ~w13605 & w13936 ) | ( w13935 & w13936 ) ;
  assign w13938 = w13936 | w13937 ;
  assign w13939 = \pi102 ^ w13592 ;
  assign w13940 = ( ~w13599 & w13938 ) | ( ~w13599 & w13939 ) | ( w13938 & w13939 ) ;
  assign w13941 = w13939 | w13940 ;
  assign w13942 = \pi103 ^ w13586 ;
  assign w13943 = ( ~w13593 & w13941 ) | ( ~w13593 & w13942 ) | ( w13941 & w13942 ) ;
  assign w13944 = w13942 | w13943 ;
  assign w13945 = \pi104 ^ w13580 ;
  assign w13946 = ( ~w13587 & w13944 ) | ( ~w13587 & w13945 ) | ( w13944 & w13945 ) ;
  assign w13947 = w13945 | w13946 ;
  assign w13948 = \pi105 ^ w13574 ;
  assign w13949 = ( ~w13581 & w13947 ) | ( ~w13581 & w13948 ) | ( w13947 & w13948 ) ;
  assign w13950 = w13948 | w13949 ;
  assign w13951 = \pi106 ^ w13568 ;
  assign w13952 = ( ~w13575 & w13950 ) | ( ~w13575 & w13951 ) | ( w13950 & w13951 ) ;
  assign w13953 = w13951 | w13952 ;
  assign w13954 = \pi107 ^ w13562 ;
  assign w13955 = ( ~w13569 & w13953 ) | ( ~w13569 & w13954 ) | ( w13953 & w13954 ) ;
  assign w13956 = w13954 | w13955 ;
  assign w13957 = \pi108 ^ w13556 ;
  assign w13958 = ( ~w13563 & w13956 ) | ( ~w13563 & w13957 ) | ( w13956 & w13957 ) ;
  assign w13959 = w13957 | w13958 ;
  assign w13960 = \pi109 ^ w13550 ;
  assign w13961 = ( ~w13557 & w13959 ) | ( ~w13557 & w13960 ) | ( w13959 & w13960 ) ;
  assign w13962 = w13960 | w13961 ;
  assign w13963 = \pi110 ^ w13544 ;
  assign w13964 = ( ~w13551 & w13962 ) | ( ~w13551 & w13963 ) | ( w13962 & w13963 ) ;
  assign w13965 = w13963 | w13964 ;
  assign w13966 = \pi111 ^ w13538 ;
  assign w13967 = ( ~w13545 & w13965 ) | ( ~w13545 & w13966 ) | ( w13965 & w13966 ) ;
  assign w13968 = w13966 | w13967 ;
  assign w13969 = \pi112 ^ w13532 ;
  assign w13970 = ( ~w13539 & w13968 ) | ( ~w13539 & w13969 ) | ( w13968 & w13969 ) ;
  assign w13971 = w13969 | w13970 ;
  assign w13972 = \pi113 ^ w13526 ;
  assign w13973 = ( ~w13533 & w13971 ) | ( ~w13533 & w13972 ) | ( w13971 & w13972 ) ;
  assign w13974 = w13972 | w13973 ;
  assign w13975 = \pi114 ^ w13520 ;
  assign w13976 = ( ~w13527 & w13974 ) | ( ~w13527 & w13975 ) | ( w13974 & w13975 ) ;
  assign w13977 = w13975 | w13976 ;
  assign w13978 = \pi115 ^ w13514 ;
  assign w13979 = ( ~w13521 & w13977 ) | ( ~w13521 & w13978 ) | ( w13977 & w13978 ) ;
  assign w13980 = w13978 | w13979 ;
  assign w13981 = w13014 & w13509 ;
  assign w13982 = ~w13015 & w13503 ;
  assign w13983 = w13504 ^ w13982 ;
  assign w13984 = ~w13509 & w13983 ;
  assign w13985 = w13981 | w13984 ;
  assign w13986 = ~\pi116 & w13985 ;
  assign w13987 = ( \pi116 & ~w13981 ) | ( \pi116 & w13984 ) | ( ~w13981 & w13984 ) ;
  assign w13988 = ~w13984 & w13987 ;
  assign w13989 = w13986 | w13988 ;
  assign w13990 = ( ~w13515 & w13980 ) | ( ~w13515 & w13989 ) | ( w13980 & w13989 ) ;
  assign w13991 = ( w448 & ~w13989 ) | ( w448 & w13990 ) | ( ~w13989 & w13990 ) ;
  assign w13992 = w13989 | w13991 ;
  assign w13993 = ~w155 & w13985 ;
  assign w13994 = w13992 & ~w13993 ;
  assign w13995 = ~w13521 & w13977 ;
  assign w13996 = w13978 ^ w13995 ;
  assign w13997 = ~w13994 & w13996 ;
  assign w13998 = ( w13514 & w13992 ) | ( w13514 & w13993 ) | ( w13992 & w13993 ) ;
  assign w13999 = ~w13993 & w13998 ;
  assign w14000 = w13997 | w13999 ;
  assign w14001 = ~\pi116 & w14000 ;
  assign w14002 = ~w13527 & w13974 ;
  assign w14003 = w13975 ^ w14002 ;
  assign w14004 = ~w13994 & w14003 ;
  assign w14005 = ( w13520 & w13992 ) | ( w13520 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14006 = ~w13993 & w14005 ;
  assign w14007 = w14004 | w14006 ;
  assign w14008 = ~\pi115 & w14007 ;
  assign w14009 = ~w13533 & w13971 ;
  assign w14010 = w13972 ^ w14009 ;
  assign w14011 = ~w13994 & w14010 ;
  assign w14012 = ( w13526 & w13992 ) | ( w13526 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14013 = ~w13993 & w14012 ;
  assign w14014 = w14011 | w14013 ;
  assign w14015 = ~\pi114 & w14014 ;
  assign w14016 = ~w13539 & w13968 ;
  assign w14017 = w13969 ^ w14016 ;
  assign w14018 = ~w13994 & w14017 ;
  assign w14019 = ( w13532 & w13992 ) | ( w13532 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14020 = ~w13993 & w14019 ;
  assign w14021 = w14018 | w14020 ;
  assign w14022 = ~\pi113 & w14021 ;
  assign w14023 = ~w13545 & w13965 ;
  assign w14024 = w13966 ^ w14023 ;
  assign w14025 = ~w13994 & w14024 ;
  assign w14026 = ( w13538 & w13992 ) | ( w13538 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14027 = ~w13993 & w14026 ;
  assign w14028 = w14025 | w14027 ;
  assign w14029 = ~\pi112 & w14028 ;
  assign w14030 = ~w13551 & w13962 ;
  assign w14031 = w13963 ^ w14030 ;
  assign w14032 = ~w13994 & w14031 ;
  assign w14033 = ( w13544 & w13992 ) | ( w13544 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14034 = ~w13993 & w14033 ;
  assign w14035 = w14032 | w14034 ;
  assign w14036 = ~\pi111 & w14035 ;
  assign w14037 = ~w13557 & w13959 ;
  assign w14038 = w13960 ^ w14037 ;
  assign w14039 = ~w13994 & w14038 ;
  assign w14040 = ( w13550 & w13992 ) | ( w13550 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14041 = ~w13993 & w14040 ;
  assign w14042 = w14039 | w14041 ;
  assign w14043 = ~\pi110 & w14042 ;
  assign w14044 = ~w13563 & w13956 ;
  assign w14045 = w13957 ^ w14044 ;
  assign w14046 = ~w13994 & w14045 ;
  assign w14047 = ( w13556 & w13992 ) | ( w13556 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14048 = ~w13993 & w14047 ;
  assign w14049 = w14046 | w14048 ;
  assign w14050 = ~\pi109 & w14049 ;
  assign w14051 = ~w13569 & w13953 ;
  assign w14052 = w13954 ^ w14051 ;
  assign w14053 = ~w13994 & w14052 ;
  assign w14054 = ( w13562 & w13992 ) | ( w13562 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14055 = ~w13993 & w14054 ;
  assign w14056 = w14053 | w14055 ;
  assign w14057 = ~\pi108 & w14056 ;
  assign w14058 = ~w13575 & w13950 ;
  assign w14059 = w13951 ^ w14058 ;
  assign w14060 = ~w13994 & w14059 ;
  assign w14061 = ( w13568 & w13992 ) | ( w13568 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14062 = ~w13993 & w14061 ;
  assign w14063 = w14060 | w14062 ;
  assign w14064 = ~\pi107 & w14063 ;
  assign w14065 = ~w13581 & w13947 ;
  assign w14066 = w13948 ^ w14065 ;
  assign w14067 = ~w13994 & w14066 ;
  assign w14068 = ( w13574 & w13992 ) | ( w13574 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14069 = ~w13993 & w14068 ;
  assign w14070 = w14067 | w14069 ;
  assign w14071 = ~\pi106 & w14070 ;
  assign w14072 = ~w13587 & w13944 ;
  assign w14073 = w13945 ^ w14072 ;
  assign w14074 = ~w13994 & w14073 ;
  assign w14075 = ( w13580 & w13992 ) | ( w13580 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14076 = ~w13993 & w14075 ;
  assign w14077 = w14074 | w14076 ;
  assign w14078 = ~\pi105 & w14077 ;
  assign w14079 = ~w13593 & w13941 ;
  assign w14080 = w13942 ^ w14079 ;
  assign w14081 = ~w13994 & w14080 ;
  assign w14082 = ( w13586 & w13992 ) | ( w13586 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14083 = ~w13993 & w14082 ;
  assign w14084 = w14081 | w14083 ;
  assign w14085 = ~\pi104 & w14084 ;
  assign w14086 = ~w13599 & w13938 ;
  assign w14087 = w13939 ^ w14086 ;
  assign w14088 = ~w13994 & w14087 ;
  assign w14089 = ( w13592 & w13992 ) | ( w13592 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14090 = ~w13993 & w14089 ;
  assign w14091 = w14088 | w14090 ;
  assign w14092 = ~\pi103 & w14091 ;
  assign w14093 = ~w13605 & w13935 ;
  assign w14094 = w13936 ^ w14093 ;
  assign w14095 = ~w13994 & w14094 ;
  assign w14096 = ( w13598 & w13992 ) | ( w13598 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14097 = ~w13993 & w14096 ;
  assign w14098 = w14095 | w14097 ;
  assign w14099 = ~\pi102 & w14098 ;
  assign w14100 = ~w13611 & w13932 ;
  assign w14101 = w13933 ^ w14100 ;
  assign w14102 = ~w13994 & w14101 ;
  assign w14103 = ( w13604 & w13992 ) | ( w13604 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14104 = ~w13993 & w14103 ;
  assign w14105 = w14102 | w14104 ;
  assign w14106 = ~\pi101 & w14105 ;
  assign w14107 = ~w13617 & w13929 ;
  assign w14108 = w13930 ^ w14107 ;
  assign w14109 = ~w13994 & w14108 ;
  assign w14110 = ( w13610 & w13992 ) | ( w13610 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14111 = ~w13993 & w14110 ;
  assign w14112 = w14109 | w14111 ;
  assign w14113 = ~\pi100 & w14112 ;
  assign w14114 = ~w13623 & w13926 ;
  assign w14115 = w13927 ^ w14114 ;
  assign w14116 = ~w13994 & w14115 ;
  assign w14117 = ( w13616 & w13992 ) | ( w13616 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14118 = ~w13993 & w14117 ;
  assign w14119 = w14116 | w14118 ;
  assign w14120 = ~\pi099 & w14119 ;
  assign w14121 = ~w13629 & w13923 ;
  assign w14122 = w13924 ^ w14121 ;
  assign w14123 = ~w13994 & w14122 ;
  assign w14124 = ( w13622 & w13992 ) | ( w13622 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14125 = ~w13993 & w14124 ;
  assign w14126 = w14123 | w14125 ;
  assign w14127 = ~\pi098 & w14126 ;
  assign w14128 = ~w13635 & w13920 ;
  assign w14129 = w13921 ^ w14128 ;
  assign w14130 = ~w13994 & w14129 ;
  assign w14131 = ( w13628 & w13992 ) | ( w13628 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14132 = ~w13993 & w14131 ;
  assign w14133 = w14130 | w14132 ;
  assign w14134 = ~\pi097 & w14133 ;
  assign w14135 = ~w13641 & w13917 ;
  assign w14136 = w13918 ^ w14135 ;
  assign w14137 = ~w13994 & w14136 ;
  assign w14138 = ( w13634 & w13992 ) | ( w13634 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14139 = ~w13993 & w14138 ;
  assign w14140 = w14137 | w14139 ;
  assign w14141 = ~\pi096 & w14140 ;
  assign w14142 = ~w13647 & w13914 ;
  assign w14143 = w13915 ^ w14142 ;
  assign w14144 = ~w13994 & w14143 ;
  assign w14145 = ( w13640 & w13992 ) | ( w13640 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14146 = ~w13993 & w14145 ;
  assign w14147 = w14144 | w14146 ;
  assign w14148 = ~\pi095 & w14147 ;
  assign w14149 = ~w13653 & w13911 ;
  assign w14150 = w13912 ^ w14149 ;
  assign w14151 = ~w13994 & w14150 ;
  assign w14152 = ( w13646 & w13992 ) | ( w13646 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14153 = ~w13993 & w14152 ;
  assign w14154 = w14151 | w14153 ;
  assign w14155 = ~\pi094 & w14154 ;
  assign w14156 = ~w13659 & w13908 ;
  assign w14157 = w13909 ^ w14156 ;
  assign w14158 = ~w13994 & w14157 ;
  assign w14159 = ( w13652 & w13992 ) | ( w13652 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14160 = ~w13993 & w14159 ;
  assign w14161 = w14158 | w14160 ;
  assign w14162 = ~\pi093 & w14161 ;
  assign w14163 = ~w13665 & w13905 ;
  assign w14164 = w13906 ^ w14163 ;
  assign w14165 = ~w13994 & w14164 ;
  assign w14166 = ( w13658 & w13992 ) | ( w13658 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14167 = ~w13993 & w14166 ;
  assign w14168 = w14165 | w14167 ;
  assign w14169 = ~\pi092 & w14168 ;
  assign w14170 = ~w13671 & w13902 ;
  assign w14171 = w13903 ^ w14170 ;
  assign w14172 = ~w13994 & w14171 ;
  assign w14173 = ( w13664 & w13992 ) | ( w13664 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14174 = ~w13993 & w14173 ;
  assign w14175 = w14172 | w14174 ;
  assign w14176 = ~\pi091 & w14175 ;
  assign w14177 = ~w13677 & w13899 ;
  assign w14178 = w13900 ^ w14177 ;
  assign w14179 = ~w13994 & w14178 ;
  assign w14180 = ( w13670 & w13992 ) | ( w13670 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14181 = ~w13993 & w14180 ;
  assign w14182 = w14179 | w14181 ;
  assign w14183 = ~\pi090 & w14182 ;
  assign w14184 = ~w13683 & w13896 ;
  assign w14185 = w13897 ^ w14184 ;
  assign w14186 = ~w13994 & w14185 ;
  assign w14187 = ( w13676 & w13992 ) | ( w13676 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14188 = ~w13993 & w14187 ;
  assign w14189 = w14186 | w14188 ;
  assign w14190 = ~\pi089 & w14189 ;
  assign w14191 = ~w13689 & w13893 ;
  assign w14192 = w13894 ^ w14191 ;
  assign w14193 = ~w13994 & w14192 ;
  assign w14194 = ( w13682 & w13992 ) | ( w13682 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14195 = ~w13993 & w14194 ;
  assign w14196 = w14193 | w14195 ;
  assign w14197 = ~\pi088 & w14196 ;
  assign w14198 = ~w13695 & w13890 ;
  assign w14199 = w13891 ^ w14198 ;
  assign w14200 = ~w13994 & w14199 ;
  assign w14201 = ( w13688 & w13992 ) | ( w13688 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14202 = ~w13993 & w14201 ;
  assign w14203 = w14200 | w14202 ;
  assign w14204 = ~\pi087 & w14203 ;
  assign w14205 = ~w13701 & w13887 ;
  assign w14206 = w13888 ^ w14205 ;
  assign w14207 = ~w13994 & w14206 ;
  assign w14208 = ( w13694 & w13992 ) | ( w13694 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14209 = ~w13993 & w14208 ;
  assign w14210 = w14207 | w14209 ;
  assign w14211 = ~\pi086 & w14210 ;
  assign w14212 = ~w13707 & w13884 ;
  assign w14213 = w13885 ^ w14212 ;
  assign w14214 = ~w13994 & w14213 ;
  assign w14215 = ( w13700 & w13992 ) | ( w13700 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14216 = ~w13993 & w14215 ;
  assign w14217 = w14214 | w14216 ;
  assign w14218 = ~\pi085 & w14217 ;
  assign w14219 = ~w13713 & w13881 ;
  assign w14220 = w13882 ^ w14219 ;
  assign w14221 = ~w13994 & w14220 ;
  assign w14222 = ( w13706 & w13992 ) | ( w13706 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14223 = ~w13993 & w14222 ;
  assign w14224 = w14221 | w14223 ;
  assign w14225 = ~\pi084 & w14224 ;
  assign w14226 = ~w13719 & w13878 ;
  assign w14227 = w13879 ^ w14226 ;
  assign w14228 = ~w13994 & w14227 ;
  assign w14229 = ( w13712 & w13992 ) | ( w13712 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14230 = ~w13993 & w14229 ;
  assign w14231 = w14228 | w14230 ;
  assign w14232 = ~\pi083 & w14231 ;
  assign w14233 = ~w13725 & w13875 ;
  assign w14234 = w13876 ^ w14233 ;
  assign w14235 = ~w13994 & w14234 ;
  assign w14236 = ( w13718 & w13992 ) | ( w13718 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14237 = ~w13993 & w14236 ;
  assign w14238 = w14235 | w14237 ;
  assign w14239 = ~\pi082 & w14238 ;
  assign w14240 = ~w13731 & w13872 ;
  assign w14241 = w13873 ^ w14240 ;
  assign w14242 = ~w13994 & w14241 ;
  assign w14243 = ( w13724 & w13992 ) | ( w13724 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14244 = ~w13993 & w14243 ;
  assign w14245 = w14242 | w14244 ;
  assign w14246 = ~\pi081 & w14245 ;
  assign w14247 = ~w13737 & w13869 ;
  assign w14248 = w13870 ^ w14247 ;
  assign w14249 = ~w13994 & w14248 ;
  assign w14250 = ( w13730 & w13992 ) | ( w13730 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14251 = ~w13993 & w14250 ;
  assign w14252 = w14249 | w14251 ;
  assign w14253 = ~\pi080 & w14252 ;
  assign w14254 = ~w13743 & w13866 ;
  assign w14255 = w13867 ^ w14254 ;
  assign w14256 = ~w13994 & w14255 ;
  assign w14257 = ( w13736 & w13992 ) | ( w13736 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14258 = ~w13993 & w14257 ;
  assign w14259 = w14256 | w14258 ;
  assign w14260 = ~\pi079 & w14259 ;
  assign w14261 = ~w13749 & w13863 ;
  assign w14262 = w13864 ^ w14261 ;
  assign w14263 = ~w13994 & w14262 ;
  assign w14264 = ( w13742 & w13992 ) | ( w13742 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14265 = ~w13993 & w14264 ;
  assign w14266 = w14263 | w14265 ;
  assign w14267 = ~\pi078 & w14266 ;
  assign w14268 = ~w13755 & w13860 ;
  assign w14269 = w13861 ^ w14268 ;
  assign w14270 = ~w13994 & w14269 ;
  assign w14271 = ( w13748 & w13992 ) | ( w13748 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14272 = ~w13993 & w14271 ;
  assign w14273 = w14270 | w14272 ;
  assign w14274 = ~\pi077 & w14273 ;
  assign w14275 = ~w13761 & w13857 ;
  assign w14276 = w13858 ^ w14275 ;
  assign w14277 = ~w13994 & w14276 ;
  assign w14278 = ( w13754 & w13992 ) | ( w13754 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14279 = ~w13993 & w14278 ;
  assign w14280 = w14277 | w14279 ;
  assign w14281 = ~\pi076 & w14280 ;
  assign w14282 = ~w13767 & w13854 ;
  assign w14283 = w13855 ^ w14282 ;
  assign w14284 = ~w13994 & w14283 ;
  assign w14285 = ( w13760 & w13992 ) | ( w13760 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14286 = ~w13993 & w14285 ;
  assign w14287 = w14284 | w14286 ;
  assign w14288 = ~\pi075 & w14287 ;
  assign w14289 = ~w13773 & w13851 ;
  assign w14290 = w13852 ^ w14289 ;
  assign w14291 = ~w13994 & w14290 ;
  assign w14292 = ( w13766 & w13992 ) | ( w13766 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14293 = ~w13993 & w14292 ;
  assign w14294 = w14291 | w14293 ;
  assign w14295 = ~\pi074 & w14294 ;
  assign w14296 = ~w13779 & w13848 ;
  assign w14297 = w13849 ^ w14296 ;
  assign w14298 = ~w13994 & w14297 ;
  assign w14299 = ( w13772 & w13992 ) | ( w13772 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14300 = ~w13993 & w14299 ;
  assign w14301 = w14298 | w14300 ;
  assign w14302 = ~\pi073 & w14301 ;
  assign w14303 = ~w13785 & w13845 ;
  assign w14304 = w13846 ^ w14303 ;
  assign w14305 = ~w13994 & w14304 ;
  assign w14306 = ( w13778 & w13992 ) | ( w13778 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14307 = ~w13993 & w14306 ;
  assign w14308 = w14305 | w14307 ;
  assign w14309 = ~\pi072 & w14308 ;
  assign w14310 = ~w13791 & w13842 ;
  assign w14311 = w13843 ^ w14310 ;
  assign w14312 = ~w13994 & w14311 ;
  assign w14313 = ( w13784 & w13992 ) | ( w13784 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14314 = ~w13993 & w14313 ;
  assign w14315 = w14312 | w14314 ;
  assign w14316 = ~\pi071 & w14315 ;
  assign w14317 = ~w13797 & w13839 ;
  assign w14318 = w13840 ^ w14317 ;
  assign w14319 = ~w13994 & w14318 ;
  assign w14320 = ( w13790 & w13992 ) | ( w13790 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14321 = ~w13993 & w14320 ;
  assign w14322 = w14319 | w14321 ;
  assign w14323 = ~\pi070 & w14322 ;
  assign w14324 = ~w13805 & w13836 ;
  assign w14325 = w13837 ^ w14324 ;
  assign w14326 = ~w13994 & w14325 ;
  assign w14327 = ( w13796 & w13992 ) | ( w13796 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14328 = ~w13993 & w14327 ;
  assign w14329 = w14326 | w14328 ;
  assign w14330 = ~\pi069 & w14329 ;
  assign w14331 = ~w13816 & w13831 ;
  assign w14332 = w13834 ^ w14331 ;
  assign w14333 = ~w13994 & w14332 ;
  assign w14334 = ( w13804 & w13992 ) | ( w13804 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14335 = ~w13993 & w14334 ;
  assign w14336 = w14333 | w14335 ;
  assign w14337 = ~\pi068 & w14336 ;
  assign w14338 = w13828 ^ w13830 ;
  assign w14339 = ~w13994 & w14338 ;
  assign w14340 = ( w13815 & w13992 ) | ( w13815 & w13993 ) | ( w13992 & w13993 ) ;
  assign w14341 = ~w13993 & w14340 ;
  assign w14342 = w14339 | w14341 ;
  assign w14343 = ~\pi067 & w14342 ;
  assign w14344 = w13825 ^ w13829 ;
  assign w14345 = \pi065 ^ w14344 ;
  assign w14346 = w13994 ^ w14345 ;
  assign w14347 = ( w13829 & w14345 ) | ( w13829 & w14346 ) | ( w14345 & w14346 ) ;
  assign w14348 = ~\pi066 & w14347 ;
  assign w14349 = w13829 ^ w13994 ;
  assign w14350 = ( w13829 & w14345 ) | ( w13829 & ~w14349 ) | ( w14345 & ~w14349 ) ;
  assign w14351 = \pi066 ^ w14350 ;
  assign w14352 = \pi064 & ~w13994 ;
  assign w14353 = \pi011 ^ w14352 ;
  assign w14354 = ( ~\pi010 & \pi064 ) | ( ~\pi010 & w14351 ) | ( \pi064 & w14351 ) ;
  assign w14355 = ( \pi065 & ~w14353 ) | ( \pi065 & w14354 ) | ( ~w14353 & w14354 ) ;
  assign w14356 = w14351 | w14355 ;
  assign w14357 = \pi067 ^ w14342 ;
  assign w14358 = ( ~w14348 & w14356 ) | ( ~w14348 & w14357 ) | ( w14356 & w14357 ) ;
  assign w14359 = w14357 | w14358 ;
  assign w14360 = \pi068 ^ w14336 ;
  assign w14361 = ( ~w14343 & w14359 ) | ( ~w14343 & w14360 ) | ( w14359 & w14360 ) ;
  assign w14362 = w14360 | w14361 ;
  assign w14363 = \pi069 ^ w14329 ;
  assign w14364 = ( ~w14337 & w14362 ) | ( ~w14337 & w14363 ) | ( w14362 & w14363 ) ;
  assign w14365 = w14363 | w14364 ;
  assign w14366 = \pi070 ^ w14322 ;
  assign w14367 = ( ~w14330 & w14365 ) | ( ~w14330 & w14366 ) | ( w14365 & w14366 ) ;
  assign w14368 = w14366 | w14367 ;
  assign w14369 = \pi071 ^ w14315 ;
  assign w14370 = ( ~w14323 & w14368 ) | ( ~w14323 & w14369 ) | ( w14368 & w14369 ) ;
  assign w14371 = w14369 | w14370 ;
  assign w14372 = \pi072 ^ w14308 ;
  assign w14373 = ( ~w14316 & w14371 ) | ( ~w14316 & w14372 ) | ( w14371 & w14372 ) ;
  assign w14374 = w14372 | w14373 ;
  assign w14375 = \pi073 ^ w14301 ;
  assign w14376 = ( ~w14309 & w14374 ) | ( ~w14309 & w14375 ) | ( w14374 & w14375 ) ;
  assign w14377 = w14375 | w14376 ;
  assign w14378 = \pi074 ^ w14294 ;
  assign w14379 = ( ~w14302 & w14377 ) | ( ~w14302 & w14378 ) | ( w14377 & w14378 ) ;
  assign w14380 = w14378 | w14379 ;
  assign w14381 = \pi075 ^ w14287 ;
  assign w14382 = ( ~w14295 & w14380 ) | ( ~w14295 & w14381 ) | ( w14380 & w14381 ) ;
  assign w14383 = w14381 | w14382 ;
  assign w14384 = \pi076 ^ w14280 ;
  assign w14385 = ( ~w14288 & w14383 ) | ( ~w14288 & w14384 ) | ( w14383 & w14384 ) ;
  assign w14386 = w14384 | w14385 ;
  assign w14387 = \pi077 ^ w14273 ;
  assign w14388 = ( ~w14281 & w14386 ) | ( ~w14281 & w14387 ) | ( w14386 & w14387 ) ;
  assign w14389 = w14387 | w14388 ;
  assign w14390 = \pi078 ^ w14266 ;
  assign w14391 = ( ~w14274 & w14389 ) | ( ~w14274 & w14390 ) | ( w14389 & w14390 ) ;
  assign w14392 = w14390 | w14391 ;
  assign w14393 = \pi079 ^ w14259 ;
  assign w14394 = ( ~w14267 & w14392 ) | ( ~w14267 & w14393 ) | ( w14392 & w14393 ) ;
  assign w14395 = w14393 | w14394 ;
  assign w14396 = \pi080 ^ w14252 ;
  assign w14397 = ( ~w14260 & w14395 ) | ( ~w14260 & w14396 ) | ( w14395 & w14396 ) ;
  assign w14398 = w14396 | w14397 ;
  assign w14399 = \pi081 ^ w14245 ;
  assign w14400 = ( ~w14253 & w14398 ) | ( ~w14253 & w14399 ) | ( w14398 & w14399 ) ;
  assign w14401 = w14399 | w14400 ;
  assign w14402 = \pi082 ^ w14238 ;
  assign w14403 = ( ~w14246 & w14401 ) | ( ~w14246 & w14402 ) | ( w14401 & w14402 ) ;
  assign w14404 = w14402 | w14403 ;
  assign w14405 = \pi083 ^ w14231 ;
  assign w14406 = ( ~w14239 & w14404 ) | ( ~w14239 & w14405 ) | ( w14404 & w14405 ) ;
  assign w14407 = w14405 | w14406 ;
  assign w14408 = \pi084 ^ w14224 ;
  assign w14409 = ( ~w14232 & w14407 ) | ( ~w14232 & w14408 ) | ( w14407 & w14408 ) ;
  assign w14410 = w14408 | w14409 ;
  assign w14411 = \pi085 ^ w14217 ;
  assign w14412 = ( ~w14225 & w14410 ) | ( ~w14225 & w14411 ) | ( w14410 & w14411 ) ;
  assign w14413 = w14411 | w14412 ;
  assign w14414 = \pi086 ^ w14210 ;
  assign w14415 = ( ~w14218 & w14413 ) | ( ~w14218 & w14414 ) | ( w14413 & w14414 ) ;
  assign w14416 = w14414 | w14415 ;
  assign w14417 = \pi087 ^ w14203 ;
  assign w14418 = ( ~w14211 & w14416 ) | ( ~w14211 & w14417 ) | ( w14416 & w14417 ) ;
  assign w14419 = w14417 | w14418 ;
  assign w14420 = \pi088 ^ w14196 ;
  assign w14421 = ( ~w14204 & w14419 ) | ( ~w14204 & w14420 ) | ( w14419 & w14420 ) ;
  assign w14422 = w14420 | w14421 ;
  assign w14423 = \pi089 ^ w14189 ;
  assign w14424 = ( ~w14197 & w14422 ) | ( ~w14197 & w14423 ) | ( w14422 & w14423 ) ;
  assign w14425 = w14423 | w14424 ;
  assign w14426 = \pi090 ^ w14182 ;
  assign w14427 = ( ~w14190 & w14425 ) | ( ~w14190 & w14426 ) | ( w14425 & w14426 ) ;
  assign w14428 = w14426 | w14427 ;
  assign w14429 = \pi091 ^ w14175 ;
  assign w14430 = ( ~w14183 & w14428 ) | ( ~w14183 & w14429 ) | ( w14428 & w14429 ) ;
  assign w14431 = w14429 | w14430 ;
  assign w14432 = \pi092 ^ w14168 ;
  assign w14433 = ( ~w14176 & w14431 ) | ( ~w14176 & w14432 ) | ( w14431 & w14432 ) ;
  assign w14434 = w14432 | w14433 ;
  assign w14435 = \pi093 ^ w14161 ;
  assign w14436 = ( ~w14169 & w14434 ) | ( ~w14169 & w14435 ) | ( w14434 & w14435 ) ;
  assign w14437 = w14435 | w14436 ;
  assign w14438 = \pi094 ^ w14154 ;
  assign w14439 = ( ~w14162 & w14437 ) | ( ~w14162 & w14438 ) | ( w14437 & w14438 ) ;
  assign w14440 = w14438 | w14439 ;
  assign w14441 = \pi095 ^ w14147 ;
  assign w14442 = ( ~w14155 & w14440 ) | ( ~w14155 & w14441 ) | ( w14440 & w14441 ) ;
  assign w14443 = w14441 | w14442 ;
  assign w14444 = \pi096 ^ w14140 ;
  assign w14445 = ( ~w14148 & w14443 ) | ( ~w14148 & w14444 ) | ( w14443 & w14444 ) ;
  assign w14446 = w14444 | w14445 ;
  assign w14447 = \pi097 ^ w14133 ;
  assign w14448 = ( ~w14141 & w14446 ) | ( ~w14141 & w14447 ) | ( w14446 & w14447 ) ;
  assign w14449 = w14447 | w14448 ;
  assign w14450 = \pi098 ^ w14126 ;
  assign w14451 = ( ~w14134 & w14449 ) | ( ~w14134 & w14450 ) | ( w14449 & w14450 ) ;
  assign w14452 = w14450 | w14451 ;
  assign w14453 = \pi099 ^ w14119 ;
  assign w14454 = ( ~w14127 & w14452 ) | ( ~w14127 & w14453 ) | ( w14452 & w14453 ) ;
  assign w14455 = w14453 | w14454 ;
  assign w14456 = \pi100 ^ w14112 ;
  assign w14457 = ( ~w14120 & w14455 ) | ( ~w14120 & w14456 ) | ( w14455 & w14456 ) ;
  assign w14458 = w14456 | w14457 ;
  assign w14459 = \pi101 ^ w14105 ;
  assign w14460 = ( ~w14113 & w14458 ) | ( ~w14113 & w14459 ) | ( w14458 & w14459 ) ;
  assign w14461 = w14459 | w14460 ;
  assign w14462 = \pi102 ^ w14098 ;
  assign w14463 = ( ~w14106 & w14461 ) | ( ~w14106 & w14462 ) | ( w14461 & w14462 ) ;
  assign w14464 = w14462 | w14463 ;
  assign w14465 = \pi103 ^ w14091 ;
  assign w14466 = ( ~w14099 & w14464 ) | ( ~w14099 & w14465 ) | ( w14464 & w14465 ) ;
  assign w14467 = w14465 | w14466 ;
  assign w14468 = \pi104 ^ w14084 ;
  assign w14469 = ( ~w14092 & w14467 ) | ( ~w14092 & w14468 ) | ( w14467 & w14468 ) ;
  assign w14470 = w14468 | w14469 ;
  assign w14471 = \pi105 ^ w14077 ;
  assign w14472 = ( ~w14085 & w14470 ) | ( ~w14085 & w14471 ) | ( w14470 & w14471 ) ;
  assign w14473 = w14471 | w14472 ;
  assign w14474 = \pi106 ^ w14070 ;
  assign w14475 = ( ~w14078 & w14473 ) | ( ~w14078 & w14474 ) | ( w14473 & w14474 ) ;
  assign w14476 = w14474 | w14475 ;
  assign w14477 = \pi107 ^ w14063 ;
  assign w14478 = ( ~w14071 & w14476 ) | ( ~w14071 & w14477 ) | ( w14476 & w14477 ) ;
  assign w14479 = w14477 | w14478 ;
  assign w14480 = \pi108 ^ w14056 ;
  assign w14481 = ( ~w14064 & w14479 ) | ( ~w14064 & w14480 ) | ( w14479 & w14480 ) ;
  assign w14482 = w14480 | w14481 ;
  assign w14483 = \pi109 ^ w14049 ;
  assign w14484 = ( ~w14057 & w14482 ) | ( ~w14057 & w14483 ) | ( w14482 & w14483 ) ;
  assign w14485 = w14483 | w14484 ;
  assign w14486 = \pi110 ^ w14042 ;
  assign w14487 = ( ~w14050 & w14485 ) | ( ~w14050 & w14486 ) | ( w14485 & w14486 ) ;
  assign w14488 = w14486 | w14487 ;
  assign w14489 = \pi111 ^ w14035 ;
  assign w14490 = ( ~w14043 & w14488 ) | ( ~w14043 & w14489 ) | ( w14488 & w14489 ) ;
  assign w14491 = w14489 | w14490 ;
  assign w14492 = \pi112 ^ w14028 ;
  assign w14493 = ( ~w14036 & w14491 ) | ( ~w14036 & w14492 ) | ( w14491 & w14492 ) ;
  assign w14494 = w14492 | w14493 ;
  assign w14495 = \pi113 ^ w14021 ;
  assign w14496 = ( ~w14029 & w14494 ) | ( ~w14029 & w14495 ) | ( w14494 & w14495 ) ;
  assign w14497 = w14495 | w14496 ;
  assign w14498 = \pi114 ^ w14014 ;
  assign w14499 = ( ~w14022 & w14497 ) | ( ~w14022 & w14498 ) | ( w14497 & w14498 ) ;
  assign w14500 = w14498 | w14499 ;
  assign w14501 = \pi115 ^ w14007 ;
  assign w14502 = ( ~w14015 & w14500 ) | ( ~w14015 & w14501 ) | ( w14500 & w14501 ) ;
  assign w14503 = w14501 | w14502 ;
  assign w14504 = \pi116 ^ w14000 ;
  assign w14505 = ( ~w14008 & w14503 ) | ( ~w14008 & w14504 ) | ( w14503 & w14504 ) ;
  assign w14506 = w14504 | w14505 ;
  assign w14507 = ( ~w13515 & w13980 ) | ( ~w13515 & w13994 ) | ( w13980 & w13994 ) ;
  assign w14508 = w13989 ^ w14507 ;
  assign w14509 = ~w13994 & w14508 ;
  assign w14510 = ( w155 & ~w13985 ) | ( w155 & w13992 ) | ( ~w13985 & w13992 ) ;
  assign w14511 = w13985 & w14510 ;
  assign w14512 = w14509 | w14511 ;
  assign w14513 = ~\pi117 & w14512 ;
  assign w14514 = ( \pi117 & ~w14509 ) | ( \pi117 & w14511 ) | ( ~w14509 & w14511 ) ;
  assign w14515 = ~w14511 & w14514 ;
  assign w14516 = \pi119 | w150 ;
  assign w14517 = ( \pi118 & w147 ) | ( \pi118 & ~w150 ) | ( w147 & ~w150 ) ;
  assign w14518 = w14516 | w14517 ;
  assign w14519 = w14513 | w14515 ;
  assign w14520 = ( ~w14001 & w14506 ) | ( ~w14001 & w14519 ) | ( w14506 & w14519 ) ;
  assign w14521 = ( w14518 & ~w14519 ) | ( w14518 & w14520 ) | ( ~w14519 & w14520 ) ;
  assign w14522 = w14519 | w14521 ;
  assign w14523 = ~w448 & w14512 ;
  assign w14524 = w14522 & ~w14523 ;
  assign w14525 = ~w14008 & w14503 ;
  assign w14526 = w14504 ^ w14525 ;
  assign w14527 = ~w14524 & w14526 ;
  assign w14528 = ( w14000 & w14522 ) | ( w14000 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14529 = ~w14523 & w14528 ;
  assign w14530 = w14527 | w14529 ;
  assign w14531 = ( ~w14001 & w14506 ) | ( ~w14001 & w14524 ) | ( w14506 & w14524 ) ;
  assign w14532 = w14519 ^ w14531 ;
  assign w14533 = ~w14524 & w14532 ;
  assign w14534 = ( w448 & ~w14512 ) | ( w448 & w14522 ) | ( ~w14512 & w14522 ) ;
  assign w14535 = w14512 & w14534 ;
  assign w14536 = w14533 | w14535 ;
  assign w14537 = ~\pi117 & w14530 ;
  assign w14538 = ~w14015 & w14500 ;
  assign w14539 = w14501 ^ w14538 ;
  assign w14540 = ~w14524 & w14539 ;
  assign w14541 = ( w14007 & w14522 ) | ( w14007 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14542 = ~w14523 & w14541 ;
  assign w14543 = w14540 | w14542 ;
  assign w14544 = ~\pi116 & w14543 ;
  assign w14545 = ~w14022 & w14497 ;
  assign w14546 = w14498 ^ w14545 ;
  assign w14547 = ~w14524 & w14546 ;
  assign w14548 = ( w14014 & w14522 ) | ( w14014 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14549 = ~w14523 & w14548 ;
  assign w14550 = w14547 | w14549 ;
  assign w14551 = ~\pi115 & w14550 ;
  assign w14552 = ~w14029 & w14494 ;
  assign w14553 = w14495 ^ w14552 ;
  assign w14554 = ~w14524 & w14553 ;
  assign w14555 = ( w14021 & w14522 ) | ( w14021 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14556 = ~w14523 & w14555 ;
  assign w14557 = w14554 | w14556 ;
  assign w14558 = ~\pi114 & w14557 ;
  assign w14559 = ~w14036 & w14491 ;
  assign w14560 = w14492 ^ w14559 ;
  assign w14561 = ~w14524 & w14560 ;
  assign w14562 = ( w14028 & w14522 ) | ( w14028 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14563 = ~w14523 & w14562 ;
  assign w14564 = w14561 | w14563 ;
  assign w14565 = ~\pi113 & w14564 ;
  assign w14566 = ~w14043 & w14488 ;
  assign w14567 = w14489 ^ w14566 ;
  assign w14568 = ~w14524 & w14567 ;
  assign w14569 = ( w14035 & w14522 ) | ( w14035 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14570 = ~w14523 & w14569 ;
  assign w14571 = w14568 | w14570 ;
  assign w14572 = ~\pi112 & w14571 ;
  assign w14573 = ~w14050 & w14485 ;
  assign w14574 = w14486 ^ w14573 ;
  assign w14575 = ~w14524 & w14574 ;
  assign w14576 = ( w14042 & w14522 ) | ( w14042 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14577 = ~w14523 & w14576 ;
  assign w14578 = w14575 | w14577 ;
  assign w14579 = ~\pi111 & w14578 ;
  assign w14580 = ~w14057 & w14482 ;
  assign w14581 = w14483 ^ w14580 ;
  assign w14582 = ~w14524 & w14581 ;
  assign w14583 = ( w14049 & w14522 ) | ( w14049 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14584 = ~w14523 & w14583 ;
  assign w14585 = w14582 | w14584 ;
  assign w14586 = ~\pi110 & w14585 ;
  assign w14587 = ~w14064 & w14479 ;
  assign w14588 = w14480 ^ w14587 ;
  assign w14589 = ~w14524 & w14588 ;
  assign w14590 = ( w14056 & w14522 ) | ( w14056 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14591 = ~w14523 & w14590 ;
  assign w14592 = w14589 | w14591 ;
  assign w14593 = ~\pi109 & w14592 ;
  assign w14594 = ~w14071 & w14476 ;
  assign w14595 = w14477 ^ w14594 ;
  assign w14596 = ~w14524 & w14595 ;
  assign w14597 = ( w14063 & w14522 ) | ( w14063 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14598 = ~w14523 & w14597 ;
  assign w14599 = w14596 | w14598 ;
  assign w14600 = ~\pi108 & w14599 ;
  assign w14601 = ~w14078 & w14473 ;
  assign w14602 = w14474 ^ w14601 ;
  assign w14603 = ~w14524 & w14602 ;
  assign w14604 = ( w14070 & w14522 ) | ( w14070 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14605 = ~w14523 & w14604 ;
  assign w14606 = w14603 | w14605 ;
  assign w14607 = ~\pi107 & w14606 ;
  assign w14608 = ~w14085 & w14470 ;
  assign w14609 = w14471 ^ w14608 ;
  assign w14610 = ~w14524 & w14609 ;
  assign w14611 = ( w14077 & w14522 ) | ( w14077 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14612 = ~w14523 & w14611 ;
  assign w14613 = w14610 | w14612 ;
  assign w14614 = ~\pi106 & w14613 ;
  assign w14615 = ~w14092 & w14467 ;
  assign w14616 = w14468 ^ w14615 ;
  assign w14617 = ~w14524 & w14616 ;
  assign w14618 = ( w14084 & w14522 ) | ( w14084 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14619 = ~w14523 & w14618 ;
  assign w14620 = w14617 | w14619 ;
  assign w14621 = ~\pi105 & w14620 ;
  assign w14622 = ~w14099 & w14464 ;
  assign w14623 = w14465 ^ w14622 ;
  assign w14624 = ~w14524 & w14623 ;
  assign w14625 = ( w14091 & w14522 ) | ( w14091 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14626 = ~w14523 & w14625 ;
  assign w14627 = w14624 | w14626 ;
  assign w14628 = ~\pi104 & w14627 ;
  assign w14629 = ~w14106 & w14461 ;
  assign w14630 = w14462 ^ w14629 ;
  assign w14631 = ~w14524 & w14630 ;
  assign w14632 = ( w14098 & w14522 ) | ( w14098 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14633 = ~w14523 & w14632 ;
  assign w14634 = w14631 | w14633 ;
  assign w14635 = ~\pi103 & w14634 ;
  assign w14636 = ~w14113 & w14458 ;
  assign w14637 = w14459 ^ w14636 ;
  assign w14638 = ~w14524 & w14637 ;
  assign w14639 = ( w14105 & w14522 ) | ( w14105 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14640 = ~w14523 & w14639 ;
  assign w14641 = w14638 | w14640 ;
  assign w14642 = ~\pi102 & w14641 ;
  assign w14643 = ~w14120 & w14455 ;
  assign w14644 = w14456 ^ w14643 ;
  assign w14645 = ~w14524 & w14644 ;
  assign w14646 = ( w14112 & w14522 ) | ( w14112 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14647 = ~w14523 & w14646 ;
  assign w14648 = w14645 | w14647 ;
  assign w14649 = ~\pi101 & w14648 ;
  assign w14650 = ~w14127 & w14452 ;
  assign w14651 = w14453 ^ w14650 ;
  assign w14652 = ~w14524 & w14651 ;
  assign w14653 = ( w14119 & w14522 ) | ( w14119 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14654 = ~w14523 & w14653 ;
  assign w14655 = w14652 | w14654 ;
  assign w14656 = ~\pi100 & w14655 ;
  assign w14657 = ~w14134 & w14449 ;
  assign w14658 = w14450 ^ w14657 ;
  assign w14659 = ~w14524 & w14658 ;
  assign w14660 = ( w14126 & w14522 ) | ( w14126 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14661 = ~w14523 & w14660 ;
  assign w14662 = w14659 | w14661 ;
  assign w14663 = ~\pi099 & w14662 ;
  assign w14664 = ~w14141 & w14446 ;
  assign w14665 = w14447 ^ w14664 ;
  assign w14666 = ~w14524 & w14665 ;
  assign w14667 = ( w14133 & w14522 ) | ( w14133 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14668 = ~w14523 & w14667 ;
  assign w14669 = w14666 | w14668 ;
  assign w14670 = ~\pi098 & w14669 ;
  assign w14671 = ~w14148 & w14443 ;
  assign w14672 = w14444 ^ w14671 ;
  assign w14673 = ~w14524 & w14672 ;
  assign w14674 = ( w14140 & w14522 ) | ( w14140 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14675 = ~w14523 & w14674 ;
  assign w14676 = w14673 | w14675 ;
  assign w14677 = ~\pi097 & w14676 ;
  assign w14678 = ~w14155 & w14440 ;
  assign w14679 = w14441 ^ w14678 ;
  assign w14680 = ~w14524 & w14679 ;
  assign w14681 = ( w14147 & w14522 ) | ( w14147 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14682 = ~w14523 & w14681 ;
  assign w14683 = w14680 | w14682 ;
  assign w14684 = ~\pi096 & w14683 ;
  assign w14685 = ~w14162 & w14437 ;
  assign w14686 = w14438 ^ w14685 ;
  assign w14687 = ~w14524 & w14686 ;
  assign w14688 = ( w14154 & w14522 ) | ( w14154 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14689 = ~w14523 & w14688 ;
  assign w14690 = w14687 | w14689 ;
  assign w14691 = ~\pi095 & w14690 ;
  assign w14692 = ~w14169 & w14434 ;
  assign w14693 = w14435 ^ w14692 ;
  assign w14694 = ~w14524 & w14693 ;
  assign w14695 = ( w14161 & w14522 ) | ( w14161 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14696 = ~w14523 & w14695 ;
  assign w14697 = w14694 | w14696 ;
  assign w14698 = ~\pi094 & w14697 ;
  assign w14699 = ~w14176 & w14431 ;
  assign w14700 = w14432 ^ w14699 ;
  assign w14701 = ~w14524 & w14700 ;
  assign w14702 = ( w14168 & w14522 ) | ( w14168 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14703 = ~w14523 & w14702 ;
  assign w14704 = w14701 | w14703 ;
  assign w14705 = ~\pi093 & w14704 ;
  assign w14706 = ~w14183 & w14428 ;
  assign w14707 = w14429 ^ w14706 ;
  assign w14708 = ~w14524 & w14707 ;
  assign w14709 = ( w14175 & w14522 ) | ( w14175 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14710 = ~w14523 & w14709 ;
  assign w14711 = w14708 | w14710 ;
  assign w14712 = ~\pi092 & w14711 ;
  assign w14713 = ~w14190 & w14425 ;
  assign w14714 = w14426 ^ w14713 ;
  assign w14715 = ~w14524 & w14714 ;
  assign w14716 = ( w14182 & w14522 ) | ( w14182 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14717 = ~w14523 & w14716 ;
  assign w14718 = w14715 | w14717 ;
  assign w14719 = ~\pi091 & w14718 ;
  assign w14720 = ~w14197 & w14422 ;
  assign w14721 = w14423 ^ w14720 ;
  assign w14722 = ~w14524 & w14721 ;
  assign w14723 = ( w14189 & w14522 ) | ( w14189 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14724 = ~w14523 & w14723 ;
  assign w14725 = w14722 | w14724 ;
  assign w14726 = ~\pi090 & w14725 ;
  assign w14727 = ~w14204 & w14419 ;
  assign w14728 = w14420 ^ w14727 ;
  assign w14729 = ~w14524 & w14728 ;
  assign w14730 = ( w14196 & w14522 ) | ( w14196 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14731 = ~w14523 & w14730 ;
  assign w14732 = w14729 | w14731 ;
  assign w14733 = ~\pi089 & w14732 ;
  assign w14734 = ~w14211 & w14416 ;
  assign w14735 = w14417 ^ w14734 ;
  assign w14736 = ~w14524 & w14735 ;
  assign w14737 = ( w14203 & w14522 ) | ( w14203 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14738 = ~w14523 & w14737 ;
  assign w14739 = w14736 | w14738 ;
  assign w14740 = ~\pi088 & w14739 ;
  assign w14741 = ~w14218 & w14413 ;
  assign w14742 = w14414 ^ w14741 ;
  assign w14743 = ~w14524 & w14742 ;
  assign w14744 = ( w14210 & w14522 ) | ( w14210 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14745 = ~w14523 & w14744 ;
  assign w14746 = w14743 | w14745 ;
  assign w14747 = ~\pi087 & w14746 ;
  assign w14748 = ~w14225 & w14410 ;
  assign w14749 = w14411 ^ w14748 ;
  assign w14750 = ~w14524 & w14749 ;
  assign w14751 = ( w14217 & w14522 ) | ( w14217 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14752 = ~w14523 & w14751 ;
  assign w14753 = w14750 | w14752 ;
  assign w14754 = ~\pi086 & w14753 ;
  assign w14755 = ~w14232 & w14407 ;
  assign w14756 = w14408 ^ w14755 ;
  assign w14757 = ~w14524 & w14756 ;
  assign w14758 = ( w14224 & w14522 ) | ( w14224 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14759 = ~w14523 & w14758 ;
  assign w14760 = w14757 | w14759 ;
  assign w14761 = ~\pi085 & w14760 ;
  assign w14762 = ~w14239 & w14404 ;
  assign w14763 = w14405 ^ w14762 ;
  assign w14764 = ~w14524 & w14763 ;
  assign w14765 = ( w14231 & w14522 ) | ( w14231 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14766 = ~w14523 & w14765 ;
  assign w14767 = w14764 | w14766 ;
  assign w14768 = ~\pi084 & w14767 ;
  assign w14769 = ~w14246 & w14401 ;
  assign w14770 = w14402 ^ w14769 ;
  assign w14771 = ~w14524 & w14770 ;
  assign w14772 = ( w14238 & w14522 ) | ( w14238 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14773 = ~w14523 & w14772 ;
  assign w14774 = w14771 | w14773 ;
  assign w14775 = ~\pi083 & w14774 ;
  assign w14776 = ~w14253 & w14398 ;
  assign w14777 = w14399 ^ w14776 ;
  assign w14778 = ~w14524 & w14777 ;
  assign w14779 = ( w14245 & w14522 ) | ( w14245 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14780 = ~w14523 & w14779 ;
  assign w14781 = w14778 | w14780 ;
  assign w14782 = ~\pi082 & w14781 ;
  assign w14783 = ~w14260 & w14395 ;
  assign w14784 = w14396 ^ w14783 ;
  assign w14785 = ~w14524 & w14784 ;
  assign w14786 = ( w14252 & w14522 ) | ( w14252 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14787 = ~w14523 & w14786 ;
  assign w14788 = w14785 | w14787 ;
  assign w14789 = ~\pi081 & w14788 ;
  assign w14790 = ~w14267 & w14392 ;
  assign w14791 = w14393 ^ w14790 ;
  assign w14792 = ~w14524 & w14791 ;
  assign w14793 = ( w14259 & w14522 ) | ( w14259 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14794 = ~w14523 & w14793 ;
  assign w14795 = w14792 | w14794 ;
  assign w14796 = ~\pi080 & w14795 ;
  assign w14797 = ~w14274 & w14389 ;
  assign w14798 = w14390 ^ w14797 ;
  assign w14799 = ~w14524 & w14798 ;
  assign w14800 = ( w14266 & w14522 ) | ( w14266 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14801 = ~w14523 & w14800 ;
  assign w14802 = w14799 | w14801 ;
  assign w14803 = ~\pi079 & w14802 ;
  assign w14804 = ~w14281 & w14386 ;
  assign w14805 = w14387 ^ w14804 ;
  assign w14806 = ~w14524 & w14805 ;
  assign w14807 = ( w14273 & w14522 ) | ( w14273 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14808 = ~w14523 & w14807 ;
  assign w14809 = w14806 | w14808 ;
  assign w14810 = ~\pi078 & w14809 ;
  assign w14811 = ~w14288 & w14383 ;
  assign w14812 = w14384 ^ w14811 ;
  assign w14813 = ~w14524 & w14812 ;
  assign w14814 = ( w14280 & w14522 ) | ( w14280 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14815 = ~w14523 & w14814 ;
  assign w14816 = w14813 | w14815 ;
  assign w14817 = ~\pi077 & w14816 ;
  assign w14818 = ~w14295 & w14380 ;
  assign w14819 = w14381 ^ w14818 ;
  assign w14820 = ~w14524 & w14819 ;
  assign w14821 = ( w14287 & w14522 ) | ( w14287 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14822 = ~w14523 & w14821 ;
  assign w14823 = w14820 | w14822 ;
  assign w14824 = ~\pi076 & w14823 ;
  assign w14825 = ~w14302 & w14377 ;
  assign w14826 = w14378 ^ w14825 ;
  assign w14827 = ~w14524 & w14826 ;
  assign w14828 = ( w14294 & w14522 ) | ( w14294 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14829 = ~w14523 & w14828 ;
  assign w14830 = w14827 | w14829 ;
  assign w14831 = ~\pi075 & w14830 ;
  assign w14832 = ~w14309 & w14374 ;
  assign w14833 = w14375 ^ w14832 ;
  assign w14834 = ~w14524 & w14833 ;
  assign w14835 = ( w14301 & w14522 ) | ( w14301 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14836 = ~w14523 & w14835 ;
  assign w14837 = w14834 | w14836 ;
  assign w14838 = ~\pi074 & w14837 ;
  assign w14839 = ~w14316 & w14371 ;
  assign w14840 = w14372 ^ w14839 ;
  assign w14841 = ~w14524 & w14840 ;
  assign w14842 = ( w14308 & w14522 ) | ( w14308 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14843 = ~w14523 & w14842 ;
  assign w14844 = w14841 | w14843 ;
  assign w14845 = ~\pi073 & w14844 ;
  assign w14846 = ~w14323 & w14368 ;
  assign w14847 = w14369 ^ w14846 ;
  assign w14848 = ~w14524 & w14847 ;
  assign w14849 = ( w14315 & w14522 ) | ( w14315 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14850 = ~w14523 & w14849 ;
  assign w14851 = w14848 | w14850 ;
  assign w14852 = ~\pi072 & w14851 ;
  assign w14853 = ~w14330 & w14365 ;
  assign w14854 = w14366 ^ w14853 ;
  assign w14855 = ~w14524 & w14854 ;
  assign w14856 = ( w14322 & w14522 ) | ( w14322 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14857 = ~w14523 & w14856 ;
  assign w14858 = w14855 | w14857 ;
  assign w14859 = ~\pi071 & w14858 ;
  assign w14860 = ~w14337 & w14362 ;
  assign w14861 = w14363 ^ w14860 ;
  assign w14862 = ~w14524 & w14861 ;
  assign w14863 = ( w14329 & w14522 ) | ( w14329 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14864 = ~w14523 & w14863 ;
  assign w14865 = w14862 | w14864 ;
  assign w14866 = ~\pi070 & w14865 ;
  assign w14867 = ~w14343 & w14359 ;
  assign w14868 = w14360 ^ w14867 ;
  assign w14869 = ~w14524 & w14868 ;
  assign w14870 = ( w14336 & w14522 ) | ( w14336 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14871 = ~w14523 & w14870 ;
  assign w14872 = w14869 | w14871 ;
  assign w14873 = ~\pi069 & w14872 ;
  assign w14874 = ~w14348 & w14356 ;
  assign w14875 = w14357 ^ w14874 ;
  assign w14876 = ~w14524 & w14875 ;
  assign w14877 = ( w14342 & w14522 ) | ( w14342 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14878 = ~w14523 & w14877 ;
  assign w14879 = w14876 | w14878 ;
  assign w14880 = ~\pi068 & w14879 ;
  assign w14881 = ~\pi010 & \pi064 ;
  assign w14882 = ( \pi065 & ~w14353 ) | ( \pi065 & w14881 ) | ( ~w14353 & w14881 ) ;
  assign w14883 = w14351 ^ w14882 ;
  assign w14884 = ~w14524 & w14883 ;
  assign w14885 = ( w14347 & w14522 ) | ( w14347 & w14523 ) | ( w14522 & w14523 ) ;
  assign w14886 = ~w14523 & w14885 ;
  assign w14887 = w14884 | w14886 ;
  assign w14888 = ~\pi067 & w14887 ;
  assign w14889 = \pi011 ^ \pi065 ;
  assign w14890 = \pi010 ^ w13994 ;
  assign w14891 = ( \pi064 & w14524 ) | ( \pi064 & w14890 ) | ( w14524 & w14890 ) ;
  assign w14892 = w14889 ^ w14891 ;
  assign w14893 = ~w14524 & w14892 ;
  assign w14894 = w14353 & w14524 ;
  assign w14895 = w14893 | w14894 ;
  assign w14896 = ~\pi066 & w14895 ;
  assign w14897 = \pi066 ^ w14895 ;
  assign w14898 = \pi064 & ~w14524 ;
  assign w14899 = \pi010 ^ w14898 ;
  assign w14900 = ( ~\pi009 & \pi064 ) | ( ~\pi009 & w14897 ) | ( \pi064 & w14897 ) ;
  assign w14901 = ( \pi065 & ~w14899 ) | ( \pi065 & w14900 ) | ( ~w14899 & w14900 ) ;
  assign w14902 = w14897 | w14901 ;
  assign w14903 = \pi067 ^ w14887 ;
  assign w14904 = ( ~w14896 & w14902 ) | ( ~w14896 & w14903 ) | ( w14902 & w14903 ) ;
  assign w14905 = w14903 | w14904 ;
  assign w14906 = \pi068 ^ w14879 ;
  assign w14907 = ( ~w14888 & w14905 ) | ( ~w14888 & w14906 ) | ( w14905 & w14906 ) ;
  assign w14908 = w14906 | w14907 ;
  assign w14909 = \pi069 ^ w14872 ;
  assign w14910 = ( ~w14880 & w14908 ) | ( ~w14880 & w14909 ) | ( w14908 & w14909 ) ;
  assign w14911 = w14909 | w14910 ;
  assign w14912 = \pi070 ^ w14865 ;
  assign w14913 = ( ~w14873 & w14911 ) | ( ~w14873 & w14912 ) | ( w14911 & w14912 ) ;
  assign w14914 = w14912 | w14913 ;
  assign w14915 = \pi071 ^ w14858 ;
  assign w14916 = ( ~w14866 & w14914 ) | ( ~w14866 & w14915 ) | ( w14914 & w14915 ) ;
  assign w14917 = w14915 | w14916 ;
  assign w14918 = \pi072 ^ w14851 ;
  assign w14919 = ( ~w14859 & w14917 ) | ( ~w14859 & w14918 ) | ( w14917 & w14918 ) ;
  assign w14920 = w14918 | w14919 ;
  assign w14921 = \pi073 ^ w14844 ;
  assign w14922 = ( ~w14852 & w14920 ) | ( ~w14852 & w14921 ) | ( w14920 & w14921 ) ;
  assign w14923 = w14921 | w14922 ;
  assign w14924 = \pi074 ^ w14837 ;
  assign w14925 = ( ~w14845 & w14923 ) | ( ~w14845 & w14924 ) | ( w14923 & w14924 ) ;
  assign w14926 = w14924 | w14925 ;
  assign w14927 = \pi075 ^ w14830 ;
  assign w14928 = ( ~w14838 & w14926 ) | ( ~w14838 & w14927 ) | ( w14926 & w14927 ) ;
  assign w14929 = w14927 | w14928 ;
  assign w14930 = \pi076 ^ w14823 ;
  assign w14931 = ( ~w14831 & w14929 ) | ( ~w14831 & w14930 ) | ( w14929 & w14930 ) ;
  assign w14932 = w14930 | w14931 ;
  assign w14933 = \pi077 ^ w14816 ;
  assign w14934 = ( ~w14824 & w14932 ) | ( ~w14824 & w14933 ) | ( w14932 & w14933 ) ;
  assign w14935 = w14933 | w14934 ;
  assign w14936 = \pi078 ^ w14809 ;
  assign w14937 = ( ~w14817 & w14935 ) | ( ~w14817 & w14936 ) | ( w14935 & w14936 ) ;
  assign w14938 = w14936 | w14937 ;
  assign w14939 = \pi079 ^ w14802 ;
  assign w14940 = ( ~w14810 & w14938 ) | ( ~w14810 & w14939 ) | ( w14938 & w14939 ) ;
  assign w14941 = w14939 | w14940 ;
  assign w14942 = \pi080 ^ w14795 ;
  assign w14943 = ( ~w14803 & w14941 ) | ( ~w14803 & w14942 ) | ( w14941 & w14942 ) ;
  assign w14944 = w14942 | w14943 ;
  assign w14945 = \pi081 ^ w14788 ;
  assign w14946 = ( ~w14796 & w14944 ) | ( ~w14796 & w14945 ) | ( w14944 & w14945 ) ;
  assign w14947 = w14945 | w14946 ;
  assign w14948 = \pi082 ^ w14781 ;
  assign w14949 = ( ~w14789 & w14947 ) | ( ~w14789 & w14948 ) | ( w14947 & w14948 ) ;
  assign w14950 = w14948 | w14949 ;
  assign w14951 = \pi083 ^ w14774 ;
  assign w14952 = ( ~w14782 & w14950 ) | ( ~w14782 & w14951 ) | ( w14950 & w14951 ) ;
  assign w14953 = w14951 | w14952 ;
  assign w14954 = \pi084 ^ w14767 ;
  assign w14955 = ( ~w14775 & w14953 ) | ( ~w14775 & w14954 ) | ( w14953 & w14954 ) ;
  assign w14956 = w14954 | w14955 ;
  assign w14957 = \pi085 ^ w14760 ;
  assign w14958 = ( ~w14768 & w14956 ) | ( ~w14768 & w14957 ) | ( w14956 & w14957 ) ;
  assign w14959 = w14957 | w14958 ;
  assign w14960 = \pi086 ^ w14753 ;
  assign w14961 = ( ~w14761 & w14959 ) | ( ~w14761 & w14960 ) | ( w14959 & w14960 ) ;
  assign w14962 = w14960 | w14961 ;
  assign w14963 = \pi087 ^ w14746 ;
  assign w14964 = ( ~w14754 & w14962 ) | ( ~w14754 & w14963 ) | ( w14962 & w14963 ) ;
  assign w14965 = w14963 | w14964 ;
  assign w14966 = \pi088 ^ w14739 ;
  assign w14967 = ( ~w14747 & w14965 ) | ( ~w14747 & w14966 ) | ( w14965 & w14966 ) ;
  assign w14968 = w14966 | w14967 ;
  assign w14969 = \pi089 ^ w14732 ;
  assign w14970 = ( ~w14740 & w14968 ) | ( ~w14740 & w14969 ) | ( w14968 & w14969 ) ;
  assign w14971 = w14969 | w14970 ;
  assign w14972 = \pi090 ^ w14725 ;
  assign w14973 = ( ~w14733 & w14971 ) | ( ~w14733 & w14972 ) | ( w14971 & w14972 ) ;
  assign w14974 = w14972 | w14973 ;
  assign w14975 = \pi091 ^ w14718 ;
  assign w14976 = ( ~w14726 & w14974 ) | ( ~w14726 & w14975 ) | ( w14974 & w14975 ) ;
  assign w14977 = w14975 | w14976 ;
  assign w14978 = \pi092 ^ w14711 ;
  assign w14979 = ( ~w14719 & w14977 ) | ( ~w14719 & w14978 ) | ( w14977 & w14978 ) ;
  assign w14980 = w14978 | w14979 ;
  assign w14981 = \pi093 ^ w14704 ;
  assign w14982 = ( ~w14712 & w14980 ) | ( ~w14712 & w14981 ) | ( w14980 & w14981 ) ;
  assign w14983 = w14981 | w14982 ;
  assign w14984 = \pi094 ^ w14697 ;
  assign w14985 = ( ~w14705 & w14983 ) | ( ~w14705 & w14984 ) | ( w14983 & w14984 ) ;
  assign w14986 = w14984 | w14985 ;
  assign w14987 = \pi095 ^ w14690 ;
  assign w14988 = ( ~w14698 & w14986 ) | ( ~w14698 & w14987 ) | ( w14986 & w14987 ) ;
  assign w14989 = w14987 | w14988 ;
  assign w14990 = \pi096 ^ w14683 ;
  assign w14991 = ( ~w14691 & w14989 ) | ( ~w14691 & w14990 ) | ( w14989 & w14990 ) ;
  assign w14992 = w14990 | w14991 ;
  assign w14993 = \pi097 ^ w14676 ;
  assign w14994 = ( ~w14684 & w14992 ) | ( ~w14684 & w14993 ) | ( w14992 & w14993 ) ;
  assign w14995 = w14993 | w14994 ;
  assign w14996 = \pi098 ^ w14669 ;
  assign w14997 = ( ~w14677 & w14995 ) | ( ~w14677 & w14996 ) | ( w14995 & w14996 ) ;
  assign w14998 = w14996 | w14997 ;
  assign w14999 = \pi099 ^ w14662 ;
  assign w15000 = ( ~w14670 & w14998 ) | ( ~w14670 & w14999 ) | ( w14998 & w14999 ) ;
  assign w15001 = w14999 | w15000 ;
  assign w15002 = \pi100 ^ w14655 ;
  assign w15003 = ( ~w14663 & w15001 ) | ( ~w14663 & w15002 ) | ( w15001 & w15002 ) ;
  assign w15004 = w15002 | w15003 ;
  assign w15005 = \pi101 ^ w14648 ;
  assign w15006 = ( ~w14656 & w15004 ) | ( ~w14656 & w15005 ) | ( w15004 & w15005 ) ;
  assign w15007 = w15005 | w15006 ;
  assign w15008 = \pi102 ^ w14641 ;
  assign w15009 = ( ~w14649 & w15007 ) | ( ~w14649 & w15008 ) | ( w15007 & w15008 ) ;
  assign w15010 = w15008 | w15009 ;
  assign w15011 = \pi103 ^ w14634 ;
  assign w15012 = ( ~w14642 & w15010 ) | ( ~w14642 & w15011 ) | ( w15010 & w15011 ) ;
  assign w15013 = w15011 | w15012 ;
  assign w15014 = \pi104 ^ w14627 ;
  assign w15015 = ( ~w14635 & w15013 ) | ( ~w14635 & w15014 ) | ( w15013 & w15014 ) ;
  assign w15016 = w15014 | w15015 ;
  assign w15017 = \pi105 ^ w14620 ;
  assign w15018 = ( ~w14628 & w15016 ) | ( ~w14628 & w15017 ) | ( w15016 & w15017 ) ;
  assign w15019 = w15017 | w15018 ;
  assign w15020 = \pi106 ^ w14613 ;
  assign w15021 = ( ~w14621 & w15019 ) | ( ~w14621 & w15020 ) | ( w15019 & w15020 ) ;
  assign w15022 = w15020 | w15021 ;
  assign w15023 = \pi107 ^ w14606 ;
  assign w15024 = ( ~w14614 & w15022 ) | ( ~w14614 & w15023 ) | ( w15022 & w15023 ) ;
  assign w15025 = w15023 | w15024 ;
  assign w15026 = \pi108 ^ w14599 ;
  assign w15027 = ( ~w14607 & w15025 ) | ( ~w14607 & w15026 ) | ( w15025 & w15026 ) ;
  assign w15028 = w15026 | w15027 ;
  assign w15029 = \pi109 ^ w14592 ;
  assign w15030 = ( ~w14600 & w15028 ) | ( ~w14600 & w15029 ) | ( w15028 & w15029 ) ;
  assign w15031 = w15029 | w15030 ;
  assign w15032 = \pi110 ^ w14585 ;
  assign w15033 = ( ~w14593 & w15031 ) | ( ~w14593 & w15032 ) | ( w15031 & w15032 ) ;
  assign w15034 = w15032 | w15033 ;
  assign w15035 = \pi111 ^ w14578 ;
  assign w15036 = ( ~w14586 & w15034 ) | ( ~w14586 & w15035 ) | ( w15034 & w15035 ) ;
  assign w15037 = w15035 | w15036 ;
  assign w15038 = \pi112 ^ w14571 ;
  assign w15039 = ( ~w14579 & w15037 ) | ( ~w14579 & w15038 ) | ( w15037 & w15038 ) ;
  assign w15040 = w15038 | w15039 ;
  assign w15041 = \pi113 ^ w14564 ;
  assign w15042 = ( ~w14572 & w15040 ) | ( ~w14572 & w15041 ) | ( w15040 & w15041 ) ;
  assign w15043 = w15041 | w15042 ;
  assign w15044 = \pi114 ^ w14557 ;
  assign w15045 = ( ~w14565 & w15043 ) | ( ~w14565 & w15044 ) | ( w15043 & w15044 ) ;
  assign w15046 = w15044 | w15045 ;
  assign w15047 = \pi115 ^ w14550 ;
  assign w15048 = ( ~w14558 & w15046 ) | ( ~w14558 & w15047 ) | ( w15046 & w15047 ) ;
  assign w15049 = w15047 | w15048 ;
  assign w15050 = \pi116 ^ w14543 ;
  assign w15051 = ( ~w14551 & w15049 ) | ( ~w14551 & w15050 ) | ( w15049 & w15050 ) ;
  assign w15052 = w15050 | w15051 ;
  assign w15053 = \pi117 ^ w14530 ;
  assign w15054 = ( ~w14544 & w15052 ) | ( ~w14544 & w15053 ) | ( w15052 & w15053 ) ;
  assign w15055 = w15053 | w15054 ;
  assign w15056 = \pi118 ^ w14536 ;
  assign w15057 = w14537 & ~w15056 ;
  assign w15058 = ( w15055 & w15056 ) | ( w15055 & ~w15057 ) | ( w15056 & ~w15057 ) ;
  assign w15059 = ~\pi118 & w14536 ;
  assign w15060 = w15058 & ~w15059 ;
  assign w15061 = \pi120 | w269 ;
  assign w15062 = ( \pi119 & ~w269 ) | ( \pi119 & w272 ) | ( ~w269 & w272 ) ;
  assign w15063 = w15061 | w15062 ;
  assign w15064 = w15060 | w15063 ;
  assign w15065 = w14530 & w15064 ;
  assign w15066 = ~w14544 & w15052 ;
  assign w15067 = w15053 ^ w15066 ;
  assign w15068 = ~w15064 & w15067 ;
  assign w15069 = w15065 | w15068 ;
  assign w15070 = ~\pi118 & w15069 ;
  assign w15071 = w14543 & w15064 ;
  assign w15072 = ~w14551 & w15049 ;
  assign w15073 = w15050 ^ w15072 ;
  assign w15074 = ~w15064 & w15073 ;
  assign w15075 = w15071 | w15074 ;
  assign w15076 = ~\pi117 & w15075 ;
  assign w15077 = w14550 & w15064 ;
  assign w15078 = ~w14558 & w15046 ;
  assign w15079 = w15047 ^ w15078 ;
  assign w15080 = ~w15064 & w15079 ;
  assign w15081 = w15077 | w15080 ;
  assign w15082 = ~\pi116 & w15081 ;
  assign w15083 = w14557 & w15064 ;
  assign w15084 = ~w14565 & w15043 ;
  assign w15085 = w15044 ^ w15084 ;
  assign w15086 = ~w15064 & w15085 ;
  assign w15087 = w15083 | w15086 ;
  assign w15088 = ~\pi115 & w15087 ;
  assign w15089 = w14564 & w15064 ;
  assign w15090 = ~w14572 & w15040 ;
  assign w15091 = w15041 ^ w15090 ;
  assign w15092 = ~w15064 & w15091 ;
  assign w15093 = w15089 | w15092 ;
  assign w15094 = ~\pi114 & w15093 ;
  assign w15095 = w14571 & w15064 ;
  assign w15096 = ~w14579 & w15037 ;
  assign w15097 = w15038 ^ w15096 ;
  assign w15098 = ~w15064 & w15097 ;
  assign w15099 = w15095 | w15098 ;
  assign w15100 = ~\pi113 & w15099 ;
  assign w15101 = w14578 & w15064 ;
  assign w15102 = ~w14586 & w15034 ;
  assign w15103 = w15035 ^ w15102 ;
  assign w15104 = ~w15064 & w15103 ;
  assign w15105 = w15101 | w15104 ;
  assign w15106 = ~\pi112 & w15105 ;
  assign w15107 = w14585 & w15064 ;
  assign w15108 = ~w14593 & w15031 ;
  assign w15109 = w15032 ^ w15108 ;
  assign w15110 = ~w15064 & w15109 ;
  assign w15111 = w15107 | w15110 ;
  assign w15112 = ~\pi111 & w15111 ;
  assign w15113 = w14592 & w15064 ;
  assign w15114 = ~w14600 & w15028 ;
  assign w15115 = w15029 ^ w15114 ;
  assign w15116 = ~w15064 & w15115 ;
  assign w15117 = w15113 | w15116 ;
  assign w15118 = ~\pi110 & w15117 ;
  assign w15119 = w14599 & w15064 ;
  assign w15120 = ~w14607 & w15025 ;
  assign w15121 = w15026 ^ w15120 ;
  assign w15122 = ~w15064 & w15121 ;
  assign w15123 = w15119 | w15122 ;
  assign w15124 = ~\pi109 & w15123 ;
  assign w15125 = w14606 & w15064 ;
  assign w15126 = ~w14614 & w15022 ;
  assign w15127 = w15023 ^ w15126 ;
  assign w15128 = ~w15064 & w15127 ;
  assign w15129 = w15125 | w15128 ;
  assign w15130 = ~\pi108 & w15129 ;
  assign w15131 = w14613 & w15064 ;
  assign w15132 = ~w14621 & w15019 ;
  assign w15133 = w15020 ^ w15132 ;
  assign w15134 = ~w15064 & w15133 ;
  assign w15135 = w15131 | w15134 ;
  assign w15136 = ~\pi107 & w15135 ;
  assign w15137 = w14620 & w15064 ;
  assign w15138 = ~w14628 & w15016 ;
  assign w15139 = w15017 ^ w15138 ;
  assign w15140 = ~w15064 & w15139 ;
  assign w15141 = w15137 | w15140 ;
  assign w15142 = ~\pi106 & w15141 ;
  assign w15143 = w14627 & w15064 ;
  assign w15144 = ~w14635 & w15013 ;
  assign w15145 = w15014 ^ w15144 ;
  assign w15146 = ~w15064 & w15145 ;
  assign w15147 = w15143 | w15146 ;
  assign w15148 = ~\pi105 & w15147 ;
  assign w15149 = w14634 & w15064 ;
  assign w15150 = ~w14642 & w15010 ;
  assign w15151 = w15011 ^ w15150 ;
  assign w15152 = ~w15064 & w15151 ;
  assign w15153 = w15149 | w15152 ;
  assign w15154 = ~\pi104 & w15153 ;
  assign w15155 = w14641 & w15064 ;
  assign w15156 = ~w14649 & w15007 ;
  assign w15157 = w15008 ^ w15156 ;
  assign w15158 = ~w15064 & w15157 ;
  assign w15159 = w15155 | w15158 ;
  assign w15160 = ~\pi103 & w15159 ;
  assign w15161 = w14648 & w15064 ;
  assign w15162 = ~w14656 & w15004 ;
  assign w15163 = w15005 ^ w15162 ;
  assign w15164 = ~w15064 & w15163 ;
  assign w15165 = w15161 | w15164 ;
  assign w15166 = ~\pi102 & w15165 ;
  assign w15167 = w14655 & w15064 ;
  assign w15168 = ~w14663 & w15001 ;
  assign w15169 = w15002 ^ w15168 ;
  assign w15170 = ~w15064 & w15169 ;
  assign w15171 = w15167 | w15170 ;
  assign w15172 = ~\pi101 & w15171 ;
  assign w15173 = w14662 & w15064 ;
  assign w15174 = ~w14670 & w14998 ;
  assign w15175 = w14999 ^ w15174 ;
  assign w15176 = ~w15064 & w15175 ;
  assign w15177 = w15173 | w15176 ;
  assign w15178 = ~\pi100 & w15177 ;
  assign w15179 = w14669 & w15064 ;
  assign w15180 = ~w14677 & w14995 ;
  assign w15181 = w14996 ^ w15180 ;
  assign w15182 = ~w15064 & w15181 ;
  assign w15183 = w15179 | w15182 ;
  assign w15184 = ~\pi099 & w15183 ;
  assign w15185 = w14676 & w15064 ;
  assign w15186 = ~w14684 & w14992 ;
  assign w15187 = w14993 ^ w15186 ;
  assign w15188 = ~w15064 & w15187 ;
  assign w15189 = w15185 | w15188 ;
  assign w15190 = ~\pi098 & w15189 ;
  assign w15191 = w14683 & w15064 ;
  assign w15192 = ~w14691 & w14989 ;
  assign w15193 = w14990 ^ w15192 ;
  assign w15194 = ~w15064 & w15193 ;
  assign w15195 = w15191 | w15194 ;
  assign w15196 = ~\pi097 & w15195 ;
  assign w15197 = w14690 & w15064 ;
  assign w15198 = ~w14698 & w14986 ;
  assign w15199 = w14987 ^ w15198 ;
  assign w15200 = ~w15064 & w15199 ;
  assign w15201 = w15197 | w15200 ;
  assign w15202 = ~\pi096 & w15201 ;
  assign w15203 = w14697 & w15064 ;
  assign w15204 = ~w14705 & w14983 ;
  assign w15205 = w14984 ^ w15204 ;
  assign w15206 = ~w15064 & w15205 ;
  assign w15207 = w15203 | w15206 ;
  assign w15208 = ~\pi095 & w15207 ;
  assign w15209 = w14704 & w15064 ;
  assign w15210 = ~w14712 & w14980 ;
  assign w15211 = w14981 ^ w15210 ;
  assign w15212 = ~w15064 & w15211 ;
  assign w15213 = w15209 | w15212 ;
  assign w15214 = ~\pi094 & w15213 ;
  assign w15215 = w14711 & w15064 ;
  assign w15216 = ~w14719 & w14977 ;
  assign w15217 = w14978 ^ w15216 ;
  assign w15218 = ~w15064 & w15217 ;
  assign w15219 = w15215 | w15218 ;
  assign w15220 = ~\pi093 & w15219 ;
  assign w15221 = w14718 & w15064 ;
  assign w15222 = ~w14726 & w14974 ;
  assign w15223 = w14975 ^ w15222 ;
  assign w15224 = ~w15064 & w15223 ;
  assign w15225 = w15221 | w15224 ;
  assign w15226 = ~\pi092 & w15225 ;
  assign w15227 = w14725 & w15064 ;
  assign w15228 = ~w14733 & w14971 ;
  assign w15229 = w14972 ^ w15228 ;
  assign w15230 = ~w15064 & w15229 ;
  assign w15231 = w15227 | w15230 ;
  assign w15232 = ~\pi091 & w15231 ;
  assign w15233 = w14732 & w15064 ;
  assign w15234 = ~w14740 & w14968 ;
  assign w15235 = w14969 ^ w15234 ;
  assign w15236 = ~w15064 & w15235 ;
  assign w15237 = w15233 | w15236 ;
  assign w15238 = ~\pi090 & w15237 ;
  assign w15239 = w14739 & w15064 ;
  assign w15240 = ~w14747 & w14965 ;
  assign w15241 = w14966 ^ w15240 ;
  assign w15242 = ~w15064 & w15241 ;
  assign w15243 = w15239 | w15242 ;
  assign w15244 = ~\pi089 & w15243 ;
  assign w15245 = w14746 & w15064 ;
  assign w15246 = ~w14754 & w14962 ;
  assign w15247 = w14963 ^ w15246 ;
  assign w15248 = ~w15064 & w15247 ;
  assign w15249 = w15245 | w15248 ;
  assign w15250 = ~\pi088 & w15249 ;
  assign w15251 = w14753 & w15064 ;
  assign w15252 = ~w14761 & w14959 ;
  assign w15253 = w14960 ^ w15252 ;
  assign w15254 = ~w15064 & w15253 ;
  assign w15255 = w15251 | w15254 ;
  assign w15256 = ~\pi087 & w15255 ;
  assign w15257 = w14760 & w15064 ;
  assign w15258 = ~w14768 & w14956 ;
  assign w15259 = w14957 ^ w15258 ;
  assign w15260 = ~w15064 & w15259 ;
  assign w15261 = w15257 | w15260 ;
  assign w15262 = ~\pi086 & w15261 ;
  assign w15263 = w14767 & w15064 ;
  assign w15264 = ~w14775 & w14953 ;
  assign w15265 = w14954 ^ w15264 ;
  assign w15266 = ~w15064 & w15265 ;
  assign w15267 = w15263 | w15266 ;
  assign w15268 = ~\pi085 & w15267 ;
  assign w15269 = w14774 & w15064 ;
  assign w15270 = ~w14782 & w14950 ;
  assign w15271 = w14951 ^ w15270 ;
  assign w15272 = ~w15064 & w15271 ;
  assign w15273 = w15269 | w15272 ;
  assign w15274 = ~\pi084 & w15273 ;
  assign w15275 = w14781 & w15064 ;
  assign w15276 = ~w14789 & w14947 ;
  assign w15277 = w14948 ^ w15276 ;
  assign w15278 = ~w15064 & w15277 ;
  assign w15279 = w15275 | w15278 ;
  assign w15280 = ~\pi083 & w15279 ;
  assign w15281 = w14788 & w15064 ;
  assign w15282 = ~w14796 & w14944 ;
  assign w15283 = w14945 ^ w15282 ;
  assign w15284 = ~w15064 & w15283 ;
  assign w15285 = w15281 | w15284 ;
  assign w15286 = ~\pi082 & w15285 ;
  assign w15287 = w14795 & w15064 ;
  assign w15288 = ~w14803 & w14941 ;
  assign w15289 = w14942 ^ w15288 ;
  assign w15290 = ~w15064 & w15289 ;
  assign w15291 = w15287 | w15290 ;
  assign w15292 = ~\pi081 & w15291 ;
  assign w15293 = w14802 & w15064 ;
  assign w15294 = ~w14810 & w14938 ;
  assign w15295 = w14939 ^ w15294 ;
  assign w15296 = ~w15064 & w15295 ;
  assign w15297 = w15293 | w15296 ;
  assign w15298 = ~\pi080 & w15297 ;
  assign w15299 = w14809 & w15064 ;
  assign w15300 = ~w14817 & w14935 ;
  assign w15301 = w14936 ^ w15300 ;
  assign w15302 = ~w15064 & w15301 ;
  assign w15303 = w15299 | w15302 ;
  assign w15304 = ~\pi079 & w15303 ;
  assign w15305 = w14816 & w15064 ;
  assign w15306 = ~w14824 & w14932 ;
  assign w15307 = w14933 ^ w15306 ;
  assign w15308 = ~w15064 & w15307 ;
  assign w15309 = w15305 | w15308 ;
  assign w15310 = ~\pi078 & w15309 ;
  assign w15311 = w14823 & w15064 ;
  assign w15312 = ~w14831 & w14929 ;
  assign w15313 = w14930 ^ w15312 ;
  assign w15314 = ~w15064 & w15313 ;
  assign w15315 = w15311 | w15314 ;
  assign w15316 = ~\pi077 & w15315 ;
  assign w15317 = w14830 & w15064 ;
  assign w15318 = ~w14838 & w14926 ;
  assign w15319 = w14927 ^ w15318 ;
  assign w15320 = ~w15064 & w15319 ;
  assign w15321 = w15317 | w15320 ;
  assign w15322 = ~\pi076 & w15321 ;
  assign w15323 = w14837 & w15064 ;
  assign w15324 = ~w14845 & w14923 ;
  assign w15325 = w14924 ^ w15324 ;
  assign w15326 = ~w15064 & w15325 ;
  assign w15327 = w15323 | w15326 ;
  assign w15328 = ~\pi075 & w15327 ;
  assign w15329 = w14844 & w15064 ;
  assign w15330 = ~w14852 & w14920 ;
  assign w15331 = w14921 ^ w15330 ;
  assign w15332 = ~w15064 & w15331 ;
  assign w15333 = w15329 | w15332 ;
  assign w15334 = ~\pi074 & w15333 ;
  assign w15335 = w14851 & w15064 ;
  assign w15336 = ~w14859 & w14917 ;
  assign w15337 = w14918 ^ w15336 ;
  assign w15338 = ~w15064 & w15337 ;
  assign w15339 = w15335 | w15338 ;
  assign w15340 = ~\pi073 & w15339 ;
  assign w15341 = w14858 & w15064 ;
  assign w15342 = ~w14866 & w14914 ;
  assign w15343 = w14915 ^ w15342 ;
  assign w15344 = ~w15064 & w15343 ;
  assign w15345 = w15341 | w15344 ;
  assign w15346 = ~\pi072 & w15345 ;
  assign w15347 = w14865 & w15064 ;
  assign w15348 = ~w14873 & w14911 ;
  assign w15349 = w14912 ^ w15348 ;
  assign w15350 = ~w15064 & w15349 ;
  assign w15351 = w15347 | w15350 ;
  assign w15352 = ~\pi071 & w15351 ;
  assign w15353 = w14872 & w15064 ;
  assign w15354 = ~w14880 & w14908 ;
  assign w15355 = w14909 ^ w15354 ;
  assign w15356 = ~w15064 & w15355 ;
  assign w15357 = w15353 | w15356 ;
  assign w15358 = ~\pi070 & w15357 ;
  assign w15359 = w14879 & w15064 ;
  assign w15360 = ~w14888 & w14905 ;
  assign w15361 = w14906 ^ w15360 ;
  assign w15362 = ~w15064 & w15361 ;
  assign w15363 = w15359 | w15362 ;
  assign w15364 = ~\pi069 & w15363 ;
  assign w15365 = w14887 & w15064 ;
  assign w15366 = ~w14896 & w14902 ;
  assign w15367 = w14903 ^ w15366 ;
  assign w15368 = ~w15064 & w15367 ;
  assign w15369 = w15365 | w15368 ;
  assign w15370 = ~\pi068 & w15369 ;
  assign w15371 = ~\pi009 & \pi064 ;
  assign w15372 = ( \pi065 & ~w14899 ) | ( \pi065 & w15371 ) | ( ~w14899 & w15371 ) ;
  assign w15373 = w14897 ^ w15372 ;
  assign w15374 = ( w15060 & w15063 ) | ( w15060 & w15373 ) | ( w15063 & w15373 ) ;
  assign w15375 = w15373 & ~w15374 ;
  assign w15376 = ( w14895 & w15064 ) | ( w14895 & w15375 ) | ( w15064 & w15375 ) ;
  assign w15377 = w15375 | w15376 ;
  assign w15378 = ~\pi067 & w15377 ;
  assign w15379 = \pi010 ^ \pi065 ;
  assign w15380 = \pi009 ^ w14524 ;
  assign w15381 = ( \pi064 & w15063 ) | ( \pi064 & w15380 ) | ( w15063 & w15380 ) ;
  assign w15382 = w15379 ^ w15381 ;
  assign w15383 = ~w15063 & w15382 ;
  assign w15384 = ~w15060 & w15383 ;
  assign w15385 = ( ~\pi064 & w14524 ) | ( ~\pi064 & w15064 ) | ( w14524 & w15064 ) ;
  assign w15386 = \pi010 ^ w15385 ;
  assign w15387 = w15064 & ~w15386 ;
  assign w15388 = w15384 | w15387 ;
  assign w15389 = ~\pi066 & w15388 ;
  assign w15390 = ( \pi064 & w147 ) | ( \pi064 & w150 ) | ( w147 & w150 ) ;
  assign w15391 = \pi009 & \pi119 ;
  assign w15392 = ( \pi009 & w15390 ) | ( \pi009 & w15391 ) | ( w15390 & w15391 ) ;
  assign w15393 = ( \pi064 & w15060 ) | ( \pi064 & w15392 ) | ( w15060 & w15392 ) ;
  assign w15394 = ( \pi009 & ~\pi064 ) | ( \pi009 & w15393 ) | ( ~\pi064 & w15393 ) ;
  assign w15395 = ( ~\pi009 & \pi064 ) | ( ~\pi009 & \pi119 ) | ( \pi064 & \pi119 ) ;
  assign w15396 = ( \pi119 & \pi120 ) | ( \pi119 & ~w269 ) | ( \pi120 & ~w269 ) ;
  assign w15397 = w273 | w15396 ;
  assign w15398 = w15395 & ~w15397 ;
  assign w15399 = ~w15060 & w15398 ;
  assign w15400 = ~\pi008 & \pi064 ;
  assign w15401 = w15064 | w15384 ;
  assign w15402 = ( w14899 & w15384 ) | ( w14899 & w15401 ) | ( w15384 & w15401 ) ;
  assign w15403 = \pi066 ^ w15402 ;
  assign w15404 = w15394 | w15399 ;
  assign w15405 = ( \pi065 & w15400 ) | ( \pi065 & ~w15404 ) | ( w15400 & ~w15404 ) ;
  assign w15406 = w15403 | w15405 ;
  assign w15407 = ~w14895 & w15064 ;
  assign w15408 = ( w15064 & w15375 ) | ( w15064 & ~w15407 ) | ( w15375 & ~w15407 ) ;
  assign w15409 = \pi067 ^ w15408 ;
  assign w15410 = ( ~w15389 & w15406 ) | ( ~w15389 & w15409 ) | ( w15406 & w15409 ) ;
  assign w15411 = w15409 | w15410 ;
  assign w15412 = \pi068 ^ w15369 ;
  assign w15413 = ( ~w15378 & w15411 ) | ( ~w15378 & w15412 ) | ( w15411 & w15412 ) ;
  assign w15414 = w15412 | w15413 ;
  assign w15415 = \pi069 ^ w15363 ;
  assign w15416 = ( ~w15370 & w15414 ) | ( ~w15370 & w15415 ) | ( w15414 & w15415 ) ;
  assign w15417 = w15415 | w15416 ;
  assign w15418 = \pi070 ^ w15357 ;
  assign w15419 = ( ~w15364 & w15417 ) | ( ~w15364 & w15418 ) | ( w15417 & w15418 ) ;
  assign w15420 = w15418 | w15419 ;
  assign w15421 = \pi071 ^ w15351 ;
  assign w15422 = ( ~w15358 & w15420 ) | ( ~w15358 & w15421 ) | ( w15420 & w15421 ) ;
  assign w15423 = w15421 | w15422 ;
  assign w15424 = \pi072 ^ w15345 ;
  assign w15425 = ( ~w15352 & w15423 ) | ( ~w15352 & w15424 ) | ( w15423 & w15424 ) ;
  assign w15426 = w15424 | w15425 ;
  assign w15427 = \pi073 ^ w15339 ;
  assign w15428 = ( ~w15346 & w15426 ) | ( ~w15346 & w15427 ) | ( w15426 & w15427 ) ;
  assign w15429 = w15427 | w15428 ;
  assign w15430 = \pi074 ^ w15333 ;
  assign w15431 = ( ~w15340 & w15429 ) | ( ~w15340 & w15430 ) | ( w15429 & w15430 ) ;
  assign w15432 = w15430 | w15431 ;
  assign w15433 = \pi075 ^ w15327 ;
  assign w15434 = ( ~w15334 & w15432 ) | ( ~w15334 & w15433 ) | ( w15432 & w15433 ) ;
  assign w15435 = w15433 | w15434 ;
  assign w15436 = \pi076 ^ w15321 ;
  assign w15437 = ( ~w15328 & w15435 ) | ( ~w15328 & w15436 ) | ( w15435 & w15436 ) ;
  assign w15438 = w15436 | w15437 ;
  assign w15439 = \pi077 ^ w15315 ;
  assign w15440 = ( ~w15322 & w15438 ) | ( ~w15322 & w15439 ) | ( w15438 & w15439 ) ;
  assign w15441 = w15439 | w15440 ;
  assign w15442 = \pi078 ^ w15309 ;
  assign w15443 = ( ~w15316 & w15441 ) | ( ~w15316 & w15442 ) | ( w15441 & w15442 ) ;
  assign w15444 = w15442 | w15443 ;
  assign w15445 = \pi079 ^ w15303 ;
  assign w15446 = ( ~w15310 & w15444 ) | ( ~w15310 & w15445 ) | ( w15444 & w15445 ) ;
  assign w15447 = w15445 | w15446 ;
  assign w15448 = \pi080 ^ w15297 ;
  assign w15449 = ( ~w15304 & w15447 ) | ( ~w15304 & w15448 ) | ( w15447 & w15448 ) ;
  assign w15450 = w15448 | w15449 ;
  assign w15451 = \pi081 ^ w15291 ;
  assign w15452 = ( ~w15298 & w15450 ) | ( ~w15298 & w15451 ) | ( w15450 & w15451 ) ;
  assign w15453 = w15451 | w15452 ;
  assign w15454 = \pi082 ^ w15285 ;
  assign w15455 = ( ~w15292 & w15453 ) | ( ~w15292 & w15454 ) | ( w15453 & w15454 ) ;
  assign w15456 = w15454 | w15455 ;
  assign w15457 = \pi083 ^ w15279 ;
  assign w15458 = ( ~w15286 & w15456 ) | ( ~w15286 & w15457 ) | ( w15456 & w15457 ) ;
  assign w15459 = w15457 | w15458 ;
  assign w15460 = \pi084 ^ w15273 ;
  assign w15461 = ( ~w15280 & w15459 ) | ( ~w15280 & w15460 ) | ( w15459 & w15460 ) ;
  assign w15462 = w15460 | w15461 ;
  assign w15463 = \pi085 ^ w15267 ;
  assign w15464 = ( ~w15274 & w15462 ) | ( ~w15274 & w15463 ) | ( w15462 & w15463 ) ;
  assign w15465 = w15463 | w15464 ;
  assign w15466 = \pi086 ^ w15261 ;
  assign w15467 = ( ~w15268 & w15465 ) | ( ~w15268 & w15466 ) | ( w15465 & w15466 ) ;
  assign w15468 = w15466 | w15467 ;
  assign w15469 = \pi087 ^ w15255 ;
  assign w15470 = ( ~w15262 & w15468 ) | ( ~w15262 & w15469 ) | ( w15468 & w15469 ) ;
  assign w15471 = w15469 | w15470 ;
  assign w15472 = \pi088 ^ w15249 ;
  assign w15473 = ( ~w15256 & w15471 ) | ( ~w15256 & w15472 ) | ( w15471 & w15472 ) ;
  assign w15474 = w15472 | w15473 ;
  assign w15475 = \pi089 ^ w15243 ;
  assign w15476 = ( ~w15250 & w15474 ) | ( ~w15250 & w15475 ) | ( w15474 & w15475 ) ;
  assign w15477 = w15475 | w15476 ;
  assign w15478 = \pi090 ^ w15237 ;
  assign w15479 = ( ~w15244 & w15477 ) | ( ~w15244 & w15478 ) | ( w15477 & w15478 ) ;
  assign w15480 = w15478 | w15479 ;
  assign w15481 = \pi091 ^ w15231 ;
  assign w15482 = ( ~w15238 & w15480 ) | ( ~w15238 & w15481 ) | ( w15480 & w15481 ) ;
  assign w15483 = w15481 | w15482 ;
  assign w15484 = \pi092 ^ w15225 ;
  assign w15485 = ( ~w15232 & w15483 ) | ( ~w15232 & w15484 ) | ( w15483 & w15484 ) ;
  assign w15486 = w15484 | w15485 ;
  assign w15487 = \pi093 ^ w15219 ;
  assign w15488 = ( ~w15226 & w15486 ) | ( ~w15226 & w15487 ) | ( w15486 & w15487 ) ;
  assign w15489 = w15487 | w15488 ;
  assign w15490 = \pi094 ^ w15213 ;
  assign w15491 = ( ~w15220 & w15489 ) | ( ~w15220 & w15490 ) | ( w15489 & w15490 ) ;
  assign w15492 = w15490 | w15491 ;
  assign w15493 = \pi095 ^ w15207 ;
  assign w15494 = ( ~w15214 & w15492 ) | ( ~w15214 & w15493 ) | ( w15492 & w15493 ) ;
  assign w15495 = w15493 | w15494 ;
  assign w15496 = \pi096 ^ w15201 ;
  assign w15497 = ( ~w15208 & w15495 ) | ( ~w15208 & w15496 ) | ( w15495 & w15496 ) ;
  assign w15498 = w15496 | w15497 ;
  assign w15499 = \pi097 ^ w15195 ;
  assign w15500 = ( ~w15202 & w15498 ) | ( ~w15202 & w15499 ) | ( w15498 & w15499 ) ;
  assign w15501 = w15499 | w15500 ;
  assign w15502 = \pi098 ^ w15189 ;
  assign w15503 = ( ~w15196 & w15501 ) | ( ~w15196 & w15502 ) | ( w15501 & w15502 ) ;
  assign w15504 = w15502 | w15503 ;
  assign w15505 = \pi099 ^ w15183 ;
  assign w15506 = ( ~w15190 & w15504 ) | ( ~w15190 & w15505 ) | ( w15504 & w15505 ) ;
  assign w15507 = w15505 | w15506 ;
  assign w15508 = \pi100 ^ w15177 ;
  assign w15509 = ( ~w15184 & w15507 ) | ( ~w15184 & w15508 ) | ( w15507 & w15508 ) ;
  assign w15510 = w15508 | w15509 ;
  assign w15511 = \pi101 ^ w15171 ;
  assign w15512 = ( ~w15178 & w15510 ) | ( ~w15178 & w15511 ) | ( w15510 & w15511 ) ;
  assign w15513 = w15511 | w15512 ;
  assign w15514 = \pi102 ^ w15165 ;
  assign w15515 = ( ~w15172 & w15513 ) | ( ~w15172 & w15514 ) | ( w15513 & w15514 ) ;
  assign w15516 = w15514 | w15515 ;
  assign w15517 = \pi103 ^ w15159 ;
  assign w15518 = ( ~w15166 & w15516 ) | ( ~w15166 & w15517 ) | ( w15516 & w15517 ) ;
  assign w15519 = w15517 | w15518 ;
  assign w15520 = \pi104 ^ w15153 ;
  assign w15521 = ( ~w15160 & w15519 ) | ( ~w15160 & w15520 ) | ( w15519 & w15520 ) ;
  assign w15522 = w15520 | w15521 ;
  assign w15523 = \pi105 ^ w15147 ;
  assign w15524 = ( ~w15154 & w15522 ) | ( ~w15154 & w15523 ) | ( w15522 & w15523 ) ;
  assign w15525 = w15523 | w15524 ;
  assign w15526 = \pi106 ^ w15141 ;
  assign w15527 = ( ~w15148 & w15525 ) | ( ~w15148 & w15526 ) | ( w15525 & w15526 ) ;
  assign w15528 = w15526 | w15527 ;
  assign w15529 = \pi107 ^ w15135 ;
  assign w15530 = ( ~w15142 & w15528 ) | ( ~w15142 & w15529 ) | ( w15528 & w15529 ) ;
  assign w15531 = w15529 | w15530 ;
  assign w15532 = \pi108 ^ w15129 ;
  assign w15533 = ( ~w15136 & w15531 ) | ( ~w15136 & w15532 ) | ( w15531 & w15532 ) ;
  assign w15534 = w15532 | w15533 ;
  assign w15535 = \pi109 ^ w15123 ;
  assign w15536 = ( ~w15130 & w15534 ) | ( ~w15130 & w15535 ) | ( w15534 & w15535 ) ;
  assign w15537 = w15535 | w15536 ;
  assign w15538 = \pi110 ^ w15117 ;
  assign w15539 = ( ~w15124 & w15537 ) | ( ~w15124 & w15538 ) | ( w15537 & w15538 ) ;
  assign w15540 = w15538 | w15539 ;
  assign w15541 = \pi111 ^ w15111 ;
  assign w15542 = ( ~w15118 & w15540 ) | ( ~w15118 & w15541 ) | ( w15540 & w15541 ) ;
  assign w15543 = w15541 | w15542 ;
  assign w15544 = \pi112 ^ w15105 ;
  assign w15545 = ( ~w15112 & w15543 ) | ( ~w15112 & w15544 ) | ( w15543 & w15544 ) ;
  assign w15546 = w15544 | w15545 ;
  assign w15547 = \pi113 ^ w15099 ;
  assign w15548 = ( ~w15106 & w15546 ) | ( ~w15106 & w15547 ) | ( w15546 & w15547 ) ;
  assign w15549 = w15547 | w15548 ;
  assign w15550 = \pi114 ^ w15093 ;
  assign w15551 = ( ~w15100 & w15549 ) | ( ~w15100 & w15550 ) | ( w15549 & w15550 ) ;
  assign w15552 = w15550 | w15551 ;
  assign w15553 = \pi115 ^ w15087 ;
  assign w15554 = ( ~w15094 & w15552 ) | ( ~w15094 & w15553 ) | ( w15552 & w15553 ) ;
  assign w15555 = w15553 | w15554 ;
  assign w15556 = \pi116 ^ w15081 ;
  assign w15557 = ( ~w15088 & w15555 ) | ( ~w15088 & w15556 ) | ( w15555 & w15556 ) ;
  assign w15558 = w15556 | w15557 ;
  assign w15559 = \pi117 ^ w15075 ;
  assign w15560 = ( ~w15082 & w15558 ) | ( ~w15082 & w15559 ) | ( w15558 & w15559 ) ;
  assign w15561 = w15559 | w15560 ;
  assign w15562 = \pi118 ^ w15069 ;
  assign w15563 = ( ~w15076 & w15561 ) | ( ~w15076 & w15562 ) | ( w15561 & w15562 ) ;
  assign w15564 = w15562 | w15563 ;
  assign w15565 = w14536 & w15064 ;
  assign w15566 = ~w14537 & w15055 ;
  assign w15567 = w15056 ^ w15566 ;
  assign w15568 = ~w15064 & w15567 ;
  assign w15569 = w15565 | w15568 ;
  assign w15570 = ~\pi119 & w15569 ;
  assign w15571 = ( \pi119 & ~w15565 ) | ( \pi119 & w15568 ) | ( ~w15565 & w15568 ) ;
  assign w15572 = ~w15568 & w15571 ;
  assign w15573 = w15570 | w15572 ;
  assign w15574 = ( ~w15070 & w15564 ) | ( ~w15070 & w15573 ) | ( w15564 & w15573 ) ;
  assign w15575 = ( w199 & ~w15573 ) | ( w199 & w15574 ) | ( ~w15573 & w15574 ) ;
  assign w15576 = w15573 | w15575 ;
  assign w15577 = ~w15063 & w15569 ;
  assign w15578 = w15576 & ~w15577 ;
  assign w15579 = ~w15076 & w15561 ;
  assign w15580 = w15562 ^ w15579 ;
  assign w15581 = ~w15578 & w15580 ;
  assign w15582 = ( w15069 & w15576 ) | ( w15069 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15583 = ~w15577 & w15582 ;
  assign w15584 = w15581 | w15583 ;
  assign w15585 = ~\pi119 & w15584 ;
  assign w15586 = ~w15082 & w15558 ;
  assign w15587 = w15559 ^ w15586 ;
  assign w15588 = ~w15578 & w15587 ;
  assign w15589 = ( w15075 & w15576 ) | ( w15075 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15590 = ~w15577 & w15589 ;
  assign w15591 = w15588 | w15590 ;
  assign w15592 = ~\pi118 & w15591 ;
  assign w15593 = ~w15088 & w15555 ;
  assign w15594 = w15556 ^ w15593 ;
  assign w15595 = ~w15578 & w15594 ;
  assign w15596 = ( w15081 & w15576 ) | ( w15081 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15597 = ~w15577 & w15596 ;
  assign w15598 = w15595 | w15597 ;
  assign w15599 = ~\pi117 & w15598 ;
  assign w15600 = ~w15094 & w15552 ;
  assign w15601 = w15553 ^ w15600 ;
  assign w15602 = ~w15578 & w15601 ;
  assign w15603 = ( w15087 & w15576 ) | ( w15087 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15604 = ~w15577 & w15603 ;
  assign w15605 = w15602 | w15604 ;
  assign w15606 = ~\pi116 & w15605 ;
  assign w15607 = ~w15100 & w15549 ;
  assign w15608 = w15550 ^ w15607 ;
  assign w15609 = ~w15578 & w15608 ;
  assign w15610 = ( w15093 & w15576 ) | ( w15093 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15611 = ~w15577 & w15610 ;
  assign w15612 = w15609 | w15611 ;
  assign w15613 = ~\pi115 & w15612 ;
  assign w15614 = ~w15106 & w15546 ;
  assign w15615 = w15547 ^ w15614 ;
  assign w15616 = ~w15578 & w15615 ;
  assign w15617 = ( w15099 & w15576 ) | ( w15099 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15618 = ~w15577 & w15617 ;
  assign w15619 = w15616 | w15618 ;
  assign w15620 = ~\pi114 & w15619 ;
  assign w15621 = ~w15112 & w15543 ;
  assign w15622 = w15544 ^ w15621 ;
  assign w15623 = ~w15578 & w15622 ;
  assign w15624 = ( w15105 & w15576 ) | ( w15105 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15625 = ~w15577 & w15624 ;
  assign w15626 = w15623 | w15625 ;
  assign w15627 = ~\pi113 & w15626 ;
  assign w15628 = ~w15118 & w15540 ;
  assign w15629 = w15541 ^ w15628 ;
  assign w15630 = ~w15578 & w15629 ;
  assign w15631 = ( w15111 & w15576 ) | ( w15111 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15632 = ~w15577 & w15631 ;
  assign w15633 = w15630 | w15632 ;
  assign w15634 = ~\pi112 & w15633 ;
  assign w15635 = ~w15124 & w15537 ;
  assign w15636 = w15538 ^ w15635 ;
  assign w15637 = ~w15578 & w15636 ;
  assign w15638 = ( w15117 & w15576 ) | ( w15117 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15639 = ~w15577 & w15638 ;
  assign w15640 = w15637 | w15639 ;
  assign w15641 = ~\pi111 & w15640 ;
  assign w15642 = ~w15130 & w15534 ;
  assign w15643 = w15535 ^ w15642 ;
  assign w15644 = ~w15578 & w15643 ;
  assign w15645 = ( w15123 & w15576 ) | ( w15123 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15646 = ~w15577 & w15645 ;
  assign w15647 = w15644 | w15646 ;
  assign w15648 = ~\pi110 & w15647 ;
  assign w15649 = ~w15136 & w15531 ;
  assign w15650 = w15532 ^ w15649 ;
  assign w15651 = ~w15578 & w15650 ;
  assign w15652 = ( w15129 & w15576 ) | ( w15129 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15653 = ~w15577 & w15652 ;
  assign w15654 = w15651 | w15653 ;
  assign w15655 = ~\pi109 & w15654 ;
  assign w15656 = ~w15142 & w15528 ;
  assign w15657 = w15529 ^ w15656 ;
  assign w15658 = ~w15578 & w15657 ;
  assign w15659 = ( w15135 & w15576 ) | ( w15135 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15660 = ~w15577 & w15659 ;
  assign w15661 = w15658 | w15660 ;
  assign w15662 = ~\pi108 & w15661 ;
  assign w15663 = ~w15148 & w15525 ;
  assign w15664 = w15526 ^ w15663 ;
  assign w15665 = ~w15578 & w15664 ;
  assign w15666 = ( w15141 & w15576 ) | ( w15141 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15667 = ~w15577 & w15666 ;
  assign w15668 = w15665 | w15667 ;
  assign w15669 = ~\pi107 & w15668 ;
  assign w15670 = ~w15154 & w15522 ;
  assign w15671 = w15523 ^ w15670 ;
  assign w15672 = ~w15578 & w15671 ;
  assign w15673 = ( w15147 & w15576 ) | ( w15147 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15674 = ~w15577 & w15673 ;
  assign w15675 = w15672 | w15674 ;
  assign w15676 = ~\pi106 & w15675 ;
  assign w15677 = ~w15160 & w15519 ;
  assign w15678 = w15520 ^ w15677 ;
  assign w15679 = ~w15578 & w15678 ;
  assign w15680 = ( w15153 & w15576 ) | ( w15153 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15681 = ~w15577 & w15680 ;
  assign w15682 = w15679 | w15681 ;
  assign w15683 = ~\pi105 & w15682 ;
  assign w15684 = ~w15166 & w15516 ;
  assign w15685 = w15517 ^ w15684 ;
  assign w15686 = ~w15578 & w15685 ;
  assign w15687 = ( w15159 & w15576 ) | ( w15159 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15688 = ~w15577 & w15687 ;
  assign w15689 = w15686 | w15688 ;
  assign w15690 = ~\pi104 & w15689 ;
  assign w15691 = ~w15172 & w15513 ;
  assign w15692 = w15514 ^ w15691 ;
  assign w15693 = ~w15578 & w15692 ;
  assign w15694 = ( w15165 & w15576 ) | ( w15165 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15695 = ~w15577 & w15694 ;
  assign w15696 = w15693 | w15695 ;
  assign w15697 = ~\pi103 & w15696 ;
  assign w15698 = ~w15178 & w15510 ;
  assign w15699 = w15511 ^ w15698 ;
  assign w15700 = ~w15578 & w15699 ;
  assign w15701 = ( w15171 & w15576 ) | ( w15171 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15702 = ~w15577 & w15701 ;
  assign w15703 = w15700 | w15702 ;
  assign w15704 = ~\pi102 & w15703 ;
  assign w15705 = ~w15184 & w15507 ;
  assign w15706 = w15508 ^ w15705 ;
  assign w15707 = ~w15578 & w15706 ;
  assign w15708 = ( w15177 & w15576 ) | ( w15177 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15709 = ~w15577 & w15708 ;
  assign w15710 = w15707 | w15709 ;
  assign w15711 = ~\pi101 & w15710 ;
  assign w15712 = ~w15190 & w15504 ;
  assign w15713 = w15505 ^ w15712 ;
  assign w15714 = ~w15578 & w15713 ;
  assign w15715 = ( w15183 & w15576 ) | ( w15183 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15716 = ~w15577 & w15715 ;
  assign w15717 = w15714 | w15716 ;
  assign w15718 = ~\pi100 & w15717 ;
  assign w15719 = ~w15196 & w15501 ;
  assign w15720 = w15502 ^ w15719 ;
  assign w15721 = ~w15578 & w15720 ;
  assign w15722 = ( w15189 & w15576 ) | ( w15189 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15723 = ~w15577 & w15722 ;
  assign w15724 = w15721 | w15723 ;
  assign w15725 = ~\pi099 & w15724 ;
  assign w15726 = ~w15202 & w15498 ;
  assign w15727 = w15499 ^ w15726 ;
  assign w15728 = ~w15578 & w15727 ;
  assign w15729 = ( w15195 & w15576 ) | ( w15195 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15730 = ~w15577 & w15729 ;
  assign w15731 = w15728 | w15730 ;
  assign w15732 = ~\pi098 & w15731 ;
  assign w15733 = ~w15208 & w15495 ;
  assign w15734 = w15496 ^ w15733 ;
  assign w15735 = ~w15578 & w15734 ;
  assign w15736 = ( w15201 & w15576 ) | ( w15201 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15737 = ~w15577 & w15736 ;
  assign w15738 = w15735 | w15737 ;
  assign w15739 = ~\pi097 & w15738 ;
  assign w15740 = ~w15214 & w15492 ;
  assign w15741 = w15493 ^ w15740 ;
  assign w15742 = ~w15578 & w15741 ;
  assign w15743 = ( w15207 & w15576 ) | ( w15207 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15744 = ~w15577 & w15743 ;
  assign w15745 = w15742 | w15744 ;
  assign w15746 = ~\pi096 & w15745 ;
  assign w15747 = ~w15220 & w15489 ;
  assign w15748 = w15490 ^ w15747 ;
  assign w15749 = ~w15578 & w15748 ;
  assign w15750 = ( w15213 & w15576 ) | ( w15213 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15751 = ~w15577 & w15750 ;
  assign w15752 = w15749 | w15751 ;
  assign w15753 = ~\pi095 & w15752 ;
  assign w15754 = ~w15226 & w15486 ;
  assign w15755 = w15487 ^ w15754 ;
  assign w15756 = ~w15578 & w15755 ;
  assign w15757 = ( w15219 & w15576 ) | ( w15219 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15758 = ~w15577 & w15757 ;
  assign w15759 = w15756 | w15758 ;
  assign w15760 = ~\pi094 & w15759 ;
  assign w15761 = ~w15232 & w15483 ;
  assign w15762 = w15484 ^ w15761 ;
  assign w15763 = ~w15578 & w15762 ;
  assign w15764 = ( w15225 & w15576 ) | ( w15225 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15765 = ~w15577 & w15764 ;
  assign w15766 = w15763 | w15765 ;
  assign w15767 = ~\pi093 & w15766 ;
  assign w15768 = ~w15238 & w15480 ;
  assign w15769 = w15481 ^ w15768 ;
  assign w15770 = ~w15578 & w15769 ;
  assign w15771 = ( w15231 & w15576 ) | ( w15231 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15772 = ~w15577 & w15771 ;
  assign w15773 = w15770 | w15772 ;
  assign w15774 = ~\pi092 & w15773 ;
  assign w15775 = ~w15244 & w15477 ;
  assign w15776 = w15478 ^ w15775 ;
  assign w15777 = ~w15578 & w15776 ;
  assign w15778 = ( w15237 & w15576 ) | ( w15237 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15779 = ~w15577 & w15778 ;
  assign w15780 = w15777 | w15779 ;
  assign w15781 = ~\pi091 & w15780 ;
  assign w15782 = ~w15250 & w15474 ;
  assign w15783 = w15475 ^ w15782 ;
  assign w15784 = ~w15578 & w15783 ;
  assign w15785 = ( w15243 & w15576 ) | ( w15243 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15786 = ~w15577 & w15785 ;
  assign w15787 = w15784 | w15786 ;
  assign w15788 = ~\pi090 & w15787 ;
  assign w15789 = ~w15256 & w15471 ;
  assign w15790 = w15472 ^ w15789 ;
  assign w15791 = ~w15578 & w15790 ;
  assign w15792 = ( w15249 & w15576 ) | ( w15249 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15793 = ~w15577 & w15792 ;
  assign w15794 = w15791 | w15793 ;
  assign w15795 = ~\pi089 & w15794 ;
  assign w15796 = ~w15262 & w15468 ;
  assign w15797 = w15469 ^ w15796 ;
  assign w15798 = ~w15578 & w15797 ;
  assign w15799 = ( w15255 & w15576 ) | ( w15255 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15800 = ~w15577 & w15799 ;
  assign w15801 = w15798 | w15800 ;
  assign w15802 = ~\pi088 & w15801 ;
  assign w15803 = ~w15268 & w15465 ;
  assign w15804 = w15466 ^ w15803 ;
  assign w15805 = ~w15578 & w15804 ;
  assign w15806 = ( w15261 & w15576 ) | ( w15261 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15807 = ~w15577 & w15806 ;
  assign w15808 = w15805 | w15807 ;
  assign w15809 = ~\pi087 & w15808 ;
  assign w15810 = ~w15274 & w15462 ;
  assign w15811 = w15463 ^ w15810 ;
  assign w15812 = ~w15578 & w15811 ;
  assign w15813 = ( w15267 & w15576 ) | ( w15267 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15814 = ~w15577 & w15813 ;
  assign w15815 = w15812 | w15814 ;
  assign w15816 = ~\pi086 & w15815 ;
  assign w15817 = ~w15280 & w15459 ;
  assign w15818 = w15460 ^ w15817 ;
  assign w15819 = ~w15578 & w15818 ;
  assign w15820 = ( w15273 & w15576 ) | ( w15273 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15821 = ~w15577 & w15820 ;
  assign w15822 = w15819 | w15821 ;
  assign w15823 = ~\pi085 & w15822 ;
  assign w15824 = ~w15286 & w15456 ;
  assign w15825 = w15457 ^ w15824 ;
  assign w15826 = ~w15578 & w15825 ;
  assign w15827 = ( w15279 & w15576 ) | ( w15279 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15828 = ~w15577 & w15827 ;
  assign w15829 = w15826 | w15828 ;
  assign w15830 = ~\pi084 & w15829 ;
  assign w15831 = ~w15292 & w15453 ;
  assign w15832 = w15454 ^ w15831 ;
  assign w15833 = ~w15578 & w15832 ;
  assign w15834 = ( w15285 & w15576 ) | ( w15285 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15835 = ~w15577 & w15834 ;
  assign w15836 = w15833 | w15835 ;
  assign w15837 = ~\pi083 & w15836 ;
  assign w15838 = ~w15298 & w15450 ;
  assign w15839 = w15451 ^ w15838 ;
  assign w15840 = ~w15578 & w15839 ;
  assign w15841 = ( w15291 & w15576 ) | ( w15291 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15842 = ~w15577 & w15841 ;
  assign w15843 = w15840 | w15842 ;
  assign w15844 = ~\pi082 & w15843 ;
  assign w15845 = ~w15304 & w15447 ;
  assign w15846 = w15448 ^ w15845 ;
  assign w15847 = ~w15578 & w15846 ;
  assign w15848 = ( w15297 & w15576 ) | ( w15297 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15849 = ~w15577 & w15848 ;
  assign w15850 = w15847 | w15849 ;
  assign w15851 = ~\pi081 & w15850 ;
  assign w15852 = ~w15310 & w15444 ;
  assign w15853 = w15445 ^ w15852 ;
  assign w15854 = ~w15578 & w15853 ;
  assign w15855 = ( w15303 & w15576 ) | ( w15303 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15856 = ~w15577 & w15855 ;
  assign w15857 = w15854 | w15856 ;
  assign w15858 = ~\pi080 & w15857 ;
  assign w15859 = ~w15316 & w15441 ;
  assign w15860 = w15442 ^ w15859 ;
  assign w15861 = ~w15578 & w15860 ;
  assign w15862 = ( w15309 & w15576 ) | ( w15309 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15863 = ~w15577 & w15862 ;
  assign w15864 = w15861 | w15863 ;
  assign w15865 = ~\pi079 & w15864 ;
  assign w15866 = ~w15322 & w15438 ;
  assign w15867 = w15439 ^ w15866 ;
  assign w15868 = ~w15578 & w15867 ;
  assign w15869 = ( w15315 & w15576 ) | ( w15315 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15870 = ~w15577 & w15869 ;
  assign w15871 = w15868 | w15870 ;
  assign w15872 = ~\pi078 & w15871 ;
  assign w15873 = ~w15328 & w15435 ;
  assign w15874 = w15436 ^ w15873 ;
  assign w15875 = ~w15578 & w15874 ;
  assign w15876 = ( w15321 & w15576 ) | ( w15321 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15877 = ~w15577 & w15876 ;
  assign w15878 = w15875 | w15877 ;
  assign w15879 = ~\pi077 & w15878 ;
  assign w15880 = ~w15334 & w15432 ;
  assign w15881 = w15433 ^ w15880 ;
  assign w15882 = ~w15578 & w15881 ;
  assign w15883 = ( w15327 & w15576 ) | ( w15327 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15884 = ~w15577 & w15883 ;
  assign w15885 = w15882 | w15884 ;
  assign w15886 = ~\pi076 & w15885 ;
  assign w15887 = ~w15340 & w15429 ;
  assign w15888 = w15430 ^ w15887 ;
  assign w15889 = ~w15578 & w15888 ;
  assign w15890 = ( w15333 & w15576 ) | ( w15333 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15891 = ~w15577 & w15890 ;
  assign w15892 = w15889 | w15891 ;
  assign w15893 = ~\pi075 & w15892 ;
  assign w15894 = ~w15346 & w15426 ;
  assign w15895 = w15427 ^ w15894 ;
  assign w15896 = ~w15578 & w15895 ;
  assign w15897 = ( w15339 & w15576 ) | ( w15339 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15898 = ~w15577 & w15897 ;
  assign w15899 = w15896 | w15898 ;
  assign w15900 = ~\pi074 & w15899 ;
  assign w15901 = ~w15352 & w15423 ;
  assign w15902 = w15424 ^ w15901 ;
  assign w15903 = ~w15578 & w15902 ;
  assign w15904 = ( w15345 & w15576 ) | ( w15345 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15905 = ~w15577 & w15904 ;
  assign w15906 = w15903 | w15905 ;
  assign w15907 = ~\pi073 & w15906 ;
  assign w15908 = ~w15358 & w15420 ;
  assign w15909 = w15421 ^ w15908 ;
  assign w15910 = ~w15578 & w15909 ;
  assign w15911 = ( w15351 & w15576 ) | ( w15351 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15912 = ~w15577 & w15911 ;
  assign w15913 = w15910 | w15912 ;
  assign w15914 = ~\pi072 & w15913 ;
  assign w15915 = ~w15364 & w15417 ;
  assign w15916 = w15418 ^ w15915 ;
  assign w15917 = ~w15578 & w15916 ;
  assign w15918 = ( w15357 & w15576 ) | ( w15357 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15919 = ~w15577 & w15918 ;
  assign w15920 = w15917 | w15919 ;
  assign w15921 = ~\pi071 & w15920 ;
  assign w15922 = ~w15370 & w15414 ;
  assign w15923 = w15415 ^ w15922 ;
  assign w15924 = ~w15578 & w15923 ;
  assign w15925 = ( w15363 & w15576 ) | ( w15363 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15926 = ~w15577 & w15925 ;
  assign w15927 = w15924 | w15926 ;
  assign w15928 = ~\pi070 & w15927 ;
  assign w15929 = ~w15378 & w15411 ;
  assign w15930 = w15412 ^ w15929 ;
  assign w15931 = ~w15578 & w15930 ;
  assign w15932 = ( w15369 & w15576 ) | ( w15369 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15933 = ~w15577 & w15932 ;
  assign w15934 = w15931 | w15933 ;
  assign w15935 = ~\pi069 & w15934 ;
  assign w15936 = ~w15389 & w15406 ;
  assign w15937 = w15409 ^ w15936 ;
  assign w15938 = ~w15578 & w15937 ;
  assign w15939 = ( w15377 & w15576 ) | ( w15377 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15940 = ~w15577 & w15939 ;
  assign w15941 = w15938 | w15940 ;
  assign w15942 = ~\pi068 & w15941 ;
  assign w15943 = w15403 ^ w15405 ;
  assign w15944 = ~w15578 & w15943 ;
  assign w15945 = ( w15388 & w15576 ) | ( w15388 & w15577 ) | ( w15576 & w15577 ) ;
  assign w15946 = ~w15577 & w15945 ;
  assign w15947 = w15944 | w15946 ;
  assign w15948 = ~\pi067 & w15947 ;
  assign w15949 = w15400 ^ w15404 ;
  assign w15950 = \pi065 ^ w15949 ;
  assign w15951 = ~w15578 & w15950 ;
  assign w15952 = ( w15394 & w15399 ) | ( w15394 & ~w15577 ) | ( w15399 & ~w15577 ) ;
  assign w15953 = w15577 & w15952 ;
  assign w15954 = ( ~w15576 & w15952 ) | ( ~w15576 & w15953 ) | ( w15952 & w15953 ) ;
  assign w15955 = ( w15951 & w15952 ) | ( w15951 & ~w15954 ) | ( w15952 & ~w15954 ) ;
  assign w15956 = ~\pi066 & w15955 ;
  assign w15957 = w15576 | w15577 ;
  assign w15958 = ( w15951 & w15952 ) | ( w15951 & w15957 ) | ( w15952 & w15957 ) ;
  assign w15959 = ( ~w15577 & w15951 ) | ( ~w15577 & w15958 ) | ( w15951 & w15958 ) ;
  assign w15960 = \pi066 ^ w15959 ;
  assign w15961 = \pi064 & ~w15578 ;
  assign w15962 = \pi008 ^ w15961 ;
  assign w15963 = ( ~\pi007 & \pi064 ) | ( ~\pi007 & w15960 ) | ( \pi064 & w15960 ) ;
  assign w15964 = ( \pi065 & ~w15962 ) | ( \pi065 & w15963 ) | ( ~w15962 & w15963 ) ;
  assign w15965 = w15960 | w15964 ;
  assign w15966 = \pi067 ^ w15947 ;
  assign w15967 = ( ~w15956 & w15965 ) | ( ~w15956 & w15966 ) | ( w15965 & w15966 ) ;
  assign w15968 = w15966 | w15967 ;
  assign w15969 = \pi068 ^ w15941 ;
  assign w15970 = ( ~w15948 & w15968 ) | ( ~w15948 & w15969 ) | ( w15968 & w15969 ) ;
  assign w15971 = w15969 | w15970 ;
  assign w15972 = \pi069 ^ w15934 ;
  assign w15973 = ( ~w15942 & w15971 ) | ( ~w15942 & w15972 ) | ( w15971 & w15972 ) ;
  assign w15974 = w15972 | w15973 ;
  assign w15975 = \pi070 ^ w15927 ;
  assign w15976 = ( ~w15935 & w15974 ) | ( ~w15935 & w15975 ) | ( w15974 & w15975 ) ;
  assign w15977 = w15975 | w15976 ;
  assign w15978 = \pi071 ^ w15920 ;
  assign w15979 = ( ~w15928 & w15977 ) | ( ~w15928 & w15978 ) | ( w15977 & w15978 ) ;
  assign w15980 = w15978 | w15979 ;
  assign w15981 = \pi072 ^ w15913 ;
  assign w15982 = ( ~w15921 & w15980 ) | ( ~w15921 & w15981 ) | ( w15980 & w15981 ) ;
  assign w15983 = w15981 | w15982 ;
  assign w15984 = \pi073 ^ w15906 ;
  assign w15985 = ( ~w15914 & w15983 ) | ( ~w15914 & w15984 ) | ( w15983 & w15984 ) ;
  assign w15986 = w15984 | w15985 ;
  assign w15987 = \pi074 ^ w15899 ;
  assign w15988 = ( ~w15907 & w15986 ) | ( ~w15907 & w15987 ) | ( w15986 & w15987 ) ;
  assign w15989 = w15987 | w15988 ;
  assign w15990 = \pi075 ^ w15892 ;
  assign w15991 = ( ~w15900 & w15989 ) | ( ~w15900 & w15990 ) | ( w15989 & w15990 ) ;
  assign w15992 = w15990 | w15991 ;
  assign w15993 = \pi076 ^ w15885 ;
  assign w15994 = ( ~w15893 & w15992 ) | ( ~w15893 & w15993 ) | ( w15992 & w15993 ) ;
  assign w15995 = w15993 | w15994 ;
  assign w15996 = \pi077 ^ w15878 ;
  assign w15997 = ( ~w15886 & w15995 ) | ( ~w15886 & w15996 ) | ( w15995 & w15996 ) ;
  assign w15998 = w15996 | w15997 ;
  assign w15999 = \pi078 ^ w15871 ;
  assign w16000 = ( ~w15879 & w15998 ) | ( ~w15879 & w15999 ) | ( w15998 & w15999 ) ;
  assign w16001 = w15999 | w16000 ;
  assign w16002 = \pi079 ^ w15864 ;
  assign w16003 = ( ~w15872 & w16001 ) | ( ~w15872 & w16002 ) | ( w16001 & w16002 ) ;
  assign w16004 = w16002 | w16003 ;
  assign w16005 = \pi080 ^ w15857 ;
  assign w16006 = ( ~w15865 & w16004 ) | ( ~w15865 & w16005 ) | ( w16004 & w16005 ) ;
  assign w16007 = w16005 | w16006 ;
  assign w16008 = \pi081 ^ w15850 ;
  assign w16009 = ( ~w15858 & w16007 ) | ( ~w15858 & w16008 ) | ( w16007 & w16008 ) ;
  assign w16010 = w16008 | w16009 ;
  assign w16011 = \pi082 ^ w15843 ;
  assign w16012 = ( ~w15851 & w16010 ) | ( ~w15851 & w16011 ) | ( w16010 & w16011 ) ;
  assign w16013 = w16011 | w16012 ;
  assign w16014 = \pi083 ^ w15836 ;
  assign w16015 = ( ~w15844 & w16013 ) | ( ~w15844 & w16014 ) | ( w16013 & w16014 ) ;
  assign w16016 = w16014 | w16015 ;
  assign w16017 = \pi084 ^ w15829 ;
  assign w16018 = ( ~w15837 & w16016 ) | ( ~w15837 & w16017 ) | ( w16016 & w16017 ) ;
  assign w16019 = w16017 | w16018 ;
  assign w16020 = \pi085 ^ w15822 ;
  assign w16021 = ( ~w15830 & w16019 ) | ( ~w15830 & w16020 ) | ( w16019 & w16020 ) ;
  assign w16022 = w16020 | w16021 ;
  assign w16023 = \pi086 ^ w15815 ;
  assign w16024 = ( ~w15823 & w16022 ) | ( ~w15823 & w16023 ) | ( w16022 & w16023 ) ;
  assign w16025 = w16023 | w16024 ;
  assign w16026 = \pi087 ^ w15808 ;
  assign w16027 = ( ~w15816 & w16025 ) | ( ~w15816 & w16026 ) | ( w16025 & w16026 ) ;
  assign w16028 = w16026 | w16027 ;
  assign w16029 = \pi088 ^ w15801 ;
  assign w16030 = ( ~w15809 & w16028 ) | ( ~w15809 & w16029 ) | ( w16028 & w16029 ) ;
  assign w16031 = w16029 | w16030 ;
  assign w16032 = \pi089 ^ w15794 ;
  assign w16033 = ( ~w15802 & w16031 ) | ( ~w15802 & w16032 ) | ( w16031 & w16032 ) ;
  assign w16034 = w16032 | w16033 ;
  assign w16035 = \pi090 ^ w15787 ;
  assign w16036 = ( ~w15795 & w16034 ) | ( ~w15795 & w16035 ) | ( w16034 & w16035 ) ;
  assign w16037 = w16035 | w16036 ;
  assign w16038 = \pi091 ^ w15780 ;
  assign w16039 = ( ~w15788 & w16037 ) | ( ~w15788 & w16038 ) | ( w16037 & w16038 ) ;
  assign w16040 = w16038 | w16039 ;
  assign w16041 = \pi092 ^ w15773 ;
  assign w16042 = ( ~w15781 & w16040 ) | ( ~w15781 & w16041 ) | ( w16040 & w16041 ) ;
  assign w16043 = w16041 | w16042 ;
  assign w16044 = \pi093 ^ w15766 ;
  assign w16045 = ( ~w15774 & w16043 ) | ( ~w15774 & w16044 ) | ( w16043 & w16044 ) ;
  assign w16046 = w16044 | w16045 ;
  assign w16047 = \pi094 ^ w15759 ;
  assign w16048 = ( ~w15767 & w16046 ) | ( ~w15767 & w16047 ) | ( w16046 & w16047 ) ;
  assign w16049 = w16047 | w16048 ;
  assign w16050 = \pi095 ^ w15752 ;
  assign w16051 = ( ~w15760 & w16049 ) | ( ~w15760 & w16050 ) | ( w16049 & w16050 ) ;
  assign w16052 = w16050 | w16051 ;
  assign w16053 = \pi096 ^ w15745 ;
  assign w16054 = ( ~w15753 & w16052 ) | ( ~w15753 & w16053 ) | ( w16052 & w16053 ) ;
  assign w16055 = w16053 | w16054 ;
  assign w16056 = \pi097 ^ w15738 ;
  assign w16057 = ( ~w15746 & w16055 ) | ( ~w15746 & w16056 ) | ( w16055 & w16056 ) ;
  assign w16058 = w16056 | w16057 ;
  assign w16059 = \pi098 ^ w15731 ;
  assign w16060 = ( ~w15739 & w16058 ) | ( ~w15739 & w16059 ) | ( w16058 & w16059 ) ;
  assign w16061 = w16059 | w16060 ;
  assign w16062 = \pi099 ^ w15724 ;
  assign w16063 = ( ~w15732 & w16061 ) | ( ~w15732 & w16062 ) | ( w16061 & w16062 ) ;
  assign w16064 = w16062 | w16063 ;
  assign w16065 = \pi100 ^ w15717 ;
  assign w16066 = ( ~w15725 & w16064 ) | ( ~w15725 & w16065 ) | ( w16064 & w16065 ) ;
  assign w16067 = w16065 | w16066 ;
  assign w16068 = \pi101 ^ w15710 ;
  assign w16069 = ( ~w15718 & w16067 ) | ( ~w15718 & w16068 ) | ( w16067 & w16068 ) ;
  assign w16070 = w16068 | w16069 ;
  assign w16071 = \pi102 ^ w15703 ;
  assign w16072 = ( ~w15711 & w16070 ) | ( ~w15711 & w16071 ) | ( w16070 & w16071 ) ;
  assign w16073 = w16071 | w16072 ;
  assign w16074 = \pi103 ^ w15696 ;
  assign w16075 = ( ~w15704 & w16073 ) | ( ~w15704 & w16074 ) | ( w16073 & w16074 ) ;
  assign w16076 = w16074 | w16075 ;
  assign w16077 = \pi104 ^ w15689 ;
  assign w16078 = ( ~w15697 & w16076 ) | ( ~w15697 & w16077 ) | ( w16076 & w16077 ) ;
  assign w16079 = w16077 | w16078 ;
  assign w16080 = \pi105 ^ w15682 ;
  assign w16081 = ( ~w15690 & w16079 ) | ( ~w15690 & w16080 ) | ( w16079 & w16080 ) ;
  assign w16082 = w16080 | w16081 ;
  assign w16083 = \pi106 ^ w15675 ;
  assign w16084 = ( ~w15683 & w16082 ) | ( ~w15683 & w16083 ) | ( w16082 & w16083 ) ;
  assign w16085 = w16083 | w16084 ;
  assign w16086 = \pi107 ^ w15668 ;
  assign w16087 = ( ~w15676 & w16085 ) | ( ~w15676 & w16086 ) | ( w16085 & w16086 ) ;
  assign w16088 = w16086 | w16087 ;
  assign w16089 = \pi108 ^ w15661 ;
  assign w16090 = ( ~w15669 & w16088 ) | ( ~w15669 & w16089 ) | ( w16088 & w16089 ) ;
  assign w16091 = w16089 | w16090 ;
  assign w16092 = \pi109 ^ w15654 ;
  assign w16093 = ( ~w15662 & w16091 ) | ( ~w15662 & w16092 ) | ( w16091 & w16092 ) ;
  assign w16094 = w16092 | w16093 ;
  assign w16095 = \pi110 ^ w15647 ;
  assign w16096 = ( ~w15655 & w16094 ) | ( ~w15655 & w16095 ) | ( w16094 & w16095 ) ;
  assign w16097 = w16095 | w16096 ;
  assign w16098 = \pi111 ^ w15640 ;
  assign w16099 = ( ~w15648 & w16097 ) | ( ~w15648 & w16098 ) | ( w16097 & w16098 ) ;
  assign w16100 = w16098 | w16099 ;
  assign w16101 = \pi112 ^ w15633 ;
  assign w16102 = ( ~w15641 & w16100 ) | ( ~w15641 & w16101 ) | ( w16100 & w16101 ) ;
  assign w16103 = w16101 | w16102 ;
  assign w16104 = \pi113 ^ w15626 ;
  assign w16105 = ( ~w15634 & w16103 ) | ( ~w15634 & w16104 ) | ( w16103 & w16104 ) ;
  assign w16106 = w16104 | w16105 ;
  assign w16107 = \pi114 ^ w15619 ;
  assign w16108 = ( ~w15627 & w16106 ) | ( ~w15627 & w16107 ) | ( w16106 & w16107 ) ;
  assign w16109 = w16107 | w16108 ;
  assign w16110 = \pi115 ^ w15612 ;
  assign w16111 = ( ~w15620 & w16109 ) | ( ~w15620 & w16110 ) | ( w16109 & w16110 ) ;
  assign w16112 = w16110 | w16111 ;
  assign w16113 = \pi116 ^ w15605 ;
  assign w16114 = ( ~w15613 & w16112 ) | ( ~w15613 & w16113 ) | ( w16112 & w16113 ) ;
  assign w16115 = w16113 | w16114 ;
  assign w16116 = \pi117 ^ w15598 ;
  assign w16117 = ( ~w15606 & w16115 ) | ( ~w15606 & w16116 ) | ( w16115 & w16116 ) ;
  assign w16118 = w16116 | w16117 ;
  assign w16119 = \pi118 ^ w15591 ;
  assign w16120 = ( ~w15599 & w16118 ) | ( ~w15599 & w16119 ) | ( w16118 & w16119 ) ;
  assign w16121 = w16119 | w16120 ;
  assign w16122 = \pi119 ^ w15584 ;
  assign w16123 = ( ~w15592 & w16121 ) | ( ~w15592 & w16122 ) | ( w16121 & w16122 ) ;
  assign w16124 = w16122 | w16123 ;
  assign w16125 = ( ~w15070 & w15564 ) | ( ~w15070 & w15578 ) | ( w15564 & w15578 ) ;
  assign w16126 = w15573 ^ w16125 ;
  assign w16127 = ~w15578 & w16126 ;
  assign w16128 = ( w15063 & ~w15569 ) | ( w15063 & w15576 ) | ( ~w15569 & w15576 ) ;
  assign w16129 = w15569 & w16128 ;
  assign w16130 = w16127 | w16129 ;
  assign w16131 = ~\pi120 & w16130 ;
  assign w16132 = ( \pi120 & ~w16127 ) | ( \pi120 & w16129 ) | ( ~w16127 & w16129 ) ;
  assign w16133 = ~w16129 & w16132 ;
  assign w16134 = w16131 | w16133 ;
  assign w16135 = ( ~w15585 & w16124 ) | ( ~w15585 & w16134 ) | ( w16124 & w16134 ) ;
  assign w16136 = ( w273 & ~w16134 ) | ( w273 & w16135 ) | ( ~w16134 & w16135 ) ;
  assign w16137 = w16134 | w16136 ;
  assign w16138 = ~w199 & w16130 ;
  assign w16139 = w16137 & ~w16138 ;
  assign w16140 = ~w15592 & w16121 ;
  assign w16141 = w16122 ^ w16140 ;
  assign w16142 = ~w16139 & w16141 ;
  assign w16143 = ( w15584 & w16137 ) | ( w15584 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16144 = ~w16138 & w16143 ;
  assign w16145 = w16142 | w16144 ;
  assign w16146 = ( ~w15585 & w16124 ) | ( ~w15585 & w16139 ) | ( w16124 & w16139 ) ;
  assign w16147 = w16134 ^ w16146 ;
  assign w16148 = ~w16139 & w16147 ;
  assign w16149 = ( w199 & ~w16130 ) | ( w199 & w16137 ) | ( ~w16130 & w16137 ) ;
  assign w16150 = w16130 & w16149 ;
  assign w16151 = w16148 | w16150 ;
  assign w16152 = ~\pi120 & w16145 ;
  assign w16153 = ~w15599 & w16118 ;
  assign w16154 = w16119 ^ w16153 ;
  assign w16155 = ~w16139 & w16154 ;
  assign w16156 = ( w15591 & w16137 ) | ( w15591 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16157 = ~w16138 & w16156 ;
  assign w16158 = w16155 | w16157 ;
  assign w16159 = ~\pi119 & w16158 ;
  assign w16160 = ~w15606 & w16115 ;
  assign w16161 = w16116 ^ w16160 ;
  assign w16162 = ~w16139 & w16161 ;
  assign w16163 = ( w15598 & w16137 ) | ( w15598 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16164 = ~w16138 & w16163 ;
  assign w16165 = w16162 | w16164 ;
  assign w16166 = ~\pi118 & w16165 ;
  assign w16167 = ~w15613 & w16112 ;
  assign w16168 = w16113 ^ w16167 ;
  assign w16169 = ~w16139 & w16168 ;
  assign w16170 = ( w15605 & w16137 ) | ( w15605 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16171 = ~w16138 & w16170 ;
  assign w16172 = w16169 | w16171 ;
  assign w16173 = ~\pi117 & w16172 ;
  assign w16174 = ~w15620 & w16109 ;
  assign w16175 = w16110 ^ w16174 ;
  assign w16176 = ~w16139 & w16175 ;
  assign w16177 = ( w15612 & w16137 ) | ( w15612 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16178 = ~w16138 & w16177 ;
  assign w16179 = w16176 | w16178 ;
  assign w16180 = ~\pi116 & w16179 ;
  assign w16181 = ~w15627 & w16106 ;
  assign w16182 = w16107 ^ w16181 ;
  assign w16183 = ~w16139 & w16182 ;
  assign w16184 = ( w15619 & w16137 ) | ( w15619 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16185 = ~w16138 & w16184 ;
  assign w16186 = w16183 | w16185 ;
  assign w16187 = ~\pi115 & w16186 ;
  assign w16188 = ~w15634 & w16103 ;
  assign w16189 = w16104 ^ w16188 ;
  assign w16190 = ~w16139 & w16189 ;
  assign w16191 = ( w15626 & w16137 ) | ( w15626 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16192 = ~w16138 & w16191 ;
  assign w16193 = w16190 | w16192 ;
  assign w16194 = ~\pi114 & w16193 ;
  assign w16195 = ~w15641 & w16100 ;
  assign w16196 = w16101 ^ w16195 ;
  assign w16197 = ~w16139 & w16196 ;
  assign w16198 = ( w15633 & w16137 ) | ( w15633 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16199 = ~w16138 & w16198 ;
  assign w16200 = w16197 | w16199 ;
  assign w16201 = ~\pi113 & w16200 ;
  assign w16202 = ~w15648 & w16097 ;
  assign w16203 = w16098 ^ w16202 ;
  assign w16204 = ~w16139 & w16203 ;
  assign w16205 = ( w15640 & w16137 ) | ( w15640 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16206 = ~w16138 & w16205 ;
  assign w16207 = w16204 | w16206 ;
  assign w16208 = ~\pi112 & w16207 ;
  assign w16209 = ~w15655 & w16094 ;
  assign w16210 = w16095 ^ w16209 ;
  assign w16211 = ~w16139 & w16210 ;
  assign w16212 = ( w15647 & w16137 ) | ( w15647 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16213 = ~w16138 & w16212 ;
  assign w16214 = w16211 | w16213 ;
  assign w16215 = ~\pi111 & w16214 ;
  assign w16216 = ~w15662 & w16091 ;
  assign w16217 = w16092 ^ w16216 ;
  assign w16218 = ~w16139 & w16217 ;
  assign w16219 = ( w15654 & w16137 ) | ( w15654 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16220 = ~w16138 & w16219 ;
  assign w16221 = w16218 | w16220 ;
  assign w16222 = ~\pi110 & w16221 ;
  assign w16223 = ~w15669 & w16088 ;
  assign w16224 = w16089 ^ w16223 ;
  assign w16225 = ~w16139 & w16224 ;
  assign w16226 = ( w15661 & w16137 ) | ( w15661 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16227 = ~w16138 & w16226 ;
  assign w16228 = w16225 | w16227 ;
  assign w16229 = ~\pi109 & w16228 ;
  assign w16230 = ~w15676 & w16085 ;
  assign w16231 = w16086 ^ w16230 ;
  assign w16232 = ~w16139 & w16231 ;
  assign w16233 = ( w15668 & w16137 ) | ( w15668 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16234 = ~w16138 & w16233 ;
  assign w16235 = w16232 | w16234 ;
  assign w16236 = ~\pi108 & w16235 ;
  assign w16237 = ~w15683 & w16082 ;
  assign w16238 = w16083 ^ w16237 ;
  assign w16239 = ~w16139 & w16238 ;
  assign w16240 = ( w15675 & w16137 ) | ( w15675 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16241 = ~w16138 & w16240 ;
  assign w16242 = w16239 | w16241 ;
  assign w16243 = ~\pi107 & w16242 ;
  assign w16244 = ~w15690 & w16079 ;
  assign w16245 = w16080 ^ w16244 ;
  assign w16246 = ~w16139 & w16245 ;
  assign w16247 = ( w15682 & w16137 ) | ( w15682 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16248 = ~w16138 & w16247 ;
  assign w16249 = w16246 | w16248 ;
  assign w16250 = ~\pi106 & w16249 ;
  assign w16251 = ~w15697 & w16076 ;
  assign w16252 = w16077 ^ w16251 ;
  assign w16253 = ~w16139 & w16252 ;
  assign w16254 = ( w15689 & w16137 ) | ( w15689 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16255 = ~w16138 & w16254 ;
  assign w16256 = w16253 | w16255 ;
  assign w16257 = ~\pi105 & w16256 ;
  assign w16258 = ~w15704 & w16073 ;
  assign w16259 = w16074 ^ w16258 ;
  assign w16260 = ~w16139 & w16259 ;
  assign w16261 = ( w15696 & w16137 ) | ( w15696 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16262 = ~w16138 & w16261 ;
  assign w16263 = w16260 | w16262 ;
  assign w16264 = ~\pi104 & w16263 ;
  assign w16265 = ~w15711 & w16070 ;
  assign w16266 = w16071 ^ w16265 ;
  assign w16267 = ~w16139 & w16266 ;
  assign w16268 = ( w15703 & w16137 ) | ( w15703 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16269 = ~w16138 & w16268 ;
  assign w16270 = w16267 | w16269 ;
  assign w16271 = ~\pi103 & w16270 ;
  assign w16272 = ~w15718 & w16067 ;
  assign w16273 = w16068 ^ w16272 ;
  assign w16274 = ~w16139 & w16273 ;
  assign w16275 = ( w15710 & w16137 ) | ( w15710 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16276 = ~w16138 & w16275 ;
  assign w16277 = w16274 | w16276 ;
  assign w16278 = ~\pi102 & w16277 ;
  assign w16279 = ~w15725 & w16064 ;
  assign w16280 = w16065 ^ w16279 ;
  assign w16281 = ~w16139 & w16280 ;
  assign w16282 = ( w15717 & w16137 ) | ( w15717 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16283 = ~w16138 & w16282 ;
  assign w16284 = w16281 | w16283 ;
  assign w16285 = ~\pi101 & w16284 ;
  assign w16286 = ~w15732 & w16061 ;
  assign w16287 = w16062 ^ w16286 ;
  assign w16288 = ~w16139 & w16287 ;
  assign w16289 = ( w15724 & w16137 ) | ( w15724 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16290 = ~w16138 & w16289 ;
  assign w16291 = w16288 | w16290 ;
  assign w16292 = ~\pi100 & w16291 ;
  assign w16293 = ~w15739 & w16058 ;
  assign w16294 = w16059 ^ w16293 ;
  assign w16295 = ~w16139 & w16294 ;
  assign w16296 = ( w15731 & w16137 ) | ( w15731 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16297 = ~w16138 & w16296 ;
  assign w16298 = w16295 | w16297 ;
  assign w16299 = ~\pi099 & w16298 ;
  assign w16300 = ~w15746 & w16055 ;
  assign w16301 = w16056 ^ w16300 ;
  assign w16302 = ~w16139 & w16301 ;
  assign w16303 = ( w15738 & w16137 ) | ( w15738 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16304 = ~w16138 & w16303 ;
  assign w16305 = w16302 | w16304 ;
  assign w16306 = ~\pi098 & w16305 ;
  assign w16307 = ~w15753 & w16052 ;
  assign w16308 = w16053 ^ w16307 ;
  assign w16309 = ~w16139 & w16308 ;
  assign w16310 = ( w15745 & w16137 ) | ( w15745 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16311 = ~w16138 & w16310 ;
  assign w16312 = w16309 | w16311 ;
  assign w16313 = ~\pi097 & w16312 ;
  assign w16314 = ~w15760 & w16049 ;
  assign w16315 = w16050 ^ w16314 ;
  assign w16316 = ~w16139 & w16315 ;
  assign w16317 = ( w15752 & w16137 ) | ( w15752 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16318 = ~w16138 & w16317 ;
  assign w16319 = w16316 | w16318 ;
  assign w16320 = ~\pi096 & w16319 ;
  assign w16321 = ~w15767 & w16046 ;
  assign w16322 = w16047 ^ w16321 ;
  assign w16323 = ~w16139 & w16322 ;
  assign w16324 = ( w15759 & w16137 ) | ( w15759 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16325 = ~w16138 & w16324 ;
  assign w16326 = w16323 | w16325 ;
  assign w16327 = ~\pi095 & w16326 ;
  assign w16328 = ~w15774 & w16043 ;
  assign w16329 = w16044 ^ w16328 ;
  assign w16330 = ~w16139 & w16329 ;
  assign w16331 = ( w15766 & w16137 ) | ( w15766 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16332 = ~w16138 & w16331 ;
  assign w16333 = w16330 | w16332 ;
  assign w16334 = ~\pi094 & w16333 ;
  assign w16335 = ~w15781 & w16040 ;
  assign w16336 = w16041 ^ w16335 ;
  assign w16337 = ~w16139 & w16336 ;
  assign w16338 = ( w15773 & w16137 ) | ( w15773 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16339 = ~w16138 & w16338 ;
  assign w16340 = w16337 | w16339 ;
  assign w16341 = ~\pi093 & w16340 ;
  assign w16342 = ~w15788 & w16037 ;
  assign w16343 = w16038 ^ w16342 ;
  assign w16344 = ~w16139 & w16343 ;
  assign w16345 = ( w15780 & w16137 ) | ( w15780 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16346 = ~w16138 & w16345 ;
  assign w16347 = w16344 | w16346 ;
  assign w16348 = ~\pi092 & w16347 ;
  assign w16349 = ~w15795 & w16034 ;
  assign w16350 = w16035 ^ w16349 ;
  assign w16351 = ~w16139 & w16350 ;
  assign w16352 = ( w15787 & w16137 ) | ( w15787 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16353 = ~w16138 & w16352 ;
  assign w16354 = w16351 | w16353 ;
  assign w16355 = ~\pi091 & w16354 ;
  assign w16356 = ~w15802 & w16031 ;
  assign w16357 = w16032 ^ w16356 ;
  assign w16358 = ~w16139 & w16357 ;
  assign w16359 = ( w15794 & w16137 ) | ( w15794 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16360 = ~w16138 & w16359 ;
  assign w16361 = w16358 | w16360 ;
  assign w16362 = ~\pi090 & w16361 ;
  assign w16363 = ~w15809 & w16028 ;
  assign w16364 = w16029 ^ w16363 ;
  assign w16365 = ~w16139 & w16364 ;
  assign w16366 = ( w15801 & w16137 ) | ( w15801 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16367 = ~w16138 & w16366 ;
  assign w16368 = w16365 | w16367 ;
  assign w16369 = ~\pi089 & w16368 ;
  assign w16370 = ~w15816 & w16025 ;
  assign w16371 = w16026 ^ w16370 ;
  assign w16372 = ~w16139 & w16371 ;
  assign w16373 = ( w15808 & w16137 ) | ( w15808 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16374 = ~w16138 & w16373 ;
  assign w16375 = w16372 | w16374 ;
  assign w16376 = ~\pi088 & w16375 ;
  assign w16377 = ~w15823 & w16022 ;
  assign w16378 = w16023 ^ w16377 ;
  assign w16379 = ~w16139 & w16378 ;
  assign w16380 = ( w15815 & w16137 ) | ( w15815 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16381 = ~w16138 & w16380 ;
  assign w16382 = w16379 | w16381 ;
  assign w16383 = ~\pi087 & w16382 ;
  assign w16384 = ~w15830 & w16019 ;
  assign w16385 = w16020 ^ w16384 ;
  assign w16386 = ~w16139 & w16385 ;
  assign w16387 = ( w15822 & w16137 ) | ( w15822 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16388 = ~w16138 & w16387 ;
  assign w16389 = w16386 | w16388 ;
  assign w16390 = ~\pi086 & w16389 ;
  assign w16391 = ~w15837 & w16016 ;
  assign w16392 = w16017 ^ w16391 ;
  assign w16393 = ~w16139 & w16392 ;
  assign w16394 = ( w15829 & w16137 ) | ( w15829 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16395 = ~w16138 & w16394 ;
  assign w16396 = w16393 | w16395 ;
  assign w16397 = ~\pi085 & w16396 ;
  assign w16398 = ~w15844 & w16013 ;
  assign w16399 = w16014 ^ w16398 ;
  assign w16400 = ~w16139 & w16399 ;
  assign w16401 = ( w15836 & w16137 ) | ( w15836 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16402 = ~w16138 & w16401 ;
  assign w16403 = w16400 | w16402 ;
  assign w16404 = ~\pi084 & w16403 ;
  assign w16405 = ~w15851 & w16010 ;
  assign w16406 = w16011 ^ w16405 ;
  assign w16407 = ~w16139 & w16406 ;
  assign w16408 = ( w15843 & w16137 ) | ( w15843 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16409 = ~w16138 & w16408 ;
  assign w16410 = w16407 | w16409 ;
  assign w16411 = ~\pi083 & w16410 ;
  assign w16412 = ~w15858 & w16007 ;
  assign w16413 = w16008 ^ w16412 ;
  assign w16414 = ~w16139 & w16413 ;
  assign w16415 = ( w15850 & w16137 ) | ( w15850 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16416 = ~w16138 & w16415 ;
  assign w16417 = w16414 | w16416 ;
  assign w16418 = ~\pi082 & w16417 ;
  assign w16419 = ~w15865 & w16004 ;
  assign w16420 = w16005 ^ w16419 ;
  assign w16421 = ~w16139 & w16420 ;
  assign w16422 = ( w15857 & w16137 ) | ( w15857 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16423 = ~w16138 & w16422 ;
  assign w16424 = w16421 | w16423 ;
  assign w16425 = ~\pi081 & w16424 ;
  assign w16426 = ~w15872 & w16001 ;
  assign w16427 = w16002 ^ w16426 ;
  assign w16428 = ~w16139 & w16427 ;
  assign w16429 = ( w15864 & w16137 ) | ( w15864 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16430 = ~w16138 & w16429 ;
  assign w16431 = w16428 | w16430 ;
  assign w16432 = ~\pi080 & w16431 ;
  assign w16433 = ~w15879 & w15998 ;
  assign w16434 = w15999 ^ w16433 ;
  assign w16435 = ~w16139 & w16434 ;
  assign w16436 = ( w15871 & w16137 ) | ( w15871 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16437 = ~w16138 & w16436 ;
  assign w16438 = w16435 | w16437 ;
  assign w16439 = ~\pi079 & w16438 ;
  assign w16440 = ~w15886 & w15995 ;
  assign w16441 = w15996 ^ w16440 ;
  assign w16442 = ~w16139 & w16441 ;
  assign w16443 = ( w15878 & w16137 ) | ( w15878 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16444 = ~w16138 & w16443 ;
  assign w16445 = w16442 | w16444 ;
  assign w16446 = ~\pi078 & w16445 ;
  assign w16447 = ~w15893 & w15992 ;
  assign w16448 = w15993 ^ w16447 ;
  assign w16449 = ~w16139 & w16448 ;
  assign w16450 = ( w15885 & w16137 ) | ( w15885 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16451 = ~w16138 & w16450 ;
  assign w16452 = w16449 | w16451 ;
  assign w16453 = ~\pi077 & w16452 ;
  assign w16454 = ~w15900 & w15989 ;
  assign w16455 = w15990 ^ w16454 ;
  assign w16456 = ~w16139 & w16455 ;
  assign w16457 = ( w15892 & w16137 ) | ( w15892 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16458 = ~w16138 & w16457 ;
  assign w16459 = w16456 | w16458 ;
  assign w16460 = ~\pi076 & w16459 ;
  assign w16461 = ~w15907 & w15986 ;
  assign w16462 = w15987 ^ w16461 ;
  assign w16463 = ~w16139 & w16462 ;
  assign w16464 = ( w15899 & w16137 ) | ( w15899 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16465 = ~w16138 & w16464 ;
  assign w16466 = w16463 | w16465 ;
  assign w16467 = ~\pi075 & w16466 ;
  assign w16468 = ~w15914 & w15983 ;
  assign w16469 = w15984 ^ w16468 ;
  assign w16470 = ~w16139 & w16469 ;
  assign w16471 = ( w15906 & w16137 ) | ( w15906 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16472 = ~w16138 & w16471 ;
  assign w16473 = w16470 | w16472 ;
  assign w16474 = ~\pi074 & w16473 ;
  assign w16475 = ~w15921 & w15980 ;
  assign w16476 = w15981 ^ w16475 ;
  assign w16477 = ~w16139 & w16476 ;
  assign w16478 = ( w15913 & w16137 ) | ( w15913 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16479 = ~w16138 & w16478 ;
  assign w16480 = w16477 | w16479 ;
  assign w16481 = ~\pi073 & w16480 ;
  assign w16482 = ~w15928 & w15977 ;
  assign w16483 = w15978 ^ w16482 ;
  assign w16484 = ~w16139 & w16483 ;
  assign w16485 = ( w15920 & w16137 ) | ( w15920 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16486 = ~w16138 & w16485 ;
  assign w16487 = w16484 | w16486 ;
  assign w16488 = ~\pi072 & w16487 ;
  assign w16489 = ~w15935 & w15974 ;
  assign w16490 = w15975 ^ w16489 ;
  assign w16491 = ~w16139 & w16490 ;
  assign w16492 = ( w15927 & w16137 ) | ( w15927 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16493 = ~w16138 & w16492 ;
  assign w16494 = w16491 | w16493 ;
  assign w16495 = ~\pi071 & w16494 ;
  assign w16496 = ~w15942 & w15971 ;
  assign w16497 = w15972 ^ w16496 ;
  assign w16498 = ~w16139 & w16497 ;
  assign w16499 = ( w15934 & w16137 ) | ( w15934 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16500 = ~w16138 & w16499 ;
  assign w16501 = w16498 | w16500 ;
  assign w16502 = ~\pi070 & w16501 ;
  assign w16503 = ~w15948 & w15968 ;
  assign w16504 = w15969 ^ w16503 ;
  assign w16505 = ~w16139 & w16504 ;
  assign w16506 = ( w15941 & w16137 ) | ( w15941 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16507 = ~w16138 & w16506 ;
  assign w16508 = w16505 | w16507 ;
  assign w16509 = ~\pi069 & w16508 ;
  assign w16510 = ~w15956 & w15965 ;
  assign w16511 = w15966 ^ w16510 ;
  assign w16512 = ~w16139 & w16511 ;
  assign w16513 = ( w15947 & w16137 ) | ( w15947 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16514 = ~w16138 & w16513 ;
  assign w16515 = w16512 | w16514 ;
  assign w16516 = ~\pi068 & w16515 ;
  assign w16517 = ~\pi007 & \pi064 ;
  assign w16518 = ( \pi065 & ~w15962 ) | ( \pi065 & w16517 ) | ( ~w15962 & w16517 ) ;
  assign w16519 = w15960 ^ w16518 ;
  assign w16520 = ~w16139 & w16519 ;
  assign w16521 = ( w15955 & w16137 ) | ( w15955 & w16138 ) | ( w16137 & w16138 ) ;
  assign w16522 = ~w16138 & w16521 ;
  assign w16523 = w16520 | w16522 ;
  assign w16524 = ~\pi067 & w16523 ;
  assign w16525 = \pi008 ^ \pi065 ;
  assign w16526 = \pi007 ^ w15578 ;
  assign w16527 = ( \pi064 & w16139 ) | ( \pi064 & w16526 ) | ( w16139 & w16526 ) ;
  assign w16528 = w16525 ^ w16527 ;
  assign w16529 = ~w16139 & w16528 ;
  assign w16530 = w15962 & w16139 ;
  assign w16531 = w16529 | w16530 ;
  assign w16532 = ~\pi066 & w16531 ;
  assign w16533 = \pi066 ^ w16531 ;
  assign w16534 = \pi064 & ~w16139 ;
  assign w16535 = \pi007 ^ w16534 ;
  assign w16536 = ( ~\pi006 & \pi064 ) | ( ~\pi006 & w16533 ) | ( \pi064 & w16533 ) ;
  assign w16537 = ( \pi065 & ~w16535 ) | ( \pi065 & w16536 ) | ( ~w16535 & w16536 ) ;
  assign w16538 = w16533 | w16537 ;
  assign w16539 = \pi067 ^ w16523 ;
  assign w16540 = ( ~w16532 & w16538 ) | ( ~w16532 & w16539 ) | ( w16538 & w16539 ) ;
  assign w16541 = w16539 | w16540 ;
  assign w16542 = \pi068 ^ w16515 ;
  assign w16543 = ( ~w16524 & w16541 ) | ( ~w16524 & w16542 ) | ( w16541 & w16542 ) ;
  assign w16544 = w16542 | w16543 ;
  assign w16545 = \pi069 ^ w16508 ;
  assign w16546 = ( ~w16516 & w16544 ) | ( ~w16516 & w16545 ) | ( w16544 & w16545 ) ;
  assign w16547 = w16545 | w16546 ;
  assign w16548 = \pi070 ^ w16501 ;
  assign w16549 = ( ~w16509 & w16547 ) | ( ~w16509 & w16548 ) | ( w16547 & w16548 ) ;
  assign w16550 = w16548 | w16549 ;
  assign w16551 = \pi071 ^ w16494 ;
  assign w16552 = ( ~w16502 & w16550 ) | ( ~w16502 & w16551 ) | ( w16550 & w16551 ) ;
  assign w16553 = w16551 | w16552 ;
  assign w16554 = \pi072 ^ w16487 ;
  assign w16555 = ( ~w16495 & w16553 ) | ( ~w16495 & w16554 ) | ( w16553 & w16554 ) ;
  assign w16556 = w16554 | w16555 ;
  assign w16557 = \pi073 ^ w16480 ;
  assign w16558 = ( ~w16488 & w16556 ) | ( ~w16488 & w16557 ) | ( w16556 & w16557 ) ;
  assign w16559 = w16557 | w16558 ;
  assign w16560 = \pi074 ^ w16473 ;
  assign w16561 = ( ~w16481 & w16559 ) | ( ~w16481 & w16560 ) | ( w16559 & w16560 ) ;
  assign w16562 = w16560 | w16561 ;
  assign w16563 = \pi075 ^ w16466 ;
  assign w16564 = ( ~w16474 & w16562 ) | ( ~w16474 & w16563 ) | ( w16562 & w16563 ) ;
  assign w16565 = w16563 | w16564 ;
  assign w16566 = \pi076 ^ w16459 ;
  assign w16567 = ( ~w16467 & w16565 ) | ( ~w16467 & w16566 ) | ( w16565 & w16566 ) ;
  assign w16568 = w16566 | w16567 ;
  assign w16569 = \pi077 ^ w16452 ;
  assign w16570 = ( ~w16460 & w16568 ) | ( ~w16460 & w16569 ) | ( w16568 & w16569 ) ;
  assign w16571 = w16569 | w16570 ;
  assign w16572 = \pi078 ^ w16445 ;
  assign w16573 = ( ~w16453 & w16571 ) | ( ~w16453 & w16572 ) | ( w16571 & w16572 ) ;
  assign w16574 = w16572 | w16573 ;
  assign w16575 = \pi079 ^ w16438 ;
  assign w16576 = ( ~w16446 & w16574 ) | ( ~w16446 & w16575 ) | ( w16574 & w16575 ) ;
  assign w16577 = w16575 | w16576 ;
  assign w16578 = \pi080 ^ w16431 ;
  assign w16579 = ( ~w16439 & w16577 ) | ( ~w16439 & w16578 ) | ( w16577 & w16578 ) ;
  assign w16580 = w16578 | w16579 ;
  assign w16581 = \pi081 ^ w16424 ;
  assign w16582 = ( ~w16432 & w16580 ) | ( ~w16432 & w16581 ) | ( w16580 & w16581 ) ;
  assign w16583 = w16581 | w16582 ;
  assign w16584 = \pi082 ^ w16417 ;
  assign w16585 = ( ~w16425 & w16583 ) | ( ~w16425 & w16584 ) | ( w16583 & w16584 ) ;
  assign w16586 = w16584 | w16585 ;
  assign w16587 = \pi083 ^ w16410 ;
  assign w16588 = ( ~w16418 & w16586 ) | ( ~w16418 & w16587 ) | ( w16586 & w16587 ) ;
  assign w16589 = w16587 | w16588 ;
  assign w16590 = \pi084 ^ w16403 ;
  assign w16591 = ( ~w16411 & w16589 ) | ( ~w16411 & w16590 ) | ( w16589 & w16590 ) ;
  assign w16592 = w16590 | w16591 ;
  assign w16593 = \pi085 ^ w16396 ;
  assign w16594 = ( ~w16404 & w16592 ) | ( ~w16404 & w16593 ) | ( w16592 & w16593 ) ;
  assign w16595 = w16593 | w16594 ;
  assign w16596 = \pi086 ^ w16389 ;
  assign w16597 = ( ~w16397 & w16595 ) | ( ~w16397 & w16596 ) | ( w16595 & w16596 ) ;
  assign w16598 = w16596 | w16597 ;
  assign w16599 = \pi087 ^ w16382 ;
  assign w16600 = ( ~w16390 & w16598 ) | ( ~w16390 & w16599 ) | ( w16598 & w16599 ) ;
  assign w16601 = w16599 | w16600 ;
  assign w16602 = \pi088 ^ w16375 ;
  assign w16603 = ( ~w16383 & w16601 ) | ( ~w16383 & w16602 ) | ( w16601 & w16602 ) ;
  assign w16604 = w16602 | w16603 ;
  assign w16605 = \pi089 ^ w16368 ;
  assign w16606 = ( ~w16376 & w16604 ) | ( ~w16376 & w16605 ) | ( w16604 & w16605 ) ;
  assign w16607 = w16605 | w16606 ;
  assign w16608 = \pi090 ^ w16361 ;
  assign w16609 = ( ~w16369 & w16607 ) | ( ~w16369 & w16608 ) | ( w16607 & w16608 ) ;
  assign w16610 = w16608 | w16609 ;
  assign w16611 = \pi091 ^ w16354 ;
  assign w16612 = ( ~w16362 & w16610 ) | ( ~w16362 & w16611 ) | ( w16610 & w16611 ) ;
  assign w16613 = w16611 | w16612 ;
  assign w16614 = \pi092 ^ w16347 ;
  assign w16615 = ( ~w16355 & w16613 ) | ( ~w16355 & w16614 ) | ( w16613 & w16614 ) ;
  assign w16616 = w16614 | w16615 ;
  assign w16617 = \pi093 ^ w16340 ;
  assign w16618 = ( ~w16348 & w16616 ) | ( ~w16348 & w16617 ) | ( w16616 & w16617 ) ;
  assign w16619 = w16617 | w16618 ;
  assign w16620 = \pi094 ^ w16333 ;
  assign w16621 = ( ~w16341 & w16619 ) | ( ~w16341 & w16620 ) | ( w16619 & w16620 ) ;
  assign w16622 = w16620 | w16621 ;
  assign w16623 = \pi095 ^ w16326 ;
  assign w16624 = ( ~w16334 & w16622 ) | ( ~w16334 & w16623 ) | ( w16622 & w16623 ) ;
  assign w16625 = w16623 | w16624 ;
  assign w16626 = \pi096 ^ w16319 ;
  assign w16627 = ( ~w16327 & w16625 ) | ( ~w16327 & w16626 ) | ( w16625 & w16626 ) ;
  assign w16628 = w16626 | w16627 ;
  assign w16629 = \pi097 ^ w16312 ;
  assign w16630 = ( ~w16320 & w16628 ) | ( ~w16320 & w16629 ) | ( w16628 & w16629 ) ;
  assign w16631 = w16629 | w16630 ;
  assign w16632 = \pi098 ^ w16305 ;
  assign w16633 = ( ~w16313 & w16631 ) | ( ~w16313 & w16632 ) | ( w16631 & w16632 ) ;
  assign w16634 = w16632 | w16633 ;
  assign w16635 = \pi099 ^ w16298 ;
  assign w16636 = ( ~w16306 & w16634 ) | ( ~w16306 & w16635 ) | ( w16634 & w16635 ) ;
  assign w16637 = w16635 | w16636 ;
  assign w16638 = \pi100 ^ w16291 ;
  assign w16639 = ( ~w16299 & w16637 ) | ( ~w16299 & w16638 ) | ( w16637 & w16638 ) ;
  assign w16640 = w16638 | w16639 ;
  assign w16641 = \pi101 ^ w16284 ;
  assign w16642 = ( ~w16292 & w16640 ) | ( ~w16292 & w16641 ) | ( w16640 & w16641 ) ;
  assign w16643 = w16641 | w16642 ;
  assign w16644 = \pi102 ^ w16277 ;
  assign w16645 = ( ~w16285 & w16643 ) | ( ~w16285 & w16644 ) | ( w16643 & w16644 ) ;
  assign w16646 = w16644 | w16645 ;
  assign w16647 = \pi103 ^ w16270 ;
  assign w16648 = ( ~w16278 & w16646 ) | ( ~w16278 & w16647 ) | ( w16646 & w16647 ) ;
  assign w16649 = w16647 | w16648 ;
  assign w16650 = \pi104 ^ w16263 ;
  assign w16651 = ( ~w16271 & w16649 ) | ( ~w16271 & w16650 ) | ( w16649 & w16650 ) ;
  assign w16652 = w16650 | w16651 ;
  assign w16653 = \pi105 ^ w16256 ;
  assign w16654 = ( ~w16264 & w16652 ) | ( ~w16264 & w16653 ) | ( w16652 & w16653 ) ;
  assign w16655 = w16653 | w16654 ;
  assign w16656 = \pi106 ^ w16249 ;
  assign w16657 = ( ~w16257 & w16655 ) | ( ~w16257 & w16656 ) | ( w16655 & w16656 ) ;
  assign w16658 = w16656 | w16657 ;
  assign w16659 = \pi107 ^ w16242 ;
  assign w16660 = ( ~w16250 & w16658 ) | ( ~w16250 & w16659 ) | ( w16658 & w16659 ) ;
  assign w16661 = w16659 | w16660 ;
  assign w16662 = \pi108 ^ w16235 ;
  assign w16663 = ( ~w16243 & w16661 ) | ( ~w16243 & w16662 ) | ( w16661 & w16662 ) ;
  assign w16664 = w16662 | w16663 ;
  assign w16665 = \pi109 ^ w16228 ;
  assign w16666 = ( ~w16236 & w16664 ) | ( ~w16236 & w16665 ) | ( w16664 & w16665 ) ;
  assign w16667 = w16665 | w16666 ;
  assign w16668 = \pi110 ^ w16221 ;
  assign w16669 = ( ~w16229 & w16667 ) | ( ~w16229 & w16668 ) | ( w16667 & w16668 ) ;
  assign w16670 = w16668 | w16669 ;
  assign w16671 = \pi111 ^ w16214 ;
  assign w16672 = ( ~w16222 & w16670 ) | ( ~w16222 & w16671 ) | ( w16670 & w16671 ) ;
  assign w16673 = w16671 | w16672 ;
  assign w16674 = \pi112 ^ w16207 ;
  assign w16675 = ( ~w16215 & w16673 ) | ( ~w16215 & w16674 ) | ( w16673 & w16674 ) ;
  assign w16676 = w16674 | w16675 ;
  assign w16677 = \pi113 ^ w16200 ;
  assign w16678 = ( ~w16208 & w16676 ) | ( ~w16208 & w16677 ) | ( w16676 & w16677 ) ;
  assign w16679 = w16677 | w16678 ;
  assign w16680 = \pi114 ^ w16193 ;
  assign w16681 = ( ~w16201 & w16679 ) | ( ~w16201 & w16680 ) | ( w16679 & w16680 ) ;
  assign w16682 = w16680 | w16681 ;
  assign w16683 = \pi115 ^ w16186 ;
  assign w16684 = ( ~w16194 & w16682 ) | ( ~w16194 & w16683 ) | ( w16682 & w16683 ) ;
  assign w16685 = w16683 | w16684 ;
  assign w16686 = \pi116 ^ w16179 ;
  assign w16687 = ( ~w16187 & w16685 ) | ( ~w16187 & w16686 ) | ( w16685 & w16686 ) ;
  assign w16688 = w16686 | w16687 ;
  assign w16689 = \pi117 ^ w16172 ;
  assign w16690 = ( ~w16180 & w16688 ) | ( ~w16180 & w16689 ) | ( w16688 & w16689 ) ;
  assign w16691 = w16689 | w16690 ;
  assign w16692 = \pi118 ^ w16165 ;
  assign w16693 = ( ~w16173 & w16691 ) | ( ~w16173 & w16692 ) | ( w16691 & w16692 ) ;
  assign w16694 = w16692 | w16693 ;
  assign w16695 = \pi119 ^ w16158 ;
  assign w16696 = ( ~w16166 & w16694 ) | ( ~w16166 & w16695 ) | ( w16694 & w16695 ) ;
  assign w16697 = w16695 | w16696 ;
  assign w16698 = \pi120 ^ w16145 ;
  assign w16699 = ( ~w16159 & w16697 ) | ( ~w16159 & w16698 ) | ( w16697 & w16698 ) ;
  assign w16700 = w16698 | w16699 ;
  assign w16701 = \pi121 ^ w16151 ;
  assign w16702 = w16152 & ~w16701 ;
  assign w16703 = ( w16700 & w16701 ) | ( w16700 & ~w16702 ) | ( w16701 & ~w16702 ) ;
  assign w16704 = ~\pi121 & w16151 ;
  assign w16705 = w16703 & ~w16704 ;
  assign w16706 = ( ~\pi122 & \pi123 ) | ( ~\pi122 & w147 ) | ( \pi123 & w147 ) ;
  assign w16707 = \pi122 | w16706 ;
  assign w16708 = w16705 | w16707 ;
  assign w16709 = w16145 & w16708 ;
  assign w16710 = ~w16159 & w16697 ;
  assign w16711 = w16698 ^ w16710 ;
  assign w16712 = ~w16708 & w16711 ;
  assign w16713 = w16709 | w16712 ;
  assign w16714 = ~\pi121 & w16713 ;
  assign w16715 = w16158 & w16708 ;
  assign w16716 = ~w16166 & w16694 ;
  assign w16717 = w16695 ^ w16716 ;
  assign w16718 = ~w16708 & w16717 ;
  assign w16719 = w16715 | w16718 ;
  assign w16720 = ~\pi120 & w16719 ;
  assign w16721 = w16165 & w16708 ;
  assign w16722 = ~w16173 & w16691 ;
  assign w16723 = w16692 ^ w16722 ;
  assign w16724 = ~w16708 & w16723 ;
  assign w16725 = w16721 | w16724 ;
  assign w16726 = ~\pi119 & w16725 ;
  assign w16727 = w16172 & w16708 ;
  assign w16728 = ~w16180 & w16688 ;
  assign w16729 = w16689 ^ w16728 ;
  assign w16730 = ~w16708 & w16729 ;
  assign w16731 = w16727 | w16730 ;
  assign w16732 = ~\pi118 & w16731 ;
  assign w16733 = w16179 & w16708 ;
  assign w16734 = ~w16187 & w16685 ;
  assign w16735 = w16686 ^ w16734 ;
  assign w16736 = ~w16708 & w16735 ;
  assign w16737 = w16733 | w16736 ;
  assign w16738 = ~\pi117 & w16737 ;
  assign w16739 = w16186 & w16708 ;
  assign w16740 = ~w16194 & w16682 ;
  assign w16741 = w16683 ^ w16740 ;
  assign w16742 = ~w16708 & w16741 ;
  assign w16743 = w16739 | w16742 ;
  assign w16744 = ~\pi116 & w16743 ;
  assign w16745 = w16193 & w16708 ;
  assign w16746 = ~w16201 & w16679 ;
  assign w16747 = w16680 ^ w16746 ;
  assign w16748 = ~w16708 & w16747 ;
  assign w16749 = w16745 | w16748 ;
  assign w16750 = ~\pi115 & w16749 ;
  assign w16751 = w16200 & w16708 ;
  assign w16752 = ~w16208 & w16676 ;
  assign w16753 = w16677 ^ w16752 ;
  assign w16754 = ~w16708 & w16753 ;
  assign w16755 = w16751 | w16754 ;
  assign w16756 = ~\pi114 & w16755 ;
  assign w16757 = w16207 & w16708 ;
  assign w16758 = ~w16215 & w16673 ;
  assign w16759 = w16674 ^ w16758 ;
  assign w16760 = ~w16708 & w16759 ;
  assign w16761 = w16757 | w16760 ;
  assign w16762 = ~\pi113 & w16761 ;
  assign w16763 = w16214 & w16708 ;
  assign w16764 = ~w16222 & w16670 ;
  assign w16765 = w16671 ^ w16764 ;
  assign w16766 = ~w16708 & w16765 ;
  assign w16767 = w16763 | w16766 ;
  assign w16768 = ~\pi112 & w16767 ;
  assign w16769 = w16221 & w16708 ;
  assign w16770 = ~w16229 & w16667 ;
  assign w16771 = w16668 ^ w16770 ;
  assign w16772 = ~w16708 & w16771 ;
  assign w16773 = w16769 | w16772 ;
  assign w16774 = ~\pi111 & w16773 ;
  assign w16775 = w16228 & w16708 ;
  assign w16776 = ~w16236 & w16664 ;
  assign w16777 = w16665 ^ w16776 ;
  assign w16778 = ~w16708 & w16777 ;
  assign w16779 = w16775 | w16778 ;
  assign w16780 = ~\pi110 & w16779 ;
  assign w16781 = w16235 & w16708 ;
  assign w16782 = ~w16243 & w16661 ;
  assign w16783 = w16662 ^ w16782 ;
  assign w16784 = ~w16708 & w16783 ;
  assign w16785 = w16781 | w16784 ;
  assign w16786 = ~\pi109 & w16785 ;
  assign w16787 = w16242 & w16708 ;
  assign w16788 = ~w16250 & w16658 ;
  assign w16789 = w16659 ^ w16788 ;
  assign w16790 = ~w16708 & w16789 ;
  assign w16791 = w16787 | w16790 ;
  assign w16792 = ~\pi108 & w16791 ;
  assign w16793 = w16249 & w16708 ;
  assign w16794 = ~w16257 & w16655 ;
  assign w16795 = w16656 ^ w16794 ;
  assign w16796 = ~w16708 & w16795 ;
  assign w16797 = w16793 | w16796 ;
  assign w16798 = ~\pi107 & w16797 ;
  assign w16799 = w16256 & w16708 ;
  assign w16800 = ~w16264 & w16652 ;
  assign w16801 = w16653 ^ w16800 ;
  assign w16802 = ~w16708 & w16801 ;
  assign w16803 = w16799 | w16802 ;
  assign w16804 = ~\pi106 & w16803 ;
  assign w16805 = w16263 & w16708 ;
  assign w16806 = ~w16271 & w16649 ;
  assign w16807 = w16650 ^ w16806 ;
  assign w16808 = ~w16708 & w16807 ;
  assign w16809 = w16805 | w16808 ;
  assign w16810 = ~\pi105 & w16809 ;
  assign w16811 = w16270 & w16708 ;
  assign w16812 = ~w16278 & w16646 ;
  assign w16813 = w16647 ^ w16812 ;
  assign w16814 = ~w16708 & w16813 ;
  assign w16815 = w16811 | w16814 ;
  assign w16816 = ~\pi104 & w16815 ;
  assign w16817 = w16277 & w16708 ;
  assign w16818 = ~w16285 & w16643 ;
  assign w16819 = w16644 ^ w16818 ;
  assign w16820 = ~w16708 & w16819 ;
  assign w16821 = w16817 | w16820 ;
  assign w16822 = ~\pi103 & w16821 ;
  assign w16823 = w16284 & w16708 ;
  assign w16824 = ~w16292 & w16640 ;
  assign w16825 = w16641 ^ w16824 ;
  assign w16826 = ~w16708 & w16825 ;
  assign w16827 = w16823 | w16826 ;
  assign w16828 = ~\pi102 & w16827 ;
  assign w16829 = w16291 & w16708 ;
  assign w16830 = ~w16299 & w16637 ;
  assign w16831 = w16638 ^ w16830 ;
  assign w16832 = ~w16708 & w16831 ;
  assign w16833 = w16829 | w16832 ;
  assign w16834 = ~\pi101 & w16833 ;
  assign w16835 = w16298 & w16708 ;
  assign w16836 = ~w16306 & w16634 ;
  assign w16837 = w16635 ^ w16836 ;
  assign w16838 = ~w16708 & w16837 ;
  assign w16839 = w16835 | w16838 ;
  assign w16840 = ~\pi100 & w16839 ;
  assign w16841 = w16305 & w16708 ;
  assign w16842 = ~w16313 & w16631 ;
  assign w16843 = w16632 ^ w16842 ;
  assign w16844 = ~w16708 & w16843 ;
  assign w16845 = w16841 | w16844 ;
  assign w16846 = ~\pi099 & w16845 ;
  assign w16847 = w16312 & w16708 ;
  assign w16848 = ~w16320 & w16628 ;
  assign w16849 = w16629 ^ w16848 ;
  assign w16850 = ~w16708 & w16849 ;
  assign w16851 = w16847 | w16850 ;
  assign w16852 = ~\pi098 & w16851 ;
  assign w16853 = w16319 & w16708 ;
  assign w16854 = ~w16327 & w16625 ;
  assign w16855 = w16626 ^ w16854 ;
  assign w16856 = ~w16708 & w16855 ;
  assign w16857 = w16853 | w16856 ;
  assign w16858 = ~\pi097 & w16857 ;
  assign w16859 = w16326 & w16708 ;
  assign w16860 = ~w16334 & w16622 ;
  assign w16861 = w16623 ^ w16860 ;
  assign w16862 = ~w16708 & w16861 ;
  assign w16863 = w16859 | w16862 ;
  assign w16864 = ~\pi096 & w16863 ;
  assign w16865 = w16333 & w16708 ;
  assign w16866 = ~w16341 & w16619 ;
  assign w16867 = w16620 ^ w16866 ;
  assign w16868 = ~w16708 & w16867 ;
  assign w16869 = w16865 | w16868 ;
  assign w16870 = ~\pi095 & w16869 ;
  assign w16871 = w16340 & w16708 ;
  assign w16872 = ~w16348 & w16616 ;
  assign w16873 = w16617 ^ w16872 ;
  assign w16874 = ~w16708 & w16873 ;
  assign w16875 = w16871 | w16874 ;
  assign w16876 = ~\pi094 & w16875 ;
  assign w16877 = w16347 & w16708 ;
  assign w16878 = ~w16355 & w16613 ;
  assign w16879 = w16614 ^ w16878 ;
  assign w16880 = ~w16708 & w16879 ;
  assign w16881 = w16877 | w16880 ;
  assign w16882 = ~\pi093 & w16881 ;
  assign w16883 = w16354 & w16708 ;
  assign w16884 = ~w16362 & w16610 ;
  assign w16885 = w16611 ^ w16884 ;
  assign w16886 = ~w16708 & w16885 ;
  assign w16887 = w16883 | w16886 ;
  assign w16888 = ~\pi092 & w16887 ;
  assign w16889 = w16361 & w16708 ;
  assign w16890 = ~w16369 & w16607 ;
  assign w16891 = w16608 ^ w16890 ;
  assign w16892 = ~w16708 & w16891 ;
  assign w16893 = w16889 | w16892 ;
  assign w16894 = ~\pi091 & w16893 ;
  assign w16895 = w16368 & w16708 ;
  assign w16896 = ~w16376 & w16604 ;
  assign w16897 = w16605 ^ w16896 ;
  assign w16898 = ~w16708 & w16897 ;
  assign w16899 = w16895 | w16898 ;
  assign w16900 = ~\pi090 & w16899 ;
  assign w16901 = w16375 & w16708 ;
  assign w16902 = ~w16383 & w16601 ;
  assign w16903 = w16602 ^ w16902 ;
  assign w16904 = ~w16708 & w16903 ;
  assign w16905 = w16901 | w16904 ;
  assign w16906 = ~\pi089 & w16905 ;
  assign w16907 = w16382 & w16708 ;
  assign w16908 = ~w16390 & w16598 ;
  assign w16909 = w16599 ^ w16908 ;
  assign w16910 = ~w16708 & w16909 ;
  assign w16911 = w16907 | w16910 ;
  assign w16912 = ~\pi088 & w16911 ;
  assign w16913 = w16389 & w16708 ;
  assign w16914 = ~w16397 & w16595 ;
  assign w16915 = w16596 ^ w16914 ;
  assign w16916 = ~w16708 & w16915 ;
  assign w16917 = w16913 | w16916 ;
  assign w16918 = ~\pi087 & w16917 ;
  assign w16919 = w16396 & w16708 ;
  assign w16920 = ~w16404 & w16592 ;
  assign w16921 = w16593 ^ w16920 ;
  assign w16922 = ~w16708 & w16921 ;
  assign w16923 = w16919 | w16922 ;
  assign w16924 = ~\pi086 & w16923 ;
  assign w16925 = w16403 & w16708 ;
  assign w16926 = ~w16411 & w16589 ;
  assign w16927 = w16590 ^ w16926 ;
  assign w16928 = ~w16708 & w16927 ;
  assign w16929 = w16925 | w16928 ;
  assign w16930 = ~\pi085 & w16929 ;
  assign w16931 = w16410 & w16708 ;
  assign w16932 = ~w16418 & w16586 ;
  assign w16933 = w16587 ^ w16932 ;
  assign w16934 = ~w16708 & w16933 ;
  assign w16935 = w16931 | w16934 ;
  assign w16936 = ~\pi084 & w16935 ;
  assign w16937 = w16417 & w16708 ;
  assign w16938 = ~w16425 & w16583 ;
  assign w16939 = w16584 ^ w16938 ;
  assign w16940 = ~w16708 & w16939 ;
  assign w16941 = w16937 | w16940 ;
  assign w16942 = ~\pi083 & w16941 ;
  assign w16943 = w16424 & w16708 ;
  assign w16944 = ~w16432 & w16580 ;
  assign w16945 = w16581 ^ w16944 ;
  assign w16946 = ~w16708 & w16945 ;
  assign w16947 = w16943 | w16946 ;
  assign w16948 = ~\pi082 & w16947 ;
  assign w16949 = w16431 & w16708 ;
  assign w16950 = ~w16439 & w16577 ;
  assign w16951 = w16578 ^ w16950 ;
  assign w16952 = ~w16708 & w16951 ;
  assign w16953 = w16949 | w16952 ;
  assign w16954 = ~\pi081 & w16953 ;
  assign w16955 = w16438 & w16708 ;
  assign w16956 = ~w16446 & w16574 ;
  assign w16957 = w16575 ^ w16956 ;
  assign w16958 = ~w16708 & w16957 ;
  assign w16959 = w16955 | w16958 ;
  assign w16960 = ~\pi080 & w16959 ;
  assign w16961 = w16445 & w16708 ;
  assign w16962 = ~w16453 & w16571 ;
  assign w16963 = w16572 ^ w16962 ;
  assign w16964 = ~w16708 & w16963 ;
  assign w16965 = w16961 | w16964 ;
  assign w16966 = ~\pi079 & w16965 ;
  assign w16967 = w16452 & w16708 ;
  assign w16968 = ~w16460 & w16568 ;
  assign w16969 = w16569 ^ w16968 ;
  assign w16970 = ~w16708 & w16969 ;
  assign w16971 = w16967 | w16970 ;
  assign w16972 = ~\pi078 & w16971 ;
  assign w16973 = w16459 & w16708 ;
  assign w16974 = ~w16467 & w16565 ;
  assign w16975 = w16566 ^ w16974 ;
  assign w16976 = ~w16708 & w16975 ;
  assign w16977 = w16973 | w16976 ;
  assign w16978 = ~\pi077 & w16977 ;
  assign w16979 = w16466 & w16708 ;
  assign w16980 = ~w16474 & w16562 ;
  assign w16981 = w16563 ^ w16980 ;
  assign w16982 = ~w16708 & w16981 ;
  assign w16983 = w16979 | w16982 ;
  assign w16984 = ~\pi076 & w16983 ;
  assign w16985 = w16473 & w16708 ;
  assign w16986 = ~w16481 & w16559 ;
  assign w16987 = w16560 ^ w16986 ;
  assign w16988 = ~w16708 & w16987 ;
  assign w16989 = w16985 | w16988 ;
  assign w16990 = ~\pi075 & w16989 ;
  assign w16991 = w16480 & w16708 ;
  assign w16992 = ~w16488 & w16556 ;
  assign w16993 = w16557 ^ w16992 ;
  assign w16994 = ~w16708 & w16993 ;
  assign w16995 = w16991 | w16994 ;
  assign w16996 = ~\pi074 & w16995 ;
  assign w16997 = w16487 & w16708 ;
  assign w16998 = ~w16495 & w16553 ;
  assign w16999 = w16554 ^ w16998 ;
  assign w17000 = ~w16708 & w16999 ;
  assign w17001 = w16997 | w17000 ;
  assign w17002 = ~\pi073 & w17001 ;
  assign w17003 = w16494 & w16708 ;
  assign w17004 = ~w16502 & w16550 ;
  assign w17005 = w16551 ^ w17004 ;
  assign w17006 = ~w16708 & w17005 ;
  assign w17007 = w17003 | w17006 ;
  assign w17008 = ~\pi072 & w17007 ;
  assign w17009 = w16501 & w16708 ;
  assign w17010 = ~w16509 & w16547 ;
  assign w17011 = w16548 ^ w17010 ;
  assign w17012 = ~w16708 & w17011 ;
  assign w17013 = w17009 | w17012 ;
  assign w17014 = ~\pi071 & w17013 ;
  assign w17015 = w16508 & w16708 ;
  assign w17016 = ~w16516 & w16544 ;
  assign w17017 = w16545 ^ w17016 ;
  assign w17018 = ~w16708 & w17017 ;
  assign w17019 = w17015 | w17018 ;
  assign w17020 = ~\pi070 & w17019 ;
  assign w17021 = w16515 & w16708 ;
  assign w17022 = ~w16524 & w16541 ;
  assign w17023 = w16542 ^ w17022 ;
  assign w17024 = ~w16708 & w17023 ;
  assign w17025 = w17021 | w17024 ;
  assign w17026 = ~\pi069 & w17025 ;
  assign w17027 = w16523 & w16708 ;
  assign w17028 = ~w16532 & w16538 ;
  assign w17029 = w16539 ^ w17028 ;
  assign w17030 = ~w16708 & w17029 ;
  assign w17031 = w17027 | w17030 ;
  assign w17032 = ~\pi068 & w17031 ;
  assign w17033 = ~\pi006 & \pi064 ;
  assign w17034 = ( \pi065 & ~w16535 ) | ( \pi065 & w17033 ) | ( ~w16535 & w17033 ) ;
  assign w17035 = w16533 ^ w17034 ;
  assign w17036 = ( w16705 & w16707 ) | ( w16705 & w17035 ) | ( w16707 & w17035 ) ;
  assign w17037 = w17035 & ~w17036 ;
  assign w17038 = ( w16531 & w16708 ) | ( w16531 & w17037 ) | ( w16708 & w17037 ) ;
  assign w17039 = w17037 | w17038 ;
  assign w17040 = ~\pi067 & w17039 ;
  assign w17041 = \pi007 ^ \pi065 ;
  assign w17042 = \pi006 ^ w16139 ;
  assign w17043 = ( \pi064 & w16707 ) | ( \pi064 & w17042 ) | ( w16707 & w17042 ) ;
  assign w17044 = w17041 ^ w17043 ;
  assign w17045 = ~w16707 & w17044 ;
  assign w17046 = ~w16705 & w17045 ;
  assign w17047 = ( ~\pi064 & w16139 ) | ( ~\pi064 & w16708 ) | ( w16139 & w16708 ) ;
  assign w17048 = \pi007 ^ w17047 ;
  assign w17049 = w16708 & ~w17048 ;
  assign w17050 = w17046 | w17049 ;
  assign w17051 = ~\pi066 & w17050 ;
  assign w17052 = ( \pi064 & w269 ) | ( \pi064 & w270 ) | ( w269 & w270 ) ;
  assign w17053 = \pi006 & \pi122 ;
  assign w17054 = ( \pi006 & w17052 ) | ( \pi006 & w17053 ) | ( w17052 & w17053 ) ;
  assign w17055 = ( \pi064 & w16705 ) | ( \pi064 & w17054 ) | ( w16705 & w17054 ) ;
  assign w17056 = ( \pi006 & ~\pi064 ) | ( \pi006 & w17055 ) | ( ~\pi064 & w17055 ) ;
  assign w17057 = ( ~\pi006 & \pi064 ) | ( ~\pi006 & \pi122 ) | ( \pi064 & \pi122 ) ;
  assign w17058 = w147 | w16705 ;
  assign w17059 = ( \pi122 & \pi123 ) | ( \pi122 & ~w147 ) | ( \pi123 & ~w147 ) ;
  assign w17060 = w17058 | w17059 ;
  assign w17061 = w17057 & ~w17060 ;
  assign w17062 = ~\pi005 & \pi064 ;
  assign w17063 = w16708 | w17046 ;
  assign w17064 = ( w16535 & w17046 ) | ( w16535 & w17063 ) | ( w17046 & w17063 ) ;
  assign w17065 = \pi066 ^ w17064 ;
  assign w17066 = w17056 | w17061 ;
  assign w17067 = ( \pi065 & w17062 ) | ( \pi065 & ~w17066 ) | ( w17062 & ~w17066 ) ;
  assign w17068 = w17065 | w17067 ;
  assign w17069 = ~w16531 & w16708 ;
  assign w17070 = ( w16708 & w17037 ) | ( w16708 & ~w17069 ) | ( w17037 & ~w17069 ) ;
  assign w17071 = \pi067 ^ w17070 ;
  assign w17072 = ( ~w17051 & w17068 ) | ( ~w17051 & w17071 ) | ( w17068 & w17071 ) ;
  assign w17073 = w17071 | w17072 ;
  assign w17074 = \pi068 ^ w17031 ;
  assign w17075 = ( ~w17040 & w17073 ) | ( ~w17040 & w17074 ) | ( w17073 & w17074 ) ;
  assign w17076 = w17074 | w17075 ;
  assign w17077 = \pi069 ^ w17025 ;
  assign w17078 = ( ~w17032 & w17076 ) | ( ~w17032 & w17077 ) | ( w17076 & w17077 ) ;
  assign w17079 = w17077 | w17078 ;
  assign w17080 = \pi070 ^ w17019 ;
  assign w17081 = ( ~w17026 & w17079 ) | ( ~w17026 & w17080 ) | ( w17079 & w17080 ) ;
  assign w17082 = w17080 | w17081 ;
  assign w17083 = \pi071 ^ w17013 ;
  assign w17084 = ( ~w17020 & w17082 ) | ( ~w17020 & w17083 ) | ( w17082 & w17083 ) ;
  assign w17085 = w17083 | w17084 ;
  assign w17086 = \pi072 ^ w17007 ;
  assign w17087 = ( ~w17014 & w17085 ) | ( ~w17014 & w17086 ) | ( w17085 & w17086 ) ;
  assign w17088 = w17086 | w17087 ;
  assign w17089 = \pi073 ^ w17001 ;
  assign w17090 = ( ~w17008 & w17088 ) | ( ~w17008 & w17089 ) | ( w17088 & w17089 ) ;
  assign w17091 = w17089 | w17090 ;
  assign w17092 = \pi074 ^ w16995 ;
  assign w17093 = ( ~w17002 & w17091 ) | ( ~w17002 & w17092 ) | ( w17091 & w17092 ) ;
  assign w17094 = w17092 | w17093 ;
  assign w17095 = \pi075 ^ w16989 ;
  assign w17096 = ( ~w16996 & w17094 ) | ( ~w16996 & w17095 ) | ( w17094 & w17095 ) ;
  assign w17097 = w17095 | w17096 ;
  assign w17098 = \pi076 ^ w16983 ;
  assign w17099 = ( ~w16990 & w17097 ) | ( ~w16990 & w17098 ) | ( w17097 & w17098 ) ;
  assign w17100 = w17098 | w17099 ;
  assign w17101 = \pi077 ^ w16977 ;
  assign w17102 = ( ~w16984 & w17100 ) | ( ~w16984 & w17101 ) | ( w17100 & w17101 ) ;
  assign w17103 = w17101 | w17102 ;
  assign w17104 = \pi078 ^ w16971 ;
  assign w17105 = ( ~w16978 & w17103 ) | ( ~w16978 & w17104 ) | ( w17103 & w17104 ) ;
  assign w17106 = w17104 | w17105 ;
  assign w17107 = \pi079 ^ w16965 ;
  assign w17108 = ( ~w16972 & w17106 ) | ( ~w16972 & w17107 ) | ( w17106 & w17107 ) ;
  assign w17109 = w17107 | w17108 ;
  assign w17110 = \pi080 ^ w16959 ;
  assign w17111 = ( ~w16966 & w17109 ) | ( ~w16966 & w17110 ) | ( w17109 & w17110 ) ;
  assign w17112 = w17110 | w17111 ;
  assign w17113 = \pi081 ^ w16953 ;
  assign w17114 = ( ~w16960 & w17112 ) | ( ~w16960 & w17113 ) | ( w17112 & w17113 ) ;
  assign w17115 = w17113 | w17114 ;
  assign w17116 = \pi082 ^ w16947 ;
  assign w17117 = ( ~w16954 & w17115 ) | ( ~w16954 & w17116 ) | ( w17115 & w17116 ) ;
  assign w17118 = w17116 | w17117 ;
  assign w17119 = \pi083 ^ w16941 ;
  assign w17120 = ( ~w16948 & w17118 ) | ( ~w16948 & w17119 ) | ( w17118 & w17119 ) ;
  assign w17121 = w17119 | w17120 ;
  assign w17122 = \pi084 ^ w16935 ;
  assign w17123 = ( ~w16942 & w17121 ) | ( ~w16942 & w17122 ) | ( w17121 & w17122 ) ;
  assign w17124 = w17122 | w17123 ;
  assign w17125 = \pi085 ^ w16929 ;
  assign w17126 = ( ~w16936 & w17124 ) | ( ~w16936 & w17125 ) | ( w17124 & w17125 ) ;
  assign w17127 = w17125 | w17126 ;
  assign w17128 = \pi086 ^ w16923 ;
  assign w17129 = ( ~w16930 & w17127 ) | ( ~w16930 & w17128 ) | ( w17127 & w17128 ) ;
  assign w17130 = w17128 | w17129 ;
  assign w17131 = \pi087 ^ w16917 ;
  assign w17132 = ( ~w16924 & w17130 ) | ( ~w16924 & w17131 ) | ( w17130 & w17131 ) ;
  assign w17133 = w17131 | w17132 ;
  assign w17134 = \pi088 ^ w16911 ;
  assign w17135 = ( ~w16918 & w17133 ) | ( ~w16918 & w17134 ) | ( w17133 & w17134 ) ;
  assign w17136 = w17134 | w17135 ;
  assign w17137 = \pi089 ^ w16905 ;
  assign w17138 = ( ~w16912 & w17136 ) | ( ~w16912 & w17137 ) | ( w17136 & w17137 ) ;
  assign w17139 = w17137 | w17138 ;
  assign w17140 = \pi090 ^ w16899 ;
  assign w17141 = ( ~w16906 & w17139 ) | ( ~w16906 & w17140 ) | ( w17139 & w17140 ) ;
  assign w17142 = w17140 | w17141 ;
  assign w17143 = \pi091 ^ w16893 ;
  assign w17144 = ( ~w16900 & w17142 ) | ( ~w16900 & w17143 ) | ( w17142 & w17143 ) ;
  assign w17145 = w17143 | w17144 ;
  assign w17146 = \pi092 ^ w16887 ;
  assign w17147 = ( ~w16894 & w17145 ) | ( ~w16894 & w17146 ) | ( w17145 & w17146 ) ;
  assign w17148 = w17146 | w17147 ;
  assign w17149 = \pi093 ^ w16881 ;
  assign w17150 = ( ~w16888 & w17148 ) | ( ~w16888 & w17149 ) | ( w17148 & w17149 ) ;
  assign w17151 = w17149 | w17150 ;
  assign w17152 = \pi094 ^ w16875 ;
  assign w17153 = ( ~w16882 & w17151 ) | ( ~w16882 & w17152 ) | ( w17151 & w17152 ) ;
  assign w17154 = w17152 | w17153 ;
  assign w17155 = \pi095 ^ w16869 ;
  assign w17156 = ( ~w16876 & w17154 ) | ( ~w16876 & w17155 ) | ( w17154 & w17155 ) ;
  assign w17157 = w17155 | w17156 ;
  assign w17158 = \pi096 ^ w16863 ;
  assign w17159 = ( ~w16870 & w17157 ) | ( ~w16870 & w17158 ) | ( w17157 & w17158 ) ;
  assign w17160 = w17158 | w17159 ;
  assign w17161 = \pi097 ^ w16857 ;
  assign w17162 = ( ~w16864 & w17160 ) | ( ~w16864 & w17161 ) | ( w17160 & w17161 ) ;
  assign w17163 = w17161 | w17162 ;
  assign w17164 = \pi098 ^ w16851 ;
  assign w17165 = ( ~w16858 & w17163 ) | ( ~w16858 & w17164 ) | ( w17163 & w17164 ) ;
  assign w17166 = w17164 | w17165 ;
  assign w17167 = \pi099 ^ w16845 ;
  assign w17168 = ( ~w16852 & w17166 ) | ( ~w16852 & w17167 ) | ( w17166 & w17167 ) ;
  assign w17169 = w17167 | w17168 ;
  assign w17170 = \pi100 ^ w16839 ;
  assign w17171 = ( ~w16846 & w17169 ) | ( ~w16846 & w17170 ) | ( w17169 & w17170 ) ;
  assign w17172 = w17170 | w17171 ;
  assign w17173 = \pi101 ^ w16833 ;
  assign w17174 = ( ~w16840 & w17172 ) | ( ~w16840 & w17173 ) | ( w17172 & w17173 ) ;
  assign w17175 = w17173 | w17174 ;
  assign w17176 = \pi102 ^ w16827 ;
  assign w17177 = ( ~w16834 & w17175 ) | ( ~w16834 & w17176 ) | ( w17175 & w17176 ) ;
  assign w17178 = w17176 | w17177 ;
  assign w17179 = \pi103 ^ w16821 ;
  assign w17180 = ( ~w16828 & w17178 ) | ( ~w16828 & w17179 ) | ( w17178 & w17179 ) ;
  assign w17181 = w17179 | w17180 ;
  assign w17182 = \pi104 ^ w16815 ;
  assign w17183 = ( ~w16822 & w17181 ) | ( ~w16822 & w17182 ) | ( w17181 & w17182 ) ;
  assign w17184 = w17182 | w17183 ;
  assign w17185 = \pi105 ^ w16809 ;
  assign w17186 = ( ~w16816 & w17184 ) | ( ~w16816 & w17185 ) | ( w17184 & w17185 ) ;
  assign w17187 = w17185 | w17186 ;
  assign w17188 = \pi106 ^ w16803 ;
  assign w17189 = ( ~w16810 & w17187 ) | ( ~w16810 & w17188 ) | ( w17187 & w17188 ) ;
  assign w17190 = w17188 | w17189 ;
  assign w17191 = \pi107 ^ w16797 ;
  assign w17192 = ( ~w16804 & w17190 ) | ( ~w16804 & w17191 ) | ( w17190 & w17191 ) ;
  assign w17193 = w17191 | w17192 ;
  assign w17194 = \pi108 ^ w16791 ;
  assign w17195 = ( ~w16798 & w17193 ) | ( ~w16798 & w17194 ) | ( w17193 & w17194 ) ;
  assign w17196 = w17194 | w17195 ;
  assign w17197 = \pi109 ^ w16785 ;
  assign w17198 = ( ~w16792 & w17196 ) | ( ~w16792 & w17197 ) | ( w17196 & w17197 ) ;
  assign w17199 = w17197 | w17198 ;
  assign w17200 = \pi110 ^ w16779 ;
  assign w17201 = ( ~w16786 & w17199 ) | ( ~w16786 & w17200 ) | ( w17199 & w17200 ) ;
  assign w17202 = w17200 | w17201 ;
  assign w17203 = \pi111 ^ w16773 ;
  assign w17204 = ( ~w16780 & w17202 ) | ( ~w16780 & w17203 ) | ( w17202 & w17203 ) ;
  assign w17205 = w17203 | w17204 ;
  assign w17206 = \pi112 ^ w16767 ;
  assign w17207 = ( ~w16774 & w17205 ) | ( ~w16774 & w17206 ) | ( w17205 & w17206 ) ;
  assign w17208 = w17206 | w17207 ;
  assign w17209 = \pi113 ^ w16761 ;
  assign w17210 = ( ~w16768 & w17208 ) | ( ~w16768 & w17209 ) | ( w17208 & w17209 ) ;
  assign w17211 = w17209 | w17210 ;
  assign w17212 = \pi114 ^ w16755 ;
  assign w17213 = ( ~w16762 & w17211 ) | ( ~w16762 & w17212 ) | ( w17211 & w17212 ) ;
  assign w17214 = w17212 | w17213 ;
  assign w17215 = \pi115 ^ w16749 ;
  assign w17216 = ( ~w16756 & w17214 ) | ( ~w16756 & w17215 ) | ( w17214 & w17215 ) ;
  assign w17217 = w17215 | w17216 ;
  assign w17218 = \pi116 ^ w16743 ;
  assign w17219 = ( ~w16750 & w17217 ) | ( ~w16750 & w17218 ) | ( w17217 & w17218 ) ;
  assign w17220 = w17218 | w17219 ;
  assign w17221 = \pi117 ^ w16737 ;
  assign w17222 = ( ~w16744 & w17220 ) | ( ~w16744 & w17221 ) | ( w17220 & w17221 ) ;
  assign w17223 = w17221 | w17222 ;
  assign w17224 = \pi118 ^ w16731 ;
  assign w17225 = ( ~w16738 & w17223 ) | ( ~w16738 & w17224 ) | ( w17223 & w17224 ) ;
  assign w17226 = w17224 | w17225 ;
  assign w17227 = \pi119 ^ w16725 ;
  assign w17228 = ( ~w16732 & w17226 ) | ( ~w16732 & w17227 ) | ( w17226 & w17227 ) ;
  assign w17229 = w17227 | w17228 ;
  assign w17230 = \pi120 ^ w16719 ;
  assign w17231 = ( ~w16726 & w17229 ) | ( ~w16726 & w17230 ) | ( w17229 & w17230 ) ;
  assign w17232 = w17230 | w17231 ;
  assign w17233 = \pi121 ^ w16713 ;
  assign w17234 = ( ~w16720 & w17232 ) | ( ~w16720 & w17233 ) | ( w17232 & w17233 ) ;
  assign w17235 = w17233 | w17234 ;
  assign w17236 = w16151 & w16708 ;
  assign w17237 = ~w16152 & w16700 ;
  assign w17238 = w16701 ^ w17237 ;
  assign w17239 = ~w16708 & w17238 ;
  assign w17240 = w17236 | w17239 ;
  assign w17241 = ~\pi122 & w17240 ;
  assign w17242 = ( \pi122 & ~w17236 ) | ( \pi122 & w17239 ) | ( ~w17236 & w17239 ) ;
  assign w17243 = ~w17239 & w17242 ;
  assign w17244 = ( ~w16714 & w17235 ) | ( ~w16714 & w17241 ) | ( w17235 & w17241 ) ;
  assign w17245 = ( w270 & w17241 ) | ( w270 & ~w17244 ) | ( w17241 & ~w17244 ) ;
  assign w17246 = ( w269 & w17243 ) | ( w269 & ~w17244 ) | ( w17243 & ~w17244 ) ;
  assign w17247 = ( w17244 & ~w17245 ) | ( w17244 & w17246 ) | ( ~w17245 & w17246 ) ;
  assign w17248 = w17245 | w17247 ;
  assign w17249 = ~w16707 & w17240 ;
  assign w17250 = w17248 & ~w17249 ;
  assign w17251 = ~w16720 & w17232 ;
  assign w17252 = w17233 ^ w17251 ;
  assign w17253 = ~w17250 & w17252 ;
  assign w17254 = ( w16713 & w17248 ) | ( w16713 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17255 = ~w17249 & w17254 ;
  assign w17256 = w17253 | w17255 ;
  assign w17257 = ~\pi122 & w17256 ;
  assign w17258 = ~w16726 & w17229 ;
  assign w17259 = w17230 ^ w17258 ;
  assign w17260 = ~w17250 & w17259 ;
  assign w17261 = ( w16719 & w17248 ) | ( w16719 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17262 = ~w17249 & w17261 ;
  assign w17263 = w17260 | w17262 ;
  assign w17264 = ~\pi121 & w17263 ;
  assign w17265 = ~w16732 & w17226 ;
  assign w17266 = w17227 ^ w17265 ;
  assign w17267 = ~w17250 & w17266 ;
  assign w17268 = ( w16725 & w17248 ) | ( w16725 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17269 = ~w17249 & w17268 ;
  assign w17270 = w17267 | w17269 ;
  assign w17271 = ~\pi120 & w17270 ;
  assign w17272 = ~w16738 & w17223 ;
  assign w17273 = w17224 ^ w17272 ;
  assign w17274 = ~w17250 & w17273 ;
  assign w17275 = ( w16731 & w17248 ) | ( w16731 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17276 = ~w17249 & w17275 ;
  assign w17277 = w17274 | w17276 ;
  assign w17278 = ~\pi119 & w17277 ;
  assign w17279 = ~w16744 & w17220 ;
  assign w17280 = w17221 ^ w17279 ;
  assign w17281 = ~w17250 & w17280 ;
  assign w17282 = ( w16737 & w17248 ) | ( w16737 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17283 = ~w17249 & w17282 ;
  assign w17284 = w17281 | w17283 ;
  assign w17285 = ~\pi118 & w17284 ;
  assign w17286 = ~w16750 & w17217 ;
  assign w17287 = w17218 ^ w17286 ;
  assign w17288 = ~w17250 & w17287 ;
  assign w17289 = ( w16743 & w17248 ) | ( w16743 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17290 = ~w17249 & w17289 ;
  assign w17291 = w17288 | w17290 ;
  assign w17292 = ~\pi117 & w17291 ;
  assign w17293 = ~w16756 & w17214 ;
  assign w17294 = w17215 ^ w17293 ;
  assign w17295 = ~w17250 & w17294 ;
  assign w17296 = ( w16749 & w17248 ) | ( w16749 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17297 = ~w17249 & w17296 ;
  assign w17298 = w17295 | w17297 ;
  assign w17299 = ~\pi116 & w17298 ;
  assign w17300 = ~w16762 & w17211 ;
  assign w17301 = w17212 ^ w17300 ;
  assign w17302 = ~w17250 & w17301 ;
  assign w17303 = ( w16755 & w17248 ) | ( w16755 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17304 = ~w17249 & w17303 ;
  assign w17305 = w17302 | w17304 ;
  assign w17306 = ~\pi115 & w17305 ;
  assign w17307 = ~w16768 & w17208 ;
  assign w17308 = w17209 ^ w17307 ;
  assign w17309 = ~w17250 & w17308 ;
  assign w17310 = ( w16761 & w17248 ) | ( w16761 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17311 = ~w17249 & w17310 ;
  assign w17312 = w17309 | w17311 ;
  assign w17313 = ~\pi114 & w17312 ;
  assign w17314 = ~w16774 & w17205 ;
  assign w17315 = w17206 ^ w17314 ;
  assign w17316 = ~w17250 & w17315 ;
  assign w17317 = ( w16767 & w17248 ) | ( w16767 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17318 = ~w17249 & w17317 ;
  assign w17319 = w17316 | w17318 ;
  assign w17320 = ~\pi113 & w17319 ;
  assign w17321 = ~w16780 & w17202 ;
  assign w17322 = w17203 ^ w17321 ;
  assign w17323 = ~w17250 & w17322 ;
  assign w17324 = ( w16773 & w17248 ) | ( w16773 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17325 = ~w17249 & w17324 ;
  assign w17326 = w17323 | w17325 ;
  assign w17327 = ~\pi112 & w17326 ;
  assign w17328 = ~w16786 & w17199 ;
  assign w17329 = w17200 ^ w17328 ;
  assign w17330 = ~w17250 & w17329 ;
  assign w17331 = ( w16779 & w17248 ) | ( w16779 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17332 = ~w17249 & w17331 ;
  assign w17333 = w17330 | w17332 ;
  assign w17334 = ~\pi111 & w17333 ;
  assign w17335 = ~w16792 & w17196 ;
  assign w17336 = w17197 ^ w17335 ;
  assign w17337 = ~w17250 & w17336 ;
  assign w17338 = ( w16785 & w17248 ) | ( w16785 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17339 = ~w17249 & w17338 ;
  assign w17340 = w17337 | w17339 ;
  assign w17341 = ~\pi110 & w17340 ;
  assign w17342 = ~w16798 & w17193 ;
  assign w17343 = w17194 ^ w17342 ;
  assign w17344 = ~w17250 & w17343 ;
  assign w17345 = ( w16791 & w17248 ) | ( w16791 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17346 = ~w17249 & w17345 ;
  assign w17347 = w17344 | w17346 ;
  assign w17348 = ~\pi109 & w17347 ;
  assign w17349 = ~w16804 & w17190 ;
  assign w17350 = w17191 ^ w17349 ;
  assign w17351 = ~w17250 & w17350 ;
  assign w17352 = ( w16797 & w17248 ) | ( w16797 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17353 = ~w17249 & w17352 ;
  assign w17354 = w17351 | w17353 ;
  assign w17355 = ~\pi108 & w17354 ;
  assign w17356 = ~w16810 & w17187 ;
  assign w17357 = w17188 ^ w17356 ;
  assign w17358 = ~w17250 & w17357 ;
  assign w17359 = ( w16803 & w17248 ) | ( w16803 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17360 = ~w17249 & w17359 ;
  assign w17361 = w17358 | w17360 ;
  assign w17362 = ~\pi107 & w17361 ;
  assign w17363 = ~w16816 & w17184 ;
  assign w17364 = w17185 ^ w17363 ;
  assign w17365 = ~w17250 & w17364 ;
  assign w17366 = ( w16809 & w17248 ) | ( w16809 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17367 = ~w17249 & w17366 ;
  assign w17368 = w17365 | w17367 ;
  assign w17369 = ~\pi106 & w17368 ;
  assign w17370 = ~w16822 & w17181 ;
  assign w17371 = w17182 ^ w17370 ;
  assign w17372 = ~w17250 & w17371 ;
  assign w17373 = ( w16815 & w17248 ) | ( w16815 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17374 = ~w17249 & w17373 ;
  assign w17375 = w17372 | w17374 ;
  assign w17376 = ~\pi105 & w17375 ;
  assign w17377 = ~w16828 & w17178 ;
  assign w17378 = w17179 ^ w17377 ;
  assign w17379 = ~w17250 & w17378 ;
  assign w17380 = ( w16821 & w17248 ) | ( w16821 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17381 = ~w17249 & w17380 ;
  assign w17382 = w17379 | w17381 ;
  assign w17383 = ~\pi104 & w17382 ;
  assign w17384 = ~w16834 & w17175 ;
  assign w17385 = w17176 ^ w17384 ;
  assign w17386 = ~w17250 & w17385 ;
  assign w17387 = ( w16827 & w17248 ) | ( w16827 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17388 = ~w17249 & w17387 ;
  assign w17389 = w17386 | w17388 ;
  assign w17390 = ~\pi103 & w17389 ;
  assign w17391 = ~w16840 & w17172 ;
  assign w17392 = w17173 ^ w17391 ;
  assign w17393 = ~w17250 & w17392 ;
  assign w17394 = ( w16833 & w17248 ) | ( w16833 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17395 = ~w17249 & w17394 ;
  assign w17396 = w17393 | w17395 ;
  assign w17397 = ~\pi102 & w17396 ;
  assign w17398 = ~w16846 & w17169 ;
  assign w17399 = w17170 ^ w17398 ;
  assign w17400 = ~w17250 & w17399 ;
  assign w17401 = ( w16839 & w17248 ) | ( w16839 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17402 = ~w17249 & w17401 ;
  assign w17403 = w17400 | w17402 ;
  assign w17404 = ~\pi101 & w17403 ;
  assign w17405 = ~w16852 & w17166 ;
  assign w17406 = w17167 ^ w17405 ;
  assign w17407 = ~w17250 & w17406 ;
  assign w17408 = ( w16845 & w17248 ) | ( w16845 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17409 = ~w17249 & w17408 ;
  assign w17410 = w17407 | w17409 ;
  assign w17411 = ~\pi100 & w17410 ;
  assign w17412 = ~w16858 & w17163 ;
  assign w17413 = w17164 ^ w17412 ;
  assign w17414 = ~w17250 & w17413 ;
  assign w17415 = ( w16851 & w17248 ) | ( w16851 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17416 = ~w17249 & w17415 ;
  assign w17417 = w17414 | w17416 ;
  assign w17418 = ~\pi099 & w17417 ;
  assign w17419 = ~w16864 & w17160 ;
  assign w17420 = w17161 ^ w17419 ;
  assign w17421 = ~w17250 & w17420 ;
  assign w17422 = ( w16857 & w17248 ) | ( w16857 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17423 = ~w17249 & w17422 ;
  assign w17424 = w17421 | w17423 ;
  assign w17425 = ~\pi098 & w17424 ;
  assign w17426 = ~w16870 & w17157 ;
  assign w17427 = w17158 ^ w17426 ;
  assign w17428 = ~w17250 & w17427 ;
  assign w17429 = ( w16863 & w17248 ) | ( w16863 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17430 = ~w17249 & w17429 ;
  assign w17431 = w17428 | w17430 ;
  assign w17432 = ~\pi097 & w17431 ;
  assign w17433 = ~w16876 & w17154 ;
  assign w17434 = w17155 ^ w17433 ;
  assign w17435 = ~w17250 & w17434 ;
  assign w17436 = ( w16869 & w17248 ) | ( w16869 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17437 = ~w17249 & w17436 ;
  assign w17438 = w17435 | w17437 ;
  assign w17439 = ~\pi096 & w17438 ;
  assign w17440 = ~w16882 & w17151 ;
  assign w17441 = w17152 ^ w17440 ;
  assign w17442 = ~w17250 & w17441 ;
  assign w17443 = ( w16875 & w17248 ) | ( w16875 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17444 = ~w17249 & w17443 ;
  assign w17445 = w17442 | w17444 ;
  assign w17446 = ~\pi095 & w17445 ;
  assign w17447 = ~w16888 & w17148 ;
  assign w17448 = w17149 ^ w17447 ;
  assign w17449 = ~w17250 & w17448 ;
  assign w17450 = ( w16881 & w17248 ) | ( w16881 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17451 = ~w17249 & w17450 ;
  assign w17452 = w17449 | w17451 ;
  assign w17453 = ~\pi094 & w17452 ;
  assign w17454 = ~w16894 & w17145 ;
  assign w17455 = w17146 ^ w17454 ;
  assign w17456 = ~w17250 & w17455 ;
  assign w17457 = ( w16887 & w17248 ) | ( w16887 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17458 = ~w17249 & w17457 ;
  assign w17459 = w17456 | w17458 ;
  assign w17460 = ~\pi093 & w17459 ;
  assign w17461 = ~w16900 & w17142 ;
  assign w17462 = w17143 ^ w17461 ;
  assign w17463 = ~w17250 & w17462 ;
  assign w17464 = ( w16893 & w17248 ) | ( w16893 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17465 = ~w17249 & w17464 ;
  assign w17466 = w17463 | w17465 ;
  assign w17467 = ~\pi092 & w17466 ;
  assign w17468 = ~w16906 & w17139 ;
  assign w17469 = w17140 ^ w17468 ;
  assign w17470 = ~w17250 & w17469 ;
  assign w17471 = ( w16899 & w17248 ) | ( w16899 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17472 = ~w17249 & w17471 ;
  assign w17473 = w17470 | w17472 ;
  assign w17474 = ~\pi091 & w17473 ;
  assign w17475 = ~w16912 & w17136 ;
  assign w17476 = w17137 ^ w17475 ;
  assign w17477 = ~w17250 & w17476 ;
  assign w17478 = ( w16905 & w17248 ) | ( w16905 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17479 = ~w17249 & w17478 ;
  assign w17480 = w17477 | w17479 ;
  assign w17481 = ~\pi090 & w17480 ;
  assign w17482 = ~w16918 & w17133 ;
  assign w17483 = w17134 ^ w17482 ;
  assign w17484 = ~w17250 & w17483 ;
  assign w17485 = ( w16911 & w17248 ) | ( w16911 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17486 = ~w17249 & w17485 ;
  assign w17487 = w17484 | w17486 ;
  assign w17488 = ~\pi089 & w17487 ;
  assign w17489 = ~w16924 & w17130 ;
  assign w17490 = w17131 ^ w17489 ;
  assign w17491 = ~w17250 & w17490 ;
  assign w17492 = ( w16917 & w17248 ) | ( w16917 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17493 = ~w17249 & w17492 ;
  assign w17494 = w17491 | w17493 ;
  assign w17495 = ~\pi088 & w17494 ;
  assign w17496 = ~w16930 & w17127 ;
  assign w17497 = w17128 ^ w17496 ;
  assign w17498 = ~w17250 & w17497 ;
  assign w17499 = ( w16923 & w17248 ) | ( w16923 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17500 = ~w17249 & w17499 ;
  assign w17501 = w17498 | w17500 ;
  assign w17502 = ~\pi087 & w17501 ;
  assign w17503 = ~w16936 & w17124 ;
  assign w17504 = w17125 ^ w17503 ;
  assign w17505 = ~w17250 & w17504 ;
  assign w17506 = ( w16929 & w17248 ) | ( w16929 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17507 = ~w17249 & w17506 ;
  assign w17508 = w17505 | w17507 ;
  assign w17509 = ~\pi086 & w17508 ;
  assign w17510 = ~w16942 & w17121 ;
  assign w17511 = w17122 ^ w17510 ;
  assign w17512 = ~w17250 & w17511 ;
  assign w17513 = ( w16935 & w17248 ) | ( w16935 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17514 = ~w17249 & w17513 ;
  assign w17515 = w17512 | w17514 ;
  assign w17516 = ~\pi085 & w17515 ;
  assign w17517 = ~w16948 & w17118 ;
  assign w17518 = w17119 ^ w17517 ;
  assign w17519 = ~w17250 & w17518 ;
  assign w17520 = ( w16941 & w17248 ) | ( w16941 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17521 = ~w17249 & w17520 ;
  assign w17522 = w17519 | w17521 ;
  assign w17523 = ~\pi084 & w17522 ;
  assign w17524 = ~w16954 & w17115 ;
  assign w17525 = w17116 ^ w17524 ;
  assign w17526 = ~w17250 & w17525 ;
  assign w17527 = ( w16947 & w17248 ) | ( w16947 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17528 = ~w17249 & w17527 ;
  assign w17529 = w17526 | w17528 ;
  assign w17530 = ~\pi083 & w17529 ;
  assign w17531 = ~w16960 & w17112 ;
  assign w17532 = w17113 ^ w17531 ;
  assign w17533 = ~w17250 & w17532 ;
  assign w17534 = ( w16953 & w17248 ) | ( w16953 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17535 = ~w17249 & w17534 ;
  assign w17536 = w17533 | w17535 ;
  assign w17537 = ~\pi082 & w17536 ;
  assign w17538 = ~w16966 & w17109 ;
  assign w17539 = w17110 ^ w17538 ;
  assign w17540 = ~w17250 & w17539 ;
  assign w17541 = ( w16959 & w17248 ) | ( w16959 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17542 = ~w17249 & w17541 ;
  assign w17543 = w17540 | w17542 ;
  assign w17544 = ~\pi081 & w17543 ;
  assign w17545 = ~w16972 & w17106 ;
  assign w17546 = w17107 ^ w17545 ;
  assign w17547 = ~w17250 & w17546 ;
  assign w17548 = ( w16965 & w17248 ) | ( w16965 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17549 = ~w17249 & w17548 ;
  assign w17550 = w17547 | w17549 ;
  assign w17551 = ~\pi080 & w17550 ;
  assign w17552 = ~w16978 & w17103 ;
  assign w17553 = w17104 ^ w17552 ;
  assign w17554 = ~w17250 & w17553 ;
  assign w17555 = ( w16971 & w17248 ) | ( w16971 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17556 = ~w17249 & w17555 ;
  assign w17557 = w17554 | w17556 ;
  assign w17558 = ~\pi079 & w17557 ;
  assign w17559 = ~w16984 & w17100 ;
  assign w17560 = w17101 ^ w17559 ;
  assign w17561 = ~w17250 & w17560 ;
  assign w17562 = ( w16977 & w17248 ) | ( w16977 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17563 = ~w17249 & w17562 ;
  assign w17564 = w17561 | w17563 ;
  assign w17565 = ~\pi078 & w17564 ;
  assign w17566 = ~w16990 & w17097 ;
  assign w17567 = w17098 ^ w17566 ;
  assign w17568 = ~w17250 & w17567 ;
  assign w17569 = ( w16983 & w17248 ) | ( w16983 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17570 = ~w17249 & w17569 ;
  assign w17571 = w17568 | w17570 ;
  assign w17572 = ~\pi077 & w17571 ;
  assign w17573 = ~w16996 & w17094 ;
  assign w17574 = w17095 ^ w17573 ;
  assign w17575 = ~w17250 & w17574 ;
  assign w17576 = ( w16989 & w17248 ) | ( w16989 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17577 = ~w17249 & w17576 ;
  assign w17578 = w17575 | w17577 ;
  assign w17579 = ~\pi076 & w17578 ;
  assign w17580 = ~w17002 & w17091 ;
  assign w17581 = w17092 ^ w17580 ;
  assign w17582 = ~w17250 & w17581 ;
  assign w17583 = ( w16995 & w17248 ) | ( w16995 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17584 = ~w17249 & w17583 ;
  assign w17585 = w17582 | w17584 ;
  assign w17586 = ~\pi075 & w17585 ;
  assign w17587 = ~w17008 & w17088 ;
  assign w17588 = w17089 ^ w17587 ;
  assign w17589 = ~w17250 & w17588 ;
  assign w17590 = ( w17001 & w17248 ) | ( w17001 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17591 = ~w17249 & w17590 ;
  assign w17592 = w17589 | w17591 ;
  assign w17593 = ~\pi074 & w17592 ;
  assign w17594 = ~w17014 & w17085 ;
  assign w17595 = w17086 ^ w17594 ;
  assign w17596 = ~w17250 & w17595 ;
  assign w17597 = ( w17007 & w17248 ) | ( w17007 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17598 = ~w17249 & w17597 ;
  assign w17599 = w17596 | w17598 ;
  assign w17600 = ~\pi073 & w17599 ;
  assign w17601 = ~w17020 & w17082 ;
  assign w17602 = w17083 ^ w17601 ;
  assign w17603 = ~w17250 & w17602 ;
  assign w17604 = ( w17013 & w17248 ) | ( w17013 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17605 = ~w17249 & w17604 ;
  assign w17606 = w17603 | w17605 ;
  assign w17607 = ~\pi072 & w17606 ;
  assign w17608 = ~w17026 & w17079 ;
  assign w17609 = w17080 ^ w17608 ;
  assign w17610 = ~w17250 & w17609 ;
  assign w17611 = ( w17019 & w17248 ) | ( w17019 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17612 = ~w17249 & w17611 ;
  assign w17613 = w17610 | w17612 ;
  assign w17614 = ~\pi071 & w17613 ;
  assign w17615 = ~w17032 & w17076 ;
  assign w17616 = w17077 ^ w17615 ;
  assign w17617 = ~w17250 & w17616 ;
  assign w17618 = ( w17025 & w17248 ) | ( w17025 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17619 = ~w17249 & w17618 ;
  assign w17620 = w17617 | w17619 ;
  assign w17621 = ~\pi070 & w17620 ;
  assign w17622 = ~w17040 & w17073 ;
  assign w17623 = w17074 ^ w17622 ;
  assign w17624 = ~w17250 & w17623 ;
  assign w17625 = ( w17031 & w17248 ) | ( w17031 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17626 = ~w17249 & w17625 ;
  assign w17627 = w17624 | w17626 ;
  assign w17628 = ~\pi069 & w17627 ;
  assign w17629 = ~w17051 & w17068 ;
  assign w17630 = w17071 ^ w17629 ;
  assign w17631 = ~w17250 & w17630 ;
  assign w17632 = ( w17039 & w17248 ) | ( w17039 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17633 = ~w17249 & w17632 ;
  assign w17634 = w17631 | w17633 ;
  assign w17635 = ~\pi068 & w17634 ;
  assign w17636 = w17065 ^ w17067 ;
  assign w17637 = ~w17250 & w17636 ;
  assign w17638 = ( w17050 & w17248 ) | ( w17050 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17639 = ~w17249 & w17638 ;
  assign w17640 = w17637 | w17639 ;
  assign w17641 = ~\pi067 & w17640 ;
  assign w17642 = w17062 ^ w17066 ;
  assign w17643 = \pi065 ^ w17642 ;
  assign w17644 = ~w17250 & w17643 ;
  assign w17645 = ( w17056 & w17061 ) | ( w17056 & ~w17249 ) | ( w17061 & ~w17249 ) ;
  assign w17646 = w17249 & w17645 ;
  assign w17647 = ( ~w17248 & w17645 ) | ( ~w17248 & w17646 ) | ( w17645 & w17646 ) ;
  assign w17648 = ( w17644 & w17645 ) | ( w17644 & ~w17647 ) | ( w17645 & ~w17647 ) ;
  assign w17649 = ~\pi066 & w17648 ;
  assign w17650 = w17248 | w17249 ;
  assign w17651 = ( w17644 & w17645 ) | ( w17644 & w17650 ) | ( w17645 & w17650 ) ;
  assign w17652 = ( ~w17249 & w17644 ) | ( ~w17249 & w17651 ) | ( w17644 & w17651 ) ;
  assign w17653 = \pi066 ^ w17652 ;
  assign w17654 = \pi064 & ~w17250 ;
  assign w17655 = \pi005 ^ w17654 ;
  assign w17656 = ( ~\pi004 & \pi064 ) | ( ~\pi004 & w17653 ) | ( \pi064 & w17653 ) ;
  assign w17657 = ( \pi065 & ~w17655 ) | ( \pi065 & w17656 ) | ( ~w17655 & w17656 ) ;
  assign w17658 = w17653 | w17657 ;
  assign w17659 = \pi067 ^ w17640 ;
  assign w17660 = ( ~w17649 & w17658 ) | ( ~w17649 & w17659 ) | ( w17658 & w17659 ) ;
  assign w17661 = w17659 | w17660 ;
  assign w17662 = \pi068 ^ w17634 ;
  assign w17663 = ( ~w17641 & w17661 ) | ( ~w17641 & w17662 ) | ( w17661 & w17662 ) ;
  assign w17664 = w17662 | w17663 ;
  assign w17665 = \pi069 ^ w17627 ;
  assign w17666 = ( ~w17635 & w17664 ) | ( ~w17635 & w17665 ) | ( w17664 & w17665 ) ;
  assign w17667 = w17665 | w17666 ;
  assign w17668 = \pi070 ^ w17620 ;
  assign w17669 = ( ~w17628 & w17667 ) | ( ~w17628 & w17668 ) | ( w17667 & w17668 ) ;
  assign w17670 = w17668 | w17669 ;
  assign w17671 = \pi071 ^ w17613 ;
  assign w17672 = ( ~w17621 & w17670 ) | ( ~w17621 & w17671 ) | ( w17670 & w17671 ) ;
  assign w17673 = w17671 | w17672 ;
  assign w17674 = \pi072 ^ w17606 ;
  assign w17675 = ( ~w17614 & w17673 ) | ( ~w17614 & w17674 ) | ( w17673 & w17674 ) ;
  assign w17676 = w17674 | w17675 ;
  assign w17677 = \pi073 ^ w17599 ;
  assign w17678 = ( ~w17607 & w17676 ) | ( ~w17607 & w17677 ) | ( w17676 & w17677 ) ;
  assign w17679 = w17677 | w17678 ;
  assign w17680 = \pi074 ^ w17592 ;
  assign w17681 = ( ~w17600 & w17679 ) | ( ~w17600 & w17680 ) | ( w17679 & w17680 ) ;
  assign w17682 = w17680 | w17681 ;
  assign w17683 = \pi075 ^ w17585 ;
  assign w17684 = ( ~w17593 & w17682 ) | ( ~w17593 & w17683 ) | ( w17682 & w17683 ) ;
  assign w17685 = w17683 | w17684 ;
  assign w17686 = \pi076 ^ w17578 ;
  assign w17687 = ( ~w17586 & w17685 ) | ( ~w17586 & w17686 ) | ( w17685 & w17686 ) ;
  assign w17688 = w17686 | w17687 ;
  assign w17689 = \pi077 ^ w17571 ;
  assign w17690 = ( ~w17579 & w17688 ) | ( ~w17579 & w17689 ) | ( w17688 & w17689 ) ;
  assign w17691 = w17689 | w17690 ;
  assign w17692 = \pi078 ^ w17564 ;
  assign w17693 = ( ~w17572 & w17691 ) | ( ~w17572 & w17692 ) | ( w17691 & w17692 ) ;
  assign w17694 = w17692 | w17693 ;
  assign w17695 = \pi079 ^ w17557 ;
  assign w17696 = ( ~w17565 & w17694 ) | ( ~w17565 & w17695 ) | ( w17694 & w17695 ) ;
  assign w17697 = w17695 | w17696 ;
  assign w17698 = \pi080 ^ w17550 ;
  assign w17699 = ( ~w17558 & w17697 ) | ( ~w17558 & w17698 ) | ( w17697 & w17698 ) ;
  assign w17700 = w17698 | w17699 ;
  assign w17701 = \pi081 ^ w17543 ;
  assign w17702 = ( ~w17551 & w17700 ) | ( ~w17551 & w17701 ) | ( w17700 & w17701 ) ;
  assign w17703 = w17701 | w17702 ;
  assign w17704 = \pi082 ^ w17536 ;
  assign w17705 = ( ~w17544 & w17703 ) | ( ~w17544 & w17704 ) | ( w17703 & w17704 ) ;
  assign w17706 = w17704 | w17705 ;
  assign w17707 = \pi083 ^ w17529 ;
  assign w17708 = ( ~w17537 & w17706 ) | ( ~w17537 & w17707 ) | ( w17706 & w17707 ) ;
  assign w17709 = w17707 | w17708 ;
  assign w17710 = \pi084 ^ w17522 ;
  assign w17711 = ( ~w17530 & w17709 ) | ( ~w17530 & w17710 ) | ( w17709 & w17710 ) ;
  assign w17712 = w17710 | w17711 ;
  assign w17713 = \pi085 ^ w17515 ;
  assign w17714 = ( ~w17523 & w17712 ) | ( ~w17523 & w17713 ) | ( w17712 & w17713 ) ;
  assign w17715 = w17713 | w17714 ;
  assign w17716 = \pi086 ^ w17508 ;
  assign w17717 = ( ~w17516 & w17715 ) | ( ~w17516 & w17716 ) | ( w17715 & w17716 ) ;
  assign w17718 = w17716 | w17717 ;
  assign w17719 = \pi087 ^ w17501 ;
  assign w17720 = ( ~w17509 & w17718 ) | ( ~w17509 & w17719 ) | ( w17718 & w17719 ) ;
  assign w17721 = w17719 | w17720 ;
  assign w17722 = \pi088 ^ w17494 ;
  assign w17723 = ( ~w17502 & w17721 ) | ( ~w17502 & w17722 ) | ( w17721 & w17722 ) ;
  assign w17724 = w17722 | w17723 ;
  assign w17725 = \pi089 ^ w17487 ;
  assign w17726 = ( ~w17495 & w17724 ) | ( ~w17495 & w17725 ) | ( w17724 & w17725 ) ;
  assign w17727 = w17725 | w17726 ;
  assign w17728 = \pi090 ^ w17480 ;
  assign w17729 = ( ~w17488 & w17727 ) | ( ~w17488 & w17728 ) | ( w17727 & w17728 ) ;
  assign w17730 = w17728 | w17729 ;
  assign w17731 = \pi091 ^ w17473 ;
  assign w17732 = ( ~w17481 & w17730 ) | ( ~w17481 & w17731 ) | ( w17730 & w17731 ) ;
  assign w17733 = w17731 | w17732 ;
  assign w17734 = \pi092 ^ w17466 ;
  assign w17735 = ( ~w17474 & w17733 ) | ( ~w17474 & w17734 ) | ( w17733 & w17734 ) ;
  assign w17736 = w17734 | w17735 ;
  assign w17737 = \pi093 ^ w17459 ;
  assign w17738 = ( ~w17467 & w17736 ) | ( ~w17467 & w17737 ) | ( w17736 & w17737 ) ;
  assign w17739 = w17737 | w17738 ;
  assign w17740 = \pi094 ^ w17452 ;
  assign w17741 = ( ~w17460 & w17739 ) | ( ~w17460 & w17740 ) | ( w17739 & w17740 ) ;
  assign w17742 = w17740 | w17741 ;
  assign w17743 = \pi095 ^ w17445 ;
  assign w17744 = ( ~w17453 & w17742 ) | ( ~w17453 & w17743 ) | ( w17742 & w17743 ) ;
  assign w17745 = w17743 | w17744 ;
  assign w17746 = \pi096 ^ w17438 ;
  assign w17747 = ( ~w17446 & w17745 ) | ( ~w17446 & w17746 ) | ( w17745 & w17746 ) ;
  assign w17748 = w17746 | w17747 ;
  assign w17749 = \pi097 ^ w17431 ;
  assign w17750 = ( ~w17439 & w17748 ) | ( ~w17439 & w17749 ) | ( w17748 & w17749 ) ;
  assign w17751 = w17749 | w17750 ;
  assign w17752 = \pi098 ^ w17424 ;
  assign w17753 = ( ~w17432 & w17751 ) | ( ~w17432 & w17752 ) | ( w17751 & w17752 ) ;
  assign w17754 = w17752 | w17753 ;
  assign w17755 = \pi099 ^ w17417 ;
  assign w17756 = ( ~w17425 & w17754 ) | ( ~w17425 & w17755 ) | ( w17754 & w17755 ) ;
  assign w17757 = w17755 | w17756 ;
  assign w17758 = \pi100 ^ w17410 ;
  assign w17759 = ( ~w17418 & w17757 ) | ( ~w17418 & w17758 ) | ( w17757 & w17758 ) ;
  assign w17760 = w17758 | w17759 ;
  assign w17761 = \pi101 ^ w17403 ;
  assign w17762 = ( ~w17411 & w17760 ) | ( ~w17411 & w17761 ) | ( w17760 & w17761 ) ;
  assign w17763 = w17761 | w17762 ;
  assign w17764 = \pi102 ^ w17396 ;
  assign w17765 = ( ~w17404 & w17763 ) | ( ~w17404 & w17764 ) | ( w17763 & w17764 ) ;
  assign w17766 = w17764 | w17765 ;
  assign w17767 = \pi103 ^ w17389 ;
  assign w17768 = ( ~w17397 & w17766 ) | ( ~w17397 & w17767 ) | ( w17766 & w17767 ) ;
  assign w17769 = w17767 | w17768 ;
  assign w17770 = \pi104 ^ w17382 ;
  assign w17771 = ( ~w17390 & w17769 ) | ( ~w17390 & w17770 ) | ( w17769 & w17770 ) ;
  assign w17772 = w17770 | w17771 ;
  assign w17773 = \pi105 ^ w17375 ;
  assign w17774 = ( ~w17383 & w17772 ) | ( ~w17383 & w17773 ) | ( w17772 & w17773 ) ;
  assign w17775 = w17773 | w17774 ;
  assign w17776 = \pi106 ^ w17368 ;
  assign w17777 = ( ~w17376 & w17775 ) | ( ~w17376 & w17776 ) | ( w17775 & w17776 ) ;
  assign w17778 = w17776 | w17777 ;
  assign w17779 = \pi107 ^ w17361 ;
  assign w17780 = ( ~w17369 & w17778 ) | ( ~w17369 & w17779 ) | ( w17778 & w17779 ) ;
  assign w17781 = w17779 | w17780 ;
  assign w17782 = \pi108 ^ w17354 ;
  assign w17783 = ( ~w17362 & w17781 ) | ( ~w17362 & w17782 ) | ( w17781 & w17782 ) ;
  assign w17784 = w17782 | w17783 ;
  assign w17785 = \pi109 ^ w17347 ;
  assign w17786 = ( ~w17355 & w17784 ) | ( ~w17355 & w17785 ) | ( w17784 & w17785 ) ;
  assign w17787 = w17785 | w17786 ;
  assign w17788 = \pi110 ^ w17340 ;
  assign w17789 = ( ~w17348 & w17787 ) | ( ~w17348 & w17788 ) | ( w17787 & w17788 ) ;
  assign w17790 = w17788 | w17789 ;
  assign w17791 = \pi111 ^ w17333 ;
  assign w17792 = ( ~w17341 & w17790 ) | ( ~w17341 & w17791 ) | ( w17790 & w17791 ) ;
  assign w17793 = w17791 | w17792 ;
  assign w17794 = \pi112 ^ w17326 ;
  assign w17795 = ( ~w17334 & w17793 ) | ( ~w17334 & w17794 ) | ( w17793 & w17794 ) ;
  assign w17796 = w17794 | w17795 ;
  assign w17797 = \pi113 ^ w17319 ;
  assign w17798 = ( ~w17327 & w17796 ) | ( ~w17327 & w17797 ) | ( w17796 & w17797 ) ;
  assign w17799 = w17797 | w17798 ;
  assign w17800 = \pi114 ^ w17312 ;
  assign w17801 = ( ~w17320 & w17799 ) | ( ~w17320 & w17800 ) | ( w17799 & w17800 ) ;
  assign w17802 = w17800 | w17801 ;
  assign w17803 = \pi115 ^ w17305 ;
  assign w17804 = ( ~w17313 & w17802 ) | ( ~w17313 & w17803 ) | ( w17802 & w17803 ) ;
  assign w17805 = w17803 | w17804 ;
  assign w17806 = \pi116 ^ w17298 ;
  assign w17807 = ( ~w17306 & w17805 ) | ( ~w17306 & w17806 ) | ( w17805 & w17806 ) ;
  assign w17808 = w17806 | w17807 ;
  assign w17809 = \pi117 ^ w17291 ;
  assign w17810 = ( ~w17299 & w17808 ) | ( ~w17299 & w17809 ) | ( w17808 & w17809 ) ;
  assign w17811 = w17809 | w17810 ;
  assign w17812 = \pi118 ^ w17284 ;
  assign w17813 = ( ~w17292 & w17811 ) | ( ~w17292 & w17812 ) | ( w17811 & w17812 ) ;
  assign w17814 = w17812 | w17813 ;
  assign w17815 = \pi119 ^ w17277 ;
  assign w17816 = ( ~w17285 & w17814 ) | ( ~w17285 & w17815 ) | ( w17814 & w17815 ) ;
  assign w17817 = w17815 | w17816 ;
  assign w17818 = \pi120 ^ w17270 ;
  assign w17819 = ( ~w17278 & w17817 ) | ( ~w17278 & w17818 ) | ( w17817 & w17818 ) ;
  assign w17820 = w17818 | w17819 ;
  assign w17821 = \pi121 ^ w17263 ;
  assign w17822 = ( ~w17271 & w17820 ) | ( ~w17271 & w17821 ) | ( w17820 & w17821 ) ;
  assign w17823 = w17821 | w17822 ;
  assign w17824 = \pi122 ^ w17256 ;
  assign w17825 = ( ~w17264 & w17823 ) | ( ~w17264 & w17824 ) | ( w17823 & w17824 ) ;
  assign w17826 = w17824 | w17825 ;
  assign w17827 = w17241 | w17243 ;
  assign w17828 = ( ~w16714 & w17235 ) | ( ~w16714 & w17250 ) | ( w17235 & w17250 ) ;
  assign w17829 = w17827 ^ w17828 ;
  assign w17830 = ~w17250 & w17829 ;
  assign w17831 = ( w16707 & ~w17240 ) | ( w16707 & w17248 ) | ( ~w17240 & w17248 ) ;
  assign w17832 = w17240 & w17831 ;
  assign w17833 = w17830 | w17832 ;
  assign w17834 = ~\pi123 & w17833 ;
  assign w17835 = ( \pi123 & ~w17830 ) | ( \pi123 & w17832 ) | ( ~w17830 & w17832 ) ;
  assign w17836 = ~w17832 & w17835 ;
  assign w17837 = w17834 | w17836 ;
  assign w17838 = ( ~w17257 & w17826 ) | ( ~w17257 & w17837 ) | ( w17826 & w17837 ) ;
  assign w17839 = ( w147 & ~w17837 ) | ( w147 & w17838 ) | ( ~w17837 & w17838 ) ;
  assign w17840 = w17837 | w17839 ;
  assign w17841 = ( w269 & ~w270 ) | ( w269 & w17833 ) | ( ~w270 & w17833 ) ;
  assign w17842 = ~w269 & w17841 ;
  assign w17843 = w17840 & ~w17842 ;
  assign w17844 = ~w17264 & w17823 ;
  assign w17845 = w17824 ^ w17844 ;
  assign w17846 = ~w17843 & w17845 ;
  assign w17847 = ( w17256 & w17840 ) | ( w17256 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17848 = ~w17842 & w17847 ;
  assign w17849 = w17846 | w17848 ;
  assign w17850 = ~\pi123 & w17849 ;
  assign w17851 = ~w17271 & w17820 ;
  assign w17852 = w17821 ^ w17851 ;
  assign w17853 = ~w17843 & w17852 ;
  assign w17854 = ( w17263 & w17840 ) | ( w17263 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17855 = ~w17842 & w17854 ;
  assign w17856 = w17853 | w17855 ;
  assign w17857 = ~\pi122 & w17856 ;
  assign w17858 = ~w17278 & w17817 ;
  assign w17859 = w17818 ^ w17858 ;
  assign w17860 = ~w17843 & w17859 ;
  assign w17861 = ( w17270 & w17840 ) | ( w17270 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17862 = ~w17842 & w17861 ;
  assign w17863 = w17860 | w17862 ;
  assign w17864 = ~\pi121 & w17863 ;
  assign w17865 = ~w17285 & w17814 ;
  assign w17866 = w17815 ^ w17865 ;
  assign w17867 = ~w17843 & w17866 ;
  assign w17868 = ( w17277 & w17840 ) | ( w17277 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17869 = ~w17842 & w17868 ;
  assign w17870 = w17867 | w17869 ;
  assign w17871 = ~\pi120 & w17870 ;
  assign w17872 = ~w17292 & w17811 ;
  assign w17873 = w17812 ^ w17872 ;
  assign w17874 = ~w17843 & w17873 ;
  assign w17875 = ( w17284 & w17840 ) | ( w17284 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17876 = ~w17842 & w17875 ;
  assign w17877 = w17874 | w17876 ;
  assign w17878 = ~\pi119 & w17877 ;
  assign w17879 = ~w17299 & w17808 ;
  assign w17880 = w17809 ^ w17879 ;
  assign w17881 = ~w17843 & w17880 ;
  assign w17882 = ( w17291 & w17840 ) | ( w17291 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17883 = ~w17842 & w17882 ;
  assign w17884 = w17881 | w17883 ;
  assign w17885 = ~\pi118 & w17884 ;
  assign w17886 = ~w17306 & w17805 ;
  assign w17887 = w17806 ^ w17886 ;
  assign w17888 = ~w17843 & w17887 ;
  assign w17889 = ( w17298 & w17840 ) | ( w17298 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17890 = ~w17842 & w17889 ;
  assign w17891 = w17888 | w17890 ;
  assign w17892 = ~\pi117 & w17891 ;
  assign w17893 = ~w17313 & w17802 ;
  assign w17894 = w17803 ^ w17893 ;
  assign w17895 = ~w17843 & w17894 ;
  assign w17896 = ( w17305 & w17840 ) | ( w17305 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17897 = ~w17842 & w17896 ;
  assign w17898 = w17895 | w17897 ;
  assign w17899 = ~\pi116 & w17898 ;
  assign w17900 = ~w17320 & w17799 ;
  assign w17901 = w17800 ^ w17900 ;
  assign w17902 = ~w17843 & w17901 ;
  assign w17903 = ( w17312 & w17840 ) | ( w17312 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17904 = ~w17842 & w17903 ;
  assign w17905 = w17902 | w17904 ;
  assign w17906 = ~\pi115 & w17905 ;
  assign w17907 = ~w17327 & w17796 ;
  assign w17908 = w17797 ^ w17907 ;
  assign w17909 = ~w17843 & w17908 ;
  assign w17910 = ( w17319 & w17840 ) | ( w17319 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17911 = ~w17842 & w17910 ;
  assign w17912 = w17909 | w17911 ;
  assign w17913 = ~\pi114 & w17912 ;
  assign w17914 = ~w17334 & w17793 ;
  assign w17915 = w17794 ^ w17914 ;
  assign w17916 = ~w17843 & w17915 ;
  assign w17917 = ( w17326 & w17840 ) | ( w17326 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17918 = ~w17842 & w17917 ;
  assign w17919 = w17916 | w17918 ;
  assign w17920 = ~\pi113 & w17919 ;
  assign w17921 = ~w17341 & w17790 ;
  assign w17922 = w17791 ^ w17921 ;
  assign w17923 = ~w17843 & w17922 ;
  assign w17924 = ( w17333 & w17840 ) | ( w17333 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17925 = ~w17842 & w17924 ;
  assign w17926 = w17923 | w17925 ;
  assign w17927 = ~\pi112 & w17926 ;
  assign w17928 = ~w17348 & w17787 ;
  assign w17929 = w17788 ^ w17928 ;
  assign w17930 = ~w17843 & w17929 ;
  assign w17931 = ( w17340 & w17840 ) | ( w17340 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17932 = ~w17842 & w17931 ;
  assign w17933 = w17930 | w17932 ;
  assign w17934 = ~\pi111 & w17933 ;
  assign w17935 = ~w17355 & w17784 ;
  assign w17936 = w17785 ^ w17935 ;
  assign w17937 = ~w17843 & w17936 ;
  assign w17938 = ( w17347 & w17840 ) | ( w17347 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17939 = ~w17842 & w17938 ;
  assign w17940 = w17937 | w17939 ;
  assign w17941 = ~\pi110 & w17940 ;
  assign w17942 = ~w17362 & w17781 ;
  assign w17943 = w17782 ^ w17942 ;
  assign w17944 = ~w17843 & w17943 ;
  assign w17945 = ( w17354 & w17840 ) | ( w17354 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17946 = ~w17842 & w17945 ;
  assign w17947 = w17944 | w17946 ;
  assign w17948 = ~\pi109 & w17947 ;
  assign w17949 = ~w17369 & w17778 ;
  assign w17950 = w17779 ^ w17949 ;
  assign w17951 = ~w17843 & w17950 ;
  assign w17952 = ( w17361 & w17840 ) | ( w17361 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17953 = ~w17842 & w17952 ;
  assign w17954 = w17951 | w17953 ;
  assign w17955 = ~\pi108 & w17954 ;
  assign w17956 = ~w17376 & w17775 ;
  assign w17957 = w17776 ^ w17956 ;
  assign w17958 = ~w17843 & w17957 ;
  assign w17959 = ( w17368 & w17840 ) | ( w17368 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17960 = ~w17842 & w17959 ;
  assign w17961 = w17958 | w17960 ;
  assign w17962 = ~\pi107 & w17961 ;
  assign w17963 = ~w17383 & w17772 ;
  assign w17964 = w17773 ^ w17963 ;
  assign w17965 = ~w17843 & w17964 ;
  assign w17966 = ( w17375 & w17840 ) | ( w17375 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17967 = ~w17842 & w17966 ;
  assign w17968 = w17965 | w17967 ;
  assign w17969 = ~\pi106 & w17968 ;
  assign w17970 = ~w17390 & w17769 ;
  assign w17971 = w17770 ^ w17970 ;
  assign w17972 = ~w17843 & w17971 ;
  assign w17973 = ( w17382 & w17840 ) | ( w17382 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17974 = ~w17842 & w17973 ;
  assign w17975 = w17972 | w17974 ;
  assign w17976 = ~\pi105 & w17975 ;
  assign w17977 = ~w17397 & w17766 ;
  assign w17978 = w17767 ^ w17977 ;
  assign w17979 = ~w17843 & w17978 ;
  assign w17980 = ( w17389 & w17840 ) | ( w17389 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17981 = ~w17842 & w17980 ;
  assign w17982 = w17979 | w17981 ;
  assign w17983 = ~\pi104 & w17982 ;
  assign w17984 = ~w17404 & w17763 ;
  assign w17985 = w17764 ^ w17984 ;
  assign w17986 = ~w17843 & w17985 ;
  assign w17987 = ( w17396 & w17840 ) | ( w17396 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17988 = ~w17842 & w17987 ;
  assign w17989 = w17986 | w17988 ;
  assign w17990 = ~\pi103 & w17989 ;
  assign w17991 = ~w17411 & w17760 ;
  assign w17992 = w17761 ^ w17991 ;
  assign w17993 = ~w17843 & w17992 ;
  assign w17994 = ( w17403 & w17840 ) | ( w17403 & w17842 ) | ( w17840 & w17842 ) ;
  assign w17995 = ~w17842 & w17994 ;
  assign w17996 = w17993 | w17995 ;
  assign w17997 = ~\pi102 & w17996 ;
  assign w17998 = ~w17418 & w17757 ;
  assign w17999 = w17758 ^ w17998 ;
  assign w18000 = ~w17843 & w17999 ;
  assign w18001 = ( w17410 & w17840 ) | ( w17410 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18002 = ~w17842 & w18001 ;
  assign w18003 = w18000 | w18002 ;
  assign w18004 = ~\pi101 & w18003 ;
  assign w18005 = ~w17425 & w17754 ;
  assign w18006 = w17755 ^ w18005 ;
  assign w18007 = ~w17843 & w18006 ;
  assign w18008 = ( w17417 & w17840 ) | ( w17417 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18009 = ~w17842 & w18008 ;
  assign w18010 = w18007 | w18009 ;
  assign w18011 = ~\pi100 & w18010 ;
  assign w18012 = ~w17432 & w17751 ;
  assign w18013 = w17752 ^ w18012 ;
  assign w18014 = ~w17843 & w18013 ;
  assign w18015 = ( w17424 & w17840 ) | ( w17424 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18016 = ~w17842 & w18015 ;
  assign w18017 = w18014 | w18016 ;
  assign w18018 = ~\pi099 & w18017 ;
  assign w18019 = ~w17439 & w17748 ;
  assign w18020 = w17749 ^ w18019 ;
  assign w18021 = ~w17843 & w18020 ;
  assign w18022 = ( w17431 & w17840 ) | ( w17431 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18023 = ~w17842 & w18022 ;
  assign w18024 = w18021 | w18023 ;
  assign w18025 = ~\pi098 & w18024 ;
  assign w18026 = ~w17446 & w17745 ;
  assign w18027 = w17746 ^ w18026 ;
  assign w18028 = ~w17843 & w18027 ;
  assign w18029 = ( w17438 & w17840 ) | ( w17438 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18030 = ~w17842 & w18029 ;
  assign w18031 = w18028 | w18030 ;
  assign w18032 = ~\pi097 & w18031 ;
  assign w18033 = ~w17453 & w17742 ;
  assign w18034 = w17743 ^ w18033 ;
  assign w18035 = ~w17843 & w18034 ;
  assign w18036 = ( w17445 & w17840 ) | ( w17445 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18037 = ~w17842 & w18036 ;
  assign w18038 = w18035 | w18037 ;
  assign w18039 = ~\pi096 & w18038 ;
  assign w18040 = ~w17460 & w17739 ;
  assign w18041 = w17740 ^ w18040 ;
  assign w18042 = ~w17843 & w18041 ;
  assign w18043 = ( w17452 & w17840 ) | ( w17452 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18044 = ~w17842 & w18043 ;
  assign w18045 = w18042 | w18044 ;
  assign w18046 = ~\pi095 & w18045 ;
  assign w18047 = ~w17467 & w17736 ;
  assign w18048 = w17737 ^ w18047 ;
  assign w18049 = ~w17843 & w18048 ;
  assign w18050 = ( w17459 & w17840 ) | ( w17459 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18051 = ~w17842 & w18050 ;
  assign w18052 = w18049 | w18051 ;
  assign w18053 = ~\pi094 & w18052 ;
  assign w18054 = ~w17474 & w17733 ;
  assign w18055 = w17734 ^ w18054 ;
  assign w18056 = ~w17843 & w18055 ;
  assign w18057 = ( w17466 & w17840 ) | ( w17466 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18058 = ~w17842 & w18057 ;
  assign w18059 = w18056 | w18058 ;
  assign w18060 = ~\pi093 & w18059 ;
  assign w18061 = ~w17481 & w17730 ;
  assign w18062 = w17731 ^ w18061 ;
  assign w18063 = ~w17843 & w18062 ;
  assign w18064 = ( w17473 & w17840 ) | ( w17473 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18065 = ~w17842 & w18064 ;
  assign w18066 = w18063 | w18065 ;
  assign w18067 = ~\pi092 & w18066 ;
  assign w18068 = ~w17488 & w17727 ;
  assign w18069 = w17728 ^ w18068 ;
  assign w18070 = ~w17843 & w18069 ;
  assign w18071 = ( w17480 & w17840 ) | ( w17480 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18072 = ~w17842 & w18071 ;
  assign w18073 = w18070 | w18072 ;
  assign w18074 = ~\pi091 & w18073 ;
  assign w18075 = ~w17495 & w17724 ;
  assign w18076 = w17725 ^ w18075 ;
  assign w18077 = ~w17843 & w18076 ;
  assign w18078 = ( w17487 & w17840 ) | ( w17487 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18079 = ~w17842 & w18078 ;
  assign w18080 = w18077 | w18079 ;
  assign w18081 = ~\pi090 & w18080 ;
  assign w18082 = ~w17502 & w17721 ;
  assign w18083 = w17722 ^ w18082 ;
  assign w18084 = ~w17843 & w18083 ;
  assign w18085 = ( w17494 & w17840 ) | ( w17494 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18086 = ~w17842 & w18085 ;
  assign w18087 = w18084 | w18086 ;
  assign w18088 = ~\pi089 & w18087 ;
  assign w18089 = ~w17509 & w17718 ;
  assign w18090 = w17719 ^ w18089 ;
  assign w18091 = ~w17843 & w18090 ;
  assign w18092 = ( w17501 & w17840 ) | ( w17501 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18093 = ~w17842 & w18092 ;
  assign w18094 = w18091 | w18093 ;
  assign w18095 = ~\pi088 & w18094 ;
  assign w18096 = ~w17516 & w17715 ;
  assign w18097 = w17716 ^ w18096 ;
  assign w18098 = ~w17843 & w18097 ;
  assign w18099 = ( w17508 & w17840 ) | ( w17508 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18100 = ~w17842 & w18099 ;
  assign w18101 = w18098 | w18100 ;
  assign w18102 = ~\pi087 & w18101 ;
  assign w18103 = ~w17523 & w17712 ;
  assign w18104 = w17713 ^ w18103 ;
  assign w18105 = ~w17843 & w18104 ;
  assign w18106 = ( w17515 & w17840 ) | ( w17515 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18107 = ~w17842 & w18106 ;
  assign w18108 = w18105 | w18107 ;
  assign w18109 = ~\pi086 & w18108 ;
  assign w18110 = ~w17530 & w17709 ;
  assign w18111 = w17710 ^ w18110 ;
  assign w18112 = ~w17843 & w18111 ;
  assign w18113 = ( w17522 & w17840 ) | ( w17522 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18114 = ~w17842 & w18113 ;
  assign w18115 = w18112 | w18114 ;
  assign w18116 = ~\pi085 & w18115 ;
  assign w18117 = ~w17537 & w17706 ;
  assign w18118 = w17707 ^ w18117 ;
  assign w18119 = ~w17843 & w18118 ;
  assign w18120 = ( w17529 & w17840 ) | ( w17529 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18121 = ~w17842 & w18120 ;
  assign w18122 = w18119 | w18121 ;
  assign w18123 = ~\pi084 & w18122 ;
  assign w18124 = ~w17544 & w17703 ;
  assign w18125 = w17704 ^ w18124 ;
  assign w18126 = ~w17843 & w18125 ;
  assign w18127 = ( w17536 & w17840 ) | ( w17536 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18128 = ~w17842 & w18127 ;
  assign w18129 = w18126 | w18128 ;
  assign w18130 = ~\pi083 & w18129 ;
  assign w18131 = ~w17551 & w17700 ;
  assign w18132 = w17701 ^ w18131 ;
  assign w18133 = ~w17843 & w18132 ;
  assign w18134 = ( w17543 & w17840 ) | ( w17543 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18135 = ~w17842 & w18134 ;
  assign w18136 = w18133 | w18135 ;
  assign w18137 = ~\pi082 & w18136 ;
  assign w18138 = ~w17558 & w17697 ;
  assign w18139 = w17698 ^ w18138 ;
  assign w18140 = ~w17843 & w18139 ;
  assign w18141 = ( w17550 & w17840 ) | ( w17550 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18142 = ~w17842 & w18141 ;
  assign w18143 = w18140 | w18142 ;
  assign w18144 = ~\pi081 & w18143 ;
  assign w18145 = ~w17565 & w17694 ;
  assign w18146 = w17695 ^ w18145 ;
  assign w18147 = ~w17843 & w18146 ;
  assign w18148 = ( w17557 & w17840 ) | ( w17557 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18149 = ~w17842 & w18148 ;
  assign w18150 = w18147 | w18149 ;
  assign w18151 = ~\pi080 & w18150 ;
  assign w18152 = ~w17572 & w17691 ;
  assign w18153 = w17692 ^ w18152 ;
  assign w18154 = ~w17843 & w18153 ;
  assign w18155 = ( w17564 & w17840 ) | ( w17564 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18156 = ~w17842 & w18155 ;
  assign w18157 = w18154 | w18156 ;
  assign w18158 = ~\pi079 & w18157 ;
  assign w18159 = ~w17579 & w17688 ;
  assign w18160 = w17689 ^ w18159 ;
  assign w18161 = ~w17843 & w18160 ;
  assign w18162 = ( w17571 & w17840 ) | ( w17571 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18163 = ~w17842 & w18162 ;
  assign w18164 = w18161 | w18163 ;
  assign w18165 = ~\pi078 & w18164 ;
  assign w18166 = ~w17586 & w17685 ;
  assign w18167 = w17686 ^ w18166 ;
  assign w18168 = ~w17843 & w18167 ;
  assign w18169 = ( w17578 & w17840 ) | ( w17578 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18170 = ~w17842 & w18169 ;
  assign w18171 = w18168 | w18170 ;
  assign w18172 = ~\pi077 & w18171 ;
  assign w18173 = ~w17593 & w17682 ;
  assign w18174 = w17683 ^ w18173 ;
  assign w18175 = ~w17843 & w18174 ;
  assign w18176 = ( w17585 & w17840 ) | ( w17585 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18177 = ~w17842 & w18176 ;
  assign w18178 = w18175 | w18177 ;
  assign w18179 = ~\pi076 & w18178 ;
  assign w18180 = ~w17600 & w17679 ;
  assign w18181 = w17680 ^ w18180 ;
  assign w18182 = ~w17843 & w18181 ;
  assign w18183 = ( w17592 & w17840 ) | ( w17592 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18184 = ~w17842 & w18183 ;
  assign w18185 = w18182 | w18184 ;
  assign w18186 = ~\pi075 & w18185 ;
  assign w18187 = ~w17607 & w17676 ;
  assign w18188 = w17677 ^ w18187 ;
  assign w18189 = ~w17843 & w18188 ;
  assign w18190 = ( w17599 & w17840 ) | ( w17599 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18191 = ~w17842 & w18190 ;
  assign w18192 = w18189 | w18191 ;
  assign w18193 = ~\pi074 & w18192 ;
  assign w18194 = ~w17614 & w17673 ;
  assign w18195 = w17674 ^ w18194 ;
  assign w18196 = ~w17843 & w18195 ;
  assign w18197 = ( w17606 & w17840 ) | ( w17606 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18198 = ~w17842 & w18197 ;
  assign w18199 = w18196 | w18198 ;
  assign w18200 = ~\pi073 & w18199 ;
  assign w18201 = ~w17621 & w17670 ;
  assign w18202 = w17671 ^ w18201 ;
  assign w18203 = ~w17843 & w18202 ;
  assign w18204 = ( w17613 & w17840 ) | ( w17613 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18205 = ~w17842 & w18204 ;
  assign w18206 = w18203 | w18205 ;
  assign w18207 = ~\pi072 & w18206 ;
  assign w18208 = ~w17628 & w17667 ;
  assign w18209 = w17668 ^ w18208 ;
  assign w18210 = ~w17843 & w18209 ;
  assign w18211 = ( w17620 & w17840 ) | ( w17620 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18212 = ~w17842 & w18211 ;
  assign w18213 = w18210 | w18212 ;
  assign w18214 = ~\pi071 & w18213 ;
  assign w18215 = ~w17635 & w17664 ;
  assign w18216 = w17665 ^ w18215 ;
  assign w18217 = ~w17843 & w18216 ;
  assign w18218 = ( w17627 & w17840 ) | ( w17627 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18219 = ~w17842 & w18218 ;
  assign w18220 = w18217 | w18219 ;
  assign w18221 = ~\pi070 & w18220 ;
  assign w18222 = ~w17641 & w17661 ;
  assign w18223 = w17662 ^ w18222 ;
  assign w18224 = ~w17843 & w18223 ;
  assign w18225 = ( w17634 & w17840 ) | ( w17634 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18226 = ~w17842 & w18225 ;
  assign w18227 = w18224 | w18226 ;
  assign w18228 = ~\pi069 & w18227 ;
  assign w18229 = ~w17649 & w17658 ;
  assign w18230 = w17659 ^ w18229 ;
  assign w18231 = ~w17843 & w18230 ;
  assign w18232 = ( w17640 & w17840 ) | ( w17640 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18233 = ~w17842 & w18232 ;
  assign w18234 = w18231 | w18233 ;
  assign w18235 = ~\pi068 & w18234 ;
  assign w18236 = ~\pi004 & \pi064 ;
  assign w18237 = ( \pi065 & ~w17655 ) | ( \pi065 & w18236 ) | ( ~w17655 & w18236 ) ;
  assign w18238 = w17653 ^ w18237 ;
  assign w18239 = ~w17843 & w18238 ;
  assign w18240 = ( w17648 & w17840 ) | ( w17648 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18241 = ~w17842 & w18240 ;
  assign w18242 = w18239 | w18241 ;
  assign w18243 = ~\pi067 & w18242 ;
  assign w18244 = \pi005 ^ \pi065 ;
  assign w18245 = \pi004 ^ w17250 ;
  assign w18246 = ( \pi064 & w17843 ) | ( \pi064 & w18245 ) | ( w17843 & w18245 ) ;
  assign w18247 = w18244 ^ w18246 ;
  assign w18248 = ~w17843 & w18247 ;
  assign w18249 = w17655 & w17843 ;
  assign w18250 = w18248 | w18249 ;
  assign w18251 = ~\pi066 & w18250 ;
  assign w18252 = \pi066 ^ w18250 ;
  assign w18253 = \pi064 & ~w17843 ;
  assign w18254 = \pi004 ^ w18253 ;
  assign w18255 = ( ~\pi003 & \pi064 ) | ( ~\pi003 & w18252 ) | ( \pi064 & w18252 ) ;
  assign w18256 = ( \pi065 & ~w18254 ) | ( \pi065 & w18255 ) | ( ~w18254 & w18255 ) ;
  assign w18257 = w18252 | w18256 ;
  assign w18258 = \pi067 ^ w18242 ;
  assign w18259 = ( ~w18251 & w18257 ) | ( ~w18251 & w18258 ) | ( w18257 & w18258 ) ;
  assign w18260 = w18258 | w18259 ;
  assign w18261 = \pi068 ^ w18234 ;
  assign w18262 = ( ~w18243 & w18260 ) | ( ~w18243 & w18261 ) | ( w18260 & w18261 ) ;
  assign w18263 = w18261 | w18262 ;
  assign w18264 = \pi069 ^ w18227 ;
  assign w18265 = ( ~w18235 & w18263 ) | ( ~w18235 & w18264 ) | ( w18263 & w18264 ) ;
  assign w18266 = w18264 | w18265 ;
  assign w18267 = \pi070 ^ w18220 ;
  assign w18268 = ( ~w18228 & w18266 ) | ( ~w18228 & w18267 ) | ( w18266 & w18267 ) ;
  assign w18269 = w18267 | w18268 ;
  assign w18270 = \pi071 ^ w18213 ;
  assign w18271 = ( ~w18221 & w18269 ) | ( ~w18221 & w18270 ) | ( w18269 & w18270 ) ;
  assign w18272 = w18270 | w18271 ;
  assign w18273 = \pi072 ^ w18206 ;
  assign w18274 = ( ~w18214 & w18272 ) | ( ~w18214 & w18273 ) | ( w18272 & w18273 ) ;
  assign w18275 = w18273 | w18274 ;
  assign w18276 = \pi073 ^ w18199 ;
  assign w18277 = ( ~w18207 & w18275 ) | ( ~w18207 & w18276 ) | ( w18275 & w18276 ) ;
  assign w18278 = w18276 | w18277 ;
  assign w18279 = \pi074 ^ w18192 ;
  assign w18280 = ( ~w18200 & w18278 ) | ( ~w18200 & w18279 ) | ( w18278 & w18279 ) ;
  assign w18281 = w18279 | w18280 ;
  assign w18282 = \pi075 ^ w18185 ;
  assign w18283 = ( ~w18193 & w18281 ) | ( ~w18193 & w18282 ) | ( w18281 & w18282 ) ;
  assign w18284 = w18282 | w18283 ;
  assign w18285 = \pi076 ^ w18178 ;
  assign w18286 = ( ~w18186 & w18284 ) | ( ~w18186 & w18285 ) | ( w18284 & w18285 ) ;
  assign w18287 = w18285 | w18286 ;
  assign w18288 = \pi077 ^ w18171 ;
  assign w18289 = ( ~w18179 & w18287 ) | ( ~w18179 & w18288 ) | ( w18287 & w18288 ) ;
  assign w18290 = w18288 | w18289 ;
  assign w18291 = \pi078 ^ w18164 ;
  assign w18292 = ( ~w18172 & w18290 ) | ( ~w18172 & w18291 ) | ( w18290 & w18291 ) ;
  assign w18293 = w18291 | w18292 ;
  assign w18294 = \pi079 ^ w18157 ;
  assign w18295 = ( ~w18165 & w18293 ) | ( ~w18165 & w18294 ) | ( w18293 & w18294 ) ;
  assign w18296 = w18294 | w18295 ;
  assign w18297 = \pi080 ^ w18150 ;
  assign w18298 = ( ~w18158 & w18296 ) | ( ~w18158 & w18297 ) | ( w18296 & w18297 ) ;
  assign w18299 = w18297 | w18298 ;
  assign w18300 = \pi081 ^ w18143 ;
  assign w18301 = ( ~w18151 & w18299 ) | ( ~w18151 & w18300 ) | ( w18299 & w18300 ) ;
  assign w18302 = w18300 | w18301 ;
  assign w18303 = \pi082 ^ w18136 ;
  assign w18304 = ( ~w18144 & w18302 ) | ( ~w18144 & w18303 ) | ( w18302 & w18303 ) ;
  assign w18305 = w18303 | w18304 ;
  assign w18306 = \pi083 ^ w18129 ;
  assign w18307 = ( ~w18137 & w18305 ) | ( ~w18137 & w18306 ) | ( w18305 & w18306 ) ;
  assign w18308 = w18306 | w18307 ;
  assign w18309 = \pi084 ^ w18122 ;
  assign w18310 = ( ~w18130 & w18308 ) | ( ~w18130 & w18309 ) | ( w18308 & w18309 ) ;
  assign w18311 = w18309 | w18310 ;
  assign w18312 = \pi085 ^ w18115 ;
  assign w18313 = ( ~w18123 & w18311 ) | ( ~w18123 & w18312 ) | ( w18311 & w18312 ) ;
  assign w18314 = w18312 | w18313 ;
  assign w18315 = \pi086 ^ w18108 ;
  assign w18316 = ( ~w18116 & w18314 ) | ( ~w18116 & w18315 ) | ( w18314 & w18315 ) ;
  assign w18317 = w18315 | w18316 ;
  assign w18318 = \pi087 ^ w18101 ;
  assign w18319 = ( ~w18109 & w18317 ) | ( ~w18109 & w18318 ) | ( w18317 & w18318 ) ;
  assign w18320 = w18318 | w18319 ;
  assign w18321 = \pi088 ^ w18094 ;
  assign w18322 = ( ~w18102 & w18320 ) | ( ~w18102 & w18321 ) | ( w18320 & w18321 ) ;
  assign w18323 = w18321 | w18322 ;
  assign w18324 = \pi089 ^ w18087 ;
  assign w18325 = ( ~w18095 & w18323 ) | ( ~w18095 & w18324 ) | ( w18323 & w18324 ) ;
  assign w18326 = w18324 | w18325 ;
  assign w18327 = \pi090 ^ w18080 ;
  assign w18328 = ( ~w18088 & w18326 ) | ( ~w18088 & w18327 ) | ( w18326 & w18327 ) ;
  assign w18329 = w18327 | w18328 ;
  assign w18330 = \pi091 ^ w18073 ;
  assign w18331 = ( ~w18081 & w18329 ) | ( ~w18081 & w18330 ) | ( w18329 & w18330 ) ;
  assign w18332 = w18330 | w18331 ;
  assign w18333 = \pi092 ^ w18066 ;
  assign w18334 = ( ~w18074 & w18332 ) | ( ~w18074 & w18333 ) | ( w18332 & w18333 ) ;
  assign w18335 = w18333 | w18334 ;
  assign w18336 = \pi093 ^ w18059 ;
  assign w18337 = ( ~w18067 & w18335 ) | ( ~w18067 & w18336 ) | ( w18335 & w18336 ) ;
  assign w18338 = w18336 | w18337 ;
  assign w18339 = \pi094 ^ w18052 ;
  assign w18340 = ( ~w18060 & w18338 ) | ( ~w18060 & w18339 ) | ( w18338 & w18339 ) ;
  assign w18341 = w18339 | w18340 ;
  assign w18342 = \pi095 ^ w18045 ;
  assign w18343 = ( ~w18053 & w18341 ) | ( ~w18053 & w18342 ) | ( w18341 & w18342 ) ;
  assign w18344 = w18342 | w18343 ;
  assign w18345 = \pi096 ^ w18038 ;
  assign w18346 = ( ~w18046 & w18344 ) | ( ~w18046 & w18345 ) | ( w18344 & w18345 ) ;
  assign w18347 = w18345 | w18346 ;
  assign w18348 = \pi097 ^ w18031 ;
  assign w18349 = ( ~w18039 & w18347 ) | ( ~w18039 & w18348 ) | ( w18347 & w18348 ) ;
  assign w18350 = w18348 | w18349 ;
  assign w18351 = \pi098 ^ w18024 ;
  assign w18352 = ( ~w18032 & w18350 ) | ( ~w18032 & w18351 ) | ( w18350 & w18351 ) ;
  assign w18353 = w18351 | w18352 ;
  assign w18354 = \pi099 ^ w18017 ;
  assign w18355 = ( ~w18025 & w18353 ) | ( ~w18025 & w18354 ) | ( w18353 & w18354 ) ;
  assign w18356 = w18354 | w18355 ;
  assign w18357 = \pi100 ^ w18010 ;
  assign w18358 = ( ~w18018 & w18356 ) | ( ~w18018 & w18357 ) | ( w18356 & w18357 ) ;
  assign w18359 = w18357 | w18358 ;
  assign w18360 = \pi101 ^ w18003 ;
  assign w18361 = ( ~w18011 & w18359 ) | ( ~w18011 & w18360 ) | ( w18359 & w18360 ) ;
  assign w18362 = w18360 | w18361 ;
  assign w18363 = \pi102 ^ w17996 ;
  assign w18364 = ( ~w18004 & w18362 ) | ( ~w18004 & w18363 ) | ( w18362 & w18363 ) ;
  assign w18365 = w18363 | w18364 ;
  assign w18366 = \pi103 ^ w17989 ;
  assign w18367 = ( ~w17997 & w18365 ) | ( ~w17997 & w18366 ) | ( w18365 & w18366 ) ;
  assign w18368 = w18366 | w18367 ;
  assign w18369 = \pi104 ^ w17982 ;
  assign w18370 = ( ~w17990 & w18368 ) | ( ~w17990 & w18369 ) | ( w18368 & w18369 ) ;
  assign w18371 = w18369 | w18370 ;
  assign w18372 = \pi105 ^ w17975 ;
  assign w18373 = ( ~w17983 & w18371 ) | ( ~w17983 & w18372 ) | ( w18371 & w18372 ) ;
  assign w18374 = w18372 | w18373 ;
  assign w18375 = \pi106 ^ w17968 ;
  assign w18376 = ( ~w17976 & w18374 ) | ( ~w17976 & w18375 ) | ( w18374 & w18375 ) ;
  assign w18377 = w18375 | w18376 ;
  assign w18378 = \pi107 ^ w17961 ;
  assign w18379 = ( ~w17969 & w18377 ) | ( ~w17969 & w18378 ) | ( w18377 & w18378 ) ;
  assign w18380 = w18378 | w18379 ;
  assign w18381 = \pi108 ^ w17954 ;
  assign w18382 = ( ~w17962 & w18380 ) | ( ~w17962 & w18381 ) | ( w18380 & w18381 ) ;
  assign w18383 = w18381 | w18382 ;
  assign w18384 = \pi109 ^ w17947 ;
  assign w18385 = ( ~w17955 & w18383 ) | ( ~w17955 & w18384 ) | ( w18383 & w18384 ) ;
  assign w18386 = w18384 | w18385 ;
  assign w18387 = \pi110 ^ w17940 ;
  assign w18388 = ( ~w17948 & w18386 ) | ( ~w17948 & w18387 ) | ( w18386 & w18387 ) ;
  assign w18389 = w18387 | w18388 ;
  assign w18390 = \pi111 ^ w17933 ;
  assign w18391 = ( ~w17941 & w18389 ) | ( ~w17941 & w18390 ) | ( w18389 & w18390 ) ;
  assign w18392 = w18390 | w18391 ;
  assign w18393 = \pi112 ^ w17926 ;
  assign w18394 = ( ~w17934 & w18392 ) | ( ~w17934 & w18393 ) | ( w18392 & w18393 ) ;
  assign w18395 = w18393 | w18394 ;
  assign w18396 = \pi113 ^ w17919 ;
  assign w18397 = ( ~w17927 & w18395 ) | ( ~w17927 & w18396 ) | ( w18395 & w18396 ) ;
  assign w18398 = w18396 | w18397 ;
  assign w18399 = \pi114 ^ w17912 ;
  assign w18400 = ( ~w17920 & w18398 ) | ( ~w17920 & w18399 ) | ( w18398 & w18399 ) ;
  assign w18401 = w18399 | w18400 ;
  assign w18402 = \pi115 ^ w17905 ;
  assign w18403 = ( ~w17913 & w18401 ) | ( ~w17913 & w18402 ) | ( w18401 & w18402 ) ;
  assign w18404 = w18402 | w18403 ;
  assign w18405 = \pi116 ^ w17898 ;
  assign w18406 = ( ~w17906 & w18404 ) | ( ~w17906 & w18405 ) | ( w18404 & w18405 ) ;
  assign w18407 = w18405 | w18406 ;
  assign w18408 = \pi117 ^ w17891 ;
  assign w18409 = ( ~w17899 & w18407 ) | ( ~w17899 & w18408 ) | ( w18407 & w18408 ) ;
  assign w18410 = w18408 | w18409 ;
  assign w18411 = \pi118 ^ w17884 ;
  assign w18412 = ( ~w17892 & w18410 ) | ( ~w17892 & w18411 ) | ( w18410 & w18411 ) ;
  assign w18413 = w18411 | w18412 ;
  assign w18414 = \pi119 ^ w17877 ;
  assign w18415 = ( ~w17885 & w18413 ) | ( ~w17885 & w18414 ) | ( w18413 & w18414 ) ;
  assign w18416 = w18414 | w18415 ;
  assign w18417 = \pi120 ^ w17870 ;
  assign w18418 = ( ~w17878 & w18416 ) | ( ~w17878 & w18417 ) | ( w18416 & w18417 ) ;
  assign w18419 = w18417 | w18418 ;
  assign w18420 = \pi121 ^ w17863 ;
  assign w18421 = ( ~w17871 & w18419 ) | ( ~w17871 & w18420 ) | ( w18419 & w18420 ) ;
  assign w18422 = w18420 | w18421 ;
  assign w18423 = \pi122 ^ w17856 ;
  assign w18424 = ( ~w17864 & w18422 ) | ( ~w17864 & w18423 ) | ( w18422 & w18423 ) ;
  assign w18425 = w18423 | w18424 ;
  assign w18426 = \pi123 ^ w17849 ;
  assign w18427 = ( ~w17857 & w18425 ) | ( ~w17857 & w18426 ) | ( w18425 & w18426 ) ;
  assign w18428 = w18426 | w18427 ;
  assign w18429 = ( ~w17257 & w17826 ) | ( ~w17257 & w17843 ) | ( w17826 & w17843 ) ;
  assign w18430 = w17837 ^ w18429 ;
  assign w18431 = ~w17843 & w18430 ;
  assign w18432 = ( w17833 & w17840 ) | ( w17833 & w17842 ) | ( w17840 & w17842 ) ;
  assign w18433 = ~w17842 & w18432 ;
  assign w18434 = w18431 | w18433 ;
  assign w18435 = ~\pi124 & w18434 ;
  assign w18436 = ( \pi124 & ~w18431 ) | ( \pi124 & w18433 ) | ( ~w18431 & w18433 ) ;
  assign w18437 = ~w18433 & w18436 ;
  assign w18438 = w18435 | w18437 ;
  assign w18439 = ( ~w17850 & w18428 ) | ( ~w17850 & w18438 ) | ( w18428 & w18438 ) ;
  assign w18440 = ( w269 & ~w18438 ) | ( w269 & w18439 ) | ( ~w18438 & w18439 ) ;
  assign w18441 = w18438 | w18440 ;
  assign w18442 = ~w147 & w18434 ;
  assign w18443 = w18441 & ~w18442 ;
  assign w18444 = ~w17857 & w18425 ;
  assign w18445 = w18426 ^ w18444 ;
  assign w18446 = ~w18443 & w18445 ;
  assign w18447 = ( w17849 & w18441 ) | ( w17849 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18448 = ~w18442 & w18447 ;
  assign w18449 = w18446 | w18448 ;
  assign w18450 = ~\pi124 & w18449 ;
  assign w18451 = ~w17864 & w18422 ;
  assign w18452 = w18423 ^ w18451 ;
  assign w18453 = ~w18443 & w18452 ;
  assign w18454 = ( w17856 & w18441 ) | ( w17856 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18455 = ~w18442 & w18454 ;
  assign w18456 = w18453 | w18455 ;
  assign w18457 = ~\pi123 & w18456 ;
  assign w18458 = ~w17871 & w18419 ;
  assign w18459 = w18420 ^ w18458 ;
  assign w18460 = ~w18443 & w18459 ;
  assign w18461 = ( w17863 & w18441 ) | ( w17863 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18462 = ~w18442 & w18461 ;
  assign w18463 = w18460 | w18462 ;
  assign w18464 = ~\pi122 & w18463 ;
  assign w18465 = ~w17878 & w18416 ;
  assign w18466 = w18417 ^ w18465 ;
  assign w18467 = ~w18443 & w18466 ;
  assign w18468 = ( w17870 & w18441 ) | ( w17870 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18469 = ~w18442 & w18468 ;
  assign w18470 = w18467 | w18469 ;
  assign w18471 = ~\pi121 & w18470 ;
  assign w18472 = ~w17885 & w18413 ;
  assign w18473 = w18414 ^ w18472 ;
  assign w18474 = ~w18443 & w18473 ;
  assign w18475 = ( w17877 & w18441 ) | ( w17877 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18476 = ~w18442 & w18475 ;
  assign w18477 = w18474 | w18476 ;
  assign w18478 = ~\pi120 & w18477 ;
  assign w18479 = ~w17892 & w18410 ;
  assign w18480 = w18411 ^ w18479 ;
  assign w18481 = ~w18443 & w18480 ;
  assign w18482 = ( w17884 & w18441 ) | ( w17884 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18483 = ~w18442 & w18482 ;
  assign w18484 = w18481 | w18483 ;
  assign w18485 = ~\pi119 & w18484 ;
  assign w18486 = ~w17899 & w18407 ;
  assign w18487 = w18408 ^ w18486 ;
  assign w18488 = ~w18443 & w18487 ;
  assign w18489 = ( w17891 & w18441 ) | ( w17891 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18490 = ~w18442 & w18489 ;
  assign w18491 = w18488 | w18490 ;
  assign w18492 = ~\pi118 & w18491 ;
  assign w18493 = ~w17906 & w18404 ;
  assign w18494 = w18405 ^ w18493 ;
  assign w18495 = ~w18443 & w18494 ;
  assign w18496 = ( w17898 & w18441 ) | ( w17898 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18497 = ~w18442 & w18496 ;
  assign w18498 = w18495 | w18497 ;
  assign w18499 = ~\pi117 & w18498 ;
  assign w18500 = ~w17913 & w18401 ;
  assign w18501 = w18402 ^ w18500 ;
  assign w18502 = ~w18443 & w18501 ;
  assign w18503 = ( w17905 & w18441 ) | ( w17905 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18504 = ~w18442 & w18503 ;
  assign w18505 = w18502 | w18504 ;
  assign w18506 = ~\pi116 & w18505 ;
  assign w18507 = ~w17920 & w18398 ;
  assign w18508 = w18399 ^ w18507 ;
  assign w18509 = ~w18443 & w18508 ;
  assign w18510 = ( w17912 & w18441 ) | ( w17912 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18511 = ~w18442 & w18510 ;
  assign w18512 = w18509 | w18511 ;
  assign w18513 = ~\pi115 & w18512 ;
  assign w18514 = ~w17927 & w18395 ;
  assign w18515 = w18396 ^ w18514 ;
  assign w18516 = ~w18443 & w18515 ;
  assign w18517 = ( w17919 & w18441 ) | ( w17919 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18518 = ~w18442 & w18517 ;
  assign w18519 = w18516 | w18518 ;
  assign w18520 = ~\pi114 & w18519 ;
  assign w18521 = ~w17934 & w18392 ;
  assign w18522 = w18393 ^ w18521 ;
  assign w18523 = ~w18443 & w18522 ;
  assign w18524 = ( w17926 & w18441 ) | ( w17926 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18525 = ~w18442 & w18524 ;
  assign w18526 = w18523 | w18525 ;
  assign w18527 = ~\pi113 & w18526 ;
  assign w18528 = ~w17941 & w18389 ;
  assign w18529 = w18390 ^ w18528 ;
  assign w18530 = ~w18443 & w18529 ;
  assign w18531 = ( w17933 & w18441 ) | ( w17933 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18532 = ~w18442 & w18531 ;
  assign w18533 = w18530 | w18532 ;
  assign w18534 = ~\pi112 & w18533 ;
  assign w18535 = ~w17948 & w18386 ;
  assign w18536 = w18387 ^ w18535 ;
  assign w18537 = ~w18443 & w18536 ;
  assign w18538 = ( w17940 & w18441 ) | ( w17940 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18539 = ~w18442 & w18538 ;
  assign w18540 = w18537 | w18539 ;
  assign w18541 = ~\pi111 & w18540 ;
  assign w18542 = ~w17955 & w18383 ;
  assign w18543 = w18384 ^ w18542 ;
  assign w18544 = ~w18443 & w18543 ;
  assign w18545 = ( w17947 & w18441 ) | ( w17947 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18546 = ~w18442 & w18545 ;
  assign w18547 = w18544 | w18546 ;
  assign w18548 = ~\pi110 & w18547 ;
  assign w18549 = ~w17962 & w18380 ;
  assign w18550 = w18381 ^ w18549 ;
  assign w18551 = ~w18443 & w18550 ;
  assign w18552 = ( w17954 & w18441 ) | ( w17954 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18553 = ~w18442 & w18552 ;
  assign w18554 = w18551 | w18553 ;
  assign w18555 = ~\pi109 & w18554 ;
  assign w18556 = ~w17969 & w18377 ;
  assign w18557 = w18378 ^ w18556 ;
  assign w18558 = ~w18443 & w18557 ;
  assign w18559 = ( w17961 & w18441 ) | ( w17961 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18560 = ~w18442 & w18559 ;
  assign w18561 = w18558 | w18560 ;
  assign w18562 = ~\pi108 & w18561 ;
  assign w18563 = ~w17976 & w18374 ;
  assign w18564 = w18375 ^ w18563 ;
  assign w18565 = ~w18443 & w18564 ;
  assign w18566 = ( w17968 & w18441 ) | ( w17968 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18567 = ~w18442 & w18566 ;
  assign w18568 = w18565 | w18567 ;
  assign w18569 = ~\pi107 & w18568 ;
  assign w18570 = ~w17983 & w18371 ;
  assign w18571 = w18372 ^ w18570 ;
  assign w18572 = ~w18443 & w18571 ;
  assign w18573 = ( w17975 & w18441 ) | ( w17975 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18574 = ~w18442 & w18573 ;
  assign w18575 = w18572 | w18574 ;
  assign w18576 = ~\pi106 & w18575 ;
  assign w18577 = ~w17990 & w18368 ;
  assign w18578 = w18369 ^ w18577 ;
  assign w18579 = ~w18443 & w18578 ;
  assign w18580 = ( w17982 & w18441 ) | ( w17982 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18581 = ~w18442 & w18580 ;
  assign w18582 = w18579 | w18581 ;
  assign w18583 = ~\pi105 & w18582 ;
  assign w18584 = ~w17997 & w18365 ;
  assign w18585 = w18366 ^ w18584 ;
  assign w18586 = ~w18443 & w18585 ;
  assign w18587 = ( w17989 & w18441 ) | ( w17989 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18588 = ~w18442 & w18587 ;
  assign w18589 = w18586 | w18588 ;
  assign w18590 = ~\pi104 & w18589 ;
  assign w18591 = ~w18004 & w18362 ;
  assign w18592 = w18363 ^ w18591 ;
  assign w18593 = ~w18443 & w18592 ;
  assign w18594 = ( w17996 & w18441 ) | ( w17996 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18595 = ~w18442 & w18594 ;
  assign w18596 = w18593 | w18595 ;
  assign w18597 = ~\pi103 & w18596 ;
  assign w18598 = ~w18011 & w18359 ;
  assign w18599 = w18360 ^ w18598 ;
  assign w18600 = ~w18443 & w18599 ;
  assign w18601 = ( w18003 & w18441 ) | ( w18003 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18602 = ~w18442 & w18601 ;
  assign w18603 = w18600 | w18602 ;
  assign w18604 = ~\pi102 & w18603 ;
  assign w18605 = ~w18018 & w18356 ;
  assign w18606 = w18357 ^ w18605 ;
  assign w18607 = ~w18443 & w18606 ;
  assign w18608 = ( w18010 & w18441 ) | ( w18010 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18609 = ~w18442 & w18608 ;
  assign w18610 = w18607 | w18609 ;
  assign w18611 = ~\pi101 & w18610 ;
  assign w18612 = ~w18025 & w18353 ;
  assign w18613 = w18354 ^ w18612 ;
  assign w18614 = ~w18443 & w18613 ;
  assign w18615 = ( w18017 & w18441 ) | ( w18017 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18616 = ~w18442 & w18615 ;
  assign w18617 = w18614 | w18616 ;
  assign w18618 = ~\pi100 & w18617 ;
  assign w18619 = ~w18032 & w18350 ;
  assign w18620 = w18351 ^ w18619 ;
  assign w18621 = ~w18443 & w18620 ;
  assign w18622 = ( w18024 & w18441 ) | ( w18024 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18623 = ~w18442 & w18622 ;
  assign w18624 = w18621 | w18623 ;
  assign w18625 = ~\pi099 & w18624 ;
  assign w18626 = ~w18039 & w18347 ;
  assign w18627 = w18348 ^ w18626 ;
  assign w18628 = ~w18443 & w18627 ;
  assign w18629 = ( w18031 & w18441 ) | ( w18031 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18630 = ~w18442 & w18629 ;
  assign w18631 = w18628 | w18630 ;
  assign w18632 = ~\pi098 & w18631 ;
  assign w18633 = ~w18046 & w18344 ;
  assign w18634 = w18345 ^ w18633 ;
  assign w18635 = ~w18443 & w18634 ;
  assign w18636 = ( w18038 & w18441 ) | ( w18038 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18637 = ~w18442 & w18636 ;
  assign w18638 = w18635 | w18637 ;
  assign w18639 = ~\pi097 & w18638 ;
  assign w18640 = ~w18053 & w18341 ;
  assign w18641 = w18342 ^ w18640 ;
  assign w18642 = ~w18443 & w18641 ;
  assign w18643 = ( w18045 & w18441 ) | ( w18045 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18644 = ~w18442 & w18643 ;
  assign w18645 = w18642 | w18644 ;
  assign w18646 = ~\pi096 & w18645 ;
  assign w18647 = ~w18060 & w18338 ;
  assign w18648 = w18339 ^ w18647 ;
  assign w18649 = ~w18443 & w18648 ;
  assign w18650 = ( w18052 & w18441 ) | ( w18052 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18651 = ~w18442 & w18650 ;
  assign w18652 = w18649 | w18651 ;
  assign w18653 = ~\pi095 & w18652 ;
  assign w18654 = ~w18067 & w18335 ;
  assign w18655 = w18336 ^ w18654 ;
  assign w18656 = ~w18443 & w18655 ;
  assign w18657 = ( w18059 & w18441 ) | ( w18059 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18658 = ~w18442 & w18657 ;
  assign w18659 = w18656 | w18658 ;
  assign w18660 = ~\pi094 & w18659 ;
  assign w18661 = ~w18074 & w18332 ;
  assign w18662 = w18333 ^ w18661 ;
  assign w18663 = ~w18443 & w18662 ;
  assign w18664 = ( w18066 & w18441 ) | ( w18066 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18665 = ~w18442 & w18664 ;
  assign w18666 = w18663 | w18665 ;
  assign w18667 = ~\pi093 & w18666 ;
  assign w18668 = ~w18081 & w18329 ;
  assign w18669 = w18330 ^ w18668 ;
  assign w18670 = ~w18443 & w18669 ;
  assign w18671 = ( w18073 & w18441 ) | ( w18073 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18672 = ~w18442 & w18671 ;
  assign w18673 = w18670 | w18672 ;
  assign w18674 = ~\pi092 & w18673 ;
  assign w18675 = ~w18088 & w18326 ;
  assign w18676 = w18327 ^ w18675 ;
  assign w18677 = ~w18443 & w18676 ;
  assign w18678 = ( w18080 & w18441 ) | ( w18080 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18679 = ~w18442 & w18678 ;
  assign w18680 = w18677 | w18679 ;
  assign w18681 = ~\pi091 & w18680 ;
  assign w18682 = ~w18095 & w18323 ;
  assign w18683 = w18324 ^ w18682 ;
  assign w18684 = ~w18443 & w18683 ;
  assign w18685 = ( w18087 & w18441 ) | ( w18087 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18686 = ~w18442 & w18685 ;
  assign w18687 = w18684 | w18686 ;
  assign w18688 = ~\pi090 & w18687 ;
  assign w18689 = ~w18102 & w18320 ;
  assign w18690 = w18321 ^ w18689 ;
  assign w18691 = ~w18443 & w18690 ;
  assign w18692 = ( w18094 & w18441 ) | ( w18094 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18693 = ~w18442 & w18692 ;
  assign w18694 = w18691 | w18693 ;
  assign w18695 = ~\pi089 & w18694 ;
  assign w18696 = ~w18109 & w18317 ;
  assign w18697 = w18318 ^ w18696 ;
  assign w18698 = ~w18443 & w18697 ;
  assign w18699 = ( w18101 & w18441 ) | ( w18101 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18700 = ~w18442 & w18699 ;
  assign w18701 = w18698 | w18700 ;
  assign w18702 = ~\pi088 & w18701 ;
  assign w18703 = ~w18116 & w18314 ;
  assign w18704 = w18315 ^ w18703 ;
  assign w18705 = ~w18443 & w18704 ;
  assign w18706 = ( w18108 & w18441 ) | ( w18108 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18707 = ~w18442 & w18706 ;
  assign w18708 = w18705 | w18707 ;
  assign w18709 = ~\pi087 & w18708 ;
  assign w18710 = ~w18123 & w18311 ;
  assign w18711 = w18312 ^ w18710 ;
  assign w18712 = ~w18443 & w18711 ;
  assign w18713 = ( w18115 & w18441 ) | ( w18115 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18714 = ~w18442 & w18713 ;
  assign w18715 = w18712 | w18714 ;
  assign w18716 = ~\pi086 & w18715 ;
  assign w18717 = ~w18130 & w18308 ;
  assign w18718 = w18309 ^ w18717 ;
  assign w18719 = ~w18443 & w18718 ;
  assign w18720 = ( w18122 & w18441 ) | ( w18122 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18721 = ~w18442 & w18720 ;
  assign w18722 = w18719 | w18721 ;
  assign w18723 = ~\pi085 & w18722 ;
  assign w18724 = ~w18137 & w18305 ;
  assign w18725 = w18306 ^ w18724 ;
  assign w18726 = ~w18443 & w18725 ;
  assign w18727 = ( w18129 & w18441 ) | ( w18129 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18728 = ~w18442 & w18727 ;
  assign w18729 = w18726 | w18728 ;
  assign w18730 = ~\pi084 & w18729 ;
  assign w18731 = ~w18144 & w18302 ;
  assign w18732 = w18303 ^ w18731 ;
  assign w18733 = ~w18443 & w18732 ;
  assign w18734 = ( w18136 & w18441 ) | ( w18136 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18735 = ~w18442 & w18734 ;
  assign w18736 = w18733 | w18735 ;
  assign w18737 = ~\pi083 & w18736 ;
  assign w18738 = ~w18151 & w18299 ;
  assign w18739 = w18300 ^ w18738 ;
  assign w18740 = ~w18443 & w18739 ;
  assign w18741 = ( w18143 & w18441 ) | ( w18143 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18742 = ~w18442 & w18741 ;
  assign w18743 = w18740 | w18742 ;
  assign w18744 = ~\pi082 & w18743 ;
  assign w18745 = ~w18158 & w18296 ;
  assign w18746 = w18297 ^ w18745 ;
  assign w18747 = ~w18443 & w18746 ;
  assign w18748 = ( w18150 & w18441 ) | ( w18150 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18749 = ~w18442 & w18748 ;
  assign w18750 = w18747 | w18749 ;
  assign w18751 = ~\pi081 & w18750 ;
  assign w18752 = ~w18165 & w18293 ;
  assign w18753 = w18294 ^ w18752 ;
  assign w18754 = ~w18443 & w18753 ;
  assign w18755 = ( w18157 & w18441 ) | ( w18157 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18756 = ~w18442 & w18755 ;
  assign w18757 = w18754 | w18756 ;
  assign w18758 = ~\pi080 & w18757 ;
  assign w18759 = ~w18172 & w18290 ;
  assign w18760 = w18291 ^ w18759 ;
  assign w18761 = ~w18443 & w18760 ;
  assign w18762 = ( w18164 & w18441 ) | ( w18164 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18763 = ~w18442 & w18762 ;
  assign w18764 = w18761 | w18763 ;
  assign w18765 = ~\pi079 & w18764 ;
  assign w18766 = ~w18179 & w18287 ;
  assign w18767 = w18288 ^ w18766 ;
  assign w18768 = ~w18443 & w18767 ;
  assign w18769 = ( w18171 & w18441 ) | ( w18171 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18770 = ~w18442 & w18769 ;
  assign w18771 = w18768 | w18770 ;
  assign w18772 = ~\pi078 & w18771 ;
  assign w18773 = ~w18186 & w18284 ;
  assign w18774 = w18285 ^ w18773 ;
  assign w18775 = ~w18443 & w18774 ;
  assign w18776 = ( w18178 & w18441 ) | ( w18178 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18777 = ~w18442 & w18776 ;
  assign w18778 = w18775 | w18777 ;
  assign w18779 = ~\pi077 & w18778 ;
  assign w18780 = ~w18193 & w18281 ;
  assign w18781 = w18282 ^ w18780 ;
  assign w18782 = ~w18443 & w18781 ;
  assign w18783 = ( w18185 & w18441 ) | ( w18185 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18784 = ~w18442 & w18783 ;
  assign w18785 = w18782 | w18784 ;
  assign w18786 = ~\pi076 & w18785 ;
  assign w18787 = ~w18200 & w18278 ;
  assign w18788 = w18279 ^ w18787 ;
  assign w18789 = ~w18443 & w18788 ;
  assign w18790 = ( w18192 & w18441 ) | ( w18192 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18791 = ~w18442 & w18790 ;
  assign w18792 = w18789 | w18791 ;
  assign w18793 = ~\pi075 & w18792 ;
  assign w18794 = ~w18207 & w18275 ;
  assign w18795 = w18276 ^ w18794 ;
  assign w18796 = ~w18443 & w18795 ;
  assign w18797 = ( w18199 & w18441 ) | ( w18199 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18798 = ~w18442 & w18797 ;
  assign w18799 = w18796 | w18798 ;
  assign w18800 = ~\pi074 & w18799 ;
  assign w18801 = ~w18214 & w18272 ;
  assign w18802 = w18273 ^ w18801 ;
  assign w18803 = ~w18443 & w18802 ;
  assign w18804 = ( w18206 & w18441 ) | ( w18206 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18805 = ~w18442 & w18804 ;
  assign w18806 = w18803 | w18805 ;
  assign w18807 = ~\pi073 & w18806 ;
  assign w18808 = ~w18221 & w18269 ;
  assign w18809 = w18270 ^ w18808 ;
  assign w18810 = ~w18443 & w18809 ;
  assign w18811 = ( w18213 & w18441 ) | ( w18213 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18812 = ~w18442 & w18811 ;
  assign w18813 = w18810 | w18812 ;
  assign w18814 = ~\pi072 & w18813 ;
  assign w18815 = ~w18228 & w18266 ;
  assign w18816 = w18267 ^ w18815 ;
  assign w18817 = ~w18443 & w18816 ;
  assign w18818 = ( w18220 & w18441 ) | ( w18220 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18819 = ~w18442 & w18818 ;
  assign w18820 = w18817 | w18819 ;
  assign w18821 = ~\pi071 & w18820 ;
  assign w18822 = ~w18235 & w18263 ;
  assign w18823 = w18264 ^ w18822 ;
  assign w18824 = ~w18443 & w18823 ;
  assign w18825 = ( w18227 & w18441 ) | ( w18227 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18826 = ~w18442 & w18825 ;
  assign w18827 = w18824 | w18826 ;
  assign w18828 = ~\pi070 & w18827 ;
  assign w18829 = ~w18243 & w18260 ;
  assign w18830 = w18261 ^ w18829 ;
  assign w18831 = ~w18443 & w18830 ;
  assign w18832 = ( w18234 & w18441 ) | ( w18234 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18833 = ~w18442 & w18832 ;
  assign w18834 = w18831 | w18833 ;
  assign w18835 = ~\pi069 & w18834 ;
  assign w18836 = ~w18251 & w18257 ;
  assign w18837 = w18258 ^ w18836 ;
  assign w18838 = ~w18443 & w18837 ;
  assign w18839 = ( w18242 & w18441 ) | ( w18242 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18840 = ~w18442 & w18839 ;
  assign w18841 = w18838 | w18840 ;
  assign w18842 = ~\pi068 & w18841 ;
  assign w18843 = ~\pi003 & \pi064 ;
  assign w18844 = ( \pi065 & ~w18254 ) | ( \pi065 & w18843 ) | ( ~w18254 & w18843 ) ;
  assign w18845 = w18252 ^ w18844 ;
  assign w18846 = ~w18443 & w18845 ;
  assign w18847 = ( w18250 & w18441 ) | ( w18250 & w18442 ) | ( w18441 & w18442 ) ;
  assign w18848 = ~w18442 & w18847 ;
  assign w18849 = w18846 | w18848 ;
  assign w18850 = ~\pi067 & w18849 ;
  assign w18851 = \pi004 ^ \pi065 ;
  assign w18852 = \pi003 ^ w17843 ;
  assign w18853 = ( \pi064 & w18443 ) | ( \pi064 & w18852 ) | ( w18443 & w18852 ) ;
  assign w18854 = w18851 ^ w18853 ;
  assign w18855 = ~w18443 & w18854 ;
  assign w18856 = w18254 & w18443 ;
  assign w18857 = w18855 | w18856 ;
  assign w18858 = ~\pi066 & w18857 ;
  assign w18859 = \pi066 ^ w18857 ;
  assign w18860 = \pi064 & ~w18443 ;
  assign w18861 = \pi003 ^ w18860 ;
  assign w18862 = ( ~\pi002 & \pi064 ) | ( ~\pi002 & w18859 ) | ( \pi064 & w18859 ) ;
  assign w18863 = ( \pi065 & ~w18861 ) | ( \pi065 & w18862 ) | ( ~w18861 & w18862 ) ;
  assign w18864 = w18859 | w18863 ;
  assign w18865 = \pi067 ^ w18849 ;
  assign w18866 = ( ~w18858 & w18864 ) | ( ~w18858 & w18865 ) | ( w18864 & w18865 ) ;
  assign w18867 = w18865 | w18866 ;
  assign w18868 = \pi068 ^ w18841 ;
  assign w18869 = ( ~w18850 & w18867 ) | ( ~w18850 & w18868 ) | ( w18867 & w18868 ) ;
  assign w18870 = w18868 | w18869 ;
  assign w18871 = \pi069 ^ w18834 ;
  assign w18872 = ( ~w18842 & w18870 ) | ( ~w18842 & w18871 ) | ( w18870 & w18871 ) ;
  assign w18873 = w18871 | w18872 ;
  assign w18874 = \pi070 ^ w18827 ;
  assign w18875 = ( ~w18835 & w18873 ) | ( ~w18835 & w18874 ) | ( w18873 & w18874 ) ;
  assign w18876 = w18874 | w18875 ;
  assign w18877 = \pi071 ^ w18820 ;
  assign w18878 = ( ~w18828 & w18876 ) | ( ~w18828 & w18877 ) | ( w18876 & w18877 ) ;
  assign w18879 = w18877 | w18878 ;
  assign w18880 = \pi072 ^ w18813 ;
  assign w18881 = ( ~w18821 & w18879 ) | ( ~w18821 & w18880 ) | ( w18879 & w18880 ) ;
  assign w18882 = w18880 | w18881 ;
  assign w18883 = \pi073 ^ w18806 ;
  assign w18884 = ( ~w18814 & w18882 ) | ( ~w18814 & w18883 ) | ( w18882 & w18883 ) ;
  assign w18885 = w18883 | w18884 ;
  assign w18886 = \pi074 ^ w18799 ;
  assign w18887 = ( ~w18807 & w18885 ) | ( ~w18807 & w18886 ) | ( w18885 & w18886 ) ;
  assign w18888 = w18886 | w18887 ;
  assign w18889 = \pi075 ^ w18792 ;
  assign w18890 = ( ~w18800 & w18888 ) | ( ~w18800 & w18889 ) | ( w18888 & w18889 ) ;
  assign w18891 = w18889 | w18890 ;
  assign w18892 = \pi076 ^ w18785 ;
  assign w18893 = ( ~w18793 & w18891 ) | ( ~w18793 & w18892 ) | ( w18891 & w18892 ) ;
  assign w18894 = w18892 | w18893 ;
  assign w18895 = \pi077 ^ w18778 ;
  assign w18896 = ( ~w18786 & w18894 ) | ( ~w18786 & w18895 ) | ( w18894 & w18895 ) ;
  assign w18897 = w18895 | w18896 ;
  assign w18898 = \pi078 ^ w18771 ;
  assign w18899 = ( ~w18779 & w18897 ) | ( ~w18779 & w18898 ) | ( w18897 & w18898 ) ;
  assign w18900 = w18898 | w18899 ;
  assign w18901 = \pi079 ^ w18764 ;
  assign w18902 = ( ~w18772 & w18900 ) | ( ~w18772 & w18901 ) | ( w18900 & w18901 ) ;
  assign w18903 = w18901 | w18902 ;
  assign w18904 = \pi080 ^ w18757 ;
  assign w18905 = ( ~w18765 & w18903 ) | ( ~w18765 & w18904 ) | ( w18903 & w18904 ) ;
  assign w18906 = w18904 | w18905 ;
  assign w18907 = \pi081 ^ w18750 ;
  assign w18908 = ( ~w18758 & w18906 ) | ( ~w18758 & w18907 ) | ( w18906 & w18907 ) ;
  assign w18909 = w18907 | w18908 ;
  assign w18910 = \pi082 ^ w18743 ;
  assign w18911 = ( ~w18751 & w18909 ) | ( ~w18751 & w18910 ) | ( w18909 & w18910 ) ;
  assign w18912 = w18910 | w18911 ;
  assign w18913 = \pi083 ^ w18736 ;
  assign w18914 = ( ~w18744 & w18912 ) | ( ~w18744 & w18913 ) | ( w18912 & w18913 ) ;
  assign w18915 = w18913 | w18914 ;
  assign w18916 = \pi084 ^ w18729 ;
  assign w18917 = ( ~w18737 & w18915 ) | ( ~w18737 & w18916 ) | ( w18915 & w18916 ) ;
  assign w18918 = w18916 | w18917 ;
  assign w18919 = \pi085 ^ w18722 ;
  assign w18920 = ( ~w18730 & w18918 ) | ( ~w18730 & w18919 ) | ( w18918 & w18919 ) ;
  assign w18921 = w18919 | w18920 ;
  assign w18922 = \pi086 ^ w18715 ;
  assign w18923 = ( ~w18723 & w18921 ) | ( ~w18723 & w18922 ) | ( w18921 & w18922 ) ;
  assign w18924 = w18922 | w18923 ;
  assign w18925 = \pi087 ^ w18708 ;
  assign w18926 = ( ~w18716 & w18924 ) | ( ~w18716 & w18925 ) | ( w18924 & w18925 ) ;
  assign w18927 = w18925 | w18926 ;
  assign w18928 = \pi088 ^ w18701 ;
  assign w18929 = ( ~w18709 & w18927 ) | ( ~w18709 & w18928 ) | ( w18927 & w18928 ) ;
  assign w18930 = w18928 | w18929 ;
  assign w18931 = \pi089 ^ w18694 ;
  assign w18932 = ( ~w18702 & w18930 ) | ( ~w18702 & w18931 ) | ( w18930 & w18931 ) ;
  assign w18933 = w18931 | w18932 ;
  assign w18934 = \pi090 ^ w18687 ;
  assign w18935 = ( ~w18695 & w18933 ) | ( ~w18695 & w18934 ) | ( w18933 & w18934 ) ;
  assign w18936 = w18934 | w18935 ;
  assign w18937 = \pi091 ^ w18680 ;
  assign w18938 = ( ~w18688 & w18936 ) | ( ~w18688 & w18937 ) | ( w18936 & w18937 ) ;
  assign w18939 = w18937 | w18938 ;
  assign w18940 = \pi092 ^ w18673 ;
  assign w18941 = ( ~w18681 & w18939 ) | ( ~w18681 & w18940 ) | ( w18939 & w18940 ) ;
  assign w18942 = w18940 | w18941 ;
  assign w18943 = \pi093 ^ w18666 ;
  assign w18944 = ( ~w18674 & w18942 ) | ( ~w18674 & w18943 ) | ( w18942 & w18943 ) ;
  assign w18945 = w18943 | w18944 ;
  assign w18946 = \pi094 ^ w18659 ;
  assign w18947 = ( ~w18667 & w18945 ) | ( ~w18667 & w18946 ) | ( w18945 & w18946 ) ;
  assign w18948 = w18946 | w18947 ;
  assign w18949 = \pi095 ^ w18652 ;
  assign w18950 = ( ~w18660 & w18948 ) | ( ~w18660 & w18949 ) | ( w18948 & w18949 ) ;
  assign w18951 = w18949 | w18950 ;
  assign w18952 = \pi096 ^ w18645 ;
  assign w18953 = ( ~w18653 & w18951 ) | ( ~w18653 & w18952 ) | ( w18951 & w18952 ) ;
  assign w18954 = w18952 | w18953 ;
  assign w18955 = \pi097 ^ w18638 ;
  assign w18956 = ( ~w18646 & w18954 ) | ( ~w18646 & w18955 ) | ( w18954 & w18955 ) ;
  assign w18957 = w18955 | w18956 ;
  assign w18958 = \pi098 ^ w18631 ;
  assign w18959 = ( ~w18639 & w18957 ) | ( ~w18639 & w18958 ) | ( w18957 & w18958 ) ;
  assign w18960 = w18958 | w18959 ;
  assign w18961 = \pi099 ^ w18624 ;
  assign w18962 = ( ~w18632 & w18960 ) | ( ~w18632 & w18961 ) | ( w18960 & w18961 ) ;
  assign w18963 = w18961 | w18962 ;
  assign w18964 = \pi100 ^ w18617 ;
  assign w18965 = ( ~w18625 & w18963 ) | ( ~w18625 & w18964 ) | ( w18963 & w18964 ) ;
  assign w18966 = w18964 | w18965 ;
  assign w18967 = \pi101 ^ w18610 ;
  assign w18968 = ( ~w18618 & w18966 ) | ( ~w18618 & w18967 ) | ( w18966 & w18967 ) ;
  assign w18969 = w18967 | w18968 ;
  assign w18970 = \pi102 ^ w18603 ;
  assign w18971 = ( ~w18611 & w18969 ) | ( ~w18611 & w18970 ) | ( w18969 & w18970 ) ;
  assign w18972 = w18970 | w18971 ;
  assign w18973 = \pi103 ^ w18596 ;
  assign w18974 = ( ~w18604 & w18972 ) | ( ~w18604 & w18973 ) | ( w18972 & w18973 ) ;
  assign w18975 = w18973 | w18974 ;
  assign w18976 = \pi104 ^ w18589 ;
  assign w18977 = ( ~w18597 & w18975 ) | ( ~w18597 & w18976 ) | ( w18975 & w18976 ) ;
  assign w18978 = w18976 | w18977 ;
  assign w18979 = \pi105 ^ w18582 ;
  assign w18980 = ( ~w18590 & w18978 ) | ( ~w18590 & w18979 ) | ( w18978 & w18979 ) ;
  assign w18981 = w18979 | w18980 ;
  assign w18982 = \pi106 ^ w18575 ;
  assign w18983 = ( ~w18583 & w18981 ) | ( ~w18583 & w18982 ) | ( w18981 & w18982 ) ;
  assign w18984 = w18982 | w18983 ;
  assign w18985 = \pi107 ^ w18568 ;
  assign w18986 = ( ~w18576 & w18984 ) | ( ~w18576 & w18985 ) | ( w18984 & w18985 ) ;
  assign w18987 = w18985 | w18986 ;
  assign w18988 = \pi108 ^ w18561 ;
  assign w18989 = ( ~w18569 & w18987 ) | ( ~w18569 & w18988 ) | ( w18987 & w18988 ) ;
  assign w18990 = w18988 | w18989 ;
  assign w18991 = \pi109 ^ w18554 ;
  assign w18992 = ( ~w18562 & w18990 ) | ( ~w18562 & w18991 ) | ( w18990 & w18991 ) ;
  assign w18993 = w18991 | w18992 ;
  assign w18994 = \pi110 ^ w18547 ;
  assign w18995 = ( ~w18555 & w18993 ) | ( ~w18555 & w18994 ) | ( w18993 & w18994 ) ;
  assign w18996 = w18994 | w18995 ;
  assign w18997 = \pi111 ^ w18540 ;
  assign w18998 = ( ~w18548 & w18996 ) | ( ~w18548 & w18997 ) | ( w18996 & w18997 ) ;
  assign w18999 = w18997 | w18998 ;
  assign w19000 = \pi112 ^ w18533 ;
  assign w19001 = ( ~w18541 & w18999 ) | ( ~w18541 & w19000 ) | ( w18999 & w19000 ) ;
  assign w19002 = w19000 | w19001 ;
  assign w19003 = \pi113 ^ w18526 ;
  assign w19004 = ( ~w18534 & w19002 ) | ( ~w18534 & w19003 ) | ( w19002 & w19003 ) ;
  assign w19005 = w19003 | w19004 ;
  assign w19006 = \pi114 ^ w18519 ;
  assign w19007 = ( ~w18527 & w19005 ) | ( ~w18527 & w19006 ) | ( w19005 & w19006 ) ;
  assign w19008 = w19006 | w19007 ;
  assign w19009 = \pi115 ^ w18512 ;
  assign w19010 = ( ~w18520 & w19008 ) | ( ~w18520 & w19009 ) | ( w19008 & w19009 ) ;
  assign w19011 = w19009 | w19010 ;
  assign w19012 = \pi116 ^ w18505 ;
  assign w19013 = ( ~w18513 & w19011 ) | ( ~w18513 & w19012 ) | ( w19011 & w19012 ) ;
  assign w19014 = w19012 | w19013 ;
  assign w19015 = \pi117 ^ w18498 ;
  assign w19016 = ( ~w18506 & w19014 ) | ( ~w18506 & w19015 ) | ( w19014 & w19015 ) ;
  assign w19017 = w19015 | w19016 ;
  assign w19018 = \pi118 ^ w18491 ;
  assign w19019 = ( ~w18499 & w19017 ) | ( ~w18499 & w19018 ) | ( w19017 & w19018 ) ;
  assign w19020 = w19018 | w19019 ;
  assign w19021 = \pi119 ^ w18484 ;
  assign w19022 = ( ~w18492 & w19020 ) | ( ~w18492 & w19021 ) | ( w19020 & w19021 ) ;
  assign w19023 = w19021 | w19022 ;
  assign w19024 = \pi120 ^ w18477 ;
  assign w19025 = ( ~w18485 & w19023 ) | ( ~w18485 & w19024 ) | ( w19023 & w19024 ) ;
  assign w19026 = w19024 | w19025 ;
  assign w19027 = \pi121 ^ w18470 ;
  assign w19028 = ( ~w18478 & w19026 ) | ( ~w18478 & w19027 ) | ( w19026 & w19027 ) ;
  assign w19029 = w19027 | w19028 ;
  assign w19030 = \pi122 ^ w18463 ;
  assign w19031 = ( ~w18471 & w19029 ) | ( ~w18471 & w19030 ) | ( w19029 & w19030 ) ;
  assign w19032 = w19030 | w19031 ;
  assign w19033 = \pi123 ^ w18456 ;
  assign w19034 = ( ~w18464 & w19032 ) | ( ~w18464 & w19033 ) | ( w19032 & w19033 ) ;
  assign w19035 = w19033 | w19034 ;
  assign w19036 = \pi124 ^ w18449 ;
  assign w19037 = ( ~w18457 & w19035 ) | ( ~w18457 & w19036 ) | ( w19035 & w19036 ) ;
  assign w19038 = w19036 | w19037 ;
  assign w19039 = ( ~w17850 & w18428 ) | ( ~w17850 & w18443 ) | ( w18428 & w18443 ) ;
  assign w19040 = w18438 ^ w19039 ;
  assign w19041 = ~w18443 & w19040 ;
  assign w19042 = ( w147 & ~w18434 ) | ( w147 & w18441 ) | ( ~w18434 & w18441 ) ;
  assign w19043 = w18434 & w19042 ;
  assign w19044 = w19041 | w19043 ;
  assign w19045 = ~\pi125 & w19044 ;
  assign w19046 = ( \pi125 & ~w19041 ) | ( \pi125 & w19043 ) | ( ~w19041 & w19043 ) ;
  assign w19047 = ~w19043 & w19046 ;
  assign w19048 = ( ~w18450 & w19038 ) | ( ~w18450 & w19045 ) | ( w19038 & w19045 ) ;
  assign w19049 = ( \pi127 & w19045 ) | ( \pi127 & ~w19048 ) | ( w19045 & ~w19048 ) ;
  assign w19050 = ( \pi126 & w19047 ) | ( \pi126 & ~w19048 ) | ( w19047 & ~w19048 ) ;
  assign w19051 = ( w19048 & ~w19049 ) | ( w19048 & w19050 ) | ( ~w19049 & w19050 ) ;
  assign w19052 = w19049 | w19051 ;
  assign w19053 = ~w269 & w19044 ;
  assign w19054 = w19052 & ~w19053 ;
  assign w19055 = ~w18457 & w19035 ;
  assign w19056 = w19036 ^ w19055 ;
  assign w19057 = ~w19054 & w19056 ;
  assign w19058 = ( w18449 & w19052 ) | ( w18449 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19059 = ~w19053 & w19058 ;
  assign w19060 = w19057 | w19059 ;
  assign w19061 = ~\pi125 & w19060 ;
  assign w19062 = ~w18464 & w19032 ;
  assign w19063 = w19033 ^ w19062 ;
  assign w19064 = ~w19054 & w19063 ;
  assign w19065 = ( w18456 & w19052 ) | ( w18456 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19066 = ~w19053 & w19065 ;
  assign w19067 = w19064 | w19066 ;
  assign w19068 = ~\pi124 & w19067 ;
  assign w19069 = ~w18471 & w19029 ;
  assign w19070 = w19030 ^ w19069 ;
  assign w19071 = ~w19054 & w19070 ;
  assign w19072 = ( w18463 & w19052 ) | ( w18463 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19073 = ~w19053 & w19072 ;
  assign w19074 = w19071 | w19073 ;
  assign w19075 = ~\pi123 & w19074 ;
  assign w19076 = ~w18478 & w19026 ;
  assign w19077 = w19027 ^ w19076 ;
  assign w19078 = ~w19054 & w19077 ;
  assign w19079 = ( w18470 & w19052 ) | ( w18470 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19080 = ~w19053 & w19079 ;
  assign w19081 = w19078 | w19080 ;
  assign w19082 = ~\pi122 & w19081 ;
  assign w19083 = ~w18485 & w19023 ;
  assign w19084 = w19024 ^ w19083 ;
  assign w19085 = ~w19054 & w19084 ;
  assign w19086 = ( w18477 & w19052 ) | ( w18477 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19087 = ~w19053 & w19086 ;
  assign w19088 = w19085 | w19087 ;
  assign w19089 = ~\pi121 & w19088 ;
  assign w19090 = ~w18492 & w19020 ;
  assign w19091 = w19021 ^ w19090 ;
  assign w19092 = ~w19054 & w19091 ;
  assign w19093 = ( w18484 & w19052 ) | ( w18484 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19094 = ~w19053 & w19093 ;
  assign w19095 = w19092 | w19094 ;
  assign w19096 = ~\pi120 & w19095 ;
  assign w19097 = ~w18499 & w19017 ;
  assign w19098 = w19018 ^ w19097 ;
  assign w19099 = ~w19054 & w19098 ;
  assign w19100 = ( w18491 & w19052 ) | ( w18491 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19101 = ~w19053 & w19100 ;
  assign w19102 = w19099 | w19101 ;
  assign w19103 = ~\pi119 & w19102 ;
  assign w19104 = ~w18506 & w19014 ;
  assign w19105 = w19015 ^ w19104 ;
  assign w19106 = ~w19054 & w19105 ;
  assign w19107 = ( w18498 & w19052 ) | ( w18498 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19108 = ~w19053 & w19107 ;
  assign w19109 = w19106 | w19108 ;
  assign w19110 = ~\pi118 & w19109 ;
  assign w19111 = ~w18513 & w19011 ;
  assign w19112 = w19012 ^ w19111 ;
  assign w19113 = ~w19054 & w19112 ;
  assign w19114 = ( w18505 & w19052 ) | ( w18505 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19115 = ~w19053 & w19114 ;
  assign w19116 = w19113 | w19115 ;
  assign w19117 = ~\pi117 & w19116 ;
  assign w19118 = ~w18520 & w19008 ;
  assign w19119 = w19009 ^ w19118 ;
  assign w19120 = ~w19054 & w19119 ;
  assign w19121 = ( w18512 & w19052 ) | ( w18512 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19122 = ~w19053 & w19121 ;
  assign w19123 = w19120 | w19122 ;
  assign w19124 = ~\pi116 & w19123 ;
  assign w19125 = ~w18527 & w19005 ;
  assign w19126 = w19006 ^ w19125 ;
  assign w19127 = ~w19054 & w19126 ;
  assign w19128 = ( w18519 & w19052 ) | ( w18519 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19129 = ~w19053 & w19128 ;
  assign w19130 = w19127 | w19129 ;
  assign w19131 = ~\pi115 & w19130 ;
  assign w19132 = ~w18534 & w19002 ;
  assign w19133 = w19003 ^ w19132 ;
  assign w19134 = ~w19054 & w19133 ;
  assign w19135 = ( w18526 & w19052 ) | ( w18526 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19136 = ~w19053 & w19135 ;
  assign w19137 = w19134 | w19136 ;
  assign w19138 = ~\pi114 & w19137 ;
  assign w19139 = ~w18541 & w18999 ;
  assign w19140 = w19000 ^ w19139 ;
  assign w19141 = ~w19054 & w19140 ;
  assign w19142 = ( w18533 & w19052 ) | ( w18533 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19143 = ~w19053 & w19142 ;
  assign w19144 = w19141 | w19143 ;
  assign w19145 = ~\pi113 & w19144 ;
  assign w19146 = ~w18548 & w18996 ;
  assign w19147 = w18997 ^ w19146 ;
  assign w19148 = ~w19054 & w19147 ;
  assign w19149 = ( w18540 & w19052 ) | ( w18540 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19150 = ~w19053 & w19149 ;
  assign w19151 = w19148 | w19150 ;
  assign w19152 = ~\pi112 & w19151 ;
  assign w19153 = ~w18555 & w18993 ;
  assign w19154 = w18994 ^ w19153 ;
  assign w19155 = ~w19054 & w19154 ;
  assign w19156 = ( w18547 & w19052 ) | ( w18547 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19157 = ~w19053 & w19156 ;
  assign w19158 = w19155 | w19157 ;
  assign w19159 = ~\pi111 & w19158 ;
  assign w19160 = ~w18562 & w18990 ;
  assign w19161 = w18991 ^ w19160 ;
  assign w19162 = ~w19054 & w19161 ;
  assign w19163 = ( w18554 & w19052 ) | ( w18554 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19164 = ~w19053 & w19163 ;
  assign w19165 = w19162 | w19164 ;
  assign w19166 = ~\pi110 & w19165 ;
  assign w19167 = ~w18569 & w18987 ;
  assign w19168 = w18988 ^ w19167 ;
  assign w19169 = ~w19054 & w19168 ;
  assign w19170 = ( w18561 & w19052 ) | ( w18561 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19171 = ~w19053 & w19170 ;
  assign w19172 = w19169 | w19171 ;
  assign w19173 = ~\pi109 & w19172 ;
  assign w19174 = ~w18576 & w18984 ;
  assign w19175 = w18985 ^ w19174 ;
  assign w19176 = ~w19054 & w19175 ;
  assign w19177 = ( w18568 & w19052 ) | ( w18568 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19178 = ~w19053 & w19177 ;
  assign w19179 = w19176 | w19178 ;
  assign w19180 = ~\pi108 & w19179 ;
  assign w19181 = ~w18583 & w18981 ;
  assign w19182 = w18982 ^ w19181 ;
  assign w19183 = ~w19054 & w19182 ;
  assign w19184 = ( w18575 & w19052 ) | ( w18575 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19185 = ~w19053 & w19184 ;
  assign w19186 = w19183 | w19185 ;
  assign w19187 = ~\pi107 & w19186 ;
  assign w19188 = ~w18590 & w18978 ;
  assign w19189 = w18979 ^ w19188 ;
  assign w19190 = ~w19054 & w19189 ;
  assign w19191 = ( w18582 & w19052 ) | ( w18582 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19192 = ~w19053 & w19191 ;
  assign w19193 = w19190 | w19192 ;
  assign w19194 = ~\pi106 & w19193 ;
  assign w19195 = ~w18597 & w18975 ;
  assign w19196 = w18976 ^ w19195 ;
  assign w19197 = ~w19054 & w19196 ;
  assign w19198 = ( w18589 & w19052 ) | ( w18589 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19199 = ~w19053 & w19198 ;
  assign w19200 = w19197 | w19199 ;
  assign w19201 = ~\pi105 & w19200 ;
  assign w19202 = ~w18604 & w18972 ;
  assign w19203 = w18973 ^ w19202 ;
  assign w19204 = ~w19054 & w19203 ;
  assign w19205 = ( w18596 & w19052 ) | ( w18596 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19206 = ~w19053 & w19205 ;
  assign w19207 = w19204 | w19206 ;
  assign w19208 = ~\pi104 & w19207 ;
  assign w19209 = ~w18611 & w18969 ;
  assign w19210 = w18970 ^ w19209 ;
  assign w19211 = ~w19054 & w19210 ;
  assign w19212 = ( w18603 & w19052 ) | ( w18603 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19213 = ~w19053 & w19212 ;
  assign w19214 = w19211 | w19213 ;
  assign w19215 = ~\pi103 & w19214 ;
  assign w19216 = ~w18618 & w18966 ;
  assign w19217 = w18967 ^ w19216 ;
  assign w19218 = ~w19054 & w19217 ;
  assign w19219 = ( w18610 & w19052 ) | ( w18610 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19220 = ~w19053 & w19219 ;
  assign w19221 = w19218 | w19220 ;
  assign w19222 = ~\pi102 & w19221 ;
  assign w19223 = ~w18625 & w18963 ;
  assign w19224 = w18964 ^ w19223 ;
  assign w19225 = ~w19054 & w19224 ;
  assign w19226 = ( w18617 & w19052 ) | ( w18617 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19227 = ~w19053 & w19226 ;
  assign w19228 = w19225 | w19227 ;
  assign w19229 = ~\pi101 & w19228 ;
  assign w19230 = ~w18632 & w18960 ;
  assign w19231 = w18961 ^ w19230 ;
  assign w19232 = ~w19054 & w19231 ;
  assign w19233 = ( w18624 & w19052 ) | ( w18624 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19234 = ~w19053 & w19233 ;
  assign w19235 = w19232 | w19234 ;
  assign w19236 = ~\pi100 & w19235 ;
  assign w19237 = ~w18639 & w18957 ;
  assign w19238 = w18958 ^ w19237 ;
  assign w19239 = ~w19054 & w19238 ;
  assign w19240 = ( w18631 & w19052 ) | ( w18631 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19241 = ~w19053 & w19240 ;
  assign w19242 = w19239 | w19241 ;
  assign w19243 = ~\pi099 & w19242 ;
  assign w19244 = ~w18646 & w18954 ;
  assign w19245 = w18955 ^ w19244 ;
  assign w19246 = ~w19054 & w19245 ;
  assign w19247 = ( w18638 & w19052 ) | ( w18638 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19248 = ~w19053 & w19247 ;
  assign w19249 = w19246 | w19248 ;
  assign w19250 = ~\pi098 & w19249 ;
  assign w19251 = ~w18653 & w18951 ;
  assign w19252 = w18952 ^ w19251 ;
  assign w19253 = ~w19054 & w19252 ;
  assign w19254 = ( w18645 & w19052 ) | ( w18645 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19255 = ~w19053 & w19254 ;
  assign w19256 = w19253 | w19255 ;
  assign w19257 = ~\pi097 & w19256 ;
  assign w19258 = ~w18660 & w18948 ;
  assign w19259 = w18949 ^ w19258 ;
  assign w19260 = ~w19054 & w19259 ;
  assign w19261 = ( w18652 & w19052 ) | ( w18652 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19262 = ~w19053 & w19261 ;
  assign w19263 = w19260 | w19262 ;
  assign w19264 = ~\pi096 & w19263 ;
  assign w19265 = ~w18667 & w18945 ;
  assign w19266 = w18946 ^ w19265 ;
  assign w19267 = ~w19054 & w19266 ;
  assign w19268 = ( w18659 & w19052 ) | ( w18659 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19269 = ~w19053 & w19268 ;
  assign w19270 = w19267 | w19269 ;
  assign w19271 = ~\pi095 & w19270 ;
  assign w19272 = ~w18674 & w18942 ;
  assign w19273 = w18943 ^ w19272 ;
  assign w19274 = ~w19054 & w19273 ;
  assign w19275 = ( w18666 & w19052 ) | ( w18666 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19276 = ~w19053 & w19275 ;
  assign w19277 = w19274 | w19276 ;
  assign w19278 = ~\pi094 & w19277 ;
  assign w19279 = ~w18681 & w18939 ;
  assign w19280 = w18940 ^ w19279 ;
  assign w19281 = ~w19054 & w19280 ;
  assign w19282 = ( w18673 & w19052 ) | ( w18673 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19283 = ~w19053 & w19282 ;
  assign w19284 = w19281 | w19283 ;
  assign w19285 = ~\pi093 & w19284 ;
  assign w19286 = ~w18688 & w18936 ;
  assign w19287 = w18937 ^ w19286 ;
  assign w19288 = ~w19054 & w19287 ;
  assign w19289 = ( w18680 & w19052 ) | ( w18680 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19290 = ~w19053 & w19289 ;
  assign w19291 = w19288 | w19290 ;
  assign w19292 = ~\pi092 & w19291 ;
  assign w19293 = ~w18695 & w18933 ;
  assign w19294 = w18934 ^ w19293 ;
  assign w19295 = ~w19054 & w19294 ;
  assign w19296 = ( w18687 & w19052 ) | ( w18687 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19297 = ~w19053 & w19296 ;
  assign w19298 = w19295 | w19297 ;
  assign w19299 = ~\pi091 & w19298 ;
  assign w19300 = ~w18702 & w18930 ;
  assign w19301 = w18931 ^ w19300 ;
  assign w19302 = ~w19054 & w19301 ;
  assign w19303 = ( w18694 & w19052 ) | ( w18694 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19304 = ~w19053 & w19303 ;
  assign w19305 = w19302 | w19304 ;
  assign w19306 = ~\pi090 & w19305 ;
  assign w19307 = ~w18709 & w18927 ;
  assign w19308 = w18928 ^ w19307 ;
  assign w19309 = ~w19054 & w19308 ;
  assign w19310 = ( w18701 & w19052 ) | ( w18701 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19311 = ~w19053 & w19310 ;
  assign w19312 = w19309 | w19311 ;
  assign w19313 = ~\pi089 & w19312 ;
  assign w19314 = ~w18716 & w18924 ;
  assign w19315 = w18925 ^ w19314 ;
  assign w19316 = ~w19054 & w19315 ;
  assign w19317 = ( w18708 & w19052 ) | ( w18708 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19318 = ~w19053 & w19317 ;
  assign w19319 = w19316 | w19318 ;
  assign w19320 = ~\pi088 & w19319 ;
  assign w19321 = ~w18723 & w18921 ;
  assign w19322 = w18922 ^ w19321 ;
  assign w19323 = ~w19054 & w19322 ;
  assign w19324 = ( w18715 & w19052 ) | ( w18715 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19325 = ~w19053 & w19324 ;
  assign w19326 = w19323 | w19325 ;
  assign w19327 = ~\pi087 & w19326 ;
  assign w19328 = ~w18730 & w18918 ;
  assign w19329 = w18919 ^ w19328 ;
  assign w19330 = ~w19054 & w19329 ;
  assign w19331 = ( w18722 & w19052 ) | ( w18722 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19332 = ~w19053 & w19331 ;
  assign w19333 = w19330 | w19332 ;
  assign w19334 = ~\pi086 & w19333 ;
  assign w19335 = ~w18737 & w18915 ;
  assign w19336 = w18916 ^ w19335 ;
  assign w19337 = ~w19054 & w19336 ;
  assign w19338 = ( w18729 & w19052 ) | ( w18729 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19339 = ~w19053 & w19338 ;
  assign w19340 = w19337 | w19339 ;
  assign w19341 = ~\pi085 & w19340 ;
  assign w19342 = ~w18744 & w18912 ;
  assign w19343 = w18913 ^ w19342 ;
  assign w19344 = ~w19054 & w19343 ;
  assign w19345 = ( w18736 & w19052 ) | ( w18736 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19346 = ~w19053 & w19345 ;
  assign w19347 = w19344 | w19346 ;
  assign w19348 = ~\pi084 & w19347 ;
  assign w19349 = ~w18751 & w18909 ;
  assign w19350 = w18910 ^ w19349 ;
  assign w19351 = ~w19054 & w19350 ;
  assign w19352 = ( w18743 & w19052 ) | ( w18743 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19353 = ~w19053 & w19352 ;
  assign w19354 = w19351 | w19353 ;
  assign w19355 = ~\pi083 & w19354 ;
  assign w19356 = ~w18758 & w18906 ;
  assign w19357 = w18907 ^ w19356 ;
  assign w19358 = ~w19054 & w19357 ;
  assign w19359 = ( w18750 & w19052 ) | ( w18750 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19360 = ~w19053 & w19359 ;
  assign w19361 = w19358 | w19360 ;
  assign w19362 = ~\pi082 & w19361 ;
  assign w19363 = ~w18765 & w18903 ;
  assign w19364 = w18904 ^ w19363 ;
  assign w19365 = ~w19054 & w19364 ;
  assign w19366 = ( w18757 & w19052 ) | ( w18757 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19367 = ~w19053 & w19366 ;
  assign w19368 = w19365 | w19367 ;
  assign w19369 = ~\pi081 & w19368 ;
  assign w19370 = ~w18772 & w18900 ;
  assign w19371 = w18901 ^ w19370 ;
  assign w19372 = ~w19054 & w19371 ;
  assign w19373 = ( w18764 & w19052 ) | ( w18764 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19374 = ~w19053 & w19373 ;
  assign w19375 = w19372 | w19374 ;
  assign w19376 = ~\pi080 & w19375 ;
  assign w19377 = ~w18779 & w18897 ;
  assign w19378 = w18898 ^ w19377 ;
  assign w19379 = ~w19054 & w19378 ;
  assign w19380 = ( w18771 & w19052 ) | ( w18771 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19381 = ~w19053 & w19380 ;
  assign w19382 = w19379 | w19381 ;
  assign w19383 = ~\pi079 & w19382 ;
  assign w19384 = ~w18786 & w18894 ;
  assign w19385 = w18895 ^ w19384 ;
  assign w19386 = ~w19054 & w19385 ;
  assign w19387 = ( w18778 & w19052 ) | ( w18778 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19388 = ~w19053 & w19387 ;
  assign w19389 = w19386 | w19388 ;
  assign w19390 = ~\pi078 & w19389 ;
  assign w19391 = ~w18793 & w18891 ;
  assign w19392 = w18892 ^ w19391 ;
  assign w19393 = ~w19054 & w19392 ;
  assign w19394 = ( w18785 & w19052 ) | ( w18785 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19395 = ~w19053 & w19394 ;
  assign w19396 = w19393 | w19395 ;
  assign w19397 = ~\pi077 & w19396 ;
  assign w19398 = ~w18800 & w18888 ;
  assign w19399 = w18889 ^ w19398 ;
  assign w19400 = ~w19054 & w19399 ;
  assign w19401 = ( w18792 & w19052 ) | ( w18792 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19402 = ~w19053 & w19401 ;
  assign w19403 = w19400 | w19402 ;
  assign w19404 = ~\pi076 & w19403 ;
  assign w19405 = ~w18807 & w18885 ;
  assign w19406 = w18886 ^ w19405 ;
  assign w19407 = ~w19054 & w19406 ;
  assign w19408 = ( w18799 & w19052 ) | ( w18799 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19409 = ~w19053 & w19408 ;
  assign w19410 = w19407 | w19409 ;
  assign w19411 = ~\pi075 & w19410 ;
  assign w19412 = ~w18814 & w18882 ;
  assign w19413 = w18883 ^ w19412 ;
  assign w19414 = ~w19054 & w19413 ;
  assign w19415 = ( w18806 & w19052 ) | ( w18806 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19416 = ~w19053 & w19415 ;
  assign w19417 = w19414 | w19416 ;
  assign w19418 = ~\pi074 & w19417 ;
  assign w19419 = ~w18821 & w18879 ;
  assign w19420 = w18880 ^ w19419 ;
  assign w19421 = ~w19054 & w19420 ;
  assign w19422 = ( w18813 & w19052 ) | ( w18813 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19423 = ~w19053 & w19422 ;
  assign w19424 = w19421 | w19423 ;
  assign w19425 = ~\pi073 & w19424 ;
  assign w19426 = ~w18828 & w18876 ;
  assign w19427 = w18877 ^ w19426 ;
  assign w19428 = ~w19054 & w19427 ;
  assign w19429 = ( w18820 & w19052 ) | ( w18820 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19430 = ~w19053 & w19429 ;
  assign w19431 = w19428 | w19430 ;
  assign w19432 = ~\pi072 & w19431 ;
  assign w19433 = ~w18835 & w18873 ;
  assign w19434 = w18874 ^ w19433 ;
  assign w19435 = ~w19054 & w19434 ;
  assign w19436 = ( w18827 & w19052 ) | ( w18827 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19437 = ~w19053 & w19436 ;
  assign w19438 = w19435 | w19437 ;
  assign w19439 = ~\pi071 & w19438 ;
  assign w19440 = ~w18842 & w18870 ;
  assign w19441 = w18871 ^ w19440 ;
  assign w19442 = ~w19054 & w19441 ;
  assign w19443 = ( w18834 & w19052 ) | ( w18834 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19444 = ~w19053 & w19443 ;
  assign w19445 = w19442 | w19444 ;
  assign w19446 = ~\pi070 & w19445 ;
  assign w19447 = ~w18850 & w18867 ;
  assign w19448 = w18868 ^ w19447 ;
  assign w19449 = ~w19054 & w19448 ;
  assign w19450 = ( w18841 & w19052 ) | ( w18841 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19451 = ~w19053 & w19450 ;
  assign w19452 = w19449 | w19451 ;
  assign w19453 = ~\pi069 & w19452 ;
  assign w19454 = ~w18858 & w18864 ;
  assign w19455 = w18865 ^ w19454 ;
  assign w19456 = ~w19054 & w19455 ;
  assign w19457 = ( w18849 & w19052 ) | ( w18849 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19458 = ~w19053 & w19457 ;
  assign w19459 = w19456 | w19458 ;
  assign w19460 = ~\pi068 & w19459 ;
  assign w19461 = ~\pi002 & \pi064 ;
  assign w19462 = ( \pi065 & ~w18861 ) | ( \pi065 & w19461 ) | ( ~w18861 & w19461 ) ;
  assign w19463 = w18859 ^ w19462 ;
  assign w19464 = ~w19054 & w19463 ;
  assign w19465 = ( w18857 & w19052 ) | ( w18857 & w19053 ) | ( w19052 & w19053 ) ;
  assign w19466 = ~w19053 & w19465 ;
  assign w19467 = w19464 | w19466 ;
  assign w19468 = ~\pi067 & w19467 ;
  assign w19469 = \pi003 ^ \pi065 ;
  assign w19470 = \pi002 ^ w18443 ;
  assign w19471 = ( \pi064 & w19054 ) | ( \pi064 & w19470 ) | ( w19054 & w19470 ) ;
  assign w19472 = w19469 ^ w19471 ;
  assign w19473 = ~w19054 & w19472 ;
  assign w19474 = w18861 & w19054 ;
  assign w19475 = w19473 | w19474 ;
  assign w19476 = ~\pi066 & w19475 ;
  assign w19477 = \pi066 ^ w19475 ;
  assign w19478 = \pi064 & ~w19054 ;
  assign w19479 = \pi002 ^ w19478 ;
  assign w19480 = ( ~\pi001 & \pi064 ) | ( ~\pi001 & w19477 ) | ( \pi064 & w19477 ) ;
  assign w19481 = ( \pi065 & ~w19479 ) | ( \pi065 & w19480 ) | ( ~w19479 & w19480 ) ;
  assign w19482 = w19477 | w19481 ;
  assign w19483 = \pi067 ^ w19467 ;
  assign w19484 = ( ~w19476 & w19482 ) | ( ~w19476 & w19483 ) | ( w19482 & w19483 ) ;
  assign w19485 = w19483 | w19484 ;
  assign w19486 = \pi068 ^ w19459 ;
  assign w19487 = ( ~w19468 & w19485 ) | ( ~w19468 & w19486 ) | ( w19485 & w19486 ) ;
  assign w19488 = w19486 | w19487 ;
  assign w19489 = \pi069 ^ w19452 ;
  assign w19490 = ( ~w19460 & w19488 ) | ( ~w19460 & w19489 ) | ( w19488 & w19489 ) ;
  assign w19491 = w19489 | w19490 ;
  assign w19492 = \pi070 ^ w19445 ;
  assign w19493 = ( ~w19453 & w19491 ) | ( ~w19453 & w19492 ) | ( w19491 & w19492 ) ;
  assign w19494 = w19492 | w19493 ;
  assign w19495 = \pi071 ^ w19438 ;
  assign w19496 = ( ~w19446 & w19494 ) | ( ~w19446 & w19495 ) | ( w19494 & w19495 ) ;
  assign w19497 = w19495 | w19496 ;
  assign w19498 = \pi072 ^ w19431 ;
  assign w19499 = ( ~w19439 & w19497 ) | ( ~w19439 & w19498 ) | ( w19497 & w19498 ) ;
  assign w19500 = w19498 | w19499 ;
  assign w19501 = \pi073 ^ w19424 ;
  assign w19502 = ( ~w19432 & w19500 ) | ( ~w19432 & w19501 ) | ( w19500 & w19501 ) ;
  assign w19503 = w19501 | w19502 ;
  assign w19504 = \pi074 ^ w19417 ;
  assign w19505 = ( ~w19425 & w19503 ) | ( ~w19425 & w19504 ) | ( w19503 & w19504 ) ;
  assign w19506 = w19504 | w19505 ;
  assign w19507 = \pi075 ^ w19410 ;
  assign w19508 = ( ~w19418 & w19506 ) | ( ~w19418 & w19507 ) | ( w19506 & w19507 ) ;
  assign w19509 = w19507 | w19508 ;
  assign w19510 = \pi076 ^ w19403 ;
  assign w19511 = ( ~w19411 & w19509 ) | ( ~w19411 & w19510 ) | ( w19509 & w19510 ) ;
  assign w19512 = w19510 | w19511 ;
  assign w19513 = \pi077 ^ w19396 ;
  assign w19514 = ( ~w19404 & w19512 ) | ( ~w19404 & w19513 ) | ( w19512 & w19513 ) ;
  assign w19515 = w19513 | w19514 ;
  assign w19516 = \pi078 ^ w19389 ;
  assign w19517 = ( ~w19397 & w19515 ) | ( ~w19397 & w19516 ) | ( w19515 & w19516 ) ;
  assign w19518 = w19516 | w19517 ;
  assign w19519 = \pi079 ^ w19382 ;
  assign w19520 = ( ~w19390 & w19518 ) | ( ~w19390 & w19519 ) | ( w19518 & w19519 ) ;
  assign w19521 = w19519 | w19520 ;
  assign w19522 = \pi080 ^ w19375 ;
  assign w19523 = ( ~w19383 & w19521 ) | ( ~w19383 & w19522 ) | ( w19521 & w19522 ) ;
  assign w19524 = w19522 | w19523 ;
  assign w19525 = \pi081 ^ w19368 ;
  assign w19526 = ( ~w19376 & w19524 ) | ( ~w19376 & w19525 ) | ( w19524 & w19525 ) ;
  assign w19527 = w19525 | w19526 ;
  assign w19528 = \pi082 ^ w19361 ;
  assign w19529 = ( ~w19369 & w19527 ) | ( ~w19369 & w19528 ) | ( w19527 & w19528 ) ;
  assign w19530 = w19528 | w19529 ;
  assign w19531 = \pi083 ^ w19354 ;
  assign w19532 = ( ~w19362 & w19530 ) | ( ~w19362 & w19531 ) | ( w19530 & w19531 ) ;
  assign w19533 = w19531 | w19532 ;
  assign w19534 = \pi084 ^ w19347 ;
  assign w19535 = ( ~w19355 & w19533 ) | ( ~w19355 & w19534 ) | ( w19533 & w19534 ) ;
  assign w19536 = w19534 | w19535 ;
  assign w19537 = \pi085 ^ w19340 ;
  assign w19538 = ( ~w19348 & w19536 ) | ( ~w19348 & w19537 ) | ( w19536 & w19537 ) ;
  assign w19539 = w19537 | w19538 ;
  assign w19540 = \pi086 ^ w19333 ;
  assign w19541 = ( ~w19341 & w19539 ) | ( ~w19341 & w19540 ) | ( w19539 & w19540 ) ;
  assign w19542 = w19540 | w19541 ;
  assign w19543 = \pi087 ^ w19326 ;
  assign w19544 = ( ~w19334 & w19542 ) | ( ~w19334 & w19543 ) | ( w19542 & w19543 ) ;
  assign w19545 = w19543 | w19544 ;
  assign w19546 = \pi088 ^ w19319 ;
  assign w19547 = ( ~w19327 & w19545 ) | ( ~w19327 & w19546 ) | ( w19545 & w19546 ) ;
  assign w19548 = w19546 | w19547 ;
  assign w19549 = \pi089 ^ w19312 ;
  assign w19550 = ( ~w19320 & w19548 ) | ( ~w19320 & w19549 ) | ( w19548 & w19549 ) ;
  assign w19551 = w19549 | w19550 ;
  assign w19552 = \pi090 ^ w19305 ;
  assign w19553 = ( ~w19313 & w19551 ) | ( ~w19313 & w19552 ) | ( w19551 & w19552 ) ;
  assign w19554 = w19552 | w19553 ;
  assign w19555 = \pi091 ^ w19298 ;
  assign w19556 = ( ~w19306 & w19554 ) | ( ~w19306 & w19555 ) | ( w19554 & w19555 ) ;
  assign w19557 = w19555 | w19556 ;
  assign w19558 = \pi092 ^ w19291 ;
  assign w19559 = ( ~w19299 & w19557 ) | ( ~w19299 & w19558 ) | ( w19557 & w19558 ) ;
  assign w19560 = w19558 | w19559 ;
  assign w19561 = \pi093 ^ w19284 ;
  assign w19562 = ( ~w19292 & w19560 ) | ( ~w19292 & w19561 ) | ( w19560 & w19561 ) ;
  assign w19563 = w19561 | w19562 ;
  assign w19564 = \pi094 ^ w19277 ;
  assign w19565 = ( ~w19285 & w19563 ) | ( ~w19285 & w19564 ) | ( w19563 & w19564 ) ;
  assign w19566 = w19564 | w19565 ;
  assign w19567 = \pi095 ^ w19270 ;
  assign w19568 = ( ~w19278 & w19566 ) | ( ~w19278 & w19567 ) | ( w19566 & w19567 ) ;
  assign w19569 = w19567 | w19568 ;
  assign w19570 = \pi096 ^ w19263 ;
  assign w19571 = ( ~w19271 & w19569 ) | ( ~w19271 & w19570 ) | ( w19569 & w19570 ) ;
  assign w19572 = w19570 | w19571 ;
  assign w19573 = \pi097 ^ w19256 ;
  assign w19574 = ( ~w19264 & w19572 ) | ( ~w19264 & w19573 ) | ( w19572 & w19573 ) ;
  assign w19575 = w19573 | w19574 ;
  assign w19576 = \pi098 ^ w19249 ;
  assign w19577 = ( ~w19257 & w19575 ) | ( ~w19257 & w19576 ) | ( w19575 & w19576 ) ;
  assign w19578 = w19576 | w19577 ;
  assign w19579 = \pi099 ^ w19242 ;
  assign w19580 = ( ~w19250 & w19578 ) | ( ~w19250 & w19579 ) | ( w19578 & w19579 ) ;
  assign w19581 = w19579 | w19580 ;
  assign w19582 = \pi100 ^ w19235 ;
  assign w19583 = ( ~w19243 & w19581 ) | ( ~w19243 & w19582 ) | ( w19581 & w19582 ) ;
  assign w19584 = w19582 | w19583 ;
  assign w19585 = \pi101 ^ w19228 ;
  assign w19586 = ( ~w19236 & w19584 ) | ( ~w19236 & w19585 ) | ( w19584 & w19585 ) ;
  assign w19587 = w19585 | w19586 ;
  assign w19588 = \pi102 ^ w19221 ;
  assign w19589 = ( ~w19229 & w19587 ) | ( ~w19229 & w19588 ) | ( w19587 & w19588 ) ;
  assign w19590 = w19588 | w19589 ;
  assign w19591 = \pi103 ^ w19214 ;
  assign w19592 = ( ~w19222 & w19590 ) | ( ~w19222 & w19591 ) | ( w19590 & w19591 ) ;
  assign w19593 = w19591 | w19592 ;
  assign w19594 = \pi104 ^ w19207 ;
  assign w19595 = ( ~w19215 & w19593 ) | ( ~w19215 & w19594 ) | ( w19593 & w19594 ) ;
  assign w19596 = w19594 | w19595 ;
  assign w19597 = \pi105 ^ w19200 ;
  assign w19598 = ( ~w19208 & w19596 ) | ( ~w19208 & w19597 ) | ( w19596 & w19597 ) ;
  assign w19599 = w19597 | w19598 ;
  assign w19600 = \pi106 ^ w19193 ;
  assign w19601 = ( ~w19201 & w19599 ) | ( ~w19201 & w19600 ) | ( w19599 & w19600 ) ;
  assign w19602 = w19600 | w19601 ;
  assign w19603 = \pi107 ^ w19186 ;
  assign w19604 = ( ~w19194 & w19602 ) | ( ~w19194 & w19603 ) | ( w19602 & w19603 ) ;
  assign w19605 = w19603 | w19604 ;
  assign w19606 = \pi108 ^ w19179 ;
  assign w19607 = ( ~w19187 & w19605 ) | ( ~w19187 & w19606 ) | ( w19605 & w19606 ) ;
  assign w19608 = w19606 | w19607 ;
  assign w19609 = \pi109 ^ w19172 ;
  assign w19610 = ( ~w19180 & w19608 ) | ( ~w19180 & w19609 ) | ( w19608 & w19609 ) ;
  assign w19611 = w19609 | w19610 ;
  assign w19612 = \pi110 ^ w19165 ;
  assign w19613 = ( ~w19173 & w19611 ) | ( ~w19173 & w19612 ) | ( w19611 & w19612 ) ;
  assign w19614 = w19612 | w19613 ;
  assign w19615 = \pi111 ^ w19158 ;
  assign w19616 = ( ~w19166 & w19614 ) | ( ~w19166 & w19615 ) | ( w19614 & w19615 ) ;
  assign w19617 = w19615 | w19616 ;
  assign w19618 = \pi112 ^ w19151 ;
  assign w19619 = ( ~w19159 & w19617 ) | ( ~w19159 & w19618 ) | ( w19617 & w19618 ) ;
  assign w19620 = w19618 | w19619 ;
  assign w19621 = \pi113 ^ w19144 ;
  assign w19622 = ( ~w19152 & w19620 ) | ( ~w19152 & w19621 ) | ( w19620 & w19621 ) ;
  assign w19623 = w19621 | w19622 ;
  assign w19624 = \pi114 ^ w19137 ;
  assign w19625 = ( ~w19145 & w19623 ) | ( ~w19145 & w19624 ) | ( w19623 & w19624 ) ;
  assign w19626 = w19624 | w19625 ;
  assign w19627 = \pi115 ^ w19130 ;
  assign w19628 = ( ~w19138 & w19626 ) | ( ~w19138 & w19627 ) | ( w19626 & w19627 ) ;
  assign w19629 = w19627 | w19628 ;
  assign w19630 = \pi116 ^ w19123 ;
  assign w19631 = ( ~w19131 & w19629 ) | ( ~w19131 & w19630 ) | ( w19629 & w19630 ) ;
  assign w19632 = w19630 | w19631 ;
  assign w19633 = \pi117 ^ w19116 ;
  assign w19634 = ( ~w19124 & w19632 ) | ( ~w19124 & w19633 ) | ( w19632 & w19633 ) ;
  assign w19635 = w19633 | w19634 ;
  assign w19636 = \pi118 ^ w19109 ;
  assign w19637 = ( ~w19117 & w19635 ) | ( ~w19117 & w19636 ) | ( w19635 & w19636 ) ;
  assign w19638 = w19636 | w19637 ;
  assign w19639 = \pi119 ^ w19102 ;
  assign w19640 = ( ~w19110 & w19638 ) | ( ~w19110 & w19639 ) | ( w19638 & w19639 ) ;
  assign w19641 = w19639 | w19640 ;
  assign w19642 = \pi120 ^ w19095 ;
  assign w19643 = ( ~w19103 & w19641 ) | ( ~w19103 & w19642 ) | ( w19641 & w19642 ) ;
  assign w19644 = w19642 | w19643 ;
  assign w19645 = \pi121 ^ w19088 ;
  assign w19646 = ( ~w19096 & w19644 ) | ( ~w19096 & w19645 ) | ( w19644 & w19645 ) ;
  assign w19647 = w19645 | w19646 ;
  assign w19648 = \pi122 ^ w19081 ;
  assign w19649 = ( ~w19089 & w19647 ) | ( ~w19089 & w19648 ) | ( w19647 & w19648 ) ;
  assign w19650 = w19648 | w19649 ;
  assign w19651 = \pi123 ^ w19074 ;
  assign w19652 = ( ~w19082 & w19650 ) | ( ~w19082 & w19651 ) | ( w19650 & w19651 ) ;
  assign w19653 = w19651 | w19652 ;
  assign w19654 = \pi124 ^ w19067 ;
  assign w19655 = ( ~w19075 & w19653 ) | ( ~w19075 & w19654 ) | ( w19653 & w19654 ) ;
  assign w19656 = w19654 | w19655 ;
  assign w19657 = \pi125 ^ w19060 ;
  assign w19658 = ( ~w19068 & w19656 ) | ( ~w19068 & w19657 ) | ( w19656 & w19657 ) ;
  assign w19659 = w19657 | w19658 ;
  assign w19660 = w19045 | w19047 ;
  assign w19661 = ( ~w18450 & w19038 ) | ( ~w18450 & w19054 ) | ( w19038 & w19054 ) ;
  assign w19662 = w19660 ^ w19661 ;
  assign w19663 = ~w19054 & w19662 ;
  assign w19664 = ( w269 & ~w19044 ) | ( w269 & w19052 ) | ( ~w19044 & w19052 ) ;
  assign w19665 = w19044 & w19664 ;
  assign w19666 = ( ~\pi127 & w19663 ) | ( ~\pi127 & w19665 ) | ( w19663 & w19665 ) ;
  assign w19667 = \pi126 ^ w19666 ;
  assign w19668 = ( w19061 & w19659 ) | ( w19061 & ~w19667 ) | ( w19659 & ~w19667 ) ;
  assign w19669 = ( \pi127 & ~w19061 ) | ( \pi127 & w19668 ) | ( ~w19061 & w19668 ) ;
  assign w19670 = w19667 | w19669 ;
  assign w19671 = \pi126 | \pi127 ;
  assign w19672 = w19666 & ~w19671 ;
  assign w19673 = w19670 & ~w19672 ;
  assign w19674 = ~w19075 & w19653 ;
  assign w19675 = w19654 ^ w19674 ;
  assign w19676 = w19067 ^ w19673 ;
  assign w19677 = ( w19067 & w19675 ) | ( w19067 & ~w19676 ) | ( w19675 & ~w19676 ) ;
  assign w19678 = ~w19089 & w19647 ;
  assign w19679 = w19648 ^ w19678 ;
  assign w19680 = w19081 ^ w19673 ;
  assign w19681 = ( w19081 & w19679 ) | ( w19081 & ~w19680 ) | ( w19679 & ~w19680 ) ;
  assign w19682 = ~w19103 & w19641 ;
  assign w19683 = w19642 ^ w19682 ;
  assign w19684 = w19095 ^ w19673 ;
  assign w19685 = ( w19095 & w19683 ) | ( w19095 & ~w19684 ) | ( w19683 & ~w19684 ) ;
  assign w19686 = ~w19117 & w19635 ;
  assign w19687 = w19636 ^ w19686 ;
  assign w19688 = w19109 ^ w19673 ;
  assign w19689 = ( w19109 & w19687 ) | ( w19109 & ~w19688 ) | ( w19687 & ~w19688 ) ;
  assign w19690 = ~w19131 & w19629 ;
  assign w19691 = w19630 ^ w19690 ;
  assign w19692 = w19123 ^ w19673 ;
  assign w19693 = ( w19123 & w19691 ) | ( w19123 & ~w19692 ) | ( w19691 & ~w19692 ) ;
  assign w19694 = ~w19145 & w19623 ;
  assign w19695 = w19624 ^ w19694 ;
  assign w19696 = w19137 ^ w19673 ;
  assign w19697 = ( w19137 & w19695 ) | ( w19137 & ~w19696 ) | ( w19695 & ~w19696 ) ;
  assign w19698 = ~w19159 & w19617 ;
  assign w19699 = w19618 ^ w19698 ;
  assign w19700 = w19151 ^ w19673 ;
  assign w19701 = ( w19151 & w19699 ) | ( w19151 & ~w19700 ) | ( w19699 & ~w19700 ) ;
  assign w19702 = ~w19173 & w19611 ;
  assign w19703 = w19612 ^ w19702 ;
  assign w19704 = w19165 ^ w19673 ;
  assign w19705 = ( w19165 & w19703 ) | ( w19165 & ~w19704 ) | ( w19703 & ~w19704 ) ;
  assign w19706 = ~w19187 & w19605 ;
  assign w19707 = w19606 ^ w19706 ;
  assign w19708 = w19179 ^ w19673 ;
  assign w19709 = ( w19179 & w19707 ) | ( w19179 & ~w19708 ) | ( w19707 & ~w19708 ) ;
  assign w19710 = ~w19201 & w19599 ;
  assign w19711 = w19600 ^ w19710 ;
  assign w19712 = w19193 ^ w19673 ;
  assign w19713 = ( w19193 & w19711 ) | ( w19193 & ~w19712 ) | ( w19711 & ~w19712 ) ;
  assign w19714 = ~w19215 & w19593 ;
  assign w19715 = w19594 ^ w19714 ;
  assign w19716 = w19207 ^ w19673 ;
  assign w19717 = ( w19207 & w19715 ) | ( w19207 & ~w19716 ) | ( w19715 & ~w19716 ) ;
  assign w19718 = ~w19229 & w19587 ;
  assign w19719 = w19588 ^ w19718 ;
  assign w19720 = w19221 ^ w19673 ;
  assign w19721 = ( w19221 & w19719 ) | ( w19221 & ~w19720 ) | ( w19719 & ~w19720 ) ;
  assign w19722 = ~w19243 & w19581 ;
  assign w19723 = w19582 ^ w19722 ;
  assign w19724 = w19235 ^ w19673 ;
  assign w19725 = ( w19235 & w19723 ) | ( w19235 & ~w19724 ) | ( w19723 & ~w19724 ) ;
  assign w19726 = ~w19257 & w19575 ;
  assign w19727 = w19576 ^ w19726 ;
  assign w19728 = w19249 ^ w19673 ;
  assign w19729 = ( w19249 & w19727 ) | ( w19249 & ~w19728 ) | ( w19727 & ~w19728 ) ;
  assign w19730 = ~w19271 & w19569 ;
  assign w19731 = w19570 ^ w19730 ;
  assign w19732 = w19263 ^ w19673 ;
  assign w19733 = ( w19263 & w19731 ) | ( w19263 & ~w19732 ) | ( w19731 & ~w19732 ) ;
  assign w19734 = ~w19285 & w19563 ;
  assign w19735 = w19564 ^ w19734 ;
  assign w19736 = w19277 ^ w19673 ;
  assign w19737 = ( w19277 & w19735 ) | ( w19277 & ~w19736 ) | ( w19735 & ~w19736 ) ;
  assign w19738 = ~w19299 & w19557 ;
  assign w19739 = w19558 ^ w19738 ;
  assign w19740 = w19291 ^ w19673 ;
  assign w19741 = ( w19291 & w19739 ) | ( w19291 & ~w19740 ) | ( w19739 & ~w19740 ) ;
  assign w19742 = ~w19313 & w19551 ;
  assign w19743 = w19552 ^ w19742 ;
  assign w19744 = w19305 ^ w19673 ;
  assign w19745 = ( w19305 & w19743 ) | ( w19305 & ~w19744 ) | ( w19743 & ~w19744 ) ;
  assign w19746 = ~w19327 & w19545 ;
  assign w19747 = w19546 ^ w19746 ;
  assign w19748 = w19319 ^ w19673 ;
  assign w19749 = ( w19319 & w19747 ) | ( w19319 & ~w19748 ) | ( w19747 & ~w19748 ) ;
  assign w19750 = ~w19341 & w19539 ;
  assign w19751 = w19540 ^ w19750 ;
  assign w19752 = w19333 ^ w19673 ;
  assign w19753 = ( w19333 & w19751 ) | ( w19333 & ~w19752 ) | ( w19751 & ~w19752 ) ;
  assign w19754 = ~w19355 & w19533 ;
  assign w19755 = w19534 ^ w19754 ;
  assign w19756 = w19347 ^ w19673 ;
  assign w19757 = ( w19347 & w19755 ) | ( w19347 & ~w19756 ) | ( w19755 & ~w19756 ) ;
  assign w19758 = ~w19369 & w19527 ;
  assign w19759 = w19528 ^ w19758 ;
  assign w19760 = w19361 ^ w19673 ;
  assign w19761 = ( w19361 & w19759 ) | ( w19361 & ~w19760 ) | ( w19759 & ~w19760 ) ;
  assign w19762 = ~w19383 & w19521 ;
  assign w19763 = w19522 ^ w19762 ;
  assign w19764 = w19375 ^ w19673 ;
  assign w19765 = ( w19375 & w19763 ) | ( w19375 & ~w19764 ) | ( w19763 & ~w19764 ) ;
  assign w19766 = ~w19397 & w19515 ;
  assign w19767 = w19516 ^ w19766 ;
  assign w19768 = w19389 ^ w19673 ;
  assign w19769 = ( w19389 & w19767 ) | ( w19389 & ~w19768 ) | ( w19767 & ~w19768 ) ;
  assign w19770 = ~w19411 & w19509 ;
  assign w19771 = w19510 ^ w19770 ;
  assign w19772 = w19403 ^ w19673 ;
  assign w19773 = ( w19403 & w19771 ) | ( w19403 & ~w19772 ) | ( w19771 & ~w19772 ) ;
  assign w19774 = ~w19425 & w19503 ;
  assign w19775 = w19504 ^ w19774 ;
  assign w19776 = w19417 ^ w19673 ;
  assign w19777 = ( w19417 & w19775 ) | ( w19417 & ~w19776 ) | ( w19775 & ~w19776 ) ;
  assign w19778 = ~w19439 & w19497 ;
  assign w19779 = w19498 ^ w19778 ;
  assign w19780 = w19431 ^ w19673 ;
  assign w19781 = ( w19431 & w19779 ) | ( w19431 & ~w19780 ) | ( w19779 & ~w19780 ) ;
  assign w19782 = ~w19453 & w19491 ;
  assign w19783 = w19492 ^ w19782 ;
  assign w19784 = w19445 ^ w19673 ;
  assign w19785 = ( w19445 & w19783 ) | ( w19445 & ~w19784 ) | ( w19783 & ~w19784 ) ;
  assign w19786 = ~w19468 & w19485 ;
  assign w19787 = w19486 ^ w19786 ;
  assign w19788 = w19459 ^ w19673 ;
  assign w19789 = ( w19459 & w19787 ) | ( w19459 & ~w19788 ) | ( w19787 & ~w19788 ) ;
  assign w19790 = ~\pi001 & \pi064 ;
  assign w19791 = ( \pi065 & ~w19479 ) | ( \pi065 & w19790 ) | ( ~w19479 & w19790 ) ;
  assign w19792 = w19477 ^ w19791 ;
  assign w19793 = w19673 ^ w19792 ;
  assign w19794 = ( w19475 & w19792 ) | ( w19475 & w19793 ) | ( w19792 & w19793 ) ;
  assign w19795 = \pi002 ^ \pi065 ;
  assign w19796 = \pi001 ^ w19054 ;
  assign w19797 = \pi064 & w19796 ;
  assign w19798 = w19795 ^ w19797 ;
  assign w19799 = ( ~\pi064 & w19054 ) | ( ~\pi064 & w19670 ) | ( w19054 & w19670 ) ;
  assign w19800 = \pi002 ^ w19799 ;
  assign w19801 = w19673 ^ w19800 ;
  assign w19802 = ( w19798 & ~w19800 ) | ( w19798 & w19801 ) | ( ~w19800 & w19801 ) ;
  assign w19803 = ( \pi064 & ~w19673 ) | ( \pi064 & w19802 ) | ( ~w19673 & w19802 ) ;
  assign w19804 = \pi001 ^ w19803 ;
  assign w19805 = ~\pi000 & \pi064 ;
  assign w19806 = ( \pi065 & ~w19804 ) | ( \pi065 & w19805 ) | ( ~w19804 & w19805 ) ;
  assign w19807 = ~w19802 & w19806 ;
  assign w19808 = \pi066 | w19807 ;
  assign w19809 = \pi064 & ~w19673 ;
  assign w19810 = \pi001 ^ w19809 ;
  assign w19811 = ( \pi000 & ~\pi064 ) | ( \pi000 & w19802 ) | ( ~\pi064 & w19802 ) ;
  assign w19812 = ( ~\pi065 & w19810 ) | ( ~\pi065 & w19811 ) | ( w19810 & w19811 ) ;
  assign w19813 = w19802 & w19812 ;
  assign w19814 = ~w19476 & w19482 ;
  assign w19815 = w19483 ^ w19814 ;
  assign w19816 = w19467 ^ w19673 ;
  assign w19817 = ( w19467 & w19815 ) | ( w19467 & ~w19816 ) | ( w19815 & ~w19816 ) ;
  assign w19818 = ~\pi068 & w19817 ;
  assign w19819 = ( w19808 & ~w19813 ) | ( w19808 & w19818 ) | ( ~w19813 & w19818 ) ;
  assign w19820 = ( \pi067 & ~w19794 ) | ( \pi067 & w19819 ) | ( ~w19794 & w19819 ) ;
  assign w19821 = ( \pi068 & ~w19818 ) | ( \pi068 & w19820 ) | ( ~w19818 & w19820 ) ;
  assign w19822 = w19808 & ~w19813 ;
  assign w19823 = ( \pi067 & ~w19794 ) | ( \pi067 & w19822 ) | ( ~w19794 & w19822 ) ;
  assign w19824 = w19817 & ~w19823 ;
  assign w19825 = ~w19460 & w19488 ;
  assign w19826 = w19489 ^ w19825 ;
  assign w19827 = w19452 ^ w19673 ;
  assign w19828 = ( w19452 & w19826 ) | ( w19452 & ~w19827 ) | ( w19826 & ~w19827 ) ;
  assign w19829 = ~\pi070 & w19828 ;
  assign w19830 = ( w19821 & ~w19824 ) | ( w19821 & w19829 ) | ( ~w19824 & w19829 ) ;
  assign w19831 = ( \pi069 & ~w19789 ) | ( \pi069 & w19830 ) | ( ~w19789 & w19830 ) ;
  assign w19832 = ( \pi070 & ~w19829 ) | ( \pi070 & w19831 ) | ( ~w19829 & w19831 ) ;
  assign w19833 = w19821 & ~w19824 ;
  assign w19834 = ( \pi069 & ~w19789 ) | ( \pi069 & w19833 ) | ( ~w19789 & w19833 ) ;
  assign w19835 = w19828 & ~w19834 ;
  assign w19836 = ~w19446 & w19494 ;
  assign w19837 = w19495 ^ w19836 ;
  assign w19838 = w19438 ^ w19673 ;
  assign w19839 = ( w19438 & w19837 ) | ( w19438 & ~w19838 ) | ( w19837 & ~w19838 ) ;
  assign w19840 = ~\pi072 & w19839 ;
  assign w19841 = ( w19832 & ~w19835 ) | ( w19832 & w19840 ) | ( ~w19835 & w19840 ) ;
  assign w19842 = ( \pi071 & ~w19785 ) | ( \pi071 & w19841 ) | ( ~w19785 & w19841 ) ;
  assign w19843 = ( \pi072 & ~w19840 ) | ( \pi072 & w19842 ) | ( ~w19840 & w19842 ) ;
  assign w19844 = w19832 & ~w19835 ;
  assign w19845 = ( \pi071 & ~w19785 ) | ( \pi071 & w19844 ) | ( ~w19785 & w19844 ) ;
  assign w19846 = w19839 & ~w19845 ;
  assign w19847 = ~w19432 & w19500 ;
  assign w19848 = w19501 ^ w19847 ;
  assign w19849 = w19424 ^ w19673 ;
  assign w19850 = ( w19424 & w19848 ) | ( w19424 & ~w19849 ) | ( w19848 & ~w19849 ) ;
  assign w19851 = ~\pi074 & w19850 ;
  assign w19852 = ( w19843 & ~w19846 ) | ( w19843 & w19851 ) | ( ~w19846 & w19851 ) ;
  assign w19853 = ( \pi073 & ~w19781 ) | ( \pi073 & w19852 ) | ( ~w19781 & w19852 ) ;
  assign w19854 = ( \pi074 & ~w19851 ) | ( \pi074 & w19853 ) | ( ~w19851 & w19853 ) ;
  assign w19855 = w19843 & ~w19846 ;
  assign w19856 = ( \pi073 & ~w19781 ) | ( \pi073 & w19855 ) | ( ~w19781 & w19855 ) ;
  assign w19857 = w19850 & ~w19856 ;
  assign w19858 = ~w19418 & w19506 ;
  assign w19859 = w19507 ^ w19858 ;
  assign w19860 = w19410 ^ w19673 ;
  assign w19861 = ( w19410 & w19859 ) | ( w19410 & ~w19860 ) | ( w19859 & ~w19860 ) ;
  assign w19862 = ~\pi076 & w19861 ;
  assign w19863 = ( w19854 & ~w19857 ) | ( w19854 & w19862 ) | ( ~w19857 & w19862 ) ;
  assign w19864 = ( \pi075 & ~w19777 ) | ( \pi075 & w19863 ) | ( ~w19777 & w19863 ) ;
  assign w19865 = ( \pi076 & ~w19862 ) | ( \pi076 & w19864 ) | ( ~w19862 & w19864 ) ;
  assign w19866 = w19854 & ~w19857 ;
  assign w19867 = ( \pi075 & ~w19777 ) | ( \pi075 & w19866 ) | ( ~w19777 & w19866 ) ;
  assign w19868 = w19861 & ~w19867 ;
  assign w19869 = ~w19404 & w19512 ;
  assign w19870 = w19513 ^ w19869 ;
  assign w19871 = w19396 ^ w19673 ;
  assign w19872 = ( w19396 & w19870 ) | ( w19396 & ~w19871 ) | ( w19870 & ~w19871 ) ;
  assign w19873 = ~\pi078 & w19872 ;
  assign w19874 = ( w19865 & ~w19868 ) | ( w19865 & w19873 ) | ( ~w19868 & w19873 ) ;
  assign w19875 = ( \pi077 & ~w19773 ) | ( \pi077 & w19874 ) | ( ~w19773 & w19874 ) ;
  assign w19876 = ( \pi078 & ~w19873 ) | ( \pi078 & w19875 ) | ( ~w19873 & w19875 ) ;
  assign w19877 = w19865 & ~w19868 ;
  assign w19878 = ( \pi077 & ~w19773 ) | ( \pi077 & w19877 ) | ( ~w19773 & w19877 ) ;
  assign w19879 = w19872 & ~w19878 ;
  assign w19880 = ~w19390 & w19518 ;
  assign w19881 = w19519 ^ w19880 ;
  assign w19882 = w19382 ^ w19673 ;
  assign w19883 = ( w19382 & w19881 ) | ( w19382 & ~w19882 ) | ( w19881 & ~w19882 ) ;
  assign w19884 = ~\pi080 & w19883 ;
  assign w19885 = ( w19876 & ~w19879 ) | ( w19876 & w19884 ) | ( ~w19879 & w19884 ) ;
  assign w19886 = ( \pi079 & ~w19769 ) | ( \pi079 & w19885 ) | ( ~w19769 & w19885 ) ;
  assign w19887 = ( \pi080 & ~w19884 ) | ( \pi080 & w19886 ) | ( ~w19884 & w19886 ) ;
  assign w19888 = w19876 & ~w19879 ;
  assign w19889 = ( \pi079 & ~w19769 ) | ( \pi079 & w19888 ) | ( ~w19769 & w19888 ) ;
  assign w19890 = w19883 & ~w19889 ;
  assign w19891 = ~w19376 & w19524 ;
  assign w19892 = w19525 ^ w19891 ;
  assign w19893 = w19368 ^ w19673 ;
  assign w19894 = ( w19368 & w19892 ) | ( w19368 & ~w19893 ) | ( w19892 & ~w19893 ) ;
  assign w19895 = ~\pi082 & w19894 ;
  assign w19896 = ( w19887 & ~w19890 ) | ( w19887 & w19895 ) | ( ~w19890 & w19895 ) ;
  assign w19897 = ( \pi081 & ~w19765 ) | ( \pi081 & w19896 ) | ( ~w19765 & w19896 ) ;
  assign w19898 = ( \pi082 & ~w19895 ) | ( \pi082 & w19897 ) | ( ~w19895 & w19897 ) ;
  assign w19899 = w19887 & ~w19890 ;
  assign w19900 = ( \pi081 & ~w19765 ) | ( \pi081 & w19899 ) | ( ~w19765 & w19899 ) ;
  assign w19901 = w19894 & ~w19900 ;
  assign w19902 = ~w19362 & w19530 ;
  assign w19903 = w19531 ^ w19902 ;
  assign w19904 = w19354 ^ w19673 ;
  assign w19905 = ( w19354 & w19903 ) | ( w19354 & ~w19904 ) | ( w19903 & ~w19904 ) ;
  assign w19906 = ~\pi084 & w19905 ;
  assign w19907 = ( w19898 & ~w19901 ) | ( w19898 & w19906 ) | ( ~w19901 & w19906 ) ;
  assign w19908 = ( \pi083 & ~w19761 ) | ( \pi083 & w19907 ) | ( ~w19761 & w19907 ) ;
  assign w19909 = ( \pi084 & ~w19906 ) | ( \pi084 & w19908 ) | ( ~w19906 & w19908 ) ;
  assign w19910 = w19898 & ~w19901 ;
  assign w19911 = ( \pi083 & ~w19761 ) | ( \pi083 & w19910 ) | ( ~w19761 & w19910 ) ;
  assign w19912 = w19905 & ~w19911 ;
  assign w19913 = ~w19348 & w19536 ;
  assign w19914 = w19537 ^ w19913 ;
  assign w19915 = w19340 ^ w19673 ;
  assign w19916 = ( w19340 & w19914 ) | ( w19340 & ~w19915 ) | ( w19914 & ~w19915 ) ;
  assign w19917 = ~\pi086 & w19916 ;
  assign w19918 = ( w19909 & ~w19912 ) | ( w19909 & w19917 ) | ( ~w19912 & w19917 ) ;
  assign w19919 = ( \pi085 & ~w19757 ) | ( \pi085 & w19918 ) | ( ~w19757 & w19918 ) ;
  assign w19920 = ( \pi086 & ~w19917 ) | ( \pi086 & w19919 ) | ( ~w19917 & w19919 ) ;
  assign w19921 = w19909 & ~w19912 ;
  assign w19922 = ( \pi085 & ~w19757 ) | ( \pi085 & w19921 ) | ( ~w19757 & w19921 ) ;
  assign w19923 = w19916 & ~w19922 ;
  assign w19924 = ~w19334 & w19542 ;
  assign w19925 = w19543 ^ w19924 ;
  assign w19926 = w19326 ^ w19673 ;
  assign w19927 = ( w19326 & w19925 ) | ( w19326 & ~w19926 ) | ( w19925 & ~w19926 ) ;
  assign w19928 = ~\pi088 & w19927 ;
  assign w19929 = ( w19920 & ~w19923 ) | ( w19920 & w19928 ) | ( ~w19923 & w19928 ) ;
  assign w19930 = ( \pi087 & ~w19753 ) | ( \pi087 & w19929 ) | ( ~w19753 & w19929 ) ;
  assign w19931 = ( \pi088 & ~w19928 ) | ( \pi088 & w19930 ) | ( ~w19928 & w19930 ) ;
  assign w19932 = w19920 & ~w19923 ;
  assign w19933 = ( \pi087 & ~w19753 ) | ( \pi087 & w19932 ) | ( ~w19753 & w19932 ) ;
  assign w19934 = w19927 & ~w19933 ;
  assign w19935 = ~w19320 & w19548 ;
  assign w19936 = w19549 ^ w19935 ;
  assign w19937 = w19312 ^ w19673 ;
  assign w19938 = ( w19312 & w19936 ) | ( w19312 & ~w19937 ) | ( w19936 & ~w19937 ) ;
  assign w19939 = ~\pi090 & w19938 ;
  assign w19940 = ( w19931 & ~w19934 ) | ( w19931 & w19939 ) | ( ~w19934 & w19939 ) ;
  assign w19941 = ( \pi089 & ~w19749 ) | ( \pi089 & w19940 ) | ( ~w19749 & w19940 ) ;
  assign w19942 = ( \pi090 & ~w19939 ) | ( \pi090 & w19941 ) | ( ~w19939 & w19941 ) ;
  assign w19943 = w19931 & ~w19934 ;
  assign w19944 = ( \pi089 & ~w19749 ) | ( \pi089 & w19943 ) | ( ~w19749 & w19943 ) ;
  assign w19945 = w19938 & ~w19944 ;
  assign w19946 = ~w19306 & w19554 ;
  assign w19947 = w19555 ^ w19946 ;
  assign w19948 = w19298 ^ w19673 ;
  assign w19949 = ( w19298 & w19947 ) | ( w19298 & ~w19948 ) | ( w19947 & ~w19948 ) ;
  assign w19950 = ~\pi092 & w19949 ;
  assign w19951 = ( w19942 & ~w19945 ) | ( w19942 & w19950 ) | ( ~w19945 & w19950 ) ;
  assign w19952 = ( \pi091 & ~w19745 ) | ( \pi091 & w19951 ) | ( ~w19745 & w19951 ) ;
  assign w19953 = ( \pi092 & ~w19950 ) | ( \pi092 & w19952 ) | ( ~w19950 & w19952 ) ;
  assign w19954 = w19942 & ~w19945 ;
  assign w19955 = ( \pi091 & ~w19745 ) | ( \pi091 & w19954 ) | ( ~w19745 & w19954 ) ;
  assign w19956 = w19949 & ~w19955 ;
  assign w19957 = ~w19292 & w19560 ;
  assign w19958 = w19561 ^ w19957 ;
  assign w19959 = w19284 ^ w19673 ;
  assign w19960 = ( w19284 & w19958 ) | ( w19284 & ~w19959 ) | ( w19958 & ~w19959 ) ;
  assign w19961 = ~\pi094 & w19960 ;
  assign w19962 = ( w19953 & ~w19956 ) | ( w19953 & w19961 ) | ( ~w19956 & w19961 ) ;
  assign w19963 = ( \pi093 & ~w19741 ) | ( \pi093 & w19962 ) | ( ~w19741 & w19962 ) ;
  assign w19964 = ( \pi094 & ~w19961 ) | ( \pi094 & w19963 ) | ( ~w19961 & w19963 ) ;
  assign w19965 = w19953 & ~w19956 ;
  assign w19966 = ( \pi093 & ~w19741 ) | ( \pi093 & w19965 ) | ( ~w19741 & w19965 ) ;
  assign w19967 = w19960 & ~w19966 ;
  assign w19968 = ~w19278 & w19566 ;
  assign w19969 = w19567 ^ w19968 ;
  assign w19970 = w19270 ^ w19673 ;
  assign w19971 = ( w19270 & w19969 ) | ( w19270 & ~w19970 ) | ( w19969 & ~w19970 ) ;
  assign w19972 = ~\pi096 & w19971 ;
  assign w19973 = ( w19964 & ~w19967 ) | ( w19964 & w19972 ) | ( ~w19967 & w19972 ) ;
  assign w19974 = ( \pi095 & ~w19737 ) | ( \pi095 & w19973 ) | ( ~w19737 & w19973 ) ;
  assign w19975 = ( \pi096 & ~w19972 ) | ( \pi096 & w19974 ) | ( ~w19972 & w19974 ) ;
  assign w19976 = w19964 & ~w19967 ;
  assign w19977 = ( \pi095 & ~w19737 ) | ( \pi095 & w19976 ) | ( ~w19737 & w19976 ) ;
  assign w19978 = w19971 & ~w19977 ;
  assign w19979 = ~w19264 & w19572 ;
  assign w19980 = w19573 ^ w19979 ;
  assign w19981 = w19256 ^ w19673 ;
  assign w19982 = ( w19256 & w19980 ) | ( w19256 & ~w19981 ) | ( w19980 & ~w19981 ) ;
  assign w19983 = ~\pi098 & w19982 ;
  assign w19984 = ( w19975 & ~w19978 ) | ( w19975 & w19983 ) | ( ~w19978 & w19983 ) ;
  assign w19985 = ( \pi097 & ~w19733 ) | ( \pi097 & w19984 ) | ( ~w19733 & w19984 ) ;
  assign w19986 = ( \pi098 & ~w19983 ) | ( \pi098 & w19985 ) | ( ~w19983 & w19985 ) ;
  assign w19987 = w19975 & ~w19978 ;
  assign w19988 = ( \pi097 & ~w19733 ) | ( \pi097 & w19987 ) | ( ~w19733 & w19987 ) ;
  assign w19989 = w19982 & ~w19988 ;
  assign w19990 = ~w19250 & w19578 ;
  assign w19991 = w19579 ^ w19990 ;
  assign w19992 = w19242 ^ w19673 ;
  assign w19993 = ( w19242 & w19991 ) | ( w19242 & ~w19992 ) | ( w19991 & ~w19992 ) ;
  assign w19994 = ~\pi100 & w19993 ;
  assign w19995 = ( w19986 & ~w19989 ) | ( w19986 & w19994 ) | ( ~w19989 & w19994 ) ;
  assign w19996 = ( \pi099 & ~w19729 ) | ( \pi099 & w19995 ) | ( ~w19729 & w19995 ) ;
  assign w19997 = ( \pi100 & ~w19994 ) | ( \pi100 & w19996 ) | ( ~w19994 & w19996 ) ;
  assign w19998 = w19986 & ~w19989 ;
  assign w19999 = ( \pi099 & ~w19729 ) | ( \pi099 & w19998 ) | ( ~w19729 & w19998 ) ;
  assign w20000 = w19993 & ~w19999 ;
  assign w20001 = ~w19236 & w19584 ;
  assign w20002 = w19585 ^ w20001 ;
  assign w20003 = w19228 ^ w19673 ;
  assign w20004 = ( w19228 & w20002 ) | ( w19228 & ~w20003 ) | ( w20002 & ~w20003 ) ;
  assign w20005 = ~\pi102 & w20004 ;
  assign w20006 = ( w19997 & ~w20000 ) | ( w19997 & w20005 ) | ( ~w20000 & w20005 ) ;
  assign w20007 = ( \pi101 & ~w19725 ) | ( \pi101 & w20006 ) | ( ~w19725 & w20006 ) ;
  assign w20008 = ( \pi102 & ~w20005 ) | ( \pi102 & w20007 ) | ( ~w20005 & w20007 ) ;
  assign w20009 = w19997 & ~w20000 ;
  assign w20010 = ( \pi101 & ~w19725 ) | ( \pi101 & w20009 ) | ( ~w19725 & w20009 ) ;
  assign w20011 = w20004 & ~w20010 ;
  assign w20012 = ~w19222 & w19590 ;
  assign w20013 = w19591 ^ w20012 ;
  assign w20014 = w19214 ^ w19673 ;
  assign w20015 = ( w19214 & w20013 ) | ( w19214 & ~w20014 ) | ( w20013 & ~w20014 ) ;
  assign w20016 = ~\pi104 & w20015 ;
  assign w20017 = ( w20008 & ~w20011 ) | ( w20008 & w20016 ) | ( ~w20011 & w20016 ) ;
  assign w20018 = ( \pi103 & ~w19721 ) | ( \pi103 & w20017 ) | ( ~w19721 & w20017 ) ;
  assign w20019 = ( \pi104 & ~w20016 ) | ( \pi104 & w20018 ) | ( ~w20016 & w20018 ) ;
  assign w20020 = w20008 & ~w20011 ;
  assign w20021 = ( \pi103 & ~w19721 ) | ( \pi103 & w20020 ) | ( ~w19721 & w20020 ) ;
  assign w20022 = w20015 & ~w20021 ;
  assign w20023 = ~w19208 & w19596 ;
  assign w20024 = w19597 ^ w20023 ;
  assign w20025 = w19200 ^ w19673 ;
  assign w20026 = ( w19200 & w20024 ) | ( w19200 & ~w20025 ) | ( w20024 & ~w20025 ) ;
  assign w20027 = ~\pi106 & w20026 ;
  assign w20028 = ( w20019 & ~w20022 ) | ( w20019 & w20027 ) | ( ~w20022 & w20027 ) ;
  assign w20029 = ( \pi105 & ~w19717 ) | ( \pi105 & w20028 ) | ( ~w19717 & w20028 ) ;
  assign w20030 = ( \pi106 & ~w20027 ) | ( \pi106 & w20029 ) | ( ~w20027 & w20029 ) ;
  assign w20031 = w20019 & ~w20022 ;
  assign w20032 = ( \pi105 & ~w19717 ) | ( \pi105 & w20031 ) | ( ~w19717 & w20031 ) ;
  assign w20033 = w20026 & ~w20032 ;
  assign w20034 = ~w19194 & w19602 ;
  assign w20035 = w19603 ^ w20034 ;
  assign w20036 = w19186 ^ w19673 ;
  assign w20037 = ( w19186 & w20035 ) | ( w19186 & ~w20036 ) | ( w20035 & ~w20036 ) ;
  assign w20038 = ~\pi108 & w20037 ;
  assign w20039 = ( w20030 & ~w20033 ) | ( w20030 & w20038 ) | ( ~w20033 & w20038 ) ;
  assign w20040 = ( \pi107 & ~w19713 ) | ( \pi107 & w20039 ) | ( ~w19713 & w20039 ) ;
  assign w20041 = ( \pi108 & ~w20038 ) | ( \pi108 & w20040 ) | ( ~w20038 & w20040 ) ;
  assign w20042 = w20030 & ~w20033 ;
  assign w20043 = ( \pi107 & ~w19713 ) | ( \pi107 & w20042 ) | ( ~w19713 & w20042 ) ;
  assign w20044 = w20037 & ~w20043 ;
  assign w20045 = ~w19180 & w19608 ;
  assign w20046 = w19609 ^ w20045 ;
  assign w20047 = w19172 ^ w19673 ;
  assign w20048 = ( w19172 & w20046 ) | ( w19172 & ~w20047 ) | ( w20046 & ~w20047 ) ;
  assign w20049 = ~\pi110 & w20048 ;
  assign w20050 = ( w20041 & ~w20044 ) | ( w20041 & w20049 ) | ( ~w20044 & w20049 ) ;
  assign w20051 = ( \pi109 & ~w19709 ) | ( \pi109 & w20050 ) | ( ~w19709 & w20050 ) ;
  assign w20052 = ( \pi110 & ~w20049 ) | ( \pi110 & w20051 ) | ( ~w20049 & w20051 ) ;
  assign w20053 = w20041 & ~w20044 ;
  assign w20054 = ( \pi109 & ~w19709 ) | ( \pi109 & w20053 ) | ( ~w19709 & w20053 ) ;
  assign w20055 = w20048 & ~w20054 ;
  assign w20056 = ~w19166 & w19614 ;
  assign w20057 = w19615 ^ w20056 ;
  assign w20058 = w19158 ^ w19673 ;
  assign w20059 = ( w19158 & w20057 ) | ( w19158 & ~w20058 ) | ( w20057 & ~w20058 ) ;
  assign w20060 = ~\pi112 & w20059 ;
  assign w20061 = ( w20052 & ~w20055 ) | ( w20052 & w20060 ) | ( ~w20055 & w20060 ) ;
  assign w20062 = ( \pi111 & ~w19705 ) | ( \pi111 & w20061 ) | ( ~w19705 & w20061 ) ;
  assign w20063 = ( \pi112 & ~w20060 ) | ( \pi112 & w20062 ) | ( ~w20060 & w20062 ) ;
  assign w20064 = w20052 & ~w20055 ;
  assign w20065 = ( \pi111 & ~w19705 ) | ( \pi111 & w20064 ) | ( ~w19705 & w20064 ) ;
  assign w20066 = w20059 & ~w20065 ;
  assign w20067 = ~w19152 & w19620 ;
  assign w20068 = w19621 ^ w20067 ;
  assign w20069 = w19144 ^ w19673 ;
  assign w20070 = ( w19144 & w20068 ) | ( w19144 & ~w20069 ) | ( w20068 & ~w20069 ) ;
  assign w20071 = ~\pi114 & w20070 ;
  assign w20072 = ( w20063 & ~w20066 ) | ( w20063 & w20071 ) | ( ~w20066 & w20071 ) ;
  assign w20073 = ( \pi113 & ~w19701 ) | ( \pi113 & w20072 ) | ( ~w19701 & w20072 ) ;
  assign w20074 = ( \pi114 & ~w20071 ) | ( \pi114 & w20073 ) | ( ~w20071 & w20073 ) ;
  assign w20075 = w20063 & ~w20066 ;
  assign w20076 = ( \pi113 & ~w19701 ) | ( \pi113 & w20075 ) | ( ~w19701 & w20075 ) ;
  assign w20077 = w20070 & ~w20076 ;
  assign w20078 = ~w19138 & w19626 ;
  assign w20079 = w19627 ^ w20078 ;
  assign w20080 = w19130 ^ w19673 ;
  assign w20081 = ( w19130 & w20079 ) | ( w19130 & ~w20080 ) | ( w20079 & ~w20080 ) ;
  assign w20082 = ~\pi116 & w20081 ;
  assign w20083 = ( w20074 & ~w20077 ) | ( w20074 & w20082 ) | ( ~w20077 & w20082 ) ;
  assign w20084 = ( \pi115 & ~w19697 ) | ( \pi115 & w20083 ) | ( ~w19697 & w20083 ) ;
  assign w20085 = ( \pi116 & ~w20082 ) | ( \pi116 & w20084 ) | ( ~w20082 & w20084 ) ;
  assign w20086 = w20074 & ~w20077 ;
  assign w20087 = ( \pi115 & ~w19697 ) | ( \pi115 & w20086 ) | ( ~w19697 & w20086 ) ;
  assign w20088 = w20081 & ~w20087 ;
  assign w20089 = ~w19124 & w19632 ;
  assign w20090 = w19633 ^ w20089 ;
  assign w20091 = w19116 ^ w19673 ;
  assign w20092 = ( w19116 & w20090 ) | ( w19116 & ~w20091 ) | ( w20090 & ~w20091 ) ;
  assign w20093 = ~\pi118 & w20092 ;
  assign w20094 = ( w20085 & ~w20088 ) | ( w20085 & w20093 ) | ( ~w20088 & w20093 ) ;
  assign w20095 = ( \pi117 & ~w19693 ) | ( \pi117 & w20094 ) | ( ~w19693 & w20094 ) ;
  assign w20096 = ( \pi118 & ~w20093 ) | ( \pi118 & w20095 ) | ( ~w20093 & w20095 ) ;
  assign w20097 = w20085 & ~w20088 ;
  assign w20098 = ( \pi117 & ~w19693 ) | ( \pi117 & w20097 ) | ( ~w19693 & w20097 ) ;
  assign w20099 = w20092 & ~w20098 ;
  assign w20100 = ~w19110 & w19638 ;
  assign w20101 = w19639 ^ w20100 ;
  assign w20102 = w19102 ^ w19673 ;
  assign w20103 = ( w19102 & w20101 ) | ( w19102 & ~w20102 ) | ( w20101 & ~w20102 ) ;
  assign w20104 = ~\pi120 & w20103 ;
  assign w20105 = ( w20096 & ~w20099 ) | ( w20096 & w20104 ) | ( ~w20099 & w20104 ) ;
  assign w20106 = ( \pi119 & ~w19689 ) | ( \pi119 & w20105 ) | ( ~w19689 & w20105 ) ;
  assign w20107 = ( \pi120 & ~w20104 ) | ( \pi120 & w20106 ) | ( ~w20104 & w20106 ) ;
  assign w20108 = w20096 & ~w20099 ;
  assign w20109 = ( \pi119 & ~w19689 ) | ( \pi119 & w20108 ) | ( ~w19689 & w20108 ) ;
  assign w20110 = w20103 & ~w20109 ;
  assign w20111 = ~w19096 & w19644 ;
  assign w20112 = w19645 ^ w20111 ;
  assign w20113 = w19088 ^ w19673 ;
  assign w20114 = ( w19088 & w20112 ) | ( w19088 & ~w20113 ) | ( w20112 & ~w20113 ) ;
  assign w20115 = ~\pi122 & w20114 ;
  assign w20116 = ( w20107 & ~w20110 ) | ( w20107 & w20115 ) | ( ~w20110 & w20115 ) ;
  assign w20117 = ( \pi121 & ~w19685 ) | ( \pi121 & w20116 ) | ( ~w19685 & w20116 ) ;
  assign w20118 = ( \pi122 & ~w20115 ) | ( \pi122 & w20117 ) | ( ~w20115 & w20117 ) ;
  assign w20119 = w20107 & ~w20110 ;
  assign w20120 = ( \pi121 & ~w19685 ) | ( \pi121 & w20119 ) | ( ~w19685 & w20119 ) ;
  assign w20121 = w20114 & ~w20120 ;
  assign w20122 = ~w19082 & w19650 ;
  assign w20123 = w19651 ^ w20122 ;
  assign w20124 = w19074 ^ w19673 ;
  assign w20125 = ( w19074 & w20123 ) | ( w19074 & ~w20124 ) | ( w20123 & ~w20124 ) ;
  assign w20126 = ~\pi124 & w20125 ;
  assign w20127 = ( w20118 & ~w20121 ) | ( w20118 & w20126 ) | ( ~w20121 & w20126 ) ;
  assign w20128 = ( \pi123 & ~w19681 ) | ( \pi123 & w20127 ) | ( ~w19681 & w20127 ) ;
  assign w20129 = ( \pi124 & ~w20126 ) | ( \pi124 & w20128 ) | ( ~w20126 & w20128 ) ;
  assign w20130 = w20118 & ~w20121 ;
  assign w20131 = ( \pi123 & ~w19681 ) | ( \pi123 & w20130 ) | ( ~w19681 & w20130 ) ;
  assign w20132 = w20125 & ~w20131 ;
  assign w20133 = ~w19068 & w19656 ;
  assign w20134 = w19657 ^ w20133 ;
  assign w20135 = w19060 ^ w19673 ;
  assign w20136 = ( w19060 & w20134 ) | ( w19060 & ~w20135 ) | ( w20134 & ~w20135 ) ;
  assign w20137 = ~\pi126 & w20136 ;
  assign w20138 = ( w20129 & ~w20132 ) | ( w20129 & w20137 ) | ( ~w20132 & w20137 ) ;
  assign w20139 = ( \pi125 & ~w19677 ) | ( \pi125 & w20138 ) | ( ~w19677 & w20138 ) ;
  assign w20140 = ( \pi126 & ~w20137 ) | ( \pi126 & w20139 ) | ( ~w20137 & w20139 ) ;
  assign w20141 = w20129 & ~w20132 ;
  assign w20142 = ( \pi125 & ~w19677 ) | ( \pi125 & w20141 ) | ( ~w19677 & w20141 ) ;
  assign w20143 = w20136 & ~w20142 ;
  assign w20144 = w19663 | w19665 ;
  assign w20145 = ( \pi127 & ~w19061 ) | ( \pi127 & w19659 ) | ( ~w19061 & w19659 ) ;
  assign w20146 = \pi126 ^ w20145 ;
  assign w20147 = ( \pi127 & w20144 ) | ( \pi127 & ~w20146 ) | ( w20144 & ~w20146 ) ;
  assign w20148 = w20144 & w20147 ;
  assign w20149 = w20140 & ~w20143 ;
  assign w20150 = ( \pi127 & ~w20148 ) | ( \pi127 & w20149 ) | ( ~w20148 & w20149 ) ;
  assign w20151 = w437 | w454 ;
  assign w20152 = ( w195 & w198 ) | ( w195 & ~w298 ) | ( w198 & ~w298 ) ;
  assign w20153 = w345 | w20152 ;
  assign w20154 = \pi065 | w250 ;
  assign w20155 = ( ~\pi063 & \pi064 ) | ( ~\pi063 & w20154 ) | ( \pi064 & w20154 ) ;
  assign w20156 = ( \pi066 & ~w20154 ) | ( \pi066 & w20155 ) | ( ~w20154 & w20155 ) ;
  assign w20157 = w20154 | w20156 ;
  assign w20158 = ( ~w446 & w491 ) | ( ~w446 & w20157 ) | ( w491 & w20157 ) ;
  assign w20159 = w446 | w20158 ;
  assign w20160 = \pi064 & ~\pi065 ;
  assign w20161 = ~w129 & w20160 ;
  assign w20162 = ~w197 & w20161 ;
  assign w20163 = ( w207 & ~w298 ) | ( w207 & w20162 ) | ( ~w298 & w20162 ) ;
  assign w20164 = ~w207 & w20163 ;
  assign w20165 = \pi063 & ~w20164 ;
  assign w20166 = ( \pi065 & w194 ) | ( \pi065 & ~w20165 ) | ( w194 & ~w20165 ) ;
  assign w20167 = w212 & ~w20166 ;
  assign w20168 = ( ~\pi063 & w212 ) | ( ~\pi063 & w20164 ) | ( w212 & w20164 ) ;
  assign w20169 = w20167 & w20168 ;
  assign w20170 = ( w228 & w20164 ) | ( w228 & ~w20166 ) | ( w20164 & ~w20166 ) ;
  assign w20171 = w20165 & ~w20170 ;
  assign w20172 = ( \pi062 & ~w293 ) | ( \pi062 & w20166 ) | ( ~w293 & w20166 ) ;
  assign w20173 = \pi062 & w20172 ;
  assign w20174 = w300 & ~w20166 ;
  assign w20175 = w20173 | w20174 ;
  assign w20176 = ( \pi065 & w231 ) | ( \pi065 & ~w20175 ) | ( w231 & ~w20175 ) ;
  assign w20177 = w20169 | w20171 ;
  assign w20178 = ( \pi066 & w20176 ) | ( \pi066 & ~w20177 ) | ( w20176 & ~w20177 ) ;
  assign w20179 = ( \pi067 & w20169 ) | ( \pi067 & w20171 ) | ( w20169 & w20171 ) ;
  assign w20180 = \pi067 & ~w20179 ;
  assign w20181 = \pi066 ^ w20176 ;
  assign w20182 = ( ~\pi067 & w309 ) | ( ~\pi067 & w20181 ) | ( w309 & w20181 ) ;
  assign w20183 = ( w20180 & w20181 ) | ( w20180 & ~w20182 ) | ( w20181 & ~w20182 ) ;
  assign w20184 = ( ~w327 & w20175 ) | ( ~w327 & w20178 ) | ( w20175 & w20178 ) ;
  assign w20185 = w20175 & w20184 ;
  assign w20186 = w336 & ~w20173 ;
  assign w20187 = ( ~w20173 & w20174 ) | ( ~w20173 & w20178 ) | ( w20174 & w20178 ) ;
  assign w20188 = w20186 & ~w20187 ;
  assign w20189 = w20185 | w20188 ;
  assign w20190 = ~\pi066 & w20189 ;
  assign w20191 = ( \pi066 & ~w20185 ) | ( \pi066 & w20188 ) | ( ~w20185 & w20188 ) ;
  assign w20192 = ~w20188 & w20191 ;
  assign w20193 = ( \pi061 & ~w348 ) | ( \pi061 & w20178 ) | ( ~w348 & w20178 ) ;
  assign w20194 = \pi061 & w20193 ;
  assign w20195 = w353 | w20178 ;
  assign w20196 = ( ~w20178 & w20194 ) | ( ~w20178 & w20195 ) | ( w20194 & w20195 ) ;
  assign w20197 = ( \pi065 & w358 ) | ( \pi065 & ~w20196 ) | ( w358 & ~w20196 ) ;
  assign w20198 = w20192 | w20197 ;
  assign w20199 = ~w20190 & w20198 ;
  assign w20200 = ( \pi066 & ~w309 ) | ( \pi066 & w20176 ) | ( ~w309 & w20176 ) ;
  assign w20201 = \pi066 & w20176 ;
  assign w20202 = ( w20177 & ~w20200 ) | ( w20177 & w20201 ) | ( ~w20200 & w20201 ) ;
  assign w20203 = ~\pi067 & w20202 ;
  assign w20204 = ( w20183 & w20199 ) | ( w20183 & ~w20203 ) | ( w20199 & ~w20203 ) ;
  assign w20205 = ~w20203 & w20204 ;
  assign w20206 = ~w20199 & w20203 ;
  assign w20207 = ~w370 & w20206 ;
  assign w20208 = ( w370 & w20202 ) | ( w370 & w20205 ) | ( w20202 & w20205 ) ;
  assign w20209 = w20202 & w20208 ;
  assign w20210 = ( \pi068 & w20207 ) | ( \pi068 & ~w20209 ) | ( w20207 & ~w20209 ) ;
  assign w20211 = ~w20207 & w20210 ;
  assign w20212 = ( w20190 & w20192 ) | ( w20190 & w20197 ) | ( w20192 & w20197 ) ;
  assign w20213 = w20197 & w20212 ;
  assign w20214 = w370 | w20213 ;
  assign w20215 = ( w20198 & ~w20205 ) | ( w20198 & w20213 ) | ( ~w20205 & w20213 ) ;
  assign w20216 = ~w20214 & w20215 ;
  assign w20217 = ( \pi066 & ~w370 ) | ( \pi066 & w20213 ) | ( ~w370 & w20213 ) ;
  assign w20218 = w370 & w20217 ;
  assign w20219 = ( w20205 & w20217 ) | ( w20205 & w20218 ) | ( w20217 & w20218 ) ;
  assign w20220 = ( w20189 & ~w20217 ) | ( w20189 & w20219 ) | ( ~w20217 & w20219 ) ;
  assign w20221 = w20216 | w20220 ;
  assign w20222 = ~\pi067 & w20221 ;
  assign w20223 = ( \pi067 & ~w20216 ) | ( \pi067 & w20220 ) | ( ~w20216 & w20220 ) ;
  assign w20224 = ~w20220 & w20223 ;
  assign w20225 = ( ~w402 & w20196 ) | ( ~w402 & w20205 ) | ( w20196 & w20205 ) ;
  assign w20226 = w20196 & w20225 ;
  assign w20227 = ( w406 & w20178 ) | ( w406 & w20205 ) | ( w20178 & w20205 ) ;
  assign w20228 = w348 & ~w20227 ;
  assign w20229 = ( \pi061 & w20205 ) | ( \pi061 & ~w20228 ) | ( w20205 & ~w20228 ) ;
  assign w20230 = ( ~w353 & w406 ) | ( ~w353 & w20227 ) | ( w406 & w20227 ) ;
  assign w20231 = ~w20229 & w20230 ;
  assign w20232 = w20226 | w20231 ;
  assign w20233 = ~\pi066 & w20232 ;
  assign w20234 = ( \pi066 & ~w20226 ) | ( \pi066 & w20231 ) | ( ~w20226 & w20231 ) ;
  assign w20235 = ~w20231 & w20234 ;
  assign w20236 = ( \pi060 & ~w420 ) | ( \pi060 & w20205 ) | ( ~w420 & w20205 ) ;
  assign w20237 = \pi060 & w20236 ;
  assign w20238 = w424 | w20205 ;
  assign w20239 = ( ~w20205 & w20237 ) | ( ~w20205 & w20238 ) | ( w20237 & w20238 ) ;
  assign w20240 = ( \pi065 & w416 ) | ( \pi065 & ~w20239 ) | ( w416 & ~w20239 ) ;
  assign w20241 = w20235 | w20240 ;
  assign w20242 = ( w20224 & ~w20233 ) | ( w20224 & w20241 ) | ( ~w20233 & w20241 ) ;
  assign w20243 = w20224 | w20242 ;
  assign w20244 = ( ~\pi068 & w20207 ) | ( ~\pi068 & w20209 ) | ( w20207 & w20209 ) ;
  assign w20245 = ~\pi068 & w20244 ;
  assign w20246 = ~w20222 & w20243 ;
  assign w20247 = w20211 & ~w20246 ;
  assign w20248 = ( ~w20245 & w20246 ) | ( ~w20245 & w20247 ) | ( w20246 & w20247 ) ;
  assign w20249 = ~w20233 & w20241 ;
  assign w20250 = ( w20222 & w20224 ) | ( w20222 & w20241 ) | ( w20224 & w20241 ) ;
  assign w20251 = w20249 & w20250 ;
  assign w20252 = ~w454 & w20243 ;
  assign w20253 = ( w20243 & w20248 ) | ( w20243 & w20251 ) | ( w20248 & w20251 ) ;
  assign w20254 = w20252 & ~w20253 ;
  assign w20255 = ( \pi067 & ~w454 ) | ( \pi067 & w20251 ) | ( ~w454 & w20251 ) ;
  assign w20256 = w454 & w20255 ;
  assign w20257 = ( w20248 & w20255 ) | ( w20248 & w20256 ) | ( w20255 & w20256 ) ;
  assign w20258 = ( w20221 & ~w20255 ) | ( w20221 & w20257 ) | ( ~w20255 & w20257 ) ;
  assign w20259 = w20254 | w20258 ;
  assign w20260 = \pi068 ^ w20259 ;
  assign w20261 = ( w20233 & w20235 ) | ( w20233 & w20240 ) | ( w20235 & w20240 ) ;
  assign w20262 = w20240 & w20261 ;
  assign w20263 = w454 | w20262 ;
  assign w20264 = ( w20241 & ~w20248 ) | ( w20241 & w20262 ) | ( ~w20248 & w20262 ) ;
  assign w20265 = ~w20263 & w20264 ;
  assign w20266 = ( \pi066 & ~w454 ) | ( \pi066 & w20262 ) | ( ~w454 & w20262 ) ;
  assign w20267 = w454 & w20266 ;
  assign w20268 = ( w20248 & w20266 ) | ( w20248 & w20267 ) | ( w20266 & w20267 ) ;
  assign w20269 = ( w20232 & ~w20266 ) | ( w20232 & w20268 ) | ( ~w20266 & w20268 ) ;
  assign w20270 = w20265 | w20269 ;
  assign w20271 = \pi067 ^ w20270 ;
  assign w20272 = ( ~w487 & w20239 ) | ( ~w487 & w20248 ) | ( w20239 & w20248 ) ;
  assign w20273 = w20239 & w20272 ;
  assign w20274 = ( w494 & w20205 ) | ( w494 & w20248 ) | ( w20205 & w20248 ) ;
  assign w20275 = w420 & ~w20274 ;
  assign w20276 = ( \pi060 & w20248 ) | ( \pi060 & ~w20275 ) | ( w20248 & ~w20275 ) ;
  assign w20277 = ( ~w424 & w494 ) | ( ~w424 & w20274 ) | ( w494 & w20274 ) ;
  assign w20278 = ~w20276 & w20277 ;
  assign w20279 = w20273 | w20278 ;
  assign w20280 = ~\pi066 & w20279 ;
  assign w20281 = ( \pi059 & ~w508 ) | ( \pi059 & w20248 ) | ( ~w508 & w20248 ) ;
  assign w20282 = \pi059 & w20281 ;
  assign w20283 = w291 | w20248 ;
  assign w20284 = w513 & ~w20283 ;
  assign w20285 = ~w511 & w20284 ;
  assign w20286 = w20282 | w20285 ;
  assign w20287 = ( ~w517 & w20282 ) | ( ~w517 & w20285 ) | ( w20282 & w20285 ) ;
  assign w20288 = \pi065 ^ w20287 ;
  assign w20289 = w517 | w20288 ;
  assign w20290 = ~\pi065 & w20286 ;
  assign w20291 = \pi066 ^ w20279 ;
  assign w20292 = ( w20289 & ~w20290 ) | ( w20289 & w20291 ) | ( ~w20290 & w20291 ) ;
  assign w20293 = w20291 | w20292 ;
  assign w20294 = ( w20271 & ~w20280 ) | ( w20271 & w20293 ) | ( ~w20280 & w20293 ) ;
  assign w20295 = w20271 | w20294 ;
  assign w20296 = ~\pi067 & w20270 ;
  assign w20297 = ( w20260 & w20295 ) | ( w20260 & ~w20296 ) | ( w20295 & ~w20296 ) ;
  assign w20298 = w20260 | w20297 ;
  assign w20299 = ~\pi068 & w20259 ;
  assign w20300 = w20211 & w20245 ;
  assign w20301 = ( w20222 & ~w20243 ) | ( w20222 & w20300 ) | ( ~w20243 & w20300 ) ;
  assign w20302 = ( w454 & w20300 ) | ( w454 & ~w20301 ) | ( w20300 & ~w20301 ) ;
  assign w20303 = w20300 & ~w20302 ;
  assign w20304 = w20207 | w20209 ;
  assign w20305 = ( w454 & ~w20222 ) | ( w454 & w20243 ) | ( ~w20222 & w20243 ) ;
  assign w20306 = \pi068 ^ w20305 ;
  assign w20307 = ( w454 & w20304 ) | ( w454 & ~w20306 ) | ( w20304 & ~w20306 ) ;
  assign w20308 = w20304 & w20307 ;
  assign w20309 = w20303 | w20308 ;
  assign w20310 = \pi069 ^ w20309 ;
  assign w20311 = w546 | w20310 ;
  assign w20312 = ( w546 & w20298 ) | ( w546 & ~w20299 ) | ( w20298 & ~w20299 ) ;
  assign w20313 = w20311 | w20312 ;
  assign w20314 = ~w454 & w20309 ;
  assign w20315 = w20313 & ~w20314 ;
  assign w20316 = w20295 & ~w20296 ;
  assign w20317 = w20260 ^ w20316 ;
  assign w20318 = ~w20315 & w20317 ;
  assign w20319 = ( w20259 & ~w20313 ) | ( w20259 & w20314 ) | ( ~w20313 & w20314 ) ;
  assign w20320 = w20259 & ~w20319 ;
  assign w20321 = w20318 | w20320 ;
  assign w20322 = w20298 & ~w20299 ;
  assign w20323 = w20310 ^ w20322 ;
  assign w20324 = ~w20315 & w20323 ;
  assign w20325 = ( w454 & ~w20309 ) | ( w454 & w20313 ) | ( ~w20309 & w20313 ) ;
  assign w20326 = w20309 & w20325 ;
  assign w20327 = w20324 | w20326 ;
  assign w20328 = ~\pi069 & w20321 ;
  assign w20329 = ~w20280 & w20293 ;
  assign w20330 = w20271 ^ w20329 ;
  assign w20331 = ~w20315 & w20330 ;
  assign w20332 = ( w20270 & ~w20313 ) | ( w20270 & w20314 ) | ( ~w20313 & w20314 ) ;
  assign w20333 = w20270 & ~w20332 ;
  assign w20334 = w20331 | w20333 ;
  assign w20335 = ~\pi068 & w20334 ;
  assign w20336 = w20289 & ~w20290 ;
  assign w20337 = w20291 ^ w20336 ;
  assign w20338 = ~w20315 & w20337 ;
  assign w20339 = ( w20279 & ~w20313 ) | ( w20279 & w20314 ) | ( ~w20313 & w20314 ) ;
  assign w20340 = w20279 & ~w20339 ;
  assign w20341 = w20338 | w20340 ;
  assign w20342 = ~\pi067 & w20341 ;
  assign w20343 = ( w20282 & w20285 ) | ( w20282 & ~w20315 ) | ( w20285 & ~w20315 ) ;
  assign w20344 = ( ~\pi058 & \pi064 ) | ( ~\pi058 & w20315 ) | ( \pi064 & w20315 ) ;
  assign w20345 = w20343 ^ w20344 ;
  assign w20346 = \pi065 ^ w20345 ;
  assign w20347 = ~w20315 & w20346 ;
  assign w20348 = ( w20286 & ~w20313 ) | ( w20286 & w20314 ) | ( ~w20313 & w20314 ) ;
  assign w20349 = w20286 & ~w20348 ;
  assign w20350 = w20347 | w20349 ;
  assign w20351 = ~\pi066 & w20350 ;
  assign w20352 = \pi064 & ~w20315 ;
  assign w20353 = \pi058 ^ w20352 ;
  assign w20354 = \pi066 ^ w20350 ;
  assign w20355 = ( \pi064 & ~w20315 ) | ( \pi064 & w20354 ) | ( ~w20315 & w20354 ) ;
  assign w20356 = \pi058 ^ w20355 ;
  assign w20357 = ( \pi065 & w638 ) | ( \pi065 & ~w20356 ) | ( w638 & ~w20356 ) ;
  assign w20358 = w20354 | w20357 ;
  assign w20359 = \pi067 ^ w20341 ;
  assign w20360 = ( ~w20351 & w20358 ) | ( ~w20351 & w20359 ) | ( w20358 & w20359 ) ;
  assign w20361 = w20359 | w20360 ;
  assign w20362 = \pi068 ^ w20334 ;
  assign w20363 = ( ~w20342 & w20361 ) | ( ~w20342 & w20362 ) | ( w20361 & w20362 ) ;
  assign w20364 = w20362 | w20363 ;
  assign w20365 = \pi069 ^ w20321 ;
  assign w20366 = ( ~w20335 & w20364 ) | ( ~w20335 & w20365 ) | ( w20364 & w20365 ) ;
  assign w20367 = w20365 | w20366 ;
  assign w20368 = \pi070 ^ w20327 ;
  assign w20369 = w20328 & ~w20368 ;
  assign w20370 = ( w20367 & w20368 ) | ( w20367 & ~w20369 ) | ( w20368 & ~w20369 ) ;
  assign w20371 = ~\pi070 & w20327 ;
  assign w20372 = w20370 & ~w20371 ;
  assign w20373 = w612 | w20372 ;
  assign w20374 = w20321 & w20373 ;
  assign w20375 = ~w20335 & w20364 ;
  assign w20376 = w20365 ^ w20375 ;
  assign w20377 = ~w20373 & w20376 ;
  assign w20378 = w20374 | w20377 ;
  assign w20379 = w20327 & w20373 ;
  assign w20380 = ~w20328 & w20367 ;
  assign w20381 = w20368 ^ w20380 ;
  assign w20382 = ~w20373 & w20381 ;
  assign w20383 = w20379 | w20382 ;
  assign w20384 = ~\pi070 & w20378 ;
  assign w20385 = w20334 & w20373 ;
  assign w20386 = ~w20342 & w20361 ;
  assign w20387 = w20362 ^ w20386 ;
  assign w20388 = ~w20373 & w20387 ;
  assign w20389 = w20385 | w20388 ;
  assign w20390 = ~\pi069 & w20389 ;
  assign w20391 = w20341 & w20373 ;
  assign w20392 = ~w20351 & w20358 ;
  assign w20393 = w20359 ^ w20392 ;
  assign w20394 = ~w20373 & w20393 ;
  assign w20395 = w20391 | w20394 ;
  assign w20396 = ~\pi068 & w20395 ;
  assign w20397 = w20350 & w20373 ;
  assign w20398 = ( \pi065 & w638 ) | ( \pi065 & ~w20353 ) | ( w638 & ~w20353 ) ;
  assign w20399 = w20354 ^ w20398 ;
  assign w20400 = ( w612 & w20372 ) | ( w612 & w20399 ) | ( w20372 & w20399 ) ;
  assign w20401 = w20399 & ~w20400 ;
  assign w20402 = w20397 | w20401 ;
  assign w20403 = ~\pi067 & w20402 ;
  assign w20404 = \pi057 ^ w20315 ;
  assign w20405 = ( \pi064 & w612 ) | ( \pi064 & w20404 ) | ( w612 & w20404 ) ;
  assign w20406 = w645 ^ w20405 ;
  assign w20407 = ~w612 & w20406 ;
  assign w20408 = ~w20372 & w20407 ;
  assign w20409 = ( w20353 & w20373 ) | ( w20353 & w20408 ) | ( w20373 & w20408 ) ;
  assign w20410 = w20408 | w20409 ;
  assign w20411 = ~\pi066 & w20410 ;
  assign w20412 = ( \pi057 & ~w659 ) | ( \pi057 & w20372 ) | ( ~w659 & w20372 ) ;
  assign w20413 = \pi057 & w20412 ;
  assign w20414 = w666 | w20372 ;
  assign w20415 = ( ~w20372 & w20413 ) | ( ~w20372 & w20414 ) | ( w20413 & w20414 ) ;
  assign w20416 = \pi065 & w20415 ;
  assign w20417 = ( \pi065 & w666 ) | ( \pi065 & ~w20372 ) | ( w666 & ~w20372 ) ;
  assign w20418 = w659 & ~w20372 ;
  assign w20419 = ( \pi057 & \pi065 ) | ( \pi057 & ~w20418 ) | ( \pi065 & ~w20418 ) ;
  assign w20420 = w20417 | w20419 ;
  assign w20421 = ~w20416 & w20420 ;
  assign w20422 = ( \pi064 & ~w676 ) | ( \pi064 & w20421 ) | ( ~w676 & w20421 ) ;
  assign w20423 = ~\pi065 & w20415 ;
  assign w20424 = ~w20353 & w20373 ;
  assign w20425 = ( w20373 & w20408 ) | ( w20373 & ~w20424 ) | ( w20408 & ~w20424 ) ;
  assign w20426 = \pi066 ^ w20425 ;
  assign w20427 = ( w20422 & ~w20423 ) | ( w20422 & w20426 ) | ( ~w20423 & w20426 ) ;
  assign w20428 = w20426 | w20427 ;
  assign w20429 = \pi067 ^ w20402 ;
  assign w20430 = ( ~w20411 & w20428 ) | ( ~w20411 & w20429 ) | ( w20428 & w20429 ) ;
  assign w20431 = w20429 | w20430 ;
  assign w20432 = \pi068 ^ w20395 ;
  assign w20433 = ( ~w20403 & w20431 ) | ( ~w20403 & w20432 ) | ( w20431 & w20432 ) ;
  assign w20434 = w20432 | w20433 ;
  assign w20435 = \pi069 ^ w20389 ;
  assign w20436 = ( ~w20396 & w20434 ) | ( ~w20396 & w20435 ) | ( w20434 & w20435 ) ;
  assign w20437 = w20435 | w20436 ;
  assign w20438 = \pi070 ^ w20378 ;
  assign w20439 = ( ~w20390 & w20437 ) | ( ~w20390 & w20438 ) | ( w20437 & w20438 ) ;
  assign w20440 = w20438 | w20439 ;
  assign w20441 = \pi071 ^ w20383 ;
  assign w20442 = w20384 & ~w20441 ;
  assign w20443 = ( w20440 & w20441 ) | ( w20440 & ~w20442 ) | ( w20441 & ~w20442 ) ;
  assign w20444 = ~\pi071 & w20383 ;
  assign w20445 = w20443 & ~w20444 ;
  assign w20446 = w703 | w20445 ;
  assign w20447 = w20378 & w20446 ;
  assign w20448 = ~w20390 & w20437 ;
  assign w20449 = w20438 ^ w20448 ;
  assign w20450 = ~w20446 & w20449 ;
  assign w20451 = w20447 | w20450 ;
  assign w20452 = ~\pi071 & w20451 ;
  assign w20453 = w20389 & w20446 ;
  assign w20454 = ~w20396 & w20434 ;
  assign w20455 = w20435 ^ w20454 ;
  assign w20456 = ~w20446 & w20455 ;
  assign w20457 = w20453 | w20456 ;
  assign w20458 = ~\pi070 & w20457 ;
  assign w20459 = w20395 & w20446 ;
  assign w20460 = ~w20403 & w20431 ;
  assign w20461 = w20432 ^ w20460 ;
  assign w20462 = ~w20446 & w20461 ;
  assign w20463 = w20459 | w20462 ;
  assign w20464 = ~\pi069 & w20463 ;
  assign w20465 = w20402 & w20446 ;
  assign w20466 = ~w20411 & w20428 ;
  assign w20467 = w20429 ^ w20466 ;
  assign w20468 = ~w20446 & w20467 ;
  assign w20469 = w20465 | w20468 ;
  assign w20470 = ~\pi068 & w20469 ;
  assign w20471 = w20410 & w20446 ;
  assign w20472 = w20422 & ~w20423 ;
  assign w20473 = w20426 ^ w20472 ;
  assign w20474 = ~w20446 & w20473 ;
  assign w20475 = w20471 | w20474 ;
  assign w20476 = ~\pi067 & w20475 ;
  assign w20477 = w20415 & w20446 ;
  assign w20478 = ( ~\pi056 & \pi064 ) | ( ~\pi056 & w20445 ) | ( \pi064 & w20445 ) ;
  assign w20479 = ( w703 & ~w20416 ) | ( w703 & w20420 ) | ( ~w20416 & w20420 ) ;
  assign w20480 = w20478 ^ w20479 ;
  assign w20481 = ( w703 & ~w20445 ) | ( w703 & w20480 ) | ( ~w20445 & w20480 ) ;
  assign w20482 = ~w703 & w20481 ;
  assign w20483 = w20477 | w20482 ;
  assign w20484 = ~\pi066 & w20483 ;
  assign w20485 = ( \pi056 & ~w746 ) | ( \pi056 & w20445 ) | ( ~w746 & w20445 ) ;
  assign w20486 = \pi056 & w20485 ;
  assign w20487 = w750 | w20445 ;
  assign w20488 = ( ~w20445 & w20486 ) | ( ~w20445 & w20487 ) | ( w20486 & w20487 ) ;
  assign w20489 = w746 & ~w20487 ;
  assign w20490 = \pi056 & ~w20489 ;
  assign w20491 = ( ~w20445 & w20487 ) | ( ~w20445 & w20490 ) | ( w20487 & w20490 ) ;
  assign w20492 = \pi065 ^ w20491 ;
  assign w20493 = w755 | w20492 ;
  assign w20494 = ~\pi065 & w20488 ;
  assign w20495 = \pi066 ^ w20483 ;
  assign w20496 = ( w20493 & ~w20494 ) | ( w20493 & w20495 ) | ( ~w20494 & w20495 ) ;
  assign w20497 = w20495 | w20496 ;
  assign w20498 = \pi067 ^ w20475 ;
  assign w20499 = ( ~w20484 & w20497 ) | ( ~w20484 & w20498 ) | ( w20497 & w20498 ) ;
  assign w20500 = w20498 | w20499 ;
  assign w20501 = \pi068 ^ w20469 ;
  assign w20502 = ( ~w20476 & w20500 ) | ( ~w20476 & w20501 ) | ( w20500 & w20501 ) ;
  assign w20503 = w20501 | w20502 ;
  assign w20504 = \pi069 ^ w20463 ;
  assign w20505 = ( ~w20470 & w20503 ) | ( ~w20470 & w20504 ) | ( w20503 & w20504 ) ;
  assign w20506 = w20504 | w20505 ;
  assign w20507 = \pi070 ^ w20457 ;
  assign w20508 = ( ~w20464 & w20506 ) | ( ~w20464 & w20507 ) | ( w20506 & w20507 ) ;
  assign w20509 = w20507 | w20508 ;
  assign w20510 = \pi071 ^ w20451 ;
  assign w20511 = ( ~w20458 & w20509 ) | ( ~w20458 & w20510 ) | ( w20509 & w20510 ) ;
  assign w20512 = w20510 | w20511 ;
  assign w20513 = w20383 & w20446 ;
  assign w20514 = ~w20384 & w20440 ;
  assign w20515 = w20441 ^ w20514 ;
  assign w20516 = ~w20446 & w20515 ;
  assign w20517 = w20513 | w20516 ;
  assign w20518 = ~\pi072 & w20517 ;
  assign w20519 = ( \pi072 & ~w20513 ) | ( \pi072 & w20516 ) | ( ~w20513 & w20516 ) ;
  assign w20520 = ~w20516 & w20519 ;
  assign w20521 = w788 | w20520 ;
  assign w20522 = ( w291 & w20518 ) | ( w291 & ~w20520 ) | ( w20518 & ~w20520 ) ;
  assign w20523 = w20521 | w20522 ;
  assign w20524 = ( ~w20452 & w20512 ) | ( ~w20452 & w20523 ) | ( w20512 & w20523 ) ;
  assign w20525 = w20523 | w20524 ;
  assign w20526 = ~w703 & w20517 ;
  assign w20527 = w20525 & ~w20526 ;
  assign w20528 = ~w20458 & w20509 ;
  assign w20529 = w20510 ^ w20528 ;
  assign w20530 = ~w20527 & w20529 ;
  assign w20531 = ( w20451 & w20525 ) | ( w20451 & w20526 ) | ( w20525 & w20526 ) ;
  assign w20532 = ~w20526 & w20531 ;
  assign w20533 = w20530 | w20532 ;
  assign w20534 = w20518 | w20520 ;
  assign w20535 = ( ~w20452 & w20512 ) | ( ~w20452 & w20527 ) | ( w20512 & w20527 ) ;
  assign w20536 = w20534 ^ w20535 ;
  assign w20537 = ~w20527 & w20536 ;
  assign w20538 = ( w703 & ~w20517 ) | ( w703 & w20525 ) | ( ~w20517 & w20525 ) ;
  assign w20539 = w20517 & w20538 ;
  assign w20540 = w20537 | w20539 ;
  assign w20541 = ~\pi072 & w20533 ;
  assign w20542 = ~w20464 & w20506 ;
  assign w20543 = w20507 ^ w20542 ;
  assign w20544 = ~w20527 & w20543 ;
  assign w20545 = ( w20457 & w20525 ) | ( w20457 & w20526 ) | ( w20525 & w20526 ) ;
  assign w20546 = ~w20526 & w20545 ;
  assign w20547 = w20544 | w20546 ;
  assign w20548 = ~\pi071 & w20547 ;
  assign w20549 = ~w20470 & w20503 ;
  assign w20550 = w20504 ^ w20549 ;
  assign w20551 = ~w20527 & w20550 ;
  assign w20552 = ( w20463 & w20525 ) | ( w20463 & w20526 ) | ( w20525 & w20526 ) ;
  assign w20553 = ~w20526 & w20552 ;
  assign w20554 = w20551 | w20553 ;
  assign w20555 = ~\pi070 & w20554 ;
  assign w20556 = ~w20476 & w20500 ;
  assign w20557 = w20501 ^ w20556 ;
  assign w20558 = ~w20527 & w20557 ;
  assign w20559 = ( w20469 & w20525 ) | ( w20469 & w20526 ) | ( w20525 & w20526 ) ;
  assign w20560 = ~w20526 & w20559 ;
  assign w20561 = w20558 | w20560 ;
  assign w20562 = ~\pi069 & w20561 ;
  assign w20563 = ~w20484 & w20497 ;
  assign w20564 = w20498 ^ w20563 ;
  assign w20565 = ~w20527 & w20564 ;
  assign w20566 = ( w20475 & w20525 ) | ( w20475 & w20526 ) | ( w20525 & w20526 ) ;
  assign w20567 = ~w20526 & w20566 ;
  assign w20568 = w20565 | w20567 ;
  assign w20569 = ~\pi068 & w20568 ;
  assign w20570 = w20493 & ~w20494 ;
  assign w20571 = w20495 ^ w20570 ;
  assign w20572 = ~w20527 & w20571 ;
  assign w20573 = ( w20483 & w20525 ) | ( w20483 & w20526 ) | ( w20525 & w20526 ) ;
  assign w20574 = ~w20526 & w20573 ;
  assign w20575 = w20572 | w20574 ;
  assign w20576 = ~\pi067 & w20575 ;
  assign w20577 = w750 ^ w20445 ;
  assign w20578 = ( \pi056 & ~w845 ) | ( \pi056 & w20577 ) | ( ~w845 & w20577 ) ;
  assign w20579 = ( \pi056 & w750 ) | ( \pi056 & w20578 ) | ( w750 & w20578 ) ;
  assign w20580 = w755 ^ w20579 ;
  assign w20581 = \pi065 ^ w20580 ;
  assign w20582 = ~w20527 & w20581 ;
  assign w20583 = ( w20488 & w20525 ) | ( w20488 & w20526 ) | ( w20525 & w20526 ) ;
  assign w20584 = ~w20526 & w20583 ;
  assign w20585 = w20582 | w20584 ;
  assign w20586 = ~\pi066 & w20585 ;
  assign w20587 = \pi066 ^ w20585 ;
  assign w20588 = ( \pi064 & ~w20527 ) | ( \pi064 & w20587 ) | ( ~w20527 & w20587 ) ;
  assign w20589 = \pi055 ^ w20588 ;
  assign w20590 = ( \pi065 & w856 ) | ( \pi065 & ~w20589 ) | ( w856 & ~w20589 ) ;
  assign w20591 = w20587 | w20590 ;
  assign w20592 = \pi067 ^ w20575 ;
  assign w20593 = ( ~w20586 & w20591 ) | ( ~w20586 & w20592 ) | ( w20591 & w20592 ) ;
  assign w20594 = w20592 | w20593 ;
  assign w20595 = \pi068 ^ w20568 ;
  assign w20596 = ( ~w20576 & w20594 ) | ( ~w20576 & w20595 ) | ( w20594 & w20595 ) ;
  assign w20597 = w20595 | w20596 ;
  assign w20598 = \pi069 ^ w20561 ;
  assign w20599 = ( ~w20569 & w20597 ) | ( ~w20569 & w20598 ) | ( w20597 & w20598 ) ;
  assign w20600 = w20598 | w20599 ;
  assign w20601 = \pi070 ^ w20554 ;
  assign w20602 = ( ~w20562 & w20600 ) | ( ~w20562 & w20601 ) | ( w20600 & w20601 ) ;
  assign w20603 = w20601 | w20602 ;
  assign w20604 = \pi071 ^ w20547 ;
  assign w20605 = ( ~w20555 & w20603 ) | ( ~w20555 & w20604 ) | ( w20603 & w20604 ) ;
  assign w20606 = w20604 | w20605 ;
  assign w20607 = \pi072 ^ w20533 ;
  assign w20608 = ( ~w20548 & w20606 ) | ( ~w20548 & w20607 ) | ( w20606 & w20607 ) ;
  assign w20609 = w20607 | w20608 ;
  assign w20610 = \pi073 ^ w20540 ;
  assign w20611 = w20541 & ~w20610 ;
  assign w20612 = ( w20609 & w20610 ) | ( w20609 & ~w20611 ) | ( w20610 & ~w20611 ) ;
  assign w20613 = ~\pi073 & w20540 ;
  assign w20614 = w20612 & ~w20613 ;
  assign w20615 = w889 | w20614 ;
  assign w20616 = w20533 & w20615 ;
  assign w20617 = ~w20548 & w20606 ;
  assign w20618 = w20607 ^ w20617 ;
  assign w20619 = ~w20615 & w20618 ;
  assign w20620 = w20616 | w20619 ;
  assign w20621 = w20540 & w20615 ;
  assign w20622 = ~w20541 & w20609 ;
  assign w20623 = w20610 ^ w20622 ;
  assign w20624 = ~w20615 & w20623 ;
  assign w20625 = w20621 | w20624 ;
  assign w20626 = ~\pi073 & w20620 ;
  assign w20627 = w20547 & w20615 ;
  assign w20628 = ~w20555 & w20603 ;
  assign w20629 = w20604 ^ w20628 ;
  assign w20630 = ~w20615 & w20629 ;
  assign w20631 = w20627 | w20630 ;
  assign w20632 = ~\pi072 & w20631 ;
  assign w20633 = w20554 & w20615 ;
  assign w20634 = ~w20562 & w20600 ;
  assign w20635 = w20601 ^ w20634 ;
  assign w20636 = ~w20615 & w20635 ;
  assign w20637 = w20633 | w20636 ;
  assign w20638 = ~\pi071 & w20637 ;
  assign w20639 = w20561 & w20615 ;
  assign w20640 = ~w20569 & w20597 ;
  assign w20641 = w20598 ^ w20640 ;
  assign w20642 = ~w20615 & w20641 ;
  assign w20643 = w20639 | w20642 ;
  assign w20644 = ~\pi070 & w20643 ;
  assign w20645 = w20568 & w20615 ;
  assign w20646 = ~w20576 & w20594 ;
  assign w20647 = w20595 ^ w20646 ;
  assign w20648 = ~w20615 & w20647 ;
  assign w20649 = w20645 | w20648 ;
  assign w20650 = ~\pi069 & w20649 ;
  assign w20651 = w20575 & w20615 ;
  assign w20652 = ~w20586 & w20591 ;
  assign w20653 = w20592 ^ w20652 ;
  assign w20654 = ~w20615 & w20653 ;
  assign w20655 = w20651 | w20654 ;
  assign w20656 = ~\pi068 & w20655 ;
  assign w20657 = w20585 & w20615 ;
  assign w20658 = \pi064 & ~w20527 ;
  assign w20659 = \pi055 ^ w20658 ;
  assign w20660 = ( \pi065 & w856 ) | ( \pi065 & ~w20659 ) | ( w856 & ~w20659 ) ;
  assign w20661 = w20587 ^ w20660 ;
  assign w20662 = ( w889 & w20614 ) | ( w889 & w20661 ) | ( w20614 & w20661 ) ;
  assign w20663 = w20661 & ~w20662 ;
  assign w20664 = w20657 | w20663 ;
  assign w20665 = ~\pi067 & w20664 ;
  assign w20666 = \pi054 ^ w20527 ;
  assign w20667 = ( \pi064 & w889 ) | ( \pi064 & w20666 ) | ( w889 & w20666 ) ;
  assign w20668 = w939 ^ w20667 ;
  assign w20669 = ~w889 & w20668 ;
  assign w20670 = ~w20614 & w20669 ;
  assign w20671 = ( ~\pi064 & w20527 ) | ( ~\pi064 & w20615 ) | ( w20527 & w20615 ) ;
  assign w20672 = \pi055 ^ w20671 ;
  assign w20673 = w20615 & ~w20672 ;
  assign w20674 = w20670 | w20673 ;
  assign w20675 = ~\pi066 & w20674 ;
  assign w20676 = ( \pi054 & ~w955 ) | ( \pi054 & w20614 ) | ( ~w955 & w20614 ) ;
  assign w20677 = \pi054 & w20676 ;
  assign w20678 = w959 | w20614 ;
  assign w20679 = ( ~w20614 & w20677 ) | ( ~w20614 & w20678 ) | ( w20677 & w20678 ) ;
  assign w20680 = ( \pi065 & w959 ) | ( \pi065 & ~w20614 ) | ( w959 & ~w20614 ) ;
  assign w20681 = w955 & ~w20614 ;
  assign w20682 = ( \pi054 & \pi065 ) | ( \pi054 & ~w20681 ) | ( \pi065 & ~w20681 ) ;
  assign w20683 = w20680 | w20682 ;
  assign w20684 = \pi065 & w20679 ;
  assign w20685 = w20683 | w20684 ;
  assign w20686 = ( w968 & ~w20684 ) | ( w968 & w20685 ) | ( ~w20684 & w20685 ) ;
  assign w20687 = ~\pi065 & w20679 ;
  assign w20688 = w20615 | w20670 ;
  assign w20689 = ( w20659 & w20670 ) | ( w20659 & w20688 ) | ( w20670 & w20688 ) ;
  assign w20690 = \pi066 ^ w20689 ;
  assign w20691 = ( w20686 & ~w20687 ) | ( w20686 & w20690 ) | ( ~w20687 & w20690 ) ;
  assign w20692 = w20690 | w20691 ;
  assign w20693 = \pi067 ^ w20664 ;
  assign w20694 = ( ~w20675 & w20692 ) | ( ~w20675 & w20693 ) | ( w20692 & w20693 ) ;
  assign w20695 = w20693 | w20694 ;
  assign w20696 = \pi068 ^ w20655 ;
  assign w20697 = ( ~w20665 & w20695 ) | ( ~w20665 & w20696 ) | ( w20695 & w20696 ) ;
  assign w20698 = w20696 | w20697 ;
  assign w20699 = \pi069 ^ w20649 ;
  assign w20700 = ( ~w20656 & w20698 ) | ( ~w20656 & w20699 ) | ( w20698 & w20699 ) ;
  assign w20701 = w20699 | w20700 ;
  assign w20702 = \pi070 ^ w20643 ;
  assign w20703 = ( ~w20650 & w20701 ) | ( ~w20650 & w20702 ) | ( w20701 & w20702 ) ;
  assign w20704 = w20702 | w20703 ;
  assign w20705 = \pi071 ^ w20637 ;
  assign w20706 = ( ~w20644 & w20704 ) | ( ~w20644 & w20705 ) | ( w20704 & w20705 ) ;
  assign w20707 = w20705 | w20706 ;
  assign w20708 = \pi072 ^ w20631 ;
  assign w20709 = ( ~w20638 & w20707 ) | ( ~w20638 & w20708 ) | ( w20707 & w20708 ) ;
  assign w20710 = w20708 | w20709 ;
  assign w20711 = \pi073 ^ w20620 ;
  assign w20712 = ( ~w20632 & w20710 ) | ( ~w20632 & w20711 ) | ( w20710 & w20711 ) ;
  assign w20713 = w20711 | w20712 ;
  assign w20714 = \pi074 ^ w20625 ;
  assign w20715 = w20626 & ~w20714 ;
  assign w20716 = ( w20713 & w20714 ) | ( w20713 & ~w20715 ) | ( w20714 & ~w20715 ) ;
  assign w20717 = ~\pi074 & w20625 ;
  assign w20718 = w20716 & ~w20717 ;
  assign w20719 = w1007 | w20718 ;
  assign w20720 = w20620 & w20719 ;
  assign w20721 = ~w20632 & w20710 ;
  assign w20722 = w20711 ^ w20721 ;
  assign w20723 = ~w20719 & w20722 ;
  assign w20724 = w20720 | w20723 ;
  assign w20725 = ~\pi074 & w20724 ;
  assign w20726 = w20631 & w20719 ;
  assign w20727 = ~w20638 & w20707 ;
  assign w20728 = w20708 ^ w20727 ;
  assign w20729 = ~w20719 & w20728 ;
  assign w20730 = w20726 | w20729 ;
  assign w20731 = ~\pi073 & w20730 ;
  assign w20732 = w20637 & w20719 ;
  assign w20733 = ~w20644 & w20704 ;
  assign w20734 = w20705 ^ w20733 ;
  assign w20735 = ~w20719 & w20734 ;
  assign w20736 = w20732 | w20735 ;
  assign w20737 = ~\pi072 & w20736 ;
  assign w20738 = w20643 & w20719 ;
  assign w20739 = ~w20650 & w20701 ;
  assign w20740 = w20702 ^ w20739 ;
  assign w20741 = ~w20719 & w20740 ;
  assign w20742 = w20738 | w20741 ;
  assign w20743 = ~\pi071 & w20742 ;
  assign w20744 = w20649 & w20719 ;
  assign w20745 = ~w20656 & w20698 ;
  assign w20746 = w20699 ^ w20745 ;
  assign w20747 = ~w20719 & w20746 ;
  assign w20748 = w20744 | w20747 ;
  assign w20749 = ~\pi070 & w20748 ;
  assign w20750 = w20655 & w20719 ;
  assign w20751 = ~w20665 & w20695 ;
  assign w20752 = w20696 ^ w20751 ;
  assign w20753 = ~w20719 & w20752 ;
  assign w20754 = w20750 | w20753 ;
  assign w20755 = ~\pi069 & w20754 ;
  assign w20756 = w20664 & w20719 ;
  assign w20757 = ~w20675 & w20692 ;
  assign w20758 = w20693 ^ w20757 ;
  assign w20759 = ~w20719 & w20758 ;
  assign w20760 = w20756 | w20759 ;
  assign w20761 = ~\pi068 & w20760 ;
  assign w20762 = w20674 & w20719 ;
  assign w20763 = w20686 & ~w20687 ;
  assign w20764 = w20690 ^ w20763 ;
  assign w20765 = ~w20719 & w20764 ;
  assign w20766 = w20762 | w20765 ;
  assign w20767 = ~\pi067 & w20766 ;
  assign w20768 = w20679 & w20719 ;
  assign w20769 = ~w20679 & w20683 ;
  assign w20770 = ( ~\pi065 & w20683 ) | ( ~\pi065 & w20769 ) | ( w20683 & w20769 ) ;
  assign w20771 = w968 ^ w20770 ;
  assign w20772 = ~w20719 & w20771 ;
  assign w20773 = w20768 | w20772 ;
  assign w20774 = ~\pi066 & w20773 ;
  assign w20775 = ( \pi053 & ~w1066 ) | ( \pi053 & w20718 ) | ( ~w1066 & w20718 ) ;
  assign w20776 = \pi053 & w20775 ;
  assign w20777 = w1070 | w20718 ;
  assign w20778 = ( ~w20718 & w20776 ) | ( ~w20718 & w20777 ) | ( w20776 & w20777 ) ;
  assign w20779 = w1066 & ~w20777 ;
  assign w20780 = \pi053 & ~w20779 ;
  assign w20781 = ( ~w20718 & w20777 ) | ( ~w20718 & w20780 ) | ( w20777 & w20780 ) ;
  assign w20782 = \pi065 ^ w20781 ;
  assign w20783 = w1075 | w20782 ;
  assign w20784 = ~\pi065 & w20778 ;
  assign w20785 = \pi066 ^ w20773 ;
  assign w20786 = ( w20783 & ~w20784 ) | ( w20783 & w20785 ) | ( ~w20784 & w20785 ) ;
  assign w20787 = w20785 | w20786 ;
  assign w20788 = \pi067 ^ w20766 ;
  assign w20789 = ( ~w20774 & w20787 ) | ( ~w20774 & w20788 ) | ( w20787 & w20788 ) ;
  assign w20790 = w20788 | w20789 ;
  assign w20791 = \pi068 ^ w20760 ;
  assign w20792 = ( ~w20767 & w20790 ) | ( ~w20767 & w20791 ) | ( w20790 & w20791 ) ;
  assign w20793 = w20791 | w20792 ;
  assign w20794 = \pi069 ^ w20754 ;
  assign w20795 = ( ~w20761 & w20793 ) | ( ~w20761 & w20794 ) | ( w20793 & w20794 ) ;
  assign w20796 = w20794 | w20795 ;
  assign w20797 = \pi070 ^ w20748 ;
  assign w20798 = ( ~w20755 & w20796 ) | ( ~w20755 & w20797 ) | ( w20796 & w20797 ) ;
  assign w20799 = w20797 | w20798 ;
  assign w20800 = \pi071 ^ w20742 ;
  assign w20801 = ( ~w20749 & w20799 ) | ( ~w20749 & w20800 ) | ( w20799 & w20800 ) ;
  assign w20802 = w20800 | w20801 ;
  assign w20803 = \pi072 ^ w20736 ;
  assign w20804 = ( ~w20743 & w20802 ) | ( ~w20743 & w20803 ) | ( w20802 & w20803 ) ;
  assign w20805 = w20803 | w20804 ;
  assign w20806 = \pi073 ^ w20730 ;
  assign w20807 = ( ~w20737 & w20805 ) | ( ~w20737 & w20806 ) | ( w20805 & w20806 ) ;
  assign w20808 = w20806 | w20807 ;
  assign w20809 = \pi074 ^ w20724 ;
  assign w20810 = ( ~w20731 & w20808 ) | ( ~w20731 & w20809 ) | ( w20808 & w20809 ) ;
  assign w20811 = w20809 | w20810 ;
  assign w20812 = w20625 & w20719 ;
  assign w20813 = ~w20626 & w20713 ;
  assign w20814 = w20714 ^ w20813 ;
  assign w20815 = ~w20719 & w20814 ;
  assign w20816 = w20812 | w20815 ;
  assign w20817 = ~\pi075 & w20816 ;
  assign w20818 = ( \pi075 & ~w20812 ) | ( \pi075 & w20815 ) | ( ~w20812 & w20815 ) ;
  assign w20819 = ~w20815 & w20818 ;
  assign w20820 = w1117 | w20819 ;
  assign w20821 = ( w368 & w20817 ) | ( w368 & ~w20819 ) | ( w20817 & ~w20819 ) ;
  assign w20822 = w20820 | w20821 ;
  assign w20823 = ( ~w20725 & w20811 ) | ( ~w20725 & w20822 ) | ( w20811 & w20822 ) ;
  assign w20824 = w20822 | w20823 ;
  assign w20825 = ~w1007 & w20816 ;
  assign w20826 = w20824 & ~w20825 ;
  assign w20827 = ~w20731 & w20808 ;
  assign w20828 = w20809 ^ w20827 ;
  assign w20829 = ~w20826 & w20828 ;
  assign w20830 = ( w20724 & w20824 ) | ( w20724 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20831 = ~w20825 & w20830 ;
  assign w20832 = w20829 | w20831 ;
  assign w20833 = w20817 | w20819 ;
  assign w20834 = ( ~w20725 & w20811 ) | ( ~w20725 & w20826 ) | ( w20811 & w20826 ) ;
  assign w20835 = w20833 ^ w20834 ;
  assign w20836 = ~w20826 & w20835 ;
  assign w20837 = ( w1007 & ~w20816 ) | ( w1007 & w20824 ) | ( ~w20816 & w20824 ) ;
  assign w20838 = w20816 & w20837 ;
  assign w20839 = w20836 | w20838 ;
  assign w20840 = ~\pi075 & w20832 ;
  assign w20841 = ~w20737 & w20805 ;
  assign w20842 = w20806 ^ w20841 ;
  assign w20843 = ~w20826 & w20842 ;
  assign w20844 = ( w20730 & w20824 ) | ( w20730 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20845 = ~w20825 & w20844 ;
  assign w20846 = w20843 | w20845 ;
  assign w20847 = ~\pi074 & w20846 ;
  assign w20848 = ~w20743 & w20802 ;
  assign w20849 = w20803 ^ w20848 ;
  assign w20850 = ~w20826 & w20849 ;
  assign w20851 = ( w20736 & w20824 ) | ( w20736 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20852 = ~w20825 & w20851 ;
  assign w20853 = w20850 | w20852 ;
  assign w20854 = ~\pi073 & w20853 ;
  assign w20855 = ~w20749 & w20799 ;
  assign w20856 = w20800 ^ w20855 ;
  assign w20857 = ~w20826 & w20856 ;
  assign w20858 = ( w20742 & w20824 ) | ( w20742 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20859 = ~w20825 & w20858 ;
  assign w20860 = w20857 | w20859 ;
  assign w20861 = ~\pi072 & w20860 ;
  assign w20862 = ~w20755 & w20796 ;
  assign w20863 = w20797 ^ w20862 ;
  assign w20864 = ~w20826 & w20863 ;
  assign w20865 = ( w20748 & w20824 ) | ( w20748 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20866 = ~w20825 & w20865 ;
  assign w20867 = w20864 | w20866 ;
  assign w20868 = ~\pi071 & w20867 ;
  assign w20869 = ~w20761 & w20793 ;
  assign w20870 = w20794 ^ w20869 ;
  assign w20871 = ~w20826 & w20870 ;
  assign w20872 = ( w20754 & w20824 ) | ( w20754 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20873 = ~w20825 & w20872 ;
  assign w20874 = w20871 | w20873 ;
  assign w20875 = ~\pi070 & w20874 ;
  assign w20876 = ~w20767 & w20790 ;
  assign w20877 = w20791 ^ w20876 ;
  assign w20878 = ~w20826 & w20877 ;
  assign w20879 = ( w20760 & w20824 ) | ( w20760 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20880 = ~w20825 & w20879 ;
  assign w20881 = w20878 | w20880 ;
  assign w20882 = ~\pi069 & w20881 ;
  assign w20883 = ~w20774 & w20787 ;
  assign w20884 = w20788 ^ w20883 ;
  assign w20885 = ~w20826 & w20884 ;
  assign w20886 = ( w20766 & w20824 ) | ( w20766 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20887 = ~w20825 & w20886 ;
  assign w20888 = w20885 | w20887 ;
  assign w20889 = ~\pi068 & w20888 ;
  assign w20890 = w20783 & ~w20784 ;
  assign w20891 = w20785 ^ w20890 ;
  assign w20892 = ~w20826 & w20891 ;
  assign w20893 = ( w20773 & w20824 ) | ( w20773 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20894 = ~w20825 & w20893 ;
  assign w20895 = w20892 | w20894 ;
  assign w20896 = ~\pi067 & w20895 ;
  assign w20897 = w1070 ^ w20718 ;
  assign w20898 = ( \pi053 & ~w1195 ) | ( \pi053 & w20897 ) | ( ~w1195 & w20897 ) ;
  assign w20899 = ( \pi053 & w1070 ) | ( \pi053 & w20898 ) | ( w1070 & w20898 ) ;
  assign w20900 = w1075 ^ w20899 ;
  assign w20901 = \pi065 ^ w20900 ;
  assign w20902 = ~w20826 & w20901 ;
  assign w20903 = ( w20778 & w20824 ) | ( w20778 & w20825 ) | ( w20824 & w20825 ) ;
  assign w20904 = ~w20825 & w20903 ;
  assign w20905 = w20902 | w20904 ;
  assign w20906 = ~\pi066 & w20905 ;
  assign w20907 = \pi066 ^ w20905 ;
  assign w20908 = ( \pi064 & ~w20826 ) | ( \pi064 & w20907 ) | ( ~w20826 & w20907 ) ;
  assign w20909 = \pi052 ^ w20908 ;
  assign w20910 = ( \pi065 & w1307 ) | ( \pi065 & ~w20909 ) | ( w1307 & ~w20909 ) ;
  assign w20911 = w20907 | w20910 ;
  assign w20912 = \pi067 ^ w20895 ;
  assign w20913 = ( ~w20906 & w20911 ) | ( ~w20906 & w20912 ) | ( w20911 & w20912 ) ;
  assign w20914 = w20912 | w20913 ;
  assign w20915 = \pi068 ^ w20888 ;
  assign w20916 = ( ~w20896 & w20914 ) | ( ~w20896 & w20915 ) | ( w20914 & w20915 ) ;
  assign w20917 = w20915 | w20916 ;
  assign w20918 = \pi069 ^ w20881 ;
  assign w20919 = ( ~w20889 & w20917 ) | ( ~w20889 & w20918 ) | ( w20917 & w20918 ) ;
  assign w20920 = w20918 | w20919 ;
  assign w20921 = \pi070 ^ w20874 ;
  assign w20922 = ( ~w20882 & w20920 ) | ( ~w20882 & w20921 ) | ( w20920 & w20921 ) ;
  assign w20923 = w20921 | w20922 ;
  assign w20924 = \pi071 ^ w20867 ;
  assign w20925 = ( ~w20875 & w20923 ) | ( ~w20875 & w20924 ) | ( w20923 & w20924 ) ;
  assign w20926 = w20924 | w20925 ;
  assign w20927 = \pi072 ^ w20860 ;
  assign w20928 = ( ~w20868 & w20926 ) | ( ~w20868 & w20927 ) | ( w20926 & w20927 ) ;
  assign w20929 = w20927 | w20928 ;
  assign w20930 = \pi073 ^ w20853 ;
  assign w20931 = ( ~w20861 & w20929 ) | ( ~w20861 & w20930 ) | ( w20929 & w20930 ) ;
  assign w20932 = w20930 | w20931 ;
  assign w20933 = \pi074 ^ w20846 ;
  assign w20934 = ( ~w20854 & w20932 ) | ( ~w20854 & w20933 ) | ( w20932 & w20933 ) ;
  assign w20935 = w20933 | w20934 ;
  assign w20936 = \pi075 ^ w20832 ;
  assign w20937 = ( ~w20847 & w20935 ) | ( ~w20847 & w20936 ) | ( w20935 & w20936 ) ;
  assign w20938 = w20936 | w20937 ;
  assign w20939 = \pi076 ^ w20839 ;
  assign w20940 = w20840 & ~w20939 ;
  assign w20941 = ( w20938 & w20939 ) | ( w20938 & ~w20940 ) | ( w20939 & ~w20940 ) ;
  assign w20942 = ~\pi076 & w20839 ;
  assign w20943 = w20941 & ~w20942 ;
  assign w20944 = w1245 | w20943 ;
  assign w20945 = w20832 & w20944 ;
  assign w20946 = ~w20847 & w20935 ;
  assign w20947 = w20936 ^ w20946 ;
  assign w20948 = ~w20944 & w20947 ;
  assign w20949 = w20945 | w20948 ;
  assign w20950 = w20839 & w20944 ;
  assign w20951 = ~w20840 & w20938 ;
  assign w20952 = w20939 ^ w20951 ;
  assign w20953 = ~w20944 & w20952 ;
  assign w20954 = w20950 | w20953 ;
  assign w20955 = ~\pi076 & w20949 ;
  assign w20956 = w20846 & w20944 ;
  assign w20957 = ~w20854 & w20932 ;
  assign w20958 = w20933 ^ w20957 ;
  assign w20959 = ~w20944 & w20958 ;
  assign w20960 = w20956 | w20959 ;
  assign w20961 = ~\pi075 & w20960 ;
  assign w20962 = w20853 & w20944 ;
  assign w20963 = ~w20861 & w20929 ;
  assign w20964 = w20930 ^ w20963 ;
  assign w20965 = ~w20944 & w20964 ;
  assign w20966 = w20962 | w20965 ;
  assign w20967 = ~\pi074 & w20966 ;
  assign w20968 = w20860 & w20944 ;
  assign w20969 = ~w20868 & w20926 ;
  assign w20970 = w20927 ^ w20969 ;
  assign w20971 = ~w20944 & w20970 ;
  assign w20972 = w20968 | w20971 ;
  assign w20973 = ~\pi073 & w20972 ;
  assign w20974 = w20867 & w20944 ;
  assign w20975 = ~w20875 & w20923 ;
  assign w20976 = w20924 ^ w20975 ;
  assign w20977 = ~w20944 & w20976 ;
  assign w20978 = w20974 | w20977 ;
  assign w20979 = ~\pi072 & w20978 ;
  assign w20980 = w20874 & w20944 ;
  assign w20981 = ~w20882 & w20920 ;
  assign w20982 = w20921 ^ w20981 ;
  assign w20983 = ~w20944 & w20982 ;
  assign w20984 = w20980 | w20983 ;
  assign w20985 = ~\pi071 & w20984 ;
  assign w20986 = w20881 & w20944 ;
  assign w20987 = ~w20889 & w20917 ;
  assign w20988 = w20918 ^ w20987 ;
  assign w20989 = ~w20944 & w20988 ;
  assign w20990 = w20986 | w20989 ;
  assign w20991 = ~\pi070 & w20990 ;
  assign w20992 = w20888 & w20944 ;
  assign w20993 = ~w20896 & w20914 ;
  assign w20994 = w20915 ^ w20993 ;
  assign w20995 = ~w20944 & w20994 ;
  assign w20996 = w20992 | w20995 ;
  assign w20997 = ~\pi069 & w20996 ;
  assign w20998 = w20895 & w20944 ;
  assign w20999 = ~w20906 & w20911 ;
  assign w21000 = w20912 ^ w20999 ;
  assign w21001 = ~w20944 & w21000 ;
  assign w21002 = w20998 | w21001 ;
  assign w21003 = ~\pi068 & w21002 ;
  assign w21004 = w20905 & w20944 ;
  assign w21005 = \pi064 & ~w20826 ;
  assign w21006 = \pi052 ^ w21005 ;
  assign w21007 = ( \pi065 & w1307 ) | ( \pi065 & ~w21006 ) | ( w1307 & ~w21006 ) ;
  assign w21008 = w20907 ^ w21007 ;
  assign w21009 = ( w1245 & w20943 ) | ( w1245 & w21008 ) | ( w20943 & w21008 ) ;
  assign w21010 = w21008 & ~w21009 ;
  assign w21011 = w21004 | w21010 ;
  assign w21012 = ~\pi067 & w21011 ;
  assign w21013 = \pi051 ^ w20826 ;
  assign w21014 = ( \pi064 & w1245 ) | ( \pi064 & w21013 ) | ( w1245 & w21013 ) ;
  assign w21015 = w1314 ^ w21014 ;
  assign w21016 = ~w1245 & w21015 ;
  assign w21017 = ~w20943 & w21016 ;
  assign w21018 = ( ~\pi064 & w20826 ) | ( ~\pi064 & w20944 ) | ( w20826 & w20944 ) ;
  assign w21019 = \pi052 ^ w21018 ;
  assign w21020 = w20944 & ~w21019 ;
  assign w21021 = w21017 | w21020 ;
  assign w21022 = ~\pi066 & w21021 ;
  assign w21023 = ( \pi051 & ~w1330 ) | ( \pi051 & w20943 ) | ( ~w1330 & w20943 ) ;
  assign w21024 = \pi051 & w21023 ;
  assign w21025 = w1334 & ~w20943 ;
  assign w21026 = w21024 | w21025 ;
  assign w21027 = \pi065 ^ w21026 ;
  assign w21028 = w1337 | w21027 ;
  assign w21029 = ~\pi065 & w21026 ;
  assign w21030 = w20944 | w21017 ;
  assign w21031 = ( w21006 & w21017 ) | ( w21006 & w21030 ) | ( w21017 & w21030 ) ;
  assign w21032 = \pi066 ^ w21031 ;
  assign w21033 = ( w21028 & ~w21029 ) | ( w21028 & w21032 ) | ( ~w21029 & w21032 ) ;
  assign w21034 = w21032 | w21033 ;
  assign w21035 = \pi067 ^ w21011 ;
  assign w21036 = ( ~w21022 & w21034 ) | ( ~w21022 & w21035 ) | ( w21034 & w21035 ) ;
  assign w21037 = w21035 | w21036 ;
  assign w21038 = \pi068 ^ w21002 ;
  assign w21039 = ( ~w21012 & w21037 ) | ( ~w21012 & w21038 ) | ( w21037 & w21038 ) ;
  assign w21040 = w21038 | w21039 ;
  assign w21041 = \pi069 ^ w20996 ;
  assign w21042 = ( ~w21003 & w21040 ) | ( ~w21003 & w21041 ) | ( w21040 & w21041 ) ;
  assign w21043 = w21041 | w21042 ;
  assign w21044 = \pi070 ^ w20990 ;
  assign w21045 = ( ~w20997 & w21043 ) | ( ~w20997 & w21044 ) | ( w21043 & w21044 ) ;
  assign w21046 = w21044 | w21045 ;
  assign w21047 = \pi071 ^ w20984 ;
  assign w21048 = ( ~w20991 & w21046 ) | ( ~w20991 & w21047 ) | ( w21046 & w21047 ) ;
  assign w21049 = w21047 | w21048 ;
  assign w21050 = \pi072 ^ w20978 ;
  assign w21051 = ( ~w20985 & w21049 ) | ( ~w20985 & w21050 ) | ( w21049 & w21050 ) ;
  assign w21052 = w21050 | w21051 ;
  assign w21053 = \pi073 ^ w20972 ;
  assign w21054 = ( ~w20979 & w21052 ) | ( ~w20979 & w21053 ) | ( w21052 & w21053 ) ;
  assign w21055 = w21053 | w21054 ;
  assign w21056 = \pi074 ^ w20966 ;
  assign w21057 = ( ~w20973 & w21055 ) | ( ~w20973 & w21056 ) | ( w21055 & w21056 ) ;
  assign w21058 = w21056 | w21057 ;
  assign w21059 = \pi075 ^ w20960 ;
  assign w21060 = ( ~w20967 & w21058 ) | ( ~w20967 & w21059 ) | ( w21058 & w21059 ) ;
  assign w21061 = w21059 | w21060 ;
  assign w21062 = \pi076 ^ w20949 ;
  assign w21063 = ( ~w20961 & w21061 ) | ( ~w20961 & w21062 ) | ( w21061 & w21062 ) ;
  assign w21064 = w21062 | w21063 ;
  assign w21065 = \pi077 ^ w20954 ;
  assign w21066 = w20955 & ~w21065 ;
  assign w21067 = ( w21064 & w21065 ) | ( w21064 & ~w21066 ) | ( w21065 & ~w21066 ) ;
  assign w21068 = ~\pi077 & w20954 ;
  assign w21069 = w21067 & ~w21068 ;
  assign w21070 = w1384 | w21069 ;
  assign w21071 = w20949 & w21070 ;
  assign w21072 = ~w20961 & w21061 ;
  assign w21073 = w21062 ^ w21072 ;
  assign w21074 = ~w21070 & w21073 ;
  assign w21075 = w21071 | w21074 ;
  assign w21076 = ~\pi077 & w21075 ;
  assign w21077 = w20960 & w21070 ;
  assign w21078 = ~w20967 & w21058 ;
  assign w21079 = w21059 ^ w21078 ;
  assign w21080 = ~w21070 & w21079 ;
  assign w21081 = w21077 | w21080 ;
  assign w21082 = ~\pi076 & w21081 ;
  assign w21083 = w20966 & w21070 ;
  assign w21084 = ~w20973 & w21055 ;
  assign w21085 = w21056 ^ w21084 ;
  assign w21086 = ~w21070 & w21085 ;
  assign w21087 = w21083 | w21086 ;
  assign w21088 = ~\pi075 & w21087 ;
  assign w21089 = w20972 & w21070 ;
  assign w21090 = ~w20979 & w21052 ;
  assign w21091 = w21053 ^ w21090 ;
  assign w21092 = ~w21070 & w21091 ;
  assign w21093 = w21089 | w21092 ;
  assign w21094 = ~\pi074 & w21093 ;
  assign w21095 = w20978 & w21070 ;
  assign w21096 = ~w20985 & w21049 ;
  assign w21097 = w21050 ^ w21096 ;
  assign w21098 = ~w21070 & w21097 ;
  assign w21099 = w21095 | w21098 ;
  assign w21100 = ~\pi073 & w21099 ;
  assign w21101 = w20984 & w21070 ;
  assign w21102 = ~w20991 & w21046 ;
  assign w21103 = w21047 ^ w21102 ;
  assign w21104 = ~w21070 & w21103 ;
  assign w21105 = w21101 | w21104 ;
  assign w21106 = ~\pi072 & w21105 ;
  assign w21107 = w20990 & w21070 ;
  assign w21108 = ~w20997 & w21043 ;
  assign w21109 = w21044 ^ w21108 ;
  assign w21110 = ~w21070 & w21109 ;
  assign w21111 = w21107 | w21110 ;
  assign w21112 = ~\pi071 & w21111 ;
  assign w21113 = w20996 & w21070 ;
  assign w21114 = ~w21003 & w21040 ;
  assign w21115 = w21041 ^ w21114 ;
  assign w21116 = ~w21070 & w21115 ;
  assign w21117 = w21113 | w21116 ;
  assign w21118 = ~\pi070 & w21117 ;
  assign w21119 = w21002 & w21070 ;
  assign w21120 = ~w21012 & w21037 ;
  assign w21121 = w21038 ^ w21120 ;
  assign w21122 = ~w21070 & w21121 ;
  assign w21123 = w21119 | w21122 ;
  assign w21124 = ~\pi069 & w21123 ;
  assign w21125 = w21011 & w21070 ;
  assign w21126 = ~w21022 & w21034 ;
  assign w21127 = w21035 ^ w21126 ;
  assign w21128 = ~w21070 & w21127 ;
  assign w21129 = w21125 | w21128 ;
  assign w21130 = ~\pi068 & w21129 ;
  assign w21131 = w21021 & w21070 ;
  assign w21132 = w21028 & ~w21029 ;
  assign w21133 = w21032 ^ w21132 ;
  assign w21134 = ~w21070 & w21133 ;
  assign w21135 = w21131 | w21134 ;
  assign w21136 = ~\pi067 & w21135 ;
  assign w21137 = w21026 & w21070 ;
  assign w21138 = ( ~w1384 & w21024 ) | ( ~w1384 & w21025 ) | ( w21024 & w21025 ) ;
  assign w21139 = \pi065 ^ w21138 ;
  assign w21140 = ( w1337 & ~w1384 ) | ( w1337 & w21139 ) | ( ~w1384 & w21139 ) ;
  assign w21141 = ( w1337 & w21069 ) | ( w1337 & w21139 ) | ( w21069 & w21139 ) ;
  assign w21142 = w21140 & ~w21141 ;
  assign w21143 = w21137 | w21142 ;
  assign w21144 = ~\pi066 & w21143 ;
  assign w21145 = ( \pi050 & ~w1465 ) | ( \pi050 & w21069 ) | ( ~w1465 & w21069 ) ;
  assign w21146 = \pi050 & w21145 ;
  assign w21147 = w1469 | w21069 ;
  assign w21148 = ( ~w21069 & w21146 ) | ( ~w21069 & w21147 ) | ( w21146 & w21147 ) ;
  assign w21149 = w1465 & ~w21147 ;
  assign w21150 = \pi050 & ~w21149 ;
  assign w21151 = ( ~w21069 & w21147 ) | ( ~w21069 & w21150 ) | ( w21147 & w21150 ) ;
  assign w21152 = \pi065 ^ w21151 ;
  assign w21153 = w1474 | w21152 ;
  assign w21154 = ~\pi065 & w21148 ;
  assign w21155 = \pi066 ^ w21143 ;
  assign w21156 = ( w21153 & ~w21154 ) | ( w21153 & w21155 ) | ( ~w21154 & w21155 ) ;
  assign w21157 = w21155 | w21156 ;
  assign w21158 = \pi067 ^ w21135 ;
  assign w21159 = ( ~w21144 & w21157 ) | ( ~w21144 & w21158 ) | ( w21157 & w21158 ) ;
  assign w21160 = w21158 | w21159 ;
  assign w21161 = \pi068 ^ w21129 ;
  assign w21162 = ( ~w21136 & w21160 ) | ( ~w21136 & w21161 ) | ( w21160 & w21161 ) ;
  assign w21163 = w21161 | w21162 ;
  assign w21164 = \pi069 ^ w21123 ;
  assign w21165 = ( ~w21130 & w21163 ) | ( ~w21130 & w21164 ) | ( w21163 & w21164 ) ;
  assign w21166 = w21164 | w21165 ;
  assign w21167 = \pi070 ^ w21117 ;
  assign w21168 = ( ~w21124 & w21166 ) | ( ~w21124 & w21167 ) | ( w21166 & w21167 ) ;
  assign w21169 = w21167 | w21168 ;
  assign w21170 = \pi071 ^ w21111 ;
  assign w21171 = ( ~w21118 & w21169 ) | ( ~w21118 & w21170 ) | ( w21169 & w21170 ) ;
  assign w21172 = w21170 | w21171 ;
  assign w21173 = \pi072 ^ w21105 ;
  assign w21174 = ( ~w21112 & w21172 ) | ( ~w21112 & w21173 ) | ( w21172 & w21173 ) ;
  assign w21175 = w21173 | w21174 ;
  assign w21176 = \pi073 ^ w21099 ;
  assign w21177 = ( ~w21106 & w21175 ) | ( ~w21106 & w21176 ) | ( w21175 & w21176 ) ;
  assign w21178 = w21176 | w21177 ;
  assign w21179 = \pi074 ^ w21093 ;
  assign w21180 = ( ~w21100 & w21178 ) | ( ~w21100 & w21179 ) | ( w21178 & w21179 ) ;
  assign w21181 = w21179 | w21180 ;
  assign w21182 = \pi075 ^ w21087 ;
  assign w21183 = ( ~w21094 & w21181 ) | ( ~w21094 & w21182 ) | ( w21181 & w21182 ) ;
  assign w21184 = w21182 | w21183 ;
  assign w21185 = \pi076 ^ w21081 ;
  assign w21186 = ( ~w21088 & w21184 ) | ( ~w21088 & w21185 ) | ( w21184 & w21185 ) ;
  assign w21187 = w21185 | w21186 ;
  assign w21188 = \pi077 ^ w21075 ;
  assign w21189 = ( ~w21082 & w21187 ) | ( ~w21082 & w21188 ) | ( w21187 & w21188 ) ;
  assign w21190 = w21188 | w21189 ;
  assign w21191 = w20954 & w21070 ;
  assign w21192 = ~w20955 & w21064 ;
  assign w21193 = w21065 ^ w21192 ;
  assign w21194 = ~w21070 & w21193 ;
  assign w21195 = w21191 | w21194 ;
  assign w21196 = ~\pi078 & w21195 ;
  assign w21197 = ( \pi078 & ~w21191 ) | ( \pi078 & w21194 ) | ( ~w21191 & w21194 ) ;
  assign w21198 = ~w21194 & w21197 ;
  assign w21199 = w21196 | w21198 ;
  assign w21200 = ( ~w21076 & w21190 ) | ( ~w21076 & w21199 ) | ( w21190 & w21199 ) ;
  assign w21201 = ( w1528 & ~w21199 ) | ( w1528 & w21200 ) | ( ~w21199 & w21200 ) ;
  assign w21202 = w21199 | w21201 ;
  assign w21203 = ~w1384 & w21195 ;
  assign w21204 = w21202 & ~w21203 ;
  assign w21205 = ~w21082 & w21187 ;
  assign w21206 = w21188 ^ w21205 ;
  assign w21207 = ~w21204 & w21206 ;
  assign w21208 = ( w21075 & w21202 ) | ( w21075 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21209 = ~w21203 & w21208 ;
  assign w21210 = w21207 | w21209 ;
  assign w21211 = ( ~w21076 & w21190 ) | ( ~w21076 & w21204 ) | ( w21190 & w21204 ) ;
  assign w21212 = w21199 ^ w21211 ;
  assign w21213 = ~w21204 & w21212 ;
  assign w21214 = ( w1384 & ~w21195 ) | ( w1384 & w21202 ) | ( ~w21195 & w21202 ) ;
  assign w21215 = w21195 & w21214 ;
  assign w21216 = w21213 | w21215 ;
  assign w21217 = ~\pi078 & w21210 ;
  assign w21218 = ~w21088 & w21184 ;
  assign w21219 = w21185 ^ w21218 ;
  assign w21220 = ~w21204 & w21219 ;
  assign w21221 = ( w21081 & w21202 ) | ( w21081 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21222 = ~w21203 & w21221 ;
  assign w21223 = w21220 | w21222 ;
  assign w21224 = ~\pi077 & w21223 ;
  assign w21225 = ~w21094 & w21181 ;
  assign w21226 = w21182 ^ w21225 ;
  assign w21227 = ~w21204 & w21226 ;
  assign w21228 = ( w21087 & w21202 ) | ( w21087 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21229 = ~w21203 & w21228 ;
  assign w21230 = w21227 | w21229 ;
  assign w21231 = ~\pi076 & w21230 ;
  assign w21232 = ~w21100 & w21178 ;
  assign w21233 = w21179 ^ w21232 ;
  assign w21234 = ~w21204 & w21233 ;
  assign w21235 = ( w21093 & w21202 ) | ( w21093 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21236 = ~w21203 & w21235 ;
  assign w21237 = w21234 | w21236 ;
  assign w21238 = ~\pi075 & w21237 ;
  assign w21239 = ~w21106 & w21175 ;
  assign w21240 = w21176 ^ w21239 ;
  assign w21241 = ~w21204 & w21240 ;
  assign w21242 = ( w21099 & w21202 ) | ( w21099 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21243 = ~w21203 & w21242 ;
  assign w21244 = w21241 | w21243 ;
  assign w21245 = ~\pi074 & w21244 ;
  assign w21246 = ~w21112 & w21172 ;
  assign w21247 = w21173 ^ w21246 ;
  assign w21248 = ~w21204 & w21247 ;
  assign w21249 = ( w21105 & w21202 ) | ( w21105 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21250 = ~w21203 & w21249 ;
  assign w21251 = w21248 | w21250 ;
  assign w21252 = ~\pi073 & w21251 ;
  assign w21253 = ~w21118 & w21169 ;
  assign w21254 = w21170 ^ w21253 ;
  assign w21255 = ~w21204 & w21254 ;
  assign w21256 = ( w21111 & w21202 ) | ( w21111 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21257 = ~w21203 & w21256 ;
  assign w21258 = w21255 | w21257 ;
  assign w21259 = ~\pi072 & w21258 ;
  assign w21260 = ~w21124 & w21166 ;
  assign w21261 = w21167 ^ w21260 ;
  assign w21262 = ~w21204 & w21261 ;
  assign w21263 = ( w21117 & w21202 ) | ( w21117 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21264 = ~w21203 & w21263 ;
  assign w21265 = w21262 | w21264 ;
  assign w21266 = ~\pi071 & w21265 ;
  assign w21267 = ~w21130 & w21163 ;
  assign w21268 = w21164 ^ w21267 ;
  assign w21269 = ~w21204 & w21268 ;
  assign w21270 = ( w21123 & w21202 ) | ( w21123 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21271 = ~w21203 & w21270 ;
  assign w21272 = w21269 | w21271 ;
  assign w21273 = ~\pi070 & w21272 ;
  assign w21274 = ~w21136 & w21160 ;
  assign w21275 = w21161 ^ w21274 ;
  assign w21276 = ~w21204 & w21275 ;
  assign w21277 = ( w21129 & w21202 ) | ( w21129 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21278 = ~w21203 & w21277 ;
  assign w21279 = w21276 | w21278 ;
  assign w21280 = ~\pi069 & w21279 ;
  assign w21281 = ~w21144 & w21157 ;
  assign w21282 = w21158 ^ w21281 ;
  assign w21283 = ~w21204 & w21282 ;
  assign w21284 = ( w21135 & w21202 ) | ( w21135 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21285 = ~w21203 & w21284 ;
  assign w21286 = w21283 | w21285 ;
  assign w21287 = ~\pi068 & w21286 ;
  assign w21288 = w21153 & ~w21154 ;
  assign w21289 = w21155 ^ w21288 ;
  assign w21290 = ~w21204 & w21289 ;
  assign w21291 = ( w21143 & w21202 ) | ( w21143 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21292 = ~w21203 & w21291 ;
  assign w21293 = w21290 | w21292 ;
  assign w21294 = ~\pi067 & w21293 ;
  assign w21295 = w1469 ^ w21069 ;
  assign w21296 = ( \pi050 & ~w1625 ) | ( \pi050 & w21295 ) | ( ~w1625 & w21295 ) ;
  assign w21297 = ( \pi050 & w1469 ) | ( \pi050 & w21296 ) | ( w1469 & w21296 ) ;
  assign w21298 = w1474 ^ w21297 ;
  assign w21299 = \pi065 ^ w21298 ;
  assign w21300 = ~w21204 & w21299 ;
  assign w21301 = ( w21148 & w21202 ) | ( w21148 & w21203 ) | ( w21202 & w21203 ) ;
  assign w21302 = ~w21203 & w21301 ;
  assign w21303 = w21300 | w21302 ;
  assign w21304 = ~\pi066 & w21303 ;
  assign w21305 = \pi066 ^ w21303 ;
  assign w21306 = ( \pi064 & ~w21204 ) | ( \pi064 & w21305 ) | ( ~w21204 & w21305 ) ;
  assign w21307 = \pi049 ^ w21306 ;
  assign w21308 = ( \pi065 & w1762 ) | ( \pi065 & ~w21307 ) | ( w1762 & ~w21307 ) ;
  assign w21309 = w21305 | w21308 ;
  assign w21310 = \pi067 ^ w21293 ;
  assign w21311 = ( ~w21304 & w21309 ) | ( ~w21304 & w21310 ) | ( w21309 & w21310 ) ;
  assign w21312 = w21310 | w21311 ;
  assign w21313 = \pi068 ^ w21286 ;
  assign w21314 = ( ~w21294 & w21312 ) | ( ~w21294 & w21313 ) | ( w21312 & w21313 ) ;
  assign w21315 = w21313 | w21314 ;
  assign w21316 = \pi069 ^ w21279 ;
  assign w21317 = ( ~w21287 & w21315 ) | ( ~w21287 & w21316 ) | ( w21315 & w21316 ) ;
  assign w21318 = w21316 | w21317 ;
  assign w21319 = \pi070 ^ w21272 ;
  assign w21320 = ( ~w21280 & w21318 ) | ( ~w21280 & w21319 ) | ( w21318 & w21319 ) ;
  assign w21321 = w21319 | w21320 ;
  assign w21322 = \pi071 ^ w21265 ;
  assign w21323 = ( ~w21273 & w21321 ) | ( ~w21273 & w21322 ) | ( w21321 & w21322 ) ;
  assign w21324 = w21322 | w21323 ;
  assign w21325 = \pi072 ^ w21258 ;
  assign w21326 = ( ~w21266 & w21324 ) | ( ~w21266 & w21325 ) | ( w21324 & w21325 ) ;
  assign w21327 = w21325 | w21326 ;
  assign w21328 = \pi073 ^ w21251 ;
  assign w21329 = ( ~w21259 & w21327 ) | ( ~w21259 & w21328 ) | ( w21327 & w21328 ) ;
  assign w21330 = w21328 | w21329 ;
  assign w21331 = \pi074 ^ w21244 ;
  assign w21332 = ( ~w21252 & w21330 ) | ( ~w21252 & w21331 ) | ( w21330 & w21331 ) ;
  assign w21333 = w21331 | w21332 ;
  assign w21334 = \pi075 ^ w21237 ;
  assign w21335 = ( ~w21245 & w21333 ) | ( ~w21245 & w21334 ) | ( w21333 & w21334 ) ;
  assign w21336 = w21334 | w21335 ;
  assign w21337 = \pi076 ^ w21230 ;
  assign w21338 = ( ~w21238 & w21336 ) | ( ~w21238 & w21337 ) | ( w21336 & w21337 ) ;
  assign w21339 = w21337 | w21338 ;
  assign w21340 = \pi077 ^ w21223 ;
  assign w21341 = ( ~w21231 & w21339 ) | ( ~w21231 & w21340 ) | ( w21339 & w21340 ) ;
  assign w21342 = w21340 | w21341 ;
  assign w21343 = \pi078 ^ w21210 ;
  assign w21344 = ( ~w21224 & w21342 ) | ( ~w21224 & w21343 ) | ( w21342 & w21343 ) ;
  assign w21345 = w21343 | w21344 ;
  assign w21346 = \pi079 ^ w21216 ;
  assign w21347 = w21217 & ~w21346 ;
  assign w21348 = ( w21345 & w21346 ) | ( w21345 & ~w21347 ) | ( w21346 & ~w21347 ) ;
  assign w21349 = ~\pi079 & w21216 ;
  assign w21350 = w21348 & ~w21349 ;
  assign w21351 = w209 | w21350 ;
  assign w21352 = w21210 & w21351 ;
  assign w21353 = ~w21224 & w21342 ;
  assign w21354 = w21343 ^ w21353 ;
  assign w21355 = ~w21351 & w21354 ;
  assign w21356 = w21352 | w21355 ;
  assign w21357 = w21216 & w21351 ;
  assign w21358 = ~w21217 & w21345 ;
  assign w21359 = w21346 ^ w21358 ;
  assign w21360 = ~w21351 & w21359 ;
  assign w21361 = w21357 | w21360 ;
  assign w21362 = ~\pi079 & w21356 ;
  assign w21363 = w21223 & w21351 ;
  assign w21364 = ~w21231 & w21339 ;
  assign w21365 = w21340 ^ w21364 ;
  assign w21366 = ~w21351 & w21365 ;
  assign w21367 = w21363 | w21366 ;
  assign w21368 = ~\pi078 & w21367 ;
  assign w21369 = w21230 & w21351 ;
  assign w21370 = ~w21238 & w21336 ;
  assign w21371 = w21337 ^ w21370 ;
  assign w21372 = ~w21351 & w21371 ;
  assign w21373 = w21369 | w21372 ;
  assign w21374 = ~\pi077 & w21373 ;
  assign w21375 = w21237 & w21351 ;
  assign w21376 = ~w21245 & w21333 ;
  assign w21377 = w21334 ^ w21376 ;
  assign w21378 = ~w21351 & w21377 ;
  assign w21379 = w21375 | w21378 ;
  assign w21380 = ~\pi076 & w21379 ;
  assign w21381 = w21244 & w21351 ;
  assign w21382 = ~w21252 & w21330 ;
  assign w21383 = w21331 ^ w21382 ;
  assign w21384 = ~w21351 & w21383 ;
  assign w21385 = w21381 | w21384 ;
  assign w21386 = ~\pi075 & w21385 ;
  assign w21387 = w21251 & w21351 ;
  assign w21388 = ~w21259 & w21327 ;
  assign w21389 = w21328 ^ w21388 ;
  assign w21390 = ~w21351 & w21389 ;
  assign w21391 = w21387 | w21390 ;
  assign w21392 = ~\pi074 & w21391 ;
  assign w21393 = w21258 & w21351 ;
  assign w21394 = ~w21266 & w21324 ;
  assign w21395 = w21325 ^ w21394 ;
  assign w21396 = ~w21351 & w21395 ;
  assign w21397 = w21393 | w21396 ;
  assign w21398 = ~\pi073 & w21397 ;
  assign w21399 = w21265 & w21351 ;
  assign w21400 = ~w21273 & w21321 ;
  assign w21401 = w21322 ^ w21400 ;
  assign w21402 = ~w21351 & w21401 ;
  assign w21403 = w21399 | w21402 ;
  assign w21404 = ~\pi072 & w21403 ;
  assign w21405 = w21272 & w21351 ;
  assign w21406 = ~w21280 & w21318 ;
  assign w21407 = w21319 ^ w21406 ;
  assign w21408 = ~w21351 & w21407 ;
  assign w21409 = w21405 | w21408 ;
  assign w21410 = ~\pi071 & w21409 ;
  assign w21411 = w21279 & w21351 ;
  assign w21412 = ~w21287 & w21315 ;
  assign w21413 = w21316 ^ w21412 ;
  assign w21414 = ~w21351 & w21413 ;
  assign w21415 = w21411 | w21414 ;
  assign w21416 = ~\pi070 & w21415 ;
  assign w21417 = w21286 & w21351 ;
  assign w21418 = ~w21294 & w21312 ;
  assign w21419 = w21313 ^ w21418 ;
  assign w21420 = ~w21351 & w21419 ;
  assign w21421 = w21417 | w21420 ;
  assign w21422 = ~\pi069 & w21421 ;
  assign w21423 = w21293 & w21351 ;
  assign w21424 = ~w21304 & w21309 ;
  assign w21425 = w21310 ^ w21424 ;
  assign w21426 = ~w21351 & w21425 ;
  assign w21427 = w21423 | w21426 ;
  assign w21428 = ~\pi068 & w21427 ;
  assign w21429 = w21303 & w21351 ;
  assign w21430 = \pi064 & ~w21204 ;
  assign w21431 = \pi049 ^ w21430 ;
  assign w21432 = ( \pi065 & w1762 ) | ( \pi065 & ~w21431 ) | ( w1762 & ~w21431 ) ;
  assign w21433 = w21305 ^ w21432 ;
  assign w21434 = ( w209 & w21350 ) | ( w209 & w21433 ) | ( w21350 & w21433 ) ;
  assign w21435 = w21433 & ~w21434 ;
  assign w21436 = w21429 | w21435 ;
  assign w21437 = ~\pi067 & w21436 ;
  assign w21438 = \pi048 ^ w21204 ;
  assign w21439 = ( \pi064 & w209 ) | ( \pi064 & w21438 ) | ( w209 & w21438 ) ;
  assign w21440 = w1769 ^ w21439 ;
  assign w21441 = ~w209 & w21440 ;
  assign w21442 = ~w21350 & w21441 ;
  assign w21443 = ( ~\pi064 & w21204 ) | ( ~\pi064 & w21351 ) | ( w21204 & w21351 ) ;
  assign w21444 = \pi049 ^ w21443 ;
  assign w21445 = w21351 & ~w21444 ;
  assign w21446 = w21442 | w21445 ;
  assign w21447 = ~\pi066 & w21446 ;
  assign w21448 = ( \pi048 & ~w1782 ) | ( \pi048 & w21350 ) | ( ~w1782 & w21350 ) ;
  assign w21449 = \pi048 & w21448 ;
  assign w21450 = w1786 & ~w21350 ;
  assign w21451 = w21449 | w21450 ;
  assign w21452 = \pi065 ^ w21451 ;
  assign w21453 = w1789 | w21452 ;
  assign w21454 = w21351 | w21442 ;
  assign w21455 = ( w21431 & w21442 ) | ( w21431 & w21454 ) | ( w21442 & w21454 ) ;
  assign w21456 = \pi066 ^ w21455 ;
  assign w21457 = ~\pi065 & w21451 ;
  assign w21458 = w21453 | w21457 ;
  assign w21459 = ( w21456 & ~w21457 ) | ( w21456 & w21458 ) | ( ~w21457 & w21458 ) ;
  assign w21460 = \pi067 ^ w21436 ;
  assign w21461 = ( ~w21447 & w21459 ) | ( ~w21447 & w21460 ) | ( w21459 & w21460 ) ;
  assign w21462 = w21460 | w21461 ;
  assign w21463 = \pi068 ^ w21427 ;
  assign w21464 = ( ~w21437 & w21462 ) | ( ~w21437 & w21463 ) | ( w21462 & w21463 ) ;
  assign w21465 = w21463 | w21464 ;
  assign w21466 = \pi069 ^ w21421 ;
  assign w21467 = ( ~w21428 & w21465 ) | ( ~w21428 & w21466 ) | ( w21465 & w21466 ) ;
  assign w21468 = w21466 | w21467 ;
  assign w21469 = \pi070 ^ w21415 ;
  assign w21470 = ( ~w21422 & w21468 ) | ( ~w21422 & w21469 ) | ( w21468 & w21469 ) ;
  assign w21471 = w21469 | w21470 ;
  assign w21472 = \pi071 ^ w21409 ;
  assign w21473 = ( ~w21416 & w21471 ) | ( ~w21416 & w21472 ) | ( w21471 & w21472 ) ;
  assign w21474 = w21472 | w21473 ;
  assign w21475 = \pi072 ^ w21403 ;
  assign w21476 = ( ~w21410 & w21474 ) | ( ~w21410 & w21475 ) | ( w21474 & w21475 ) ;
  assign w21477 = w21475 | w21476 ;
  assign w21478 = \pi073 ^ w21397 ;
  assign w21479 = ( ~w21404 & w21477 ) | ( ~w21404 & w21478 ) | ( w21477 & w21478 ) ;
  assign w21480 = w21478 | w21479 ;
  assign w21481 = \pi074 ^ w21391 ;
  assign w21482 = ( ~w21398 & w21480 ) | ( ~w21398 & w21481 ) | ( w21480 & w21481 ) ;
  assign w21483 = w21481 | w21482 ;
  assign w21484 = \pi075 ^ w21385 ;
  assign w21485 = ( ~w21392 & w21483 ) | ( ~w21392 & w21484 ) | ( w21483 & w21484 ) ;
  assign w21486 = w21484 | w21485 ;
  assign w21487 = \pi076 ^ w21379 ;
  assign w21488 = ( ~w21386 & w21486 ) | ( ~w21386 & w21487 ) | ( w21486 & w21487 ) ;
  assign w21489 = w21487 | w21488 ;
  assign w21490 = \pi077 ^ w21373 ;
  assign w21491 = ( ~w21380 & w21489 ) | ( ~w21380 & w21490 ) | ( w21489 & w21490 ) ;
  assign w21492 = w21490 | w21491 ;
  assign w21493 = \pi078 ^ w21367 ;
  assign w21494 = ( ~w21374 & w21492 ) | ( ~w21374 & w21493 ) | ( w21492 & w21493 ) ;
  assign w21495 = w21493 | w21494 ;
  assign w21496 = \pi079 ^ w21356 ;
  assign w21497 = ( ~w21368 & w21495 ) | ( ~w21368 & w21496 ) | ( w21495 & w21496 ) ;
  assign w21498 = w21496 | w21497 ;
  assign w21499 = \pi080 ^ w21361 ;
  assign w21500 = w21362 & ~w21499 ;
  assign w21501 = ( w21498 & w21499 ) | ( w21498 & ~w21500 ) | ( w21499 & ~w21500 ) ;
  assign w21502 = ~\pi080 & w21361 ;
  assign w21503 = w21501 & ~w21502 ;
  assign w21504 = w331 | w21503 ;
  assign w21505 = w21356 & w21504 ;
  assign w21506 = ~w21368 & w21495 ;
  assign w21507 = w21496 ^ w21506 ;
  assign w21508 = ~w21504 & w21507 ;
  assign w21509 = w21505 | w21508 ;
  assign w21510 = ~\pi080 & w21509 ;
  assign w21511 = w21367 & w21504 ;
  assign w21512 = ~w21374 & w21492 ;
  assign w21513 = w21493 ^ w21512 ;
  assign w21514 = ~w21504 & w21513 ;
  assign w21515 = w21511 | w21514 ;
  assign w21516 = ~\pi079 & w21515 ;
  assign w21517 = w21373 & w21504 ;
  assign w21518 = ~w21380 & w21489 ;
  assign w21519 = w21490 ^ w21518 ;
  assign w21520 = ~w21504 & w21519 ;
  assign w21521 = w21517 | w21520 ;
  assign w21522 = ~\pi078 & w21521 ;
  assign w21523 = w21379 & w21504 ;
  assign w21524 = ~w21386 & w21486 ;
  assign w21525 = w21487 ^ w21524 ;
  assign w21526 = ~w21504 & w21525 ;
  assign w21527 = w21523 | w21526 ;
  assign w21528 = ~\pi077 & w21527 ;
  assign w21529 = w21385 & w21504 ;
  assign w21530 = ~w21392 & w21483 ;
  assign w21531 = w21484 ^ w21530 ;
  assign w21532 = ~w21504 & w21531 ;
  assign w21533 = w21529 | w21532 ;
  assign w21534 = ~\pi076 & w21533 ;
  assign w21535 = w21391 & w21504 ;
  assign w21536 = ~w21398 & w21480 ;
  assign w21537 = w21481 ^ w21536 ;
  assign w21538 = ~w21504 & w21537 ;
  assign w21539 = w21535 | w21538 ;
  assign w21540 = ~\pi075 & w21539 ;
  assign w21541 = w21397 & w21504 ;
  assign w21542 = ~w21404 & w21477 ;
  assign w21543 = w21478 ^ w21542 ;
  assign w21544 = ~w21504 & w21543 ;
  assign w21545 = w21541 | w21544 ;
  assign w21546 = ~\pi074 & w21545 ;
  assign w21547 = w21403 & w21504 ;
  assign w21548 = ~w21410 & w21474 ;
  assign w21549 = w21475 ^ w21548 ;
  assign w21550 = ~w21504 & w21549 ;
  assign w21551 = w21547 | w21550 ;
  assign w21552 = ~\pi073 & w21551 ;
  assign w21553 = w21409 & w21504 ;
  assign w21554 = ~w21416 & w21471 ;
  assign w21555 = w21472 ^ w21554 ;
  assign w21556 = ~w21504 & w21555 ;
  assign w21557 = w21553 | w21556 ;
  assign w21558 = ~\pi072 & w21557 ;
  assign w21559 = w21415 & w21504 ;
  assign w21560 = ~w21422 & w21468 ;
  assign w21561 = w21469 ^ w21560 ;
  assign w21562 = ~w21504 & w21561 ;
  assign w21563 = w21559 | w21562 ;
  assign w21564 = ~\pi071 & w21563 ;
  assign w21565 = w21421 & w21504 ;
  assign w21566 = ~w21428 & w21465 ;
  assign w21567 = w21466 ^ w21566 ;
  assign w21568 = ~w21504 & w21567 ;
  assign w21569 = w21565 | w21568 ;
  assign w21570 = ~\pi070 & w21569 ;
  assign w21571 = w21427 & w21504 ;
  assign w21572 = ~w21437 & w21462 ;
  assign w21573 = w21463 ^ w21572 ;
  assign w21574 = ~w21504 & w21573 ;
  assign w21575 = w21571 | w21574 ;
  assign w21576 = ~\pi069 & w21575 ;
  assign w21577 = w21436 & w21504 ;
  assign w21578 = ~w21447 & w21459 ;
  assign w21579 = w21460 ^ w21578 ;
  assign w21580 = ~w21504 & w21579 ;
  assign w21581 = w21577 | w21580 ;
  assign w21582 = ~\pi068 & w21581 ;
  assign w21583 = w21446 & w21504 ;
  assign w21584 = ~w21451 & w21453 ;
  assign w21585 = ( \pi065 & w21453 ) | ( \pi065 & w21584 ) | ( w21453 & w21584 ) ;
  assign w21586 = w21456 ^ w21585 ;
  assign w21587 = ~w21504 & w21586 ;
  assign w21588 = w21583 | w21587 ;
  assign w21589 = ~\pi067 & w21588 ;
  assign w21590 = w21451 & w21504 ;
  assign w21591 = ( ~w331 & w21449 ) | ( ~w331 & w21450 ) | ( w21449 & w21450 ) ;
  assign w21592 = \pi065 ^ w21591 ;
  assign w21593 = ( ~w331 & w1789 ) | ( ~w331 & w21592 ) | ( w1789 & w21592 ) ;
  assign w21594 = ( w1789 & w21503 ) | ( w1789 & w21592 ) | ( w21503 & w21592 ) ;
  assign w21595 = w21593 & ~w21594 ;
  assign w21596 = w21590 | w21595 ;
  assign w21597 = ~\pi066 & w21596 ;
  assign w21598 = ( \pi047 & ~w1942 ) | ( \pi047 & w21503 ) | ( ~w1942 & w21503 ) ;
  assign w21599 = \pi047 & w21598 ;
  assign w21600 = ( w443 & ~w452 ) | ( w443 & w21503 ) | ( ~w452 & w21503 ) ;
  assign w21601 = w1946 & ~w21600 ;
  assign w21602 = w21599 | w21601 ;
  assign w21603 = ( ~w1950 & w21599 ) | ( ~w1950 & w21601 ) | ( w21599 & w21601 ) ;
  assign w21604 = \pi065 ^ w21603 ;
  assign w21605 = w1950 | w21604 ;
  assign w21606 = ~\pi065 & w21602 ;
  assign w21607 = \pi066 ^ w21596 ;
  assign w21608 = ( w21605 & ~w21606 ) | ( w21605 & w21607 ) | ( ~w21606 & w21607 ) ;
  assign w21609 = w21607 | w21608 ;
  assign w21610 = \pi067 ^ w21588 ;
  assign w21611 = ( ~w21597 & w21609 ) | ( ~w21597 & w21610 ) | ( w21609 & w21610 ) ;
  assign w21612 = w21610 | w21611 ;
  assign w21613 = \pi068 ^ w21581 ;
  assign w21614 = ( ~w21589 & w21612 ) | ( ~w21589 & w21613 ) | ( w21612 & w21613 ) ;
  assign w21615 = w21613 | w21614 ;
  assign w21616 = \pi069 ^ w21575 ;
  assign w21617 = ( ~w21582 & w21615 ) | ( ~w21582 & w21616 ) | ( w21615 & w21616 ) ;
  assign w21618 = w21616 | w21617 ;
  assign w21619 = \pi070 ^ w21569 ;
  assign w21620 = ( ~w21576 & w21618 ) | ( ~w21576 & w21619 ) | ( w21618 & w21619 ) ;
  assign w21621 = w21619 | w21620 ;
  assign w21622 = \pi071 ^ w21563 ;
  assign w21623 = ( ~w21570 & w21621 ) | ( ~w21570 & w21622 ) | ( w21621 & w21622 ) ;
  assign w21624 = w21622 | w21623 ;
  assign w21625 = \pi072 ^ w21557 ;
  assign w21626 = ( ~w21564 & w21624 ) | ( ~w21564 & w21625 ) | ( w21624 & w21625 ) ;
  assign w21627 = w21625 | w21626 ;
  assign w21628 = \pi073 ^ w21551 ;
  assign w21629 = ( ~w21558 & w21627 ) | ( ~w21558 & w21628 ) | ( w21627 & w21628 ) ;
  assign w21630 = w21628 | w21629 ;
  assign w21631 = \pi074 ^ w21545 ;
  assign w21632 = ( ~w21552 & w21630 ) | ( ~w21552 & w21631 ) | ( w21630 & w21631 ) ;
  assign w21633 = w21631 | w21632 ;
  assign w21634 = \pi075 ^ w21539 ;
  assign w21635 = ( ~w21546 & w21633 ) | ( ~w21546 & w21634 ) | ( w21633 & w21634 ) ;
  assign w21636 = w21634 | w21635 ;
  assign w21637 = \pi076 ^ w21533 ;
  assign w21638 = ( ~w21540 & w21636 ) | ( ~w21540 & w21637 ) | ( w21636 & w21637 ) ;
  assign w21639 = w21637 | w21638 ;
  assign w21640 = \pi077 ^ w21527 ;
  assign w21641 = ( ~w21534 & w21639 ) | ( ~w21534 & w21640 ) | ( w21639 & w21640 ) ;
  assign w21642 = w21640 | w21641 ;
  assign w21643 = \pi078 ^ w21521 ;
  assign w21644 = ( ~w21528 & w21642 ) | ( ~w21528 & w21643 ) | ( w21642 & w21643 ) ;
  assign w21645 = w21643 | w21644 ;
  assign w21646 = \pi079 ^ w21515 ;
  assign w21647 = ( ~w21522 & w21645 ) | ( ~w21522 & w21646 ) | ( w21645 & w21646 ) ;
  assign w21648 = w21646 | w21647 ;
  assign w21649 = \pi080 ^ w21509 ;
  assign w21650 = ( ~w21516 & w21648 ) | ( ~w21516 & w21649 ) | ( w21648 & w21649 ) ;
  assign w21651 = w21649 | w21650 ;
  assign w21652 = w21361 & w21504 ;
  assign w21653 = ~w21362 & w21498 ;
  assign w21654 = w21499 ^ w21653 ;
  assign w21655 = ~w21504 & w21654 ;
  assign w21656 = w21652 | w21655 ;
  assign w21657 = ~\pi081 & w21656 ;
  assign w21658 = ( \pi081 & ~w21652 ) | ( \pi081 & w21655 ) | ( ~w21652 & w21655 ) ;
  assign w21659 = ~w21655 & w21658 ;
  assign w21660 = w21657 | w21659 ;
  assign w21661 = ( ~w21510 & w21651 ) | ( ~w21510 & w21660 ) | ( w21651 & w21660 ) ;
  assign w21662 = ( w2011 & ~w21660 ) | ( w2011 & w21661 ) | ( ~w21660 & w21661 ) ;
  assign w21663 = w21660 | w21662 ;
  assign w21664 = ~w331 & w21656 ;
  assign w21665 = w21663 & ~w21664 ;
  assign w21666 = ~w21516 & w21648 ;
  assign w21667 = w21649 ^ w21666 ;
  assign w21668 = ~w21665 & w21667 ;
  assign w21669 = ( w21509 & w21663 ) | ( w21509 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21670 = ~w21664 & w21669 ;
  assign w21671 = w21668 | w21670 ;
  assign w21672 = ( ~w21510 & w21651 ) | ( ~w21510 & w21665 ) | ( w21651 & w21665 ) ;
  assign w21673 = w21660 ^ w21672 ;
  assign w21674 = ~w21665 & w21673 ;
  assign w21675 = ( w331 & ~w21656 ) | ( w331 & w21663 ) | ( ~w21656 & w21663 ) ;
  assign w21676 = w21656 & w21675 ;
  assign w21677 = w21674 | w21676 ;
  assign w21678 = ~\pi081 & w21671 ;
  assign w21679 = ~w21522 & w21645 ;
  assign w21680 = w21646 ^ w21679 ;
  assign w21681 = ~w21665 & w21680 ;
  assign w21682 = ( w21515 & w21663 ) | ( w21515 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21683 = ~w21664 & w21682 ;
  assign w21684 = w21681 | w21683 ;
  assign w21685 = ~\pi080 & w21684 ;
  assign w21686 = ~w21528 & w21642 ;
  assign w21687 = w21643 ^ w21686 ;
  assign w21688 = ~w21665 & w21687 ;
  assign w21689 = ( w21521 & w21663 ) | ( w21521 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21690 = ~w21664 & w21689 ;
  assign w21691 = w21688 | w21690 ;
  assign w21692 = ~\pi079 & w21691 ;
  assign w21693 = ~w21534 & w21639 ;
  assign w21694 = w21640 ^ w21693 ;
  assign w21695 = ~w21665 & w21694 ;
  assign w21696 = ( w21527 & w21663 ) | ( w21527 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21697 = ~w21664 & w21696 ;
  assign w21698 = w21695 | w21697 ;
  assign w21699 = ~\pi078 & w21698 ;
  assign w21700 = ~w21540 & w21636 ;
  assign w21701 = w21637 ^ w21700 ;
  assign w21702 = ~w21665 & w21701 ;
  assign w21703 = ( w21533 & w21663 ) | ( w21533 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21704 = ~w21664 & w21703 ;
  assign w21705 = w21702 | w21704 ;
  assign w21706 = ~\pi077 & w21705 ;
  assign w21707 = ~w21546 & w21633 ;
  assign w21708 = w21634 ^ w21707 ;
  assign w21709 = ~w21665 & w21708 ;
  assign w21710 = ( w21539 & w21663 ) | ( w21539 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21711 = ~w21664 & w21710 ;
  assign w21712 = w21709 | w21711 ;
  assign w21713 = ~\pi076 & w21712 ;
  assign w21714 = ~w21552 & w21630 ;
  assign w21715 = w21631 ^ w21714 ;
  assign w21716 = ~w21665 & w21715 ;
  assign w21717 = ( w21545 & w21663 ) | ( w21545 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21718 = ~w21664 & w21717 ;
  assign w21719 = w21716 | w21718 ;
  assign w21720 = ~\pi075 & w21719 ;
  assign w21721 = ~w21558 & w21627 ;
  assign w21722 = w21628 ^ w21721 ;
  assign w21723 = ~w21665 & w21722 ;
  assign w21724 = ( w21551 & w21663 ) | ( w21551 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21725 = ~w21664 & w21724 ;
  assign w21726 = w21723 | w21725 ;
  assign w21727 = ~\pi074 & w21726 ;
  assign w21728 = ~w21564 & w21624 ;
  assign w21729 = w21625 ^ w21728 ;
  assign w21730 = ~w21665 & w21729 ;
  assign w21731 = ( w21557 & w21663 ) | ( w21557 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21732 = ~w21664 & w21731 ;
  assign w21733 = w21730 | w21732 ;
  assign w21734 = ~\pi073 & w21733 ;
  assign w21735 = ~w21570 & w21621 ;
  assign w21736 = w21622 ^ w21735 ;
  assign w21737 = ~w21665 & w21736 ;
  assign w21738 = ( w21563 & w21663 ) | ( w21563 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21739 = ~w21664 & w21738 ;
  assign w21740 = w21737 | w21739 ;
  assign w21741 = ~\pi072 & w21740 ;
  assign w21742 = ~w21576 & w21618 ;
  assign w21743 = w21619 ^ w21742 ;
  assign w21744 = ~w21665 & w21743 ;
  assign w21745 = ( w21569 & w21663 ) | ( w21569 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21746 = ~w21664 & w21745 ;
  assign w21747 = w21744 | w21746 ;
  assign w21748 = ~\pi071 & w21747 ;
  assign w21749 = ~w21582 & w21615 ;
  assign w21750 = w21616 ^ w21749 ;
  assign w21751 = ~w21665 & w21750 ;
  assign w21752 = ( w21575 & w21663 ) | ( w21575 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21753 = ~w21664 & w21752 ;
  assign w21754 = w21751 | w21753 ;
  assign w21755 = ~\pi070 & w21754 ;
  assign w21756 = ~w21589 & w21612 ;
  assign w21757 = w21613 ^ w21756 ;
  assign w21758 = ~w21665 & w21757 ;
  assign w21759 = ( w21581 & w21663 ) | ( w21581 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21760 = ~w21664 & w21759 ;
  assign w21761 = w21758 | w21760 ;
  assign w21762 = ~\pi069 & w21761 ;
  assign w21763 = ~w21597 & w21609 ;
  assign w21764 = w21610 ^ w21763 ;
  assign w21765 = ~w21665 & w21764 ;
  assign w21766 = ( w21588 & w21663 ) | ( w21588 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21767 = ~w21664 & w21766 ;
  assign w21768 = w21765 | w21767 ;
  assign w21769 = ~\pi068 & w21768 ;
  assign w21770 = w21605 & ~w21606 ;
  assign w21771 = w21607 ^ w21770 ;
  assign w21772 = ~w21665 & w21771 ;
  assign w21773 = ( w21596 & w21663 ) | ( w21596 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21774 = ~w21664 & w21773 ;
  assign w21775 = w21772 | w21774 ;
  assign w21776 = ~\pi067 & w21775 ;
  assign w21777 = ( w21599 & w21601 ) | ( w21599 & ~w21665 ) | ( w21601 & ~w21665 ) ;
  assign w21778 = ( ~\pi046 & \pi064 ) | ( ~\pi046 & w21665 ) | ( \pi064 & w21665 ) ;
  assign w21779 = w21777 ^ w21778 ;
  assign w21780 = \pi065 ^ w21779 ;
  assign w21781 = ~w21665 & w21780 ;
  assign w21782 = ( w21602 & w21663 ) | ( w21602 & w21664 ) | ( w21663 & w21664 ) ;
  assign w21783 = ~w21664 & w21782 ;
  assign w21784 = w21781 | w21783 ;
  assign w21785 = ~\pi066 & w21784 ;
  assign w21786 = \pi066 ^ w21784 ;
  assign w21787 = ( \pi064 & ~w21665 ) | ( \pi064 & w21786 ) | ( ~w21665 & w21786 ) ;
  assign w21788 = \pi046 ^ w21787 ;
  assign w21789 = ( \pi065 & w2295 ) | ( \pi065 & ~w21788 ) | ( w2295 & ~w21788 ) ;
  assign w21790 = w21786 | w21789 ;
  assign w21791 = \pi067 ^ w21775 ;
  assign w21792 = ( ~w21785 & w21790 ) | ( ~w21785 & w21791 ) | ( w21790 & w21791 ) ;
  assign w21793 = w21791 | w21792 ;
  assign w21794 = \pi068 ^ w21768 ;
  assign w21795 = ( ~w21776 & w21793 ) | ( ~w21776 & w21794 ) | ( w21793 & w21794 ) ;
  assign w21796 = w21794 | w21795 ;
  assign w21797 = \pi069 ^ w21761 ;
  assign w21798 = ( ~w21769 & w21796 ) | ( ~w21769 & w21797 ) | ( w21796 & w21797 ) ;
  assign w21799 = w21797 | w21798 ;
  assign w21800 = \pi070 ^ w21754 ;
  assign w21801 = ( ~w21762 & w21799 ) | ( ~w21762 & w21800 ) | ( w21799 & w21800 ) ;
  assign w21802 = w21800 | w21801 ;
  assign w21803 = \pi071 ^ w21747 ;
  assign w21804 = ( ~w21755 & w21802 ) | ( ~w21755 & w21803 ) | ( w21802 & w21803 ) ;
  assign w21805 = w21803 | w21804 ;
  assign w21806 = \pi072 ^ w21740 ;
  assign w21807 = ( ~w21748 & w21805 ) | ( ~w21748 & w21806 ) | ( w21805 & w21806 ) ;
  assign w21808 = w21806 | w21807 ;
  assign w21809 = \pi073 ^ w21733 ;
  assign w21810 = ( ~w21741 & w21808 ) | ( ~w21741 & w21809 ) | ( w21808 & w21809 ) ;
  assign w21811 = w21809 | w21810 ;
  assign w21812 = \pi074 ^ w21726 ;
  assign w21813 = ( ~w21734 & w21811 ) | ( ~w21734 & w21812 ) | ( w21811 & w21812 ) ;
  assign w21814 = w21812 | w21813 ;
  assign w21815 = \pi075 ^ w21719 ;
  assign w21816 = ( ~w21727 & w21814 ) | ( ~w21727 & w21815 ) | ( w21814 & w21815 ) ;
  assign w21817 = w21815 | w21816 ;
  assign w21818 = \pi076 ^ w21712 ;
  assign w21819 = ( ~w21720 & w21817 ) | ( ~w21720 & w21818 ) | ( w21817 & w21818 ) ;
  assign w21820 = w21818 | w21819 ;
  assign w21821 = \pi077 ^ w21705 ;
  assign w21822 = ( ~w21713 & w21820 ) | ( ~w21713 & w21821 ) | ( w21820 & w21821 ) ;
  assign w21823 = w21821 | w21822 ;
  assign w21824 = \pi078 ^ w21698 ;
  assign w21825 = ( ~w21706 & w21823 ) | ( ~w21706 & w21824 ) | ( w21823 & w21824 ) ;
  assign w21826 = w21824 | w21825 ;
  assign w21827 = \pi079 ^ w21691 ;
  assign w21828 = ( ~w21699 & w21826 ) | ( ~w21699 & w21827 ) | ( w21826 & w21827 ) ;
  assign w21829 = w21827 | w21828 ;
  assign w21830 = \pi080 ^ w21684 ;
  assign w21831 = ( ~w21692 & w21829 ) | ( ~w21692 & w21830 ) | ( w21829 & w21830 ) ;
  assign w21832 = w21830 | w21831 ;
  assign w21833 = \pi081 ^ w21671 ;
  assign w21834 = ( ~w21685 & w21832 ) | ( ~w21685 & w21833 ) | ( w21832 & w21833 ) ;
  assign w21835 = w21833 | w21834 ;
  assign w21836 = \pi082 ^ w21677 ;
  assign w21837 = w21678 & ~w21836 ;
  assign w21838 = ( w21835 & w21836 ) | ( w21835 & ~w21837 ) | ( w21836 & ~w21837 ) ;
  assign w21839 = ~\pi082 & w21677 ;
  assign w21840 = w21838 & ~w21839 ;
  assign w21841 = w2197 | w21840 ;
  assign w21842 = w21671 & w21841 ;
  assign w21843 = ~w21685 & w21832 ;
  assign w21844 = w21833 ^ w21843 ;
  assign w21845 = ~w21841 & w21844 ;
  assign w21846 = w21842 | w21845 ;
  assign w21847 = w21677 & w21841 ;
  assign w21848 = ~w21678 & w21835 ;
  assign w21849 = w21836 ^ w21848 ;
  assign w21850 = ~w21841 & w21849 ;
  assign w21851 = w21847 | w21850 ;
  assign w21852 = ~\pi082 & w21846 ;
  assign w21853 = w21684 & w21841 ;
  assign w21854 = ~w21692 & w21829 ;
  assign w21855 = w21830 ^ w21854 ;
  assign w21856 = ~w21841 & w21855 ;
  assign w21857 = w21853 | w21856 ;
  assign w21858 = ~\pi081 & w21857 ;
  assign w21859 = w21691 & w21841 ;
  assign w21860 = ~w21699 & w21826 ;
  assign w21861 = w21827 ^ w21860 ;
  assign w21862 = ~w21841 & w21861 ;
  assign w21863 = w21859 | w21862 ;
  assign w21864 = ~\pi080 & w21863 ;
  assign w21865 = w21698 & w21841 ;
  assign w21866 = ~w21706 & w21823 ;
  assign w21867 = w21824 ^ w21866 ;
  assign w21868 = ~w21841 & w21867 ;
  assign w21869 = w21865 | w21868 ;
  assign w21870 = ~\pi079 & w21869 ;
  assign w21871 = w21705 & w21841 ;
  assign w21872 = ~w21713 & w21820 ;
  assign w21873 = w21821 ^ w21872 ;
  assign w21874 = ~w21841 & w21873 ;
  assign w21875 = w21871 | w21874 ;
  assign w21876 = ~\pi078 & w21875 ;
  assign w21877 = w21712 & w21841 ;
  assign w21878 = ~w21720 & w21817 ;
  assign w21879 = w21818 ^ w21878 ;
  assign w21880 = ~w21841 & w21879 ;
  assign w21881 = w21877 | w21880 ;
  assign w21882 = ~\pi077 & w21881 ;
  assign w21883 = w21719 & w21841 ;
  assign w21884 = ~w21727 & w21814 ;
  assign w21885 = w21815 ^ w21884 ;
  assign w21886 = ~w21841 & w21885 ;
  assign w21887 = w21883 | w21886 ;
  assign w21888 = ~\pi076 & w21887 ;
  assign w21889 = w21726 & w21841 ;
  assign w21890 = ~w21734 & w21811 ;
  assign w21891 = w21812 ^ w21890 ;
  assign w21892 = ~w21841 & w21891 ;
  assign w21893 = w21889 | w21892 ;
  assign w21894 = ~\pi075 & w21893 ;
  assign w21895 = w21733 & w21841 ;
  assign w21896 = ~w21741 & w21808 ;
  assign w21897 = w21809 ^ w21896 ;
  assign w21898 = ~w21841 & w21897 ;
  assign w21899 = w21895 | w21898 ;
  assign w21900 = ~\pi074 & w21899 ;
  assign w21901 = w21740 & w21841 ;
  assign w21902 = ~w21748 & w21805 ;
  assign w21903 = w21806 ^ w21902 ;
  assign w21904 = ~w21841 & w21903 ;
  assign w21905 = w21901 | w21904 ;
  assign w21906 = ~\pi073 & w21905 ;
  assign w21907 = w21747 & w21841 ;
  assign w21908 = ~w21755 & w21802 ;
  assign w21909 = w21803 ^ w21908 ;
  assign w21910 = ~w21841 & w21909 ;
  assign w21911 = w21907 | w21910 ;
  assign w21912 = ~\pi072 & w21911 ;
  assign w21913 = w21754 & w21841 ;
  assign w21914 = ~w21762 & w21799 ;
  assign w21915 = w21800 ^ w21914 ;
  assign w21916 = ~w21841 & w21915 ;
  assign w21917 = w21913 | w21916 ;
  assign w21918 = ~\pi071 & w21917 ;
  assign w21919 = w21761 & w21841 ;
  assign w21920 = ~w21769 & w21796 ;
  assign w21921 = w21797 ^ w21920 ;
  assign w21922 = ~w21841 & w21921 ;
  assign w21923 = w21919 | w21922 ;
  assign w21924 = ~\pi070 & w21923 ;
  assign w21925 = w21768 & w21841 ;
  assign w21926 = ~w21776 & w21793 ;
  assign w21927 = w21794 ^ w21926 ;
  assign w21928 = ~w21841 & w21927 ;
  assign w21929 = w21925 | w21928 ;
  assign w21930 = ~\pi069 & w21929 ;
  assign w21931 = w21775 & w21841 ;
  assign w21932 = ~w21785 & w21790 ;
  assign w21933 = w21791 ^ w21932 ;
  assign w21934 = ~w21841 & w21933 ;
  assign w21935 = w21931 | w21934 ;
  assign w21936 = ~\pi068 & w21935 ;
  assign w21937 = w21784 & w21841 ;
  assign w21938 = \pi064 & ~w21665 ;
  assign w21939 = \pi046 ^ w21938 ;
  assign w21940 = ( \pi065 & w2295 ) | ( \pi065 & ~w21939 ) | ( w2295 & ~w21939 ) ;
  assign w21941 = w21786 ^ w21940 ;
  assign w21942 = ( w2197 & w21840 ) | ( w2197 & w21941 ) | ( w21840 & w21941 ) ;
  assign w21943 = w21941 & ~w21942 ;
  assign w21944 = w21937 | w21943 ;
  assign w21945 = ~\pi067 & w21944 ;
  assign w21946 = \pi045 ^ w21665 ;
  assign w21947 = ( \pi064 & w2197 ) | ( \pi064 & w21946 ) | ( w2197 & w21946 ) ;
  assign w21948 = w2302 ^ w21947 ;
  assign w21949 = ~w2197 & w21948 ;
  assign w21950 = ~w21840 & w21949 ;
  assign w21951 = ( ~\pi064 & w21665 ) | ( ~\pi064 & w21841 ) | ( w21665 & w21841 ) ;
  assign w21952 = \pi046 ^ w21951 ;
  assign w21953 = w21841 & ~w21952 ;
  assign w21954 = w21950 | w21953 ;
  assign w21955 = ~\pi066 & w21954 ;
  assign w21956 = ( \pi045 & ~w2316 ) | ( \pi045 & w21840 ) | ( ~w2316 & w21840 ) ;
  assign w21957 = \pi045 & w21956 ;
  assign w21958 = w2325 & ~w21840 ;
  assign w21959 = w21957 | w21958 ;
  assign w21960 = \pi065 ^ w21959 ;
  assign w21961 = w2328 | w21960 ;
  assign w21962 = ~\pi065 & w21959 ;
  assign w21963 = w21841 | w21950 ;
  assign w21964 = ( w21939 & w21950 ) | ( w21939 & w21963 ) | ( w21950 & w21963 ) ;
  assign w21965 = \pi066 ^ w21964 ;
  assign w21966 = ( w21961 & ~w21962 ) | ( w21961 & w21965 ) | ( ~w21962 & w21965 ) ;
  assign w21967 = w21965 | w21966 ;
  assign w21968 = \pi067 ^ w21944 ;
  assign w21969 = ( ~w21955 & w21967 ) | ( ~w21955 & w21968 ) | ( w21967 & w21968 ) ;
  assign w21970 = w21968 | w21969 ;
  assign w21971 = \pi068 ^ w21935 ;
  assign w21972 = ( ~w21945 & w21970 ) | ( ~w21945 & w21971 ) | ( w21970 & w21971 ) ;
  assign w21973 = w21971 | w21972 ;
  assign w21974 = \pi069 ^ w21929 ;
  assign w21975 = ( ~w21936 & w21973 ) | ( ~w21936 & w21974 ) | ( w21973 & w21974 ) ;
  assign w21976 = w21974 | w21975 ;
  assign w21977 = \pi070 ^ w21923 ;
  assign w21978 = ( ~w21930 & w21976 ) | ( ~w21930 & w21977 ) | ( w21976 & w21977 ) ;
  assign w21979 = w21977 | w21978 ;
  assign w21980 = \pi071 ^ w21917 ;
  assign w21981 = ( ~w21924 & w21979 ) | ( ~w21924 & w21980 ) | ( w21979 & w21980 ) ;
  assign w21982 = w21980 | w21981 ;
  assign w21983 = \pi072 ^ w21911 ;
  assign w21984 = ( ~w21918 & w21982 ) | ( ~w21918 & w21983 ) | ( w21982 & w21983 ) ;
  assign w21985 = w21983 | w21984 ;
  assign w21986 = \pi073 ^ w21905 ;
  assign w21987 = ( ~w21912 & w21985 ) | ( ~w21912 & w21986 ) | ( w21985 & w21986 ) ;
  assign w21988 = w21986 | w21987 ;
  assign w21989 = \pi074 ^ w21899 ;
  assign w21990 = ( ~w21906 & w21988 ) | ( ~w21906 & w21989 ) | ( w21988 & w21989 ) ;
  assign w21991 = w21989 | w21990 ;
  assign w21992 = \pi075 ^ w21893 ;
  assign w21993 = ( ~w21900 & w21991 ) | ( ~w21900 & w21992 ) | ( w21991 & w21992 ) ;
  assign w21994 = w21992 | w21993 ;
  assign w21995 = \pi076 ^ w21887 ;
  assign w21996 = ( ~w21894 & w21994 ) | ( ~w21894 & w21995 ) | ( w21994 & w21995 ) ;
  assign w21997 = w21995 | w21996 ;
  assign w21998 = \pi077 ^ w21881 ;
  assign w21999 = ( ~w21888 & w21997 ) | ( ~w21888 & w21998 ) | ( w21997 & w21998 ) ;
  assign w22000 = w21998 | w21999 ;
  assign w22001 = \pi078 ^ w21875 ;
  assign w22002 = ( ~w21882 & w22000 ) | ( ~w21882 & w22001 ) | ( w22000 & w22001 ) ;
  assign w22003 = w22001 | w22002 ;
  assign w22004 = \pi079 ^ w21869 ;
  assign w22005 = ( ~w21876 & w22003 ) | ( ~w21876 & w22004 ) | ( w22003 & w22004 ) ;
  assign w22006 = w22004 | w22005 ;
  assign w22007 = \pi080 ^ w21863 ;
  assign w22008 = ( ~w21870 & w22006 ) | ( ~w21870 & w22007 ) | ( w22006 & w22007 ) ;
  assign w22009 = w22007 | w22008 ;
  assign w22010 = \pi081 ^ w21857 ;
  assign w22011 = ( ~w21864 & w22009 ) | ( ~w21864 & w22010 ) | ( w22009 & w22010 ) ;
  assign w22012 = w22010 | w22011 ;
  assign w22013 = \pi082 ^ w21846 ;
  assign w22014 = ( ~w21858 & w22012 ) | ( ~w21858 & w22013 ) | ( w22012 & w22013 ) ;
  assign w22015 = w22013 | w22014 ;
  assign w22016 = \pi083 ^ w21851 ;
  assign w22017 = w21852 & ~w22016 ;
  assign w22018 = ( w22015 & w22016 ) | ( w22015 & ~w22017 ) | ( w22016 & ~w22017 ) ;
  assign w22019 = ~\pi083 & w21851 ;
  assign w22020 = w22018 & ~w22019 ;
  assign w22021 = w187 | w22020 ;
  assign w22022 = w21846 & w22021 ;
  assign w22023 = ~w21858 & w22012 ;
  assign w22024 = w22013 ^ w22023 ;
  assign w22025 = ~w22021 & w22024 ;
  assign w22026 = w22022 | w22025 ;
  assign w22027 = ~\pi083 & w22026 ;
  assign w22028 = w21857 & w22021 ;
  assign w22029 = ~w21864 & w22009 ;
  assign w22030 = w22010 ^ w22029 ;
  assign w22031 = ~w22021 & w22030 ;
  assign w22032 = w22028 | w22031 ;
  assign w22033 = ~\pi082 & w22032 ;
  assign w22034 = w21863 & w22021 ;
  assign w22035 = ~w21870 & w22006 ;
  assign w22036 = w22007 ^ w22035 ;
  assign w22037 = ~w22021 & w22036 ;
  assign w22038 = w22034 | w22037 ;
  assign w22039 = ~\pi081 & w22038 ;
  assign w22040 = w21869 & w22021 ;
  assign w22041 = ~w21876 & w22003 ;
  assign w22042 = w22004 ^ w22041 ;
  assign w22043 = ~w22021 & w22042 ;
  assign w22044 = w22040 | w22043 ;
  assign w22045 = ~\pi080 & w22044 ;
  assign w22046 = w21875 & w22021 ;
  assign w22047 = ~w21882 & w22000 ;
  assign w22048 = w22001 ^ w22047 ;
  assign w22049 = ~w22021 & w22048 ;
  assign w22050 = w22046 | w22049 ;
  assign w22051 = ~\pi079 & w22050 ;
  assign w22052 = w21881 & w22021 ;
  assign w22053 = ~w21888 & w21997 ;
  assign w22054 = w21998 ^ w22053 ;
  assign w22055 = ~w22021 & w22054 ;
  assign w22056 = w22052 | w22055 ;
  assign w22057 = ~\pi078 & w22056 ;
  assign w22058 = w21887 & w22021 ;
  assign w22059 = ~w21894 & w21994 ;
  assign w22060 = w21995 ^ w22059 ;
  assign w22061 = ~w22021 & w22060 ;
  assign w22062 = w22058 | w22061 ;
  assign w22063 = ~\pi077 & w22062 ;
  assign w22064 = w21893 & w22021 ;
  assign w22065 = ~w21900 & w21991 ;
  assign w22066 = w21992 ^ w22065 ;
  assign w22067 = ~w22021 & w22066 ;
  assign w22068 = w22064 | w22067 ;
  assign w22069 = ~\pi076 & w22068 ;
  assign w22070 = w21899 & w22021 ;
  assign w22071 = ~w21906 & w21988 ;
  assign w22072 = w21989 ^ w22071 ;
  assign w22073 = ~w22021 & w22072 ;
  assign w22074 = w22070 | w22073 ;
  assign w22075 = ~\pi075 & w22074 ;
  assign w22076 = w21905 & w22021 ;
  assign w22077 = ~w21912 & w21985 ;
  assign w22078 = w21986 ^ w22077 ;
  assign w22079 = ~w22021 & w22078 ;
  assign w22080 = w22076 | w22079 ;
  assign w22081 = ~\pi074 & w22080 ;
  assign w22082 = w21911 & w22021 ;
  assign w22083 = ~w21918 & w21982 ;
  assign w22084 = w21983 ^ w22083 ;
  assign w22085 = ~w22021 & w22084 ;
  assign w22086 = w22082 | w22085 ;
  assign w22087 = ~\pi073 & w22086 ;
  assign w22088 = w21917 & w22021 ;
  assign w22089 = ~w21924 & w21979 ;
  assign w22090 = w21980 ^ w22089 ;
  assign w22091 = ~w22021 & w22090 ;
  assign w22092 = w22088 | w22091 ;
  assign w22093 = ~\pi072 & w22092 ;
  assign w22094 = w21923 & w22021 ;
  assign w22095 = ~w21930 & w21976 ;
  assign w22096 = w21977 ^ w22095 ;
  assign w22097 = ~w22021 & w22096 ;
  assign w22098 = w22094 | w22097 ;
  assign w22099 = ~\pi071 & w22098 ;
  assign w22100 = w21929 & w22021 ;
  assign w22101 = ~w21936 & w21973 ;
  assign w22102 = w21974 ^ w22101 ;
  assign w22103 = ~w22021 & w22102 ;
  assign w22104 = w22100 | w22103 ;
  assign w22105 = ~\pi070 & w22104 ;
  assign w22106 = w21935 & w22021 ;
  assign w22107 = ~w21945 & w21970 ;
  assign w22108 = w21971 ^ w22107 ;
  assign w22109 = ~w22021 & w22108 ;
  assign w22110 = w22106 | w22109 ;
  assign w22111 = ~\pi069 & w22110 ;
  assign w22112 = w21944 & w22021 ;
  assign w22113 = ~w21955 & w21967 ;
  assign w22114 = w21968 ^ w22113 ;
  assign w22115 = ~w22021 & w22114 ;
  assign w22116 = w22112 | w22115 ;
  assign w22117 = ~\pi068 & w22116 ;
  assign w22118 = w21954 & w22021 ;
  assign w22119 = w21961 & ~w21962 ;
  assign w22120 = w21965 ^ w22119 ;
  assign w22121 = ~w22021 & w22120 ;
  assign w22122 = w22118 | w22121 ;
  assign w22123 = ~\pi067 & w22122 ;
  assign w22124 = w21959 & w22021 ;
  assign w22125 = ( ~w187 & w21957 ) | ( ~w187 & w21958 ) | ( w21957 & w21958 ) ;
  assign w22126 = \pi065 ^ w22125 ;
  assign w22127 = ( ~w187 & w2328 ) | ( ~w187 & w22126 ) | ( w2328 & w22126 ) ;
  assign w22128 = ( w2328 & w22020 ) | ( w2328 & w22126 ) | ( w22020 & w22126 ) ;
  assign w22129 = w22127 & ~w22128 ;
  assign w22130 = w22124 | w22129 ;
  assign w22131 = ~\pi066 & w22130 ;
  assign w22132 = ( \pi044 & ~w2504 ) | ( \pi044 & w22020 ) | ( ~w2504 & w22020 ) ;
  assign w22133 = \pi044 & w22132 ;
  assign w22134 = w2508 | w22020 ;
  assign w22135 = ( ~w22020 & w22133 ) | ( ~w22020 & w22134 ) | ( w22133 & w22134 ) ;
  assign w22136 = w2504 & ~w22134 ;
  assign w22137 = \pi044 & ~w22136 ;
  assign w22138 = ( ~w22020 & w22134 ) | ( ~w22020 & w22137 ) | ( w22134 & w22137 ) ;
  assign w22139 = \pi065 ^ w22138 ;
  assign w22140 = w2513 | w22139 ;
  assign w22141 = ~\pi065 & w22135 ;
  assign w22142 = \pi066 ^ w22130 ;
  assign w22143 = ( w22140 & ~w22141 ) | ( w22140 & w22142 ) | ( ~w22141 & w22142 ) ;
  assign w22144 = w22142 | w22143 ;
  assign w22145 = \pi067 ^ w22122 ;
  assign w22146 = ( ~w22131 & w22144 ) | ( ~w22131 & w22145 ) | ( w22144 & w22145 ) ;
  assign w22147 = w22145 | w22146 ;
  assign w22148 = \pi068 ^ w22116 ;
  assign w22149 = ( ~w22123 & w22147 ) | ( ~w22123 & w22148 ) | ( w22147 & w22148 ) ;
  assign w22150 = w22148 | w22149 ;
  assign w22151 = \pi069 ^ w22110 ;
  assign w22152 = ( ~w22117 & w22150 ) | ( ~w22117 & w22151 ) | ( w22150 & w22151 ) ;
  assign w22153 = w22151 | w22152 ;
  assign w22154 = \pi070 ^ w22104 ;
  assign w22155 = ( ~w22111 & w22153 ) | ( ~w22111 & w22154 ) | ( w22153 & w22154 ) ;
  assign w22156 = w22154 | w22155 ;
  assign w22157 = \pi071 ^ w22098 ;
  assign w22158 = ( ~w22105 & w22156 ) | ( ~w22105 & w22157 ) | ( w22156 & w22157 ) ;
  assign w22159 = w22157 | w22158 ;
  assign w22160 = \pi072 ^ w22092 ;
  assign w22161 = ( ~w22099 & w22159 ) | ( ~w22099 & w22160 ) | ( w22159 & w22160 ) ;
  assign w22162 = w22160 | w22161 ;
  assign w22163 = \pi073 ^ w22086 ;
  assign w22164 = ( ~w22093 & w22162 ) | ( ~w22093 & w22163 ) | ( w22162 & w22163 ) ;
  assign w22165 = w22163 | w22164 ;
  assign w22166 = \pi074 ^ w22080 ;
  assign w22167 = ( ~w22087 & w22165 ) | ( ~w22087 & w22166 ) | ( w22165 & w22166 ) ;
  assign w22168 = w22166 | w22167 ;
  assign w22169 = \pi075 ^ w22074 ;
  assign w22170 = ( ~w22081 & w22168 ) | ( ~w22081 & w22169 ) | ( w22168 & w22169 ) ;
  assign w22171 = w22169 | w22170 ;
  assign w22172 = \pi076 ^ w22068 ;
  assign w22173 = ( ~w22075 & w22171 ) | ( ~w22075 & w22172 ) | ( w22171 & w22172 ) ;
  assign w22174 = w22172 | w22173 ;
  assign w22175 = \pi077 ^ w22062 ;
  assign w22176 = ( ~w22069 & w22174 ) | ( ~w22069 & w22175 ) | ( w22174 & w22175 ) ;
  assign w22177 = w22175 | w22176 ;
  assign w22178 = \pi078 ^ w22056 ;
  assign w22179 = ( ~w22063 & w22177 ) | ( ~w22063 & w22178 ) | ( w22177 & w22178 ) ;
  assign w22180 = w22178 | w22179 ;
  assign w22181 = \pi079 ^ w22050 ;
  assign w22182 = ( ~w22057 & w22180 ) | ( ~w22057 & w22181 ) | ( w22180 & w22181 ) ;
  assign w22183 = w22181 | w22182 ;
  assign w22184 = \pi080 ^ w22044 ;
  assign w22185 = ( ~w22051 & w22183 ) | ( ~w22051 & w22184 ) | ( w22183 & w22184 ) ;
  assign w22186 = w22184 | w22185 ;
  assign w22187 = \pi081 ^ w22038 ;
  assign w22188 = ( ~w22045 & w22186 ) | ( ~w22045 & w22187 ) | ( w22186 & w22187 ) ;
  assign w22189 = w22187 | w22188 ;
  assign w22190 = \pi082 ^ w22032 ;
  assign w22191 = ( ~w22039 & w22189 ) | ( ~w22039 & w22190 ) | ( w22189 & w22190 ) ;
  assign w22192 = w22190 | w22191 ;
  assign w22193 = \pi083 ^ w22026 ;
  assign w22194 = ( ~w22033 & w22192 ) | ( ~w22033 & w22193 ) | ( w22192 & w22193 ) ;
  assign w22195 = w22193 | w22194 ;
  assign w22196 = w21851 & w22021 ;
  assign w22197 = ~w21852 & w22015 ;
  assign w22198 = w22016 ^ w22197 ;
  assign w22199 = ~w22021 & w22198 ;
  assign w22200 = w22196 | w22199 ;
  assign w22201 = ~\pi084 & w22200 ;
  assign w22202 = ( \pi084 & ~w22196 ) | ( \pi084 & w22199 ) | ( ~w22196 & w22199 ) ;
  assign w22203 = ~w22199 & w22202 ;
  assign w22204 = w22201 | w22203 ;
  assign w22205 = ( ~w22027 & w22195 ) | ( ~w22027 & w22204 ) | ( w22195 & w22204 ) ;
  assign w22206 = ( w491 & ~w22204 ) | ( w491 & w22205 ) | ( ~w22204 & w22205 ) ;
  assign w22207 = w22204 | w22206 ;
  assign w22208 = ~w187 & w22200 ;
  assign w22209 = w22207 & ~w22208 ;
  assign w22210 = ~w22033 & w22192 ;
  assign w22211 = w22193 ^ w22210 ;
  assign w22212 = ~w22209 & w22211 ;
  assign w22213 = ( w22026 & w22207 ) | ( w22026 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22214 = ~w22208 & w22213 ;
  assign w22215 = w22212 | w22214 ;
  assign w22216 = ( ~w22027 & w22195 ) | ( ~w22027 & w22209 ) | ( w22195 & w22209 ) ;
  assign w22217 = w22204 ^ w22216 ;
  assign w22218 = ~w22209 & w22217 ;
  assign w22219 = ( w187 & ~w22200 ) | ( w187 & w22207 ) | ( ~w22200 & w22207 ) ;
  assign w22220 = w22200 & w22219 ;
  assign w22221 = w22218 | w22220 ;
  assign w22222 = ~\pi084 & w22215 ;
  assign w22223 = ~w22039 & w22189 ;
  assign w22224 = w22190 ^ w22223 ;
  assign w22225 = ~w22209 & w22224 ;
  assign w22226 = ( w22032 & w22207 ) | ( w22032 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22227 = ~w22208 & w22226 ;
  assign w22228 = w22225 | w22227 ;
  assign w22229 = ~\pi083 & w22228 ;
  assign w22230 = ~w22045 & w22186 ;
  assign w22231 = w22187 ^ w22230 ;
  assign w22232 = ~w22209 & w22231 ;
  assign w22233 = ( w22038 & w22207 ) | ( w22038 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22234 = ~w22208 & w22233 ;
  assign w22235 = w22232 | w22234 ;
  assign w22236 = ~\pi082 & w22235 ;
  assign w22237 = ~w22051 & w22183 ;
  assign w22238 = w22184 ^ w22237 ;
  assign w22239 = ~w22209 & w22238 ;
  assign w22240 = ( w22044 & w22207 ) | ( w22044 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22241 = ~w22208 & w22240 ;
  assign w22242 = w22239 | w22241 ;
  assign w22243 = ~\pi081 & w22242 ;
  assign w22244 = ~w22057 & w22180 ;
  assign w22245 = w22181 ^ w22244 ;
  assign w22246 = ~w22209 & w22245 ;
  assign w22247 = ( w22050 & w22207 ) | ( w22050 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22248 = ~w22208 & w22247 ;
  assign w22249 = w22246 | w22248 ;
  assign w22250 = ~\pi080 & w22249 ;
  assign w22251 = ~w22063 & w22177 ;
  assign w22252 = w22178 ^ w22251 ;
  assign w22253 = ~w22209 & w22252 ;
  assign w22254 = ( w22056 & w22207 ) | ( w22056 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22255 = ~w22208 & w22254 ;
  assign w22256 = w22253 | w22255 ;
  assign w22257 = ~\pi079 & w22256 ;
  assign w22258 = ~w22069 & w22174 ;
  assign w22259 = w22175 ^ w22258 ;
  assign w22260 = ~w22209 & w22259 ;
  assign w22261 = ( w22062 & w22207 ) | ( w22062 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22262 = ~w22208 & w22261 ;
  assign w22263 = w22260 | w22262 ;
  assign w22264 = ~\pi078 & w22263 ;
  assign w22265 = ~w22075 & w22171 ;
  assign w22266 = w22172 ^ w22265 ;
  assign w22267 = ~w22209 & w22266 ;
  assign w22268 = ( w22068 & w22207 ) | ( w22068 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22269 = ~w22208 & w22268 ;
  assign w22270 = w22267 | w22269 ;
  assign w22271 = ~\pi077 & w22270 ;
  assign w22272 = ~w22081 & w22168 ;
  assign w22273 = w22169 ^ w22272 ;
  assign w22274 = ~w22209 & w22273 ;
  assign w22275 = ( w22074 & w22207 ) | ( w22074 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22276 = ~w22208 & w22275 ;
  assign w22277 = w22274 | w22276 ;
  assign w22278 = ~\pi076 & w22277 ;
  assign w22279 = ~w22087 & w22165 ;
  assign w22280 = w22166 ^ w22279 ;
  assign w22281 = ~w22209 & w22280 ;
  assign w22282 = ( w22080 & w22207 ) | ( w22080 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22283 = ~w22208 & w22282 ;
  assign w22284 = w22281 | w22283 ;
  assign w22285 = ~\pi075 & w22284 ;
  assign w22286 = ~w22093 & w22162 ;
  assign w22287 = w22163 ^ w22286 ;
  assign w22288 = ~w22209 & w22287 ;
  assign w22289 = ( w22086 & w22207 ) | ( w22086 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22290 = ~w22208 & w22289 ;
  assign w22291 = w22288 | w22290 ;
  assign w22292 = ~\pi074 & w22291 ;
  assign w22293 = ~w22099 & w22159 ;
  assign w22294 = w22160 ^ w22293 ;
  assign w22295 = ~w22209 & w22294 ;
  assign w22296 = ( w22092 & w22207 ) | ( w22092 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22297 = ~w22208 & w22296 ;
  assign w22298 = w22295 | w22297 ;
  assign w22299 = ~\pi073 & w22298 ;
  assign w22300 = ~w22105 & w22156 ;
  assign w22301 = w22157 ^ w22300 ;
  assign w22302 = ~w22209 & w22301 ;
  assign w22303 = ( w22098 & w22207 ) | ( w22098 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22304 = ~w22208 & w22303 ;
  assign w22305 = w22302 | w22304 ;
  assign w22306 = ~\pi072 & w22305 ;
  assign w22307 = ~w22111 & w22153 ;
  assign w22308 = w22154 ^ w22307 ;
  assign w22309 = ~w22209 & w22308 ;
  assign w22310 = ( w22104 & w22207 ) | ( w22104 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22311 = ~w22208 & w22310 ;
  assign w22312 = w22309 | w22311 ;
  assign w22313 = ~\pi071 & w22312 ;
  assign w22314 = ~w22117 & w22150 ;
  assign w22315 = w22151 ^ w22314 ;
  assign w22316 = ~w22209 & w22315 ;
  assign w22317 = ( w22110 & w22207 ) | ( w22110 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22318 = ~w22208 & w22317 ;
  assign w22319 = w22316 | w22318 ;
  assign w22320 = ~\pi070 & w22319 ;
  assign w22321 = ~w22123 & w22147 ;
  assign w22322 = w22148 ^ w22321 ;
  assign w22323 = ~w22209 & w22322 ;
  assign w22324 = ( w22116 & w22207 ) | ( w22116 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22325 = ~w22208 & w22324 ;
  assign w22326 = w22323 | w22325 ;
  assign w22327 = ~\pi069 & w22326 ;
  assign w22328 = ~w22131 & w22144 ;
  assign w22329 = w22145 ^ w22328 ;
  assign w22330 = ~w22209 & w22329 ;
  assign w22331 = ( w22122 & w22207 ) | ( w22122 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22332 = ~w22208 & w22331 ;
  assign w22333 = w22330 | w22332 ;
  assign w22334 = ~\pi068 & w22333 ;
  assign w22335 = w22140 & ~w22141 ;
  assign w22336 = w22142 ^ w22335 ;
  assign w22337 = ~w22209 & w22336 ;
  assign w22338 = ( w22130 & w22207 ) | ( w22130 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22339 = ~w22208 & w22338 ;
  assign w22340 = w22337 | w22339 ;
  assign w22341 = ~\pi067 & w22340 ;
  assign w22342 = w2508 ^ w22020 ;
  assign w22343 = ( \pi044 & ~w2720 ) | ( \pi044 & w22342 ) | ( ~w2720 & w22342 ) ;
  assign w22344 = ( \pi044 & w2508 ) | ( \pi044 & w22343 ) | ( w2508 & w22343 ) ;
  assign w22345 = w2513 ^ w22344 ;
  assign w22346 = \pi065 ^ w22345 ;
  assign w22347 = ~w22209 & w22346 ;
  assign w22348 = ( w22135 & w22207 ) | ( w22135 & w22208 ) | ( w22207 & w22208 ) ;
  assign w22349 = ~w22208 & w22348 ;
  assign w22350 = w22347 | w22349 ;
  assign w22351 = ~\pi066 & w22350 ;
  assign w22352 = \pi066 ^ w22350 ;
  assign w22353 = ( \pi064 & ~w22209 ) | ( \pi064 & w22352 ) | ( ~w22209 & w22352 ) ;
  assign w22354 = \pi043 ^ w22353 ;
  assign w22355 = ( \pi065 & w2915 ) | ( \pi065 & ~w22354 ) | ( w2915 & ~w22354 ) ;
  assign w22356 = w22352 | w22355 ;
  assign w22357 = \pi067 ^ w22340 ;
  assign w22358 = ( ~w22351 & w22356 ) | ( ~w22351 & w22357 ) | ( w22356 & w22357 ) ;
  assign w22359 = w22357 | w22358 ;
  assign w22360 = \pi068 ^ w22333 ;
  assign w22361 = ( ~w22341 & w22359 ) | ( ~w22341 & w22360 ) | ( w22359 & w22360 ) ;
  assign w22362 = w22360 | w22361 ;
  assign w22363 = \pi069 ^ w22326 ;
  assign w22364 = ( ~w22334 & w22362 ) | ( ~w22334 & w22363 ) | ( w22362 & w22363 ) ;
  assign w22365 = w22363 | w22364 ;
  assign w22366 = \pi070 ^ w22319 ;
  assign w22367 = ( ~w22327 & w22365 ) | ( ~w22327 & w22366 ) | ( w22365 & w22366 ) ;
  assign w22368 = w22366 | w22367 ;
  assign w22369 = \pi071 ^ w22312 ;
  assign w22370 = ( ~w22320 & w22368 ) | ( ~w22320 & w22369 ) | ( w22368 & w22369 ) ;
  assign w22371 = w22369 | w22370 ;
  assign w22372 = \pi072 ^ w22305 ;
  assign w22373 = ( ~w22313 & w22371 ) | ( ~w22313 & w22372 ) | ( w22371 & w22372 ) ;
  assign w22374 = w22372 | w22373 ;
  assign w22375 = \pi073 ^ w22298 ;
  assign w22376 = ( ~w22306 & w22374 ) | ( ~w22306 & w22375 ) | ( w22374 & w22375 ) ;
  assign w22377 = w22375 | w22376 ;
  assign w22378 = \pi074 ^ w22291 ;
  assign w22379 = ( ~w22299 & w22377 ) | ( ~w22299 & w22378 ) | ( w22377 & w22378 ) ;
  assign w22380 = w22378 | w22379 ;
  assign w22381 = \pi075 ^ w22284 ;
  assign w22382 = ( ~w22292 & w22380 ) | ( ~w22292 & w22381 ) | ( w22380 & w22381 ) ;
  assign w22383 = w22381 | w22382 ;
  assign w22384 = \pi076 ^ w22277 ;
  assign w22385 = ( ~w22285 & w22383 ) | ( ~w22285 & w22384 ) | ( w22383 & w22384 ) ;
  assign w22386 = w22384 | w22385 ;
  assign w22387 = \pi077 ^ w22270 ;
  assign w22388 = ( ~w22278 & w22386 ) | ( ~w22278 & w22387 ) | ( w22386 & w22387 ) ;
  assign w22389 = w22387 | w22388 ;
  assign w22390 = \pi078 ^ w22263 ;
  assign w22391 = ( ~w22271 & w22389 ) | ( ~w22271 & w22390 ) | ( w22389 & w22390 ) ;
  assign w22392 = w22390 | w22391 ;
  assign w22393 = \pi079 ^ w22256 ;
  assign w22394 = ( ~w22264 & w22392 ) | ( ~w22264 & w22393 ) | ( w22392 & w22393 ) ;
  assign w22395 = w22393 | w22394 ;
  assign w22396 = \pi080 ^ w22249 ;
  assign w22397 = ( ~w22257 & w22395 ) | ( ~w22257 & w22396 ) | ( w22395 & w22396 ) ;
  assign w22398 = w22396 | w22397 ;
  assign w22399 = \pi081 ^ w22242 ;
  assign w22400 = ( ~w22250 & w22398 ) | ( ~w22250 & w22399 ) | ( w22398 & w22399 ) ;
  assign w22401 = w22399 | w22400 ;
  assign w22402 = \pi082 ^ w22235 ;
  assign w22403 = ( ~w22243 & w22401 ) | ( ~w22243 & w22402 ) | ( w22401 & w22402 ) ;
  assign w22404 = w22402 | w22403 ;
  assign w22405 = \pi083 ^ w22228 ;
  assign w22406 = ( ~w22236 & w22404 ) | ( ~w22236 & w22405 ) | ( w22404 & w22405 ) ;
  assign w22407 = w22405 | w22406 ;
  assign w22408 = \pi084 ^ w22215 ;
  assign w22409 = ( ~w22229 & w22407 ) | ( ~w22229 & w22408 ) | ( w22407 & w22408 ) ;
  assign w22410 = w22408 | w22409 ;
  assign w22411 = \pi085 ^ w22221 ;
  assign w22412 = w22222 & ~w22411 ;
  assign w22413 = ( w22410 & w22411 ) | ( w22410 & ~w22412 ) | ( w22411 & ~w22412 ) ;
  assign w22414 = ~\pi085 & w22221 ;
  assign w22415 = w22413 & ~w22414 ;
  assign w22416 = w2799 | w22415 ;
  assign w22417 = w22215 & w22416 ;
  assign w22418 = ~w22229 & w22407 ;
  assign w22419 = w22408 ^ w22418 ;
  assign w22420 = ~w22416 & w22419 ;
  assign w22421 = w22417 | w22420 ;
  assign w22422 = w22221 & w22416 ;
  assign w22423 = ~w22222 & w22410 ;
  assign w22424 = w22411 ^ w22423 ;
  assign w22425 = ~w22416 & w22424 ;
  assign w22426 = w22422 | w22425 ;
  assign w22427 = ~\pi085 & w22421 ;
  assign w22428 = w22228 & w22416 ;
  assign w22429 = ~w22236 & w22404 ;
  assign w22430 = w22405 ^ w22429 ;
  assign w22431 = ~w22416 & w22430 ;
  assign w22432 = w22428 | w22431 ;
  assign w22433 = ~\pi084 & w22432 ;
  assign w22434 = w22235 & w22416 ;
  assign w22435 = ~w22243 & w22401 ;
  assign w22436 = w22402 ^ w22435 ;
  assign w22437 = ~w22416 & w22436 ;
  assign w22438 = w22434 | w22437 ;
  assign w22439 = ~\pi083 & w22438 ;
  assign w22440 = w22242 & w22416 ;
  assign w22441 = ~w22250 & w22398 ;
  assign w22442 = w22399 ^ w22441 ;
  assign w22443 = ~w22416 & w22442 ;
  assign w22444 = w22440 | w22443 ;
  assign w22445 = ~\pi082 & w22444 ;
  assign w22446 = w22249 & w22416 ;
  assign w22447 = ~w22257 & w22395 ;
  assign w22448 = w22396 ^ w22447 ;
  assign w22449 = ~w22416 & w22448 ;
  assign w22450 = w22446 | w22449 ;
  assign w22451 = ~\pi081 & w22450 ;
  assign w22452 = w22256 & w22416 ;
  assign w22453 = ~w22264 & w22392 ;
  assign w22454 = w22393 ^ w22453 ;
  assign w22455 = ~w22416 & w22454 ;
  assign w22456 = w22452 | w22455 ;
  assign w22457 = ~\pi080 & w22456 ;
  assign w22458 = w22263 & w22416 ;
  assign w22459 = ~w22271 & w22389 ;
  assign w22460 = w22390 ^ w22459 ;
  assign w22461 = ~w22416 & w22460 ;
  assign w22462 = w22458 | w22461 ;
  assign w22463 = ~\pi079 & w22462 ;
  assign w22464 = w22270 & w22416 ;
  assign w22465 = ~w22278 & w22386 ;
  assign w22466 = w22387 ^ w22465 ;
  assign w22467 = ~w22416 & w22466 ;
  assign w22468 = w22464 | w22467 ;
  assign w22469 = ~\pi078 & w22468 ;
  assign w22470 = w22277 & w22416 ;
  assign w22471 = ~w22285 & w22383 ;
  assign w22472 = w22384 ^ w22471 ;
  assign w22473 = ~w22416 & w22472 ;
  assign w22474 = w22470 | w22473 ;
  assign w22475 = ~\pi077 & w22474 ;
  assign w22476 = w22284 & w22416 ;
  assign w22477 = ~w22292 & w22380 ;
  assign w22478 = w22381 ^ w22477 ;
  assign w22479 = ~w22416 & w22478 ;
  assign w22480 = w22476 | w22479 ;
  assign w22481 = ~\pi076 & w22480 ;
  assign w22482 = w22291 & w22416 ;
  assign w22483 = ~w22299 & w22377 ;
  assign w22484 = w22378 ^ w22483 ;
  assign w22485 = ~w22416 & w22484 ;
  assign w22486 = w22482 | w22485 ;
  assign w22487 = ~\pi075 & w22486 ;
  assign w22488 = w22298 & w22416 ;
  assign w22489 = ~w22306 & w22374 ;
  assign w22490 = w22375 ^ w22489 ;
  assign w22491 = ~w22416 & w22490 ;
  assign w22492 = w22488 | w22491 ;
  assign w22493 = ~\pi074 & w22492 ;
  assign w22494 = w22305 & w22416 ;
  assign w22495 = ~w22313 & w22371 ;
  assign w22496 = w22372 ^ w22495 ;
  assign w22497 = ~w22416 & w22496 ;
  assign w22498 = w22494 | w22497 ;
  assign w22499 = ~\pi073 & w22498 ;
  assign w22500 = w22312 & w22416 ;
  assign w22501 = ~w22320 & w22368 ;
  assign w22502 = w22369 ^ w22501 ;
  assign w22503 = ~w22416 & w22502 ;
  assign w22504 = w22500 | w22503 ;
  assign w22505 = ~\pi072 & w22504 ;
  assign w22506 = w22319 & w22416 ;
  assign w22507 = ~w22327 & w22365 ;
  assign w22508 = w22366 ^ w22507 ;
  assign w22509 = ~w22416 & w22508 ;
  assign w22510 = w22506 | w22509 ;
  assign w22511 = ~\pi071 & w22510 ;
  assign w22512 = w22326 & w22416 ;
  assign w22513 = ~w22334 & w22362 ;
  assign w22514 = w22363 ^ w22513 ;
  assign w22515 = ~w22416 & w22514 ;
  assign w22516 = w22512 | w22515 ;
  assign w22517 = ~\pi070 & w22516 ;
  assign w22518 = w22333 & w22416 ;
  assign w22519 = ~w22341 & w22359 ;
  assign w22520 = w22360 ^ w22519 ;
  assign w22521 = ~w22416 & w22520 ;
  assign w22522 = w22518 | w22521 ;
  assign w22523 = ~\pi069 & w22522 ;
  assign w22524 = w22340 & w22416 ;
  assign w22525 = ~w22351 & w22356 ;
  assign w22526 = w22357 ^ w22525 ;
  assign w22527 = ~w22416 & w22526 ;
  assign w22528 = w22524 | w22527 ;
  assign w22529 = ~\pi068 & w22528 ;
  assign w22530 = w22350 & w22416 ;
  assign w22531 = \pi064 & ~w22209 ;
  assign w22532 = \pi043 ^ w22531 ;
  assign w22533 = ( \pi065 & w2915 ) | ( \pi065 & ~w22532 ) | ( w2915 & ~w22532 ) ;
  assign w22534 = w22352 ^ w22533 ;
  assign w22535 = ( w2799 & w22415 ) | ( w2799 & w22534 ) | ( w22415 & w22534 ) ;
  assign w22536 = w22534 & ~w22535 ;
  assign w22537 = w22530 | w22536 ;
  assign w22538 = ~\pi067 & w22537 ;
  assign w22539 = \pi042 ^ w22209 ;
  assign w22540 = ( \pi064 & w2799 ) | ( \pi064 & w22539 ) | ( w2799 & w22539 ) ;
  assign w22541 = w2922 ^ w22540 ;
  assign w22542 = ~w2799 & w22541 ;
  assign w22543 = ~w22415 & w22542 ;
  assign w22544 = ( ~\pi064 & w22209 ) | ( ~\pi064 & w22416 ) | ( w22209 & w22416 ) ;
  assign w22545 = \pi043 ^ w22544 ;
  assign w22546 = w22416 & ~w22545 ;
  assign w22547 = w22543 | w22546 ;
  assign w22548 = ~\pi066 & w22547 ;
  assign w22549 = ( \pi042 & ~w2939 ) | ( \pi042 & w22415 ) | ( ~w2939 & w22415 ) ;
  assign w22550 = \pi042 & w22549 ;
  assign w22551 = w2948 & ~w22415 ;
  assign w22552 = w22550 | w22551 ;
  assign w22553 = \pi065 ^ w22552 ;
  assign w22554 = w2951 | w22553 ;
  assign w22555 = ~\pi065 & w22552 ;
  assign w22556 = w22416 | w22543 ;
  assign w22557 = ( w22532 & w22543 ) | ( w22532 & w22556 ) | ( w22543 & w22556 ) ;
  assign w22558 = \pi066 ^ w22557 ;
  assign w22559 = ( w22554 & ~w22555 ) | ( w22554 & w22558 ) | ( ~w22555 & w22558 ) ;
  assign w22560 = w22558 | w22559 ;
  assign w22561 = \pi067 ^ w22537 ;
  assign w22562 = ( ~w22548 & w22560 ) | ( ~w22548 & w22561 ) | ( w22560 & w22561 ) ;
  assign w22563 = w22561 | w22562 ;
  assign w22564 = \pi068 ^ w22528 ;
  assign w22565 = ( ~w22538 & w22563 ) | ( ~w22538 & w22564 ) | ( w22563 & w22564 ) ;
  assign w22566 = w22564 | w22565 ;
  assign w22567 = \pi069 ^ w22522 ;
  assign w22568 = ( ~w22529 & w22566 ) | ( ~w22529 & w22567 ) | ( w22566 & w22567 ) ;
  assign w22569 = w22567 | w22568 ;
  assign w22570 = \pi070 ^ w22516 ;
  assign w22571 = ( ~w22523 & w22569 ) | ( ~w22523 & w22570 ) | ( w22569 & w22570 ) ;
  assign w22572 = w22570 | w22571 ;
  assign w22573 = \pi071 ^ w22510 ;
  assign w22574 = ( ~w22517 & w22572 ) | ( ~w22517 & w22573 ) | ( w22572 & w22573 ) ;
  assign w22575 = w22573 | w22574 ;
  assign w22576 = \pi072 ^ w22504 ;
  assign w22577 = ( ~w22511 & w22575 ) | ( ~w22511 & w22576 ) | ( w22575 & w22576 ) ;
  assign w22578 = w22576 | w22577 ;
  assign w22579 = \pi073 ^ w22498 ;
  assign w22580 = ( ~w22505 & w22578 ) | ( ~w22505 & w22579 ) | ( w22578 & w22579 ) ;
  assign w22581 = w22579 | w22580 ;
  assign w22582 = \pi074 ^ w22492 ;
  assign w22583 = ( ~w22499 & w22581 ) | ( ~w22499 & w22582 ) | ( w22581 & w22582 ) ;
  assign w22584 = w22582 | w22583 ;
  assign w22585 = \pi075 ^ w22486 ;
  assign w22586 = ( ~w22493 & w22584 ) | ( ~w22493 & w22585 ) | ( w22584 & w22585 ) ;
  assign w22587 = w22585 | w22586 ;
  assign w22588 = \pi076 ^ w22480 ;
  assign w22589 = ( ~w22487 & w22587 ) | ( ~w22487 & w22588 ) | ( w22587 & w22588 ) ;
  assign w22590 = w22588 | w22589 ;
  assign w22591 = \pi077 ^ w22474 ;
  assign w22592 = ( ~w22481 & w22590 ) | ( ~w22481 & w22591 ) | ( w22590 & w22591 ) ;
  assign w22593 = w22591 | w22592 ;
  assign w22594 = \pi078 ^ w22468 ;
  assign w22595 = ( ~w22475 & w22593 ) | ( ~w22475 & w22594 ) | ( w22593 & w22594 ) ;
  assign w22596 = w22594 | w22595 ;
  assign w22597 = \pi079 ^ w22462 ;
  assign w22598 = ( ~w22469 & w22596 ) | ( ~w22469 & w22597 ) | ( w22596 & w22597 ) ;
  assign w22599 = w22597 | w22598 ;
  assign w22600 = \pi080 ^ w22456 ;
  assign w22601 = ( ~w22463 & w22599 ) | ( ~w22463 & w22600 ) | ( w22599 & w22600 ) ;
  assign w22602 = w22600 | w22601 ;
  assign w22603 = \pi081 ^ w22450 ;
  assign w22604 = ( ~w22457 & w22602 ) | ( ~w22457 & w22603 ) | ( w22602 & w22603 ) ;
  assign w22605 = w22603 | w22604 ;
  assign w22606 = \pi082 ^ w22444 ;
  assign w22607 = ( ~w22451 & w22605 ) | ( ~w22451 & w22606 ) | ( w22605 & w22606 ) ;
  assign w22608 = w22606 | w22607 ;
  assign w22609 = \pi083 ^ w22438 ;
  assign w22610 = ( ~w22445 & w22608 ) | ( ~w22445 & w22609 ) | ( w22608 & w22609 ) ;
  assign w22611 = w22609 | w22610 ;
  assign w22612 = \pi084 ^ w22432 ;
  assign w22613 = ( ~w22439 & w22611 ) | ( ~w22439 & w22612 ) | ( w22611 & w22612 ) ;
  assign w22614 = w22612 | w22613 ;
  assign w22615 = \pi085 ^ w22421 ;
  assign w22616 = ( ~w22433 & w22614 ) | ( ~w22433 & w22615 ) | ( w22614 & w22615 ) ;
  assign w22617 = w22615 | w22616 ;
  assign w22618 = \pi086 ^ w22426 ;
  assign w22619 = w22427 & ~w22618 ;
  assign w22620 = ( w22617 & w22618 ) | ( w22617 & ~w22619 ) | ( w22618 & ~w22619 ) ;
  assign w22621 = ~\pi086 & w22426 ;
  assign w22622 = w22620 & ~w22621 ;
  assign w22623 = w3025 | w22622 ;
  assign w22624 = w22421 & w22623 ;
  assign w22625 = ~w22433 & w22614 ;
  assign w22626 = w22615 ^ w22625 ;
  assign w22627 = ~w22623 & w22626 ;
  assign w22628 = w22624 | w22627 ;
  assign w22629 = ~\pi086 & w22628 ;
  assign w22630 = w22432 & w22623 ;
  assign w22631 = ~w22439 & w22611 ;
  assign w22632 = w22612 ^ w22631 ;
  assign w22633 = ~w22623 & w22632 ;
  assign w22634 = w22630 | w22633 ;
  assign w22635 = ~\pi085 & w22634 ;
  assign w22636 = w22438 & w22623 ;
  assign w22637 = ~w22445 & w22608 ;
  assign w22638 = w22609 ^ w22637 ;
  assign w22639 = ~w22623 & w22638 ;
  assign w22640 = w22636 | w22639 ;
  assign w22641 = ~\pi084 & w22640 ;
  assign w22642 = w22444 & w22623 ;
  assign w22643 = ~w22451 & w22605 ;
  assign w22644 = w22606 ^ w22643 ;
  assign w22645 = ~w22623 & w22644 ;
  assign w22646 = w22642 | w22645 ;
  assign w22647 = ~\pi083 & w22646 ;
  assign w22648 = w22450 & w22623 ;
  assign w22649 = ~w22457 & w22602 ;
  assign w22650 = w22603 ^ w22649 ;
  assign w22651 = ~w22623 & w22650 ;
  assign w22652 = w22648 | w22651 ;
  assign w22653 = ~\pi082 & w22652 ;
  assign w22654 = w22456 & w22623 ;
  assign w22655 = ~w22463 & w22599 ;
  assign w22656 = w22600 ^ w22655 ;
  assign w22657 = ~w22623 & w22656 ;
  assign w22658 = w22654 | w22657 ;
  assign w22659 = ~\pi081 & w22658 ;
  assign w22660 = w22462 & w22623 ;
  assign w22661 = ~w22469 & w22596 ;
  assign w22662 = w22597 ^ w22661 ;
  assign w22663 = ~w22623 & w22662 ;
  assign w22664 = w22660 | w22663 ;
  assign w22665 = ~\pi080 & w22664 ;
  assign w22666 = w22468 & w22623 ;
  assign w22667 = ~w22475 & w22593 ;
  assign w22668 = w22594 ^ w22667 ;
  assign w22669 = ~w22623 & w22668 ;
  assign w22670 = w22666 | w22669 ;
  assign w22671 = ~\pi079 & w22670 ;
  assign w22672 = w22474 & w22623 ;
  assign w22673 = ~w22481 & w22590 ;
  assign w22674 = w22591 ^ w22673 ;
  assign w22675 = ~w22623 & w22674 ;
  assign w22676 = w22672 | w22675 ;
  assign w22677 = ~\pi078 & w22676 ;
  assign w22678 = w22480 & w22623 ;
  assign w22679 = ~w22487 & w22587 ;
  assign w22680 = w22588 ^ w22679 ;
  assign w22681 = ~w22623 & w22680 ;
  assign w22682 = w22678 | w22681 ;
  assign w22683 = ~\pi077 & w22682 ;
  assign w22684 = w22486 & w22623 ;
  assign w22685 = ~w22493 & w22584 ;
  assign w22686 = w22585 ^ w22685 ;
  assign w22687 = ~w22623 & w22686 ;
  assign w22688 = w22684 | w22687 ;
  assign w22689 = ~\pi076 & w22688 ;
  assign w22690 = w22492 & w22623 ;
  assign w22691 = ~w22499 & w22581 ;
  assign w22692 = w22582 ^ w22691 ;
  assign w22693 = ~w22623 & w22692 ;
  assign w22694 = w22690 | w22693 ;
  assign w22695 = ~\pi075 & w22694 ;
  assign w22696 = w22498 & w22623 ;
  assign w22697 = ~w22505 & w22578 ;
  assign w22698 = w22579 ^ w22697 ;
  assign w22699 = ~w22623 & w22698 ;
  assign w22700 = w22696 | w22699 ;
  assign w22701 = ~\pi074 & w22700 ;
  assign w22702 = w22504 & w22623 ;
  assign w22703 = ~w22511 & w22575 ;
  assign w22704 = w22576 ^ w22703 ;
  assign w22705 = ~w22623 & w22704 ;
  assign w22706 = w22702 | w22705 ;
  assign w22707 = ~\pi073 & w22706 ;
  assign w22708 = w22510 & w22623 ;
  assign w22709 = ~w22517 & w22572 ;
  assign w22710 = w22573 ^ w22709 ;
  assign w22711 = ~w22623 & w22710 ;
  assign w22712 = w22708 | w22711 ;
  assign w22713 = ~\pi072 & w22712 ;
  assign w22714 = w22516 & w22623 ;
  assign w22715 = ~w22523 & w22569 ;
  assign w22716 = w22570 ^ w22715 ;
  assign w22717 = ~w22623 & w22716 ;
  assign w22718 = w22714 | w22717 ;
  assign w22719 = ~\pi071 & w22718 ;
  assign w22720 = w22522 & w22623 ;
  assign w22721 = ~w22529 & w22566 ;
  assign w22722 = w22567 ^ w22721 ;
  assign w22723 = ~w22623 & w22722 ;
  assign w22724 = w22720 | w22723 ;
  assign w22725 = ~\pi070 & w22724 ;
  assign w22726 = w22528 & w22623 ;
  assign w22727 = ~w22538 & w22563 ;
  assign w22728 = w22564 ^ w22727 ;
  assign w22729 = ~w22623 & w22728 ;
  assign w22730 = w22726 | w22729 ;
  assign w22731 = ~\pi069 & w22730 ;
  assign w22732 = w22537 & w22623 ;
  assign w22733 = ~w22548 & w22560 ;
  assign w22734 = w22561 ^ w22733 ;
  assign w22735 = ~w22623 & w22734 ;
  assign w22736 = w22732 | w22735 ;
  assign w22737 = ~\pi068 & w22736 ;
  assign w22738 = w22547 & w22623 ;
  assign w22739 = w22554 & ~w22555 ;
  assign w22740 = w22558 ^ w22739 ;
  assign w22741 = ~w22623 & w22740 ;
  assign w22742 = w22738 | w22741 ;
  assign w22743 = ~\pi067 & w22742 ;
  assign w22744 = w2951 ^ w22553 ;
  assign w22745 = ~w3025 & w22744 ;
  assign w22746 = ( w3025 & w22552 ) | ( w3025 & w22622 ) | ( w22552 & w22622 ) ;
  assign w22747 = w22552 & w22746 ;
  assign w22748 = w22622 | w22745 ;
  assign w22749 = ( ~w22622 & w22747 ) | ( ~w22622 & w22748 ) | ( w22747 & w22748 ) ;
  assign w22750 = ~\pi066 & w22749 ;
  assign w22751 = ( \pi041 & ~w3157 ) | ( \pi041 & w22622 ) | ( ~w3157 & w22622 ) ;
  assign w22752 = \pi041 & w22751 ;
  assign w22753 = w3165 & ~w22622 ;
  assign w22754 = w22752 | w22753 ;
  assign w22755 = ( ~w3168 & w22752 ) | ( ~w3168 & w22753 ) | ( w22752 & w22753 ) ;
  assign w22756 = \pi065 ^ w22755 ;
  assign w22757 = w3168 | w22756 ;
  assign w22758 = ~\pi065 & w22754 ;
  assign w22759 = ~w22622 & w22745 ;
  assign w22760 = ( w3025 & ~w22622 ) | ( w3025 & w22759 ) | ( ~w22622 & w22759 ) ;
  assign w22761 = w22552 | w22759 ;
  assign w22762 = ( w22622 & w22760 ) | ( w22622 & w22761 ) | ( w22760 & w22761 ) ;
  assign w22763 = \pi066 ^ w22762 ;
  assign w22764 = ( w22757 & ~w22758 ) | ( w22757 & w22763 ) | ( ~w22758 & w22763 ) ;
  assign w22765 = w22763 | w22764 ;
  assign w22766 = \pi067 ^ w22742 ;
  assign w22767 = ( ~w22750 & w22765 ) | ( ~w22750 & w22766 ) | ( w22765 & w22766 ) ;
  assign w22768 = w22766 | w22767 ;
  assign w22769 = \pi068 ^ w22736 ;
  assign w22770 = ( ~w22743 & w22768 ) | ( ~w22743 & w22769 ) | ( w22768 & w22769 ) ;
  assign w22771 = w22769 | w22770 ;
  assign w22772 = \pi069 ^ w22730 ;
  assign w22773 = ( ~w22737 & w22771 ) | ( ~w22737 & w22772 ) | ( w22771 & w22772 ) ;
  assign w22774 = w22772 | w22773 ;
  assign w22775 = \pi070 ^ w22724 ;
  assign w22776 = ( ~w22731 & w22774 ) | ( ~w22731 & w22775 ) | ( w22774 & w22775 ) ;
  assign w22777 = w22775 | w22776 ;
  assign w22778 = \pi071 ^ w22718 ;
  assign w22779 = ( ~w22725 & w22777 ) | ( ~w22725 & w22778 ) | ( w22777 & w22778 ) ;
  assign w22780 = w22778 | w22779 ;
  assign w22781 = \pi072 ^ w22712 ;
  assign w22782 = ( ~w22719 & w22780 ) | ( ~w22719 & w22781 ) | ( w22780 & w22781 ) ;
  assign w22783 = w22781 | w22782 ;
  assign w22784 = \pi073 ^ w22706 ;
  assign w22785 = ( ~w22713 & w22783 ) | ( ~w22713 & w22784 ) | ( w22783 & w22784 ) ;
  assign w22786 = w22784 | w22785 ;
  assign w22787 = \pi074 ^ w22700 ;
  assign w22788 = ( ~w22707 & w22786 ) | ( ~w22707 & w22787 ) | ( w22786 & w22787 ) ;
  assign w22789 = w22787 | w22788 ;
  assign w22790 = \pi075 ^ w22694 ;
  assign w22791 = ( ~w22701 & w22789 ) | ( ~w22701 & w22790 ) | ( w22789 & w22790 ) ;
  assign w22792 = w22790 | w22791 ;
  assign w22793 = \pi076 ^ w22688 ;
  assign w22794 = ( ~w22695 & w22792 ) | ( ~w22695 & w22793 ) | ( w22792 & w22793 ) ;
  assign w22795 = w22793 | w22794 ;
  assign w22796 = \pi077 ^ w22682 ;
  assign w22797 = ( ~w22689 & w22795 ) | ( ~w22689 & w22796 ) | ( w22795 & w22796 ) ;
  assign w22798 = w22796 | w22797 ;
  assign w22799 = \pi078 ^ w22676 ;
  assign w22800 = ( ~w22683 & w22798 ) | ( ~w22683 & w22799 ) | ( w22798 & w22799 ) ;
  assign w22801 = w22799 | w22800 ;
  assign w22802 = \pi079 ^ w22670 ;
  assign w22803 = ( ~w22677 & w22801 ) | ( ~w22677 & w22802 ) | ( w22801 & w22802 ) ;
  assign w22804 = w22802 | w22803 ;
  assign w22805 = \pi080 ^ w22664 ;
  assign w22806 = ( ~w22671 & w22804 ) | ( ~w22671 & w22805 ) | ( w22804 & w22805 ) ;
  assign w22807 = w22805 | w22806 ;
  assign w22808 = \pi081 ^ w22658 ;
  assign w22809 = ( ~w22665 & w22807 ) | ( ~w22665 & w22808 ) | ( w22807 & w22808 ) ;
  assign w22810 = w22808 | w22809 ;
  assign w22811 = \pi082 ^ w22652 ;
  assign w22812 = ( ~w22659 & w22810 ) | ( ~w22659 & w22811 ) | ( w22810 & w22811 ) ;
  assign w22813 = w22811 | w22812 ;
  assign w22814 = \pi083 ^ w22646 ;
  assign w22815 = ( ~w22653 & w22813 ) | ( ~w22653 & w22814 ) | ( w22813 & w22814 ) ;
  assign w22816 = w22814 | w22815 ;
  assign w22817 = \pi084 ^ w22640 ;
  assign w22818 = ( ~w22647 & w22816 ) | ( ~w22647 & w22817 ) | ( w22816 & w22817 ) ;
  assign w22819 = w22817 | w22818 ;
  assign w22820 = \pi085 ^ w22634 ;
  assign w22821 = ( ~w22641 & w22819 ) | ( ~w22641 & w22820 ) | ( w22819 & w22820 ) ;
  assign w22822 = w22820 | w22821 ;
  assign w22823 = \pi086 ^ w22628 ;
  assign w22824 = ( ~w22635 & w22822 ) | ( ~w22635 & w22823 ) | ( w22822 & w22823 ) ;
  assign w22825 = w22823 | w22824 ;
  assign w22826 = w22426 & w22623 ;
  assign w22827 = ~w22427 & w22617 ;
  assign w22828 = w22618 ^ w22827 ;
  assign w22829 = ~w22623 & w22828 ;
  assign w22830 = w22826 | w22829 ;
  assign w22831 = ~\pi087 & w22830 ;
  assign w22832 = ( \pi087 & ~w22826 ) | ( \pi087 & w22829 ) | ( ~w22826 & w22829 ) ;
  assign w22833 = ~w22829 & w22832 ;
  assign w22834 = w3248 | w22833 ;
  assign w22835 = ( w201 & w22831 ) | ( w201 & ~w22833 ) | ( w22831 & ~w22833 ) ;
  assign w22836 = w22834 | w22835 ;
  assign w22837 = ( ~w22629 & w22825 ) | ( ~w22629 & w22836 ) | ( w22825 & w22836 ) ;
  assign w22838 = w22836 | w22837 ;
  assign w22839 = ~w3025 & w22830 ;
  assign w22840 = w22838 & ~w22839 ;
  assign w22841 = ~w22635 & w22822 ;
  assign w22842 = w22823 ^ w22841 ;
  assign w22843 = ~w22840 & w22842 ;
  assign w22844 = ( w22628 & w22838 ) | ( w22628 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22845 = ~w22839 & w22844 ;
  assign w22846 = w22843 | w22845 ;
  assign w22847 = w22831 | w22833 ;
  assign w22848 = ( ~w22629 & w22825 ) | ( ~w22629 & w22840 ) | ( w22825 & w22840 ) ;
  assign w22849 = w22847 ^ w22848 ;
  assign w22850 = ~w22840 & w22849 ;
  assign w22851 = ( w3025 & ~w22830 ) | ( w3025 & w22838 ) | ( ~w22830 & w22838 ) ;
  assign w22852 = w22830 & w22851 ;
  assign w22853 = w22850 | w22852 ;
  assign w22854 = ~\pi087 & w22846 ;
  assign w22855 = ~w22641 & w22819 ;
  assign w22856 = w22820 ^ w22855 ;
  assign w22857 = ~w22840 & w22856 ;
  assign w22858 = ( w22634 & w22838 ) | ( w22634 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22859 = ~w22839 & w22858 ;
  assign w22860 = w22857 | w22859 ;
  assign w22861 = ~\pi086 & w22860 ;
  assign w22862 = ~w22647 & w22816 ;
  assign w22863 = w22817 ^ w22862 ;
  assign w22864 = ~w22840 & w22863 ;
  assign w22865 = ( w22640 & w22838 ) | ( w22640 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22866 = ~w22839 & w22865 ;
  assign w22867 = w22864 | w22866 ;
  assign w22868 = ~\pi085 & w22867 ;
  assign w22869 = ~w22653 & w22813 ;
  assign w22870 = w22814 ^ w22869 ;
  assign w22871 = ~w22840 & w22870 ;
  assign w22872 = ( w22646 & w22838 ) | ( w22646 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22873 = ~w22839 & w22872 ;
  assign w22874 = w22871 | w22873 ;
  assign w22875 = ~\pi084 & w22874 ;
  assign w22876 = ~w22659 & w22810 ;
  assign w22877 = w22811 ^ w22876 ;
  assign w22878 = ~w22840 & w22877 ;
  assign w22879 = ( w22652 & w22838 ) | ( w22652 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22880 = ~w22839 & w22879 ;
  assign w22881 = w22878 | w22880 ;
  assign w22882 = ~\pi083 & w22881 ;
  assign w22883 = ~w22665 & w22807 ;
  assign w22884 = w22808 ^ w22883 ;
  assign w22885 = ~w22840 & w22884 ;
  assign w22886 = ( w22658 & w22838 ) | ( w22658 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22887 = ~w22839 & w22886 ;
  assign w22888 = w22885 | w22887 ;
  assign w22889 = ~\pi082 & w22888 ;
  assign w22890 = ~w22671 & w22804 ;
  assign w22891 = w22805 ^ w22890 ;
  assign w22892 = ~w22840 & w22891 ;
  assign w22893 = ( w22664 & w22838 ) | ( w22664 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22894 = ~w22839 & w22893 ;
  assign w22895 = w22892 | w22894 ;
  assign w22896 = ~\pi081 & w22895 ;
  assign w22897 = ~w22677 & w22801 ;
  assign w22898 = w22802 ^ w22897 ;
  assign w22899 = ~w22840 & w22898 ;
  assign w22900 = ( w22670 & w22838 ) | ( w22670 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22901 = ~w22839 & w22900 ;
  assign w22902 = w22899 | w22901 ;
  assign w22903 = ~\pi080 & w22902 ;
  assign w22904 = ~w22683 & w22798 ;
  assign w22905 = w22799 ^ w22904 ;
  assign w22906 = ~w22840 & w22905 ;
  assign w22907 = ( w22676 & w22838 ) | ( w22676 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22908 = ~w22839 & w22907 ;
  assign w22909 = w22906 | w22908 ;
  assign w22910 = ~\pi079 & w22909 ;
  assign w22911 = ~w22689 & w22795 ;
  assign w22912 = w22796 ^ w22911 ;
  assign w22913 = ~w22840 & w22912 ;
  assign w22914 = ( w22682 & w22838 ) | ( w22682 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22915 = ~w22839 & w22914 ;
  assign w22916 = w22913 | w22915 ;
  assign w22917 = ~\pi078 & w22916 ;
  assign w22918 = ~w22695 & w22792 ;
  assign w22919 = w22793 ^ w22918 ;
  assign w22920 = ~w22840 & w22919 ;
  assign w22921 = ( w22688 & w22838 ) | ( w22688 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22922 = ~w22839 & w22921 ;
  assign w22923 = w22920 | w22922 ;
  assign w22924 = ~\pi077 & w22923 ;
  assign w22925 = ~w22701 & w22789 ;
  assign w22926 = w22790 ^ w22925 ;
  assign w22927 = ~w22840 & w22926 ;
  assign w22928 = ( w22694 & w22838 ) | ( w22694 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22929 = ~w22839 & w22928 ;
  assign w22930 = w22927 | w22929 ;
  assign w22931 = ~\pi076 & w22930 ;
  assign w22932 = ~w22707 & w22786 ;
  assign w22933 = w22787 ^ w22932 ;
  assign w22934 = ~w22840 & w22933 ;
  assign w22935 = ( w22700 & w22838 ) | ( w22700 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22936 = ~w22839 & w22935 ;
  assign w22937 = w22934 | w22936 ;
  assign w22938 = ~\pi075 & w22937 ;
  assign w22939 = ~w22713 & w22783 ;
  assign w22940 = w22784 ^ w22939 ;
  assign w22941 = ~w22840 & w22940 ;
  assign w22942 = ( w22706 & w22838 ) | ( w22706 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22943 = ~w22839 & w22942 ;
  assign w22944 = w22941 | w22943 ;
  assign w22945 = ~\pi074 & w22944 ;
  assign w22946 = ~w22719 & w22780 ;
  assign w22947 = w22781 ^ w22946 ;
  assign w22948 = ~w22840 & w22947 ;
  assign w22949 = ( w22712 & w22838 ) | ( w22712 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22950 = ~w22839 & w22949 ;
  assign w22951 = w22948 | w22950 ;
  assign w22952 = ~\pi073 & w22951 ;
  assign w22953 = ~w22725 & w22777 ;
  assign w22954 = w22778 ^ w22953 ;
  assign w22955 = ~w22840 & w22954 ;
  assign w22956 = ( w22718 & w22838 ) | ( w22718 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22957 = ~w22839 & w22956 ;
  assign w22958 = w22955 | w22957 ;
  assign w22959 = ~\pi072 & w22958 ;
  assign w22960 = ~w22731 & w22774 ;
  assign w22961 = w22775 ^ w22960 ;
  assign w22962 = ~w22840 & w22961 ;
  assign w22963 = ( w22724 & w22838 ) | ( w22724 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22964 = ~w22839 & w22963 ;
  assign w22965 = w22962 | w22964 ;
  assign w22966 = ~\pi071 & w22965 ;
  assign w22967 = ~w22737 & w22771 ;
  assign w22968 = w22772 ^ w22967 ;
  assign w22969 = ~w22840 & w22968 ;
  assign w22970 = ( w22730 & w22838 ) | ( w22730 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22971 = ~w22839 & w22970 ;
  assign w22972 = w22969 | w22971 ;
  assign w22973 = ~\pi070 & w22972 ;
  assign w22974 = ~w22743 & w22768 ;
  assign w22975 = w22769 ^ w22974 ;
  assign w22976 = ~w22840 & w22975 ;
  assign w22977 = ( w22736 & w22838 ) | ( w22736 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22978 = ~w22839 & w22977 ;
  assign w22979 = w22976 | w22978 ;
  assign w22980 = ~\pi069 & w22979 ;
  assign w22981 = ~w22750 & w22765 ;
  assign w22982 = w22766 ^ w22981 ;
  assign w22983 = ~w22840 & w22982 ;
  assign w22984 = ( w22742 & w22838 ) | ( w22742 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22985 = ~w22839 & w22984 ;
  assign w22986 = w22983 | w22985 ;
  assign w22987 = ~\pi068 & w22986 ;
  assign w22988 = w22757 & ~w22758 ;
  assign w22989 = w22763 ^ w22988 ;
  assign w22990 = ~w22840 & w22989 ;
  assign w22991 = ( w22749 & w22838 ) | ( w22749 & w22839 ) | ( w22838 & w22839 ) ;
  assign w22992 = ~w22839 & w22991 ;
  assign w22993 = w22990 | w22992 ;
  assign w22994 = ~\pi067 & w22993 ;
  assign w22995 = ( w22752 & w22753 ) | ( w22752 & ~w22840 ) | ( w22753 & ~w22840 ) ;
  assign w22996 = ( ~\pi040 & \pi064 ) | ( ~\pi040 & w22840 ) | ( \pi064 & w22840 ) ;
  assign w22997 = w22995 ^ w22996 ;
  assign w22998 = \pi065 ^ w22997 ;
  assign w22999 = ~w22840 & w22998 ;
  assign w23000 = ( w22754 & w22838 ) | ( w22754 & w22839 ) | ( w22838 & w22839 ) ;
  assign w23001 = ~w22839 & w23000 ;
  assign w23002 = w22999 | w23001 ;
  assign w23003 = ~\pi066 & w23002 ;
  assign w23004 = \pi066 ^ w23002 ;
  assign w23005 = ( \pi064 & ~w22840 ) | ( \pi064 & w23004 ) | ( ~w22840 & w23004 ) ;
  assign w23006 = \pi040 ^ w23005 ;
  assign w23007 = ( \pi065 & w3628 ) | ( \pi065 & ~w23006 ) | ( w3628 & ~w23006 ) ;
  assign w23008 = w23004 | w23007 ;
  assign w23009 = \pi067 ^ w22993 ;
  assign w23010 = ( ~w23003 & w23008 ) | ( ~w23003 & w23009 ) | ( w23008 & w23009 ) ;
  assign w23011 = w23009 | w23010 ;
  assign w23012 = \pi068 ^ w22986 ;
  assign w23013 = ( ~w22994 & w23011 ) | ( ~w22994 & w23012 ) | ( w23011 & w23012 ) ;
  assign w23014 = w23012 | w23013 ;
  assign w23015 = \pi069 ^ w22979 ;
  assign w23016 = ( ~w22987 & w23014 ) | ( ~w22987 & w23015 ) | ( w23014 & w23015 ) ;
  assign w23017 = w23015 | w23016 ;
  assign w23018 = \pi070 ^ w22972 ;
  assign w23019 = ( ~w22980 & w23017 ) | ( ~w22980 & w23018 ) | ( w23017 & w23018 ) ;
  assign w23020 = w23018 | w23019 ;
  assign w23021 = \pi071 ^ w22965 ;
  assign w23022 = ( ~w22973 & w23020 ) | ( ~w22973 & w23021 ) | ( w23020 & w23021 ) ;
  assign w23023 = w23021 | w23022 ;
  assign w23024 = \pi072 ^ w22958 ;
  assign w23025 = ( ~w22966 & w23023 ) | ( ~w22966 & w23024 ) | ( w23023 & w23024 ) ;
  assign w23026 = w23024 | w23025 ;
  assign w23027 = \pi073 ^ w22951 ;
  assign w23028 = ( ~w22959 & w23026 ) | ( ~w22959 & w23027 ) | ( w23026 & w23027 ) ;
  assign w23029 = w23027 | w23028 ;
  assign w23030 = \pi074 ^ w22944 ;
  assign w23031 = ( ~w22952 & w23029 ) | ( ~w22952 & w23030 ) | ( w23029 & w23030 ) ;
  assign w23032 = w23030 | w23031 ;
  assign w23033 = \pi075 ^ w22937 ;
  assign w23034 = ( ~w22945 & w23032 ) | ( ~w22945 & w23033 ) | ( w23032 & w23033 ) ;
  assign w23035 = w23033 | w23034 ;
  assign w23036 = \pi076 ^ w22930 ;
  assign w23037 = ( ~w22938 & w23035 ) | ( ~w22938 & w23036 ) | ( w23035 & w23036 ) ;
  assign w23038 = w23036 | w23037 ;
  assign w23039 = \pi077 ^ w22923 ;
  assign w23040 = ( ~w22931 & w23038 ) | ( ~w22931 & w23039 ) | ( w23038 & w23039 ) ;
  assign w23041 = w23039 | w23040 ;
  assign w23042 = \pi078 ^ w22916 ;
  assign w23043 = ( ~w22924 & w23041 ) | ( ~w22924 & w23042 ) | ( w23041 & w23042 ) ;
  assign w23044 = w23042 | w23043 ;
  assign w23045 = \pi079 ^ w22909 ;
  assign w23046 = ( ~w22917 & w23044 ) | ( ~w22917 & w23045 ) | ( w23044 & w23045 ) ;
  assign w23047 = w23045 | w23046 ;
  assign w23048 = \pi080 ^ w22902 ;
  assign w23049 = ( ~w22910 & w23047 ) | ( ~w22910 & w23048 ) | ( w23047 & w23048 ) ;
  assign w23050 = w23048 | w23049 ;
  assign w23051 = \pi081 ^ w22895 ;
  assign w23052 = ( ~w22903 & w23050 ) | ( ~w22903 & w23051 ) | ( w23050 & w23051 ) ;
  assign w23053 = w23051 | w23052 ;
  assign w23054 = \pi082 ^ w22888 ;
  assign w23055 = ( ~w22896 & w23053 ) | ( ~w22896 & w23054 ) | ( w23053 & w23054 ) ;
  assign w23056 = w23054 | w23055 ;
  assign w23057 = \pi083 ^ w22881 ;
  assign w23058 = ( ~w22889 & w23056 ) | ( ~w22889 & w23057 ) | ( w23056 & w23057 ) ;
  assign w23059 = w23057 | w23058 ;
  assign w23060 = \pi084 ^ w22874 ;
  assign w23061 = ( ~w22882 & w23059 ) | ( ~w22882 & w23060 ) | ( w23059 & w23060 ) ;
  assign w23062 = w23060 | w23061 ;
  assign w23063 = \pi085 ^ w22867 ;
  assign w23064 = ( ~w22875 & w23062 ) | ( ~w22875 & w23063 ) | ( w23062 & w23063 ) ;
  assign w23065 = w23063 | w23064 ;
  assign w23066 = \pi086 ^ w22860 ;
  assign w23067 = ( ~w22868 & w23065 ) | ( ~w22868 & w23066 ) | ( w23065 & w23066 ) ;
  assign w23068 = w23066 | w23067 ;
  assign w23069 = \pi087 ^ w22846 ;
  assign w23070 = ( ~w22861 & w23068 ) | ( ~w22861 & w23069 ) | ( w23068 & w23069 ) ;
  assign w23071 = w23069 | w23070 ;
  assign w23072 = \pi088 ^ w22853 ;
  assign w23073 = w22854 & ~w23072 ;
  assign w23074 = ( w23071 & w23072 ) | ( w23071 & ~w23073 ) | ( w23072 & ~w23073 ) ;
  assign w23075 = ~\pi088 & w22853 ;
  assign w23076 = w23074 & ~w23075 ;
  assign w23077 = w3494 | w23076 ;
  assign w23078 = w22846 & w23077 ;
  assign w23079 = ~w22861 & w23068 ;
  assign w23080 = w23069 ^ w23079 ;
  assign w23081 = ~w23077 & w23080 ;
  assign w23082 = w23078 | w23081 ;
  assign w23083 = w22853 & w23077 ;
  assign w23084 = ~w22854 & w23071 ;
  assign w23085 = w23072 ^ w23084 ;
  assign w23086 = ~w23077 & w23085 ;
  assign w23087 = w23083 | w23086 ;
  assign w23088 = ~\pi088 & w23082 ;
  assign w23089 = w22860 & w23077 ;
  assign w23090 = ~w22868 & w23065 ;
  assign w23091 = w23066 ^ w23090 ;
  assign w23092 = ~w23077 & w23091 ;
  assign w23093 = w23089 | w23092 ;
  assign w23094 = ~\pi087 & w23093 ;
  assign w23095 = w22867 & w23077 ;
  assign w23096 = ~w22875 & w23062 ;
  assign w23097 = w23063 ^ w23096 ;
  assign w23098 = ~w23077 & w23097 ;
  assign w23099 = w23095 | w23098 ;
  assign w23100 = ~\pi086 & w23099 ;
  assign w23101 = w22874 & w23077 ;
  assign w23102 = ~w22882 & w23059 ;
  assign w23103 = w23060 ^ w23102 ;
  assign w23104 = ~w23077 & w23103 ;
  assign w23105 = w23101 | w23104 ;
  assign w23106 = ~\pi085 & w23105 ;
  assign w23107 = w22881 & w23077 ;
  assign w23108 = ~w22889 & w23056 ;
  assign w23109 = w23057 ^ w23108 ;
  assign w23110 = ~w23077 & w23109 ;
  assign w23111 = w23107 | w23110 ;
  assign w23112 = ~\pi084 & w23111 ;
  assign w23113 = w22888 & w23077 ;
  assign w23114 = ~w22896 & w23053 ;
  assign w23115 = w23054 ^ w23114 ;
  assign w23116 = ~w23077 & w23115 ;
  assign w23117 = w23113 | w23116 ;
  assign w23118 = ~\pi083 & w23117 ;
  assign w23119 = w22895 & w23077 ;
  assign w23120 = ~w22903 & w23050 ;
  assign w23121 = w23051 ^ w23120 ;
  assign w23122 = ~w23077 & w23121 ;
  assign w23123 = w23119 | w23122 ;
  assign w23124 = ~\pi082 & w23123 ;
  assign w23125 = w22902 & w23077 ;
  assign w23126 = ~w22910 & w23047 ;
  assign w23127 = w23048 ^ w23126 ;
  assign w23128 = ~w23077 & w23127 ;
  assign w23129 = w23125 | w23128 ;
  assign w23130 = ~\pi081 & w23129 ;
  assign w23131 = w22909 & w23077 ;
  assign w23132 = ~w22917 & w23044 ;
  assign w23133 = w23045 ^ w23132 ;
  assign w23134 = ~w23077 & w23133 ;
  assign w23135 = w23131 | w23134 ;
  assign w23136 = ~\pi080 & w23135 ;
  assign w23137 = w22916 & w23077 ;
  assign w23138 = ~w22924 & w23041 ;
  assign w23139 = w23042 ^ w23138 ;
  assign w23140 = ~w23077 & w23139 ;
  assign w23141 = w23137 | w23140 ;
  assign w23142 = ~\pi079 & w23141 ;
  assign w23143 = w22923 & w23077 ;
  assign w23144 = ~w22931 & w23038 ;
  assign w23145 = w23039 ^ w23144 ;
  assign w23146 = ~w23077 & w23145 ;
  assign w23147 = w23143 | w23146 ;
  assign w23148 = ~\pi078 & w23147 ;
  assign w23149 = w22930 & w23077 ;
  assign w23150 = ~w22938 & w23035 ;
  assign w23151 = w23036 ^ w23150 ;
  assign w23152 = ~w23077 & w23151 ;
  assign w23153 = w23149 | w23152 ;
  assign w23154 = ~\pi077 & w23153 ;
  assign w23155 = w22937 & w23077 ;
  assign w23156 = ~w22945 & w23032 ;
  assign w23157 = w23033 ^ w23156 ;
  assign w23158 = ~w23077 & w23157 ;
  assign w23159 = w23155 | w23158 ;
  assign w23160 = ~\pi076 & w23159 ;
  assign w23161 = w22944 & w23077 ;
  assign w23162 = ~w22952 & w23029 ;
  assign w23163 = w23030 ^ w23162 ;
  assign w23164 = ~w23077 & w23163 ;
  assign w23165 = w23161 | w23164 ;
  assign w23166 = ~\pi075 & w23165 ;
  assign w23167 = w22951 & w23077 ;
  assign w23168 = ~w22959 & w23026 ;
  assign w23169 = w23027 ^ w23168 ;
  assign w23170 = ~w23077 & w23169 ;
  assign w23171 = w23167 | w23170 ;
  assign w23172 = ~\pi074 & w23171 ;
  assign w23173 = w22958 & w23077 ;
  assign w23174 = ~w22966 & w23023 ;
  assign w23175 = w23024 ^ w23174 ;
  assign w23176 = ~w23077 & w23175 ;
  assign w23177 = w23173 | w23176 ;
  assign w23178 = ~\pi073 & w23177 ;
  assign w23179 = w22965 & w23077 ;
  assign w23180 = ~w22973 & w23020 ;
  assign w23181 = w23021 ^ w23180 ;
  assign w23182 = ~w23077 & w23181 ;
  assign w23183 = w23179 | w23182 ;
  assign w23184 = ~\pi072 & w23183 ;
  assign w23185 = w22972 & w23077 ;
  assign w23186 = ~w22980 & w23017 ;
  assign w23187 = w23018 ^ w23186 ;
  assign w23188 = ~w23077 & w23187 ;
  assign w23189 = w23185 | w23188 ;
  assign w23190 = ~\pi071 & w23189 ;
  assign w23191 = w22979 & w23077 ;
  assign w23192 = ~w22987 & w23014 ;
  assign w23193 = w23015 ^ w23192 ;
  assign w23194 = ~w23077 & w23193 ;
  assign w23195 = w23191 | w23194 ;
  assign w23196 = ~\pi070 & w23195 ;
  assign w23197 = w22986 & w23077 ;
  assign w23198 = ~w22994 & w23011 ;
  assign w23199 = w23012 ^ w23198 ;
  assign w23200 = ~w23077 & w23199 ;
  assign w23201 = w23197 | w23200 ;
  assign w23202 = ~\pi069 & w23201 ;
  assign w23203 = w22993 & w23077 ;
  assign w23204 = ~w23003 & w23008 ;
  assign w23205 = w23009 ^ w23204 ;
  assign w23206 = ~w23077 & w23205 ;
  assign w23207 = w23203 | w23206 ;
  assign w23208 = ~\pi068 & w23207 ;
  assign w23209 = w23002 & w23077 ;
  assign w23210 = \pi064 & ~w22840 ;
  assign w23211 = \pi040 ^ w23210 ;
  assign w23212 = ( \pi065 & w3628 ) | ( \pi065 & ~w23211 ) | ( w3628 & ~w23211 ) ;
  assign w23213 = w23004 ^ w23212 ;
  assign w23214 = ( w3494 & w23076 ) | ( w3494 & w23213 ) | ( w23076 & w23213 ) ;
  assign w23215 = w23213 & ~w23214 ;
  assign w23216 = w23209 | w23215 ;
  assign w23217 = ~\pi067 & w23216 ;
  assign w23218 = \pi039 ^ w22840 ;
  assign w23219 = ( \pi064 & w3494 ) | ( \pi064 & w23218 ) | ( w3494 & w23218 ) ;
  assign w23220 = w3635 ^ w23219 ;
  assign w23221 = ~w3494 & w23220 ;
  assign w23222 = ~w23076 & w23221 ;
  assign w23223 = ( ~\pi064 & w22840 ) | ( ~\pi064 & w23077 ) | ( w22840 & w23077 ) ;
  assign w23224 = \pi040 ^ w23223 ;
  assign w23225 = w23077 & ~w23224 ;
  assign w23226 = w23222 | w23225 ;
  assign w23227 = ~\pi066 & w23226 ;
  assign w23228 = ( \pi039 & ~w3651 ) | ( \pi039 & w23076 ) | ( ~w3651 & w23076 ) ;
  assign w23229 = \pi039 & w23228 ;
  assign w23230 = w3657 & ~w23076 ;
  assign w23231 = w23229 | w23230 ;
  assign w23232 = \pi065 ^ w23231 ;
  assign w23233 = w3660 | w23232 ;
  assign w23234 = w23077 | w23222 ;
  assign w23235 = ( w23211 & w23222 ) | ( w23211 & w23234 ) | ( w23222 & w23234 ) ;
  assign w23236 = \pi066 ^ w23235 ;
  assign w23237 = ~\pi065 & w23231 ;
  assign w23238 = w23233 | w23237 ;
  assign w23239 = ( w23236 & ~w23237 ) | ( w23236 & w23238 ) | ( ~w23237 & w23238 ) ;
  assign w23240 = \pi067 ^ w23216 ;
  assign w23241 = ( ~w23227 & w23239 ) | ( ~w23227 & w23240 ) | ( w23239 & w23240 ) ;
  assign w23242 = w23240 | w23241 ;
  assign w23243 = \pi068 ^ w23207 ;
  assign w23244 = ( ~w23217 & w23242 ) | ( ~w23217 & w23243 ) | ( w23242 & w23243 ) ;
  assign w23245 = w23243 | w23244 ;
  assign w23246 = \pi069 ^ w23201 ;
  assign w23247 = ( ~w23208 & w23245 ) | ( ~w23208 & w23246 ) | ( w23245 & w23246 ) ;
  assign w23248 = w23246 | w23247 ;
  assign w23249 = \pi070 ^ w23195 ;
  assign w23250 = ( ~w23202 & w23248 ) | ( ~w23202 & w23249 ) | ( w23248 & w23249 ) ;
  assign w23251 = w23249 | w23250 ;
  assign w23252 = \pi071 ^ w23189 ;
  assign w23253 = ( ~w23196 & w23251 ) | ( ~w23196 & w23252 ) | ( w23251 & w23252 ) ;
  assign w23254 = w23252 | w23253 ;
  assign w23255 = \pi072 ^ w23183 ;
  assign w23256 = ( ~w23190 & w23254 ) | ( ~w23190 & w23255 ) | ( w23254 & w23255 ) ;
  assign w23257 = w23255 | w23256 ;
  assign w23258 = \pi073 ^ w23177 ;
  assign w23259 = ( ~w23184 & w23257 ) | ( ~w23184 & w23258 ) | ( w23257 & w23258 ) ;
  assign w23260 = w23258 | w23259 ;
  assign w23261 = \pi074 ^ w23171 ;
  assign w23262 = ( ~w23178 & w23260 ) | ( ~w23178 & w23261 ) | ( w23260 & w23261 ) ;
  assign w23263 = w23261 | w23262 ;
  assign w23264 = \pi075 ^ w23165 ;
  assign w23265 = ( ~w23172 & w23263 ) | ( ~w23172 & w23264 ) | ( w23263 & w23264 ) ;
  assign w23266 = w23264 | w23265 ;
  assign w23267 = \pi076 ^ w23159 ;
  assign w23268 = ( ~w23166 & w23266 ) | ( ~w23166 & w23267 ) | ( w23266 & w23267 ) ;
  assign w23269 = w23267 | w23268 ;
  assign w23270 = \pi077 ^ w23153 ;
  assign w23271 = ( ~w23160 & w23269 ) | ( ~w23160 & w23270 ) | ( w23269 & w23270 ) ;
  assign w23272 = w23270 | w23271 ;
  assign w23273 = \pi078 ^ w23147 ;
  assign w23274 = ( ~w23154 & w23272 ) | ( ~w23154 & w23273 ) | ( w23272 & w23273 ) ;
  assign w23275 = w23273 | w23274 ;
  assign w23276 = \pi079 ^ w23141 ;
  assign w23277 = ( ~w23148 & w23275 ) | ( ~w23148 & w23276 ) | ( w23275 & w23276 ) ;
  assign w23278 = w23276 | w23277 ;
  assign w23279 = \pi080 ^ w23135 ;
  assign w23280 = ( ~w23142 & w23278 ) | ( ~w23142 & w23279 ) | ( w23278 & w23279 ) ;
  assign w23281 = w23279 | w23280 ;
  assign w23282 = \pi081 ^ w23129 ;
  assign w23283 = ( ~w23136 & w23281 ) | ( ~w23136 & w23282 ) | ( w23281 & w23282 ) ;
  assign w23284 = w23282 | w23283 ;
  assign w23285 = \pi082 ^ w23123 ;
  assign w23286 = ( ~w23130 & w23284 ) | ( ~w23130 & w23285 ) | ( w23284 & w23285 ) ;
  assign w23287 = w23285 | w23286 ;
  assign w23288 = \pi083 ^ w23117 ;
  assign w23289 = ( ~w23124 & w23287 ) | ( ~w23124 & w23288 ) | ( w23287 & w23288 ) ;
  assign w23290 = w23288 | w23289 ;
  assign w23291 = \pi084 ^ w23111 ;
  assign w23292 = ( ~w23118 & w23290 ) | ( ~w23118 & w23291 ) | ( w23290 & w23291 ) ;
  assign w23293 = w23291 | w23292 ;
  assign w23294 = \pi085 ^ w23105 ;
  assign w23295 = ( ~w23112 & w23293 ) | ( ~w23112 & w23294 ) | ( w23293 & w23294 ) ;
  assign w23296 = w23294 | w23295 ;
  assign w23297 = \pi086 ^ w23099 ;
  assign w23298 = ( ~w23106 & w23296 ) | ( ~w23106 & w23297 ) | ( w23296 & w23297 ) ;
  assign w23299 = w23297 | w23298 ;
  assign w23300 = \pi087 ^ w23093 ;
  assign w23301 = ( ~w23100 & w23299 ) | ( ~w23100 & w23300 ) | ( w23299 & w23300 ) ;
  assign w23302 = w23300 | w23301 ;
  assign w23303 = \pi088 ^ w23082 ;
  assign w23304 = ( ~w23094 & w23302 ) | ( ~w23094 & w23303 ) | ( w23302 & w23303 ) ;
  assign w23305 = w23303 | w23304 ;
  assign w23306 = \pi089 ^ w23087 ;
  assign w23307 = w23088 & ~w23306 ;
  assign w23308 = ( w23305 & w23306 ) | ( w23305 & ~w23307 ) | ( w23306 & ~w23307 ) ;
  assign w23309 = ~\pi089 & w23087 ;
  assign w23310 = w23308 & ~w23309 ;
  assign w23311 = w3743 | w23310 ;
  assign w23312 = w23082 & w23311 ;
  assign w23313 = ~w23094 & w23302 ;
  assign w23314 = w23303 ^ w23313 ;
  assign w23315 = ~w23311 & w23314 ;
  assign w23316 = w23312 | w23315 ;
  assign w23317 = ~\pi089 & w23316 ;
  assign w23318 = w23093 & w23311 ;
  assign w23319 = ~w23100 & w23299 ;
  assign w23320 = w23300 ^ w23319 ;
  assign w23321 = ~w23311 & w23320 ;
  assign w23322 = w23318 | w23321 ;
  assign w23323 = ~\pi088 & w23322 ;
  assign w23324 = w23099 & w23311 ;
  assign w23325 = ~w23106 & w23296 ;
  assign w23326 = w23297 ^ w23325 ;
  assign w23327 = ~w23311 & w23326 ;
  assign w23328 = w23324 | w23327 ;
  assign w23329 = ~\pi087 & w23328 ;
  assign w23330 = w23105 & w23311 ;
  assign w23331 = ~w23112 & w23293 ;
  assign w23332 = w23294 ^ w23331 ;
  assign w23333 = ~w23311 & w23332 ;
  assign w23334 = w23330 | w23333 ;
  assign w23335 = ~\pi086 & w23334 ;
  assign w23336 = w23111 & w23311 ;
  assign w23337 = ~w23118 & w23290 ;
  assign w23338 = w23291 ^ w23337 ;
  assign w23339 = ~w23311 & w23338 ;
  assign w23340 = w23336 | w23339 ;
  assign w23341 = ~\pi085 & w23340 ;
  assign w23342 = w23117 & w23311 ;
  assign w23343 = ~w23124 & w23287 ;
  assign w23344 = w23288 ^ w23343 ;
  assign w23345 = ~w23311 & w23344 ;
  assign w23346 = w23342 | w23345 ;
  assign w23347 = ~\pi084 & w23346 ;
  assign w23348 = w23123 & w23311 ;
  assign w23349 = ~w23130 & w23284 ;
  assign w23350 = w23285 ^ w23349 ;
  assign w23351 = ~w23311 & w23350 ;
  assign w23352 = w23348 | w23351 ;
  assign w23353 = ~\pi083 & w23352 ;
  assign w23354 = w23129 & w23311 ;
  assign w23355 = ~w23136 & w23281 ;
  assign w23356 = w23282 ^ w23355 ;
  assign w23357 = ~w23311 & w23356 ;
  assign w23358 = w23354 | w23357 ;
  assign w23359 = ~\pi082 & w23358 ;
  assign w23360 = w23135 & w23311 ;
  assign w23361 = ~w23142 & w23278 ;
  assign w23362 = w23279 ^ w23361 ;
  assign w23363 = ~w23311 & w23362 ;
  assign w23364 = w23360 | w23363 ;
  assign w23365 = ~\pi081 & w23364 ;
  assign w23366 = w23141 & w23311 ;
  assign w23367 = ~w23148 & w23275 ;
  assign w23368 = w23276 ^ w23367 ;
  assign w23369 = ~w23311 & w23368 ;
  assign w23370 = w23366 | w23369 ;
  assign w23371 = ~\pi080 & w23370 ;
  assign w23372 = w23147 & w23311 ;
  assign w23373 = ~w23154 & w23272 ;
  assign w23374 = w23273 ^ w23373 ;
  assign w23375 = ~w23311 & w23374 ;
  assign w23376 = w23372 | w23375 ;
  assign w23377 = ~\pi079 & w23376 ;
  assign w23378 = w23153 & w23311 ;
  assign w23379 = ~w23160 & w23269 ;
  assign w23380 = w23270 ^ w23379 ;
  assign w23381 = ~w23311 & w23380 ;
  assign w23382 = w23378 | w23381 ;
  assign w23383 = ~\pi078 & w23382 ;
  assign w23384 = w23159 & w23311 ;
  assign w23385 = ~w23166 & w23266 ;
  assign w23386 = w23267 ^ w23385 ;
  assign w23387 = ~w23311 & w23386 ;
  assign w23388 = w23384 | w23387 ;
  assign w23389 = ~\pi077 & w23388 ;
  assign w23390 = w23165 & w23311 ;
  assign w23391 = ~w23172 & w23263 ;
  assign w23392 = w23264 ^ w23391 ;
  assign w23393 = ~w23311 & w23392 ;
  assign w23394 = w23390 | w23393 ;
  assign w23395 = ~\pi076 & w23394 ;
  assign w23396 = w23171 & w23311 ;
  assign w23397 = ~w23178 & w23260 ;
  assign w23398 = w23261 ^ w23397 ;
  assign w23399 = ~w23311 & w23398 ;
  assign w23400 = w23396 | w23399 ;
  assign w23401 = ~\pi075 & w23400 ;
  assign w23402 = w23177 & w23311 ;
  assign w23403 = ~w23184 & w23257 ;
  assign w23404 = w23258 ^ w23403 ;
  assign w23405 = ~w23311 & w23404 ;
  assign w23406 = w23402 | w23405 ;
  assign w23407 = ~\pi074 & w23406 ;
  assign w23408 = w23183 & w23311 ;
  assign w23409 = ~w23190 & w23254 ;
  assign w23410 = w23255 ^ w23409 ;
  assign w23411 = ~w23311 & w23410 ;
  assign w23412 = w23408 | w23411 ;
  assign w23413 = ~\pi073 & w23412 ;
  assign w23414 = w23189 & w23311 ;
  assign w23415 = ~w23196 & w23251 ;
  assign w23416 = w23252 ^ w23415 ;
  assign w23417 = ~w23311 & w23416 ;
  assign w23418 = w23414 | w23417 ;
  assign w23419 = ~\pi072 & w23418 ;
  assign w23420 = w23195 & w23311 ;
  assign w23421 = ~w23202 & w23248 ;
  assign w23422 = w23249 ^ w23421 ;
  assign w23423 = ~w23311 & w23422 ;
  assign w23424 = w23420 | w23423 ;
  assign w23425 = ~\pi071 & w23424 ;
  assign w23426 = w23201 & w23311 ;
  assign w23427 = ~w23208 & w23245 ;
  assign w23428 = w23246 ^ w23427 ;
  assign w23429 = ~w23311 & w23428 ;
  assign w23430 = w23426 | w23429 ;
  assign w23431 = ~\pi070 & w23430 ;
  assign w23432 = w23207 & w23311 ;
  assign w23433 = ~w23217 & w23242 ;
  assign w23434 = w23243 ^ w23433 ;
  assign w23435 = ~w23311 & w23434 ;
  assign w23436 = w23432 | w23435 ;
  assign w23437 = ~\pi069 & w23436 ;
  assign w23438 = w23216 & w23311 ;
  assign w23439 = ~w23227 & w23239 ;
  assign w23440 = w23240 ^ w23439 ;
  assign w23441 = ~w23311 & w23440 ;
  assign w23442 = w23438 | w23441 ;
  assign w23443 = ~\pi068 & w23442 ;
  assign w23444 = w23226 & w23311 ;
  assign w23445 = ~w23231 & w23233 ;
  assign w23446 = ( \pi065 & w23233 ) | ( \pi065 & w23445 ) | ( w23233 & w23445 ) ;
  assign w23447 = w23236 ^ w23446 ;
  assign w23448 = ~w23311 & w23447 ;
  assign w23449 = w23444 | w23448 ;
  assign w23450 = ~\pi067 & w23449 ;
  assign w23451 = w23231 & w23311 ;
  assign w23452 = ( ~w3743 & w23229 ) | ( ~w3743 & w23230 ) | ( w23229 & w23230 ) ;
  assign w23453 = \pi065 ^ w23452 ;
  assign w23454 = ( w3660 & ~w3743 ) | ( w3660 & w23453 ) | ( ~w3743 & w23453 ) ;
  assign w23455 = ( w3660 & w23310 ) | ( w3660 & w23453 ) | ( w23310 & w23453 ) ;
  assign w23456 = w23454 & ~w23455 ;
  assign w23457 = w23451 | w23456 ;
  assign w23458 = ~\pi066 & w23457 ;
  assign w23459 = ( \pi038 & ~w3897 ) | ( \pi038 & w23310 ) | ( ~w3897 & w23310 ) ;
  assign w23460 = \pi038 & w23459 ;
  assign w23461 = w3903 & ~w23310 ;
  assign w23462 = w23460 | w23461 ;
  assign w23463 = \pi065 ^ w23462 ;
  assign w23464 = w3906 | w23463 ;
  assign w23465 = \pi066 ^ w23457 ;
  assign w23466 = ~\pi065 & w23462 ;
  assign w23467 = w23464 | w23466 ;
  assign w23468 = ( w23465 & ~w23466 ) | ( w23465 & w23467 ) | ( ~w23466 & w23467 ) ;
  assign w23469 = \pi067 ^ w23449 ;
  assign w23470 = ( ~w23458 & w23468 ) | ( ~w23458 & w23469 ) | ( w23468 & w23469 ) ;
  assign w23471 = w23469 | w23470 ;
  assign w23472 = \pi068 ^ w23442 ;
  assign w23473 = ( ~w23450 & w23471 ) | ( ~w23450 & w23472 ) | ( w23471 & w23472 ) ;
  assign w23474 = w23472 | w23473 ;
  assign w23475 = \pi069 ^ w23436 ;
  assign w23476 = ( ~w23443 & w23474 ) | ( ~w23443 & w23475 ) | ( w23474 & w23475 ) ;
  assign w23477 = w23475 | w23476 ;
  assign w23478 = \pi070 ^ w23430 ;
  assign w23479 = ( ~w23437 & w23477 ) | ( ~w23437 & w23478 ) | ( w23477 & w23478 ) ;
  assign w23480 = w23478 | w23479 ;
  assign w23481 = \pi071 ^ w23424 ;
  assign w23482 = ( ~w23431 & w23480 ) | ( ~w23431 & w23481 ) | ( w23480 & w23481 ) ;
  assign w23483 = w23481 | w23482 ;
  assign w23484 = \pi072 ^ w23418 ;
  assign w23485 = ( ~w23425 & w23483 ) | ( ~w23425 & w23484 ) | ( w23483 & w23484 ) ;
  assign w23486 = w23484 | w23485 ;
  assign w23487 = \pi073 ^ w23412 ;
  assign w23488 = ( ~w23419 & w23486 ) | ( ~w23419 & w23487 ) | ( w23486 & w23487 ) ;
  assign w23489 = w23487 | w23488 ;
  assign w23490 = \pi074 ^ w23406 ;
  assign w23491 = ( ~w23413 & w23489 ) | ( ~w23413 & w23490 ) | ( w23489 & w23490 ) ;
  assign w23492 = w23490 | w23491 ;
  assign w23493 = \pi075 ^ w23400 ;
  assign w23494 = ( ~w23407 & w23492 ) | ( ~w23407 & w23493 ) | ( w23492 & w23493 ) ;
  assign w23495 = w23493 | w23494 ;
  assign w23496 = \pi076 ^ w23394 ;
  assign w23497 = ( ~w23401 & w23495 ) | ( ~w23401 & w23496 ) | ( w23495 & w23496 ) ;
  assign w23498 = w23496 | w23497 ;
  assign w23499 = \pi077 ^ w23388 ;
  assign w23500 = ( ~w23395 & w23498 ) | ( ~w23395 & w23499 ) | ( w23498 & w23499 ) ;
  assign w23501 = w23499 | w23500 ;
  assign w23502 = \pi078 ^ w23382 ;
  assign w23503 = ( ~w23389 & w23501 ) | ( ~w23389 & w23502 ) | ( w23501 & w23502 ) ;
  assign w23504 = w23502 | w23503 ;
  assign w23505 = \pi079 ^ w23376 ;
  assign w23506 = ( ~w23383 & w23504 ) | ( ~w23383 & w23505 ) | ( w23504 & w23505 ) ;
  assign w23507 = w23505 | w23506 ;
  assign w23508 = \pi080 ^ w23370 ;
  assign w23509 = ( ~w23377 & w23507 ) | ( ~w23377 & w23508 ) | ( w23507 & w23508 ) ;
  assign w23510 = w23508 | w23509 ;
  assign w23511 = \pi081 ^ w23364 ;
  assign w23512 = ( ~w23371 & w23510 ) | ( ~w23371 & w23511 ) | ( w23510 & w23511 ) ;
  assign w23513 = w23511 | w23512 ;
  assign w23514 = \pi082 ^ w23358 ;
  assign w23515 = ( ~w23365 & w23513 ) | ( ~w23365 & w23514 ) | ( w23513 & w23514 ) ;
  assign w23516 = w23514 | w23515 ;
  assign w23517 = \pi083 ^ w23352 ;
  assign w23518 = ( ~w23359 & w23516 ) | ( ~w23359 & w23517 ) | ( w23516 & w23517 ) ;
  assign w23519 = w23517 | w23518 ;
  assign w23520 = \pi084 ^ w23346 ;
  assign w23521 = ( ~w23353 & w23519 ) | ( ~w23353 & w23520 ) | ( w23519 & w23520 ) ;
  assign w23522 = w23520 | w23521 ;
  assign w23523 = \pi085 ^ w23340 ;
  assign w23524 = ( ~w23347 & w23522 ) | ( ~w23347 & w23523 ) | ( w23522 & w23523 ) ;
  assign w23525 = w23523 | w23524 ;
  assign w23526 = \pi086 ^ w23334 ;
  assign w23527 = ( ~w23341 & w23525 ) | ( ~w23341 & w23526 ) | ( w23525 & w23526 ) ;
  assign w23528 = w23526 | w23527 ;
  assign w23529 = \pi087 ^ w23328 ;
  assign w23530 = ( ~w23335 & w23528 ) | ( ~w23335 & w23529 ) | ( w23528 & w23529 ) ;
  assign w23531 = w23529 | w23530 ;
  assign w23532 = \pi088 ^ w23322 ;
  assign w23533 = ( ~w23329 & w23531 ) | ( ~w23329 & w23532 ) | ( w23531 & w23532 ) ;
  assign w23534 = w23532 | w23533 ;
  assign w23535 = \pi089 ^ w23316 ;
  assign w23536 = ( ~w23323 & w23534 ) | ( ~w23323 & w23535 ) | ( w23534 & w23535 ) ;
  assign w23537 = w23535 | w23536 ;
  assign w23538 = w23087 & w23311 ;
  assign w23539 = ~w23088 & w23305 ;
  assign w23540 = w23306 ^ w23539 ;
  assign w23541 = ~w23311 & w23540 ;
  assign w23542 = w23538 | w23541 ;
  assign w23543 = ~\pi090 & w23542 ;
  assign w23544 = ( \pi090 & ~w23538 ) | ( \pi090 & w23541 ) | ( ~w23538 & w23541 ) ;
  assign w23545 = ~w23541 & w23544 ;
  assign w23546 = w23543 | w23545 ;
  assign w23547 = ( ~w23317 & w23537 ) | ( ~w23317 & w23546 ) | ( w23537 & w23546 ) ;
  assign w23548 = ( w3993 & ~w23546 ) | ( w3993 & w23547 ) | ( ~w23546 & w23547 ) ;
  assign w23549 = w23546 | w23548 ;
  assign w23550 = ~w3743 & w23542 ;
  assign w23551 = w23549 & ~w23550 ;
  assign w23552 = ~w23323 & w23534 ;
  assign w23553 = w23535 ^ w23552 ;
  assign w23554 = ~w23551 & w23553 ;
  assign w23555 = ( w23316 & w23549 ) | ( w23316 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23556 = ~w23550 & w23555 ;
  assign w23557 = w23554 | w23556 ;
  assign w23558 = ( ~w23317 & w23537 ) | ( ~w23317 & w23551 ) | ( w23537 & w23551 ) ;
  assign w23559 = w23546 ^ w23558 ;
  assign w23560 = ~w23551 & w23559 ;
  assign w23561 = ( w3743 & ~w23542 ) | ( w3743 & w23549 ) | ( ~w23542 & w23549 ) ;
  assign w23562 = w23542 & w23561 ;
  assign w23563 = w23560 | w23562 ;
  assign w23564 = ~\pi090 & w23557 ;
  assign w23565 = ~w23329 & w23531 ;
  assign w23566 = w23532 ^ w23565 ;
  assign w23567 = ~w23551 & w23566 ;
  assign w23568 = ( w23322 & w23549 ) | ( w23322 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23569 = ~w23550 & w23568 ;
  assign w23570 = w23567 | w23569 ;
  assign w23571 = ~\pi089 & w23570 ;
  assign w23572 = ~w23335 & w23528 ;
  assign w23573 = w23529 ^ w23572 ;
  assign w23574 = ~w23551 & w23573 ;
  assign w23575 = ( w23328 & w23549 ) | ( w23328 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23576 = ~w23550 & w23575 ;
  assign w23577 = w23574 | w23576 ;
  assign w23578 = ~\pi088 & w23577 ;
  assign w23579 = ~w23341 & w23525 ;
  assign w23580 = w23526 ^ w23579 ;
  assign w23581 = ~w23551 & w23580 ;
  assign w23582 = ( w23334 & w23549 ) | ( w23334 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23583 = ~w23550 & w23582 ;
  assign w23584 = w23581 | w23583 ;
  assign w23585 = ~\pi087 & w23584 ;
  assign w23586 = ~w23347 & w23522 ;
  assign w23587 = w23523 ^ w23586 ;
  assign w23588 = ~w23551 & w23587 ;
  assign w23589 = ( w23340 & w23549 ) | ( w23340 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23590 = ~w23550 & w23589 ;
  assign w23591 = w23588 | w23590 ;
  assign w23592 = ~\pi086 & w23591 ;
  assign w23593 = ~w23353 & w23519 ;
  assign w23594 = w23520 ^ w23593 ;
  assign w23595 = ~w23551 & w23594 ;
  assign w23596 = ( w23346 & w23549 ) | ( w23346 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23597 = ~w23550 & w23596 ;
  assign w23598 = w23595 | w23597 ;
  assign w23599 = ~\pi085 & w23598 ;
  assign w23600 = ~w23359 & w23516 ;
  assign w23601 = w23517 ^ w23600 ;
  assign w23602 = ~w23551 & w23601 ;
  assign w23603 = ( w23352 & w23549 ) | ( w23352 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23604 = ~w23550 & w23603 ;
  assign w23605 = w23602 | w23604 ;
  assign w23606 = ~\pi084 & w23605 ;
  assign w23607 = ~w23365 & w23513 ;
  assign w23608 = w23514 ^ w23607 ;
  assign w23609 = ~w23551 & w23608 ;
  assign w23610 = ( w23358 & w23549 ) | ( w23358 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23611 = ~w23550 & w23610 ;
  assign w23612 = w23609 | w23611 ;
  assign w23613 = ~\pi083 & w23612 ;
  assign w23614 = ~w23371 & w23510 ;
  assign w23615 = w23511 ^ w23614 ;
  assign w23616 = ~w23551 & w23615 ;
  assign w23617 = ( w23364 & w23549 ) | ( w23364 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23618 = ~w23550 & w23617 ;
  assign w23619 = w23616 | w23618 ;
  assign w23620 = ~\pi082 & w23619 ;
  assign w23621 = ~w23377 & w23507 ;
  assign w23622 = w23508 ^ w23621 ;
  assign w23623 = ~w23551 & w23622 ;
  assign w23624 = ( w23370 & w23549 ) | ( w23370 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23625 = ~w23550 & w23624 ;
  assign w23626 = w23623 | w23625 ;
  assign w23627 = ~\pi081 & w23626 ;
  assign w23628 = ~w23383 & w23504 ;
  assign w23629 = w23505 ^ w23628 ;
  assign w23630 = ~w23551 & w23629 ;
  assign w23631 = ( w23376 & w23549 ) | ( w23376 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23632 = ~w23550 & w23631 ;
  assign w23633 = w23630 | w23632 ;
  assign w23634 = ~\pi080 & w23633 ;
  assign w23635 = ~w23389 & w23501 ;
  assign w23636 = w23502 ^ w23635 ;
  assign w23637 = ~w23551 & w23636 ;
  assign w23638 = ( w23382 & w23549 ) | ( w23382 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23639 = ~w23550 & w23638 ;
  assign w23640 = w23637 | w23639 ;
  assign w23641 = ~\pi079 & w23640 ;
  assign w23642 = ~w23395 & w23498 ;
  assign w23643 = w23499 ^ w23642 ;
  assign w23644 = ~w23551 & w23643 ;
  assign w23645 = ( w23388 & w23549 ) | ( w23388 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23646 = ~w23550 & w23645 ;
  assign w23647 = w23644 | w23646 ;
  assign w23648 = ~\pi078 & w23647 ;
  assign w23649 = ~w23401 & w23495 ;
  assign w23650 = w23496 ^ w23649 ;
  assign w23651 = ~w23551 & w23650 ;
  assign w23652 = ( w23394 & w23549 ) | ( w23394 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23653 = ~w23550 & w23652 ;
  assign w23654 = w23651 | w23653 ;
  assign w23655 = ~\pi077 & w23654 ;
  assign w23656 = ~w23407 & w23492 ;
  assign w23657 = w23493 ^ w23656 ;
  assign w23658 = ~w23551 & w23657 ;
  assign w23659 = ( w23400 & w23549 ) | ( w23400 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23660 = ~w23550 & w23659 ;
  assign w23661 = w23658 | w23660 ;
  assign w23662 = ~\pi076 & w23661 ;
  assign w23663 = ~w23413 & w23489 ;
  assign w23664 = w23490 ^ w23663 ;
  assign w23665 = ~w23551 & w23664 ;
  assign w23666 = ( w23406 & w23549 ) | ( w23406 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23667 = ~w23550 & w23666 ;
  assign w23668 = w23665 | w23667 ;
  assign w23669 = ~\pi075 & w23668 ;
  assign w23670 = ~w23419 & w23486 ;
  assign w23671 = w23487 ^ w23670 ;
  assign w23672 = ~w23551 & w23671 ;
  assign w23673 = ( w23412 & w23549 ) | ( w23412 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23674 = ~w23550 & w23673 ;
  assign w23675 = w23672 | w23674 ;
  assign w23676 = ~\pi074 & w23675 ;
  assign w23677 = ~w23425 & w23483 ;
  assign w23678 = w23484 ^ w23677 ;
  assign w23679 = ~w23551 & w23678 ;
  assign w23680 = ( w23418 & w23549 ) | ( w23418 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23681 = ~w23550 & w23680 ;
  assign w23682 = w23679 | w23681 ;
  assign w23683 = ~\pi073 & w23682 ;
  assign w23684 = ~w23431 & w23480 ;
  assign w23685 = w23481 ^ w23684 ;
  assign w23686 = ~w23551 & w23685 ;
  assign w23687 = ( w23424 & w23549 ) | ( w23424 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23688 = ~w23550 & w23687 ;
  assign w23689 = w23686 | w23688 ;
  assign w23690 = ~\pi072 & w23689 ;
  assign w23691 = ~w23437 & w23477 ;
  assign w23692 = w23478 ^ w23691 ;
  assign w23693 = ~w23551 & w23692 ;
  assign w23694 = ( w23430 & w23549 ) | ( w23430 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23695 = ~w23550 & w23694 ;
  assign w23696 = w23693 | w23695 ;
  assign w23697 = ~\pi071 & w23696 ;
  assign w23698 = ~w23443 & w23474 ;
  assign w23699 = w23475 ^ w23698 ;
  assign w23700 = ~w23551 & w23699 ;
  assign w23701 = ( w23436 & w23549 ) | ( w23436 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23702 = ~w23550 & w23701 ;
  assign w23703 = w23700 | w23702 ;
  assign w23704 = ~\pi070 & w23703 ;
  assign w23705 = ~w23450 & w23471 ;
  assign w23706 = w23472 ^ w23705 ;
  assign w23707 = ~w23551 & w23706 ;
  assign w23708 = ( w23442 & w23549 ) | ( w23442 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23709 = ~w23550 & w23708 ;
  assign w23710 = w23707 | w23709 ;
  assign w23711 = ~\pi069 & w23710 ;
  assign w23712 = ~w23458 & w23468 ;
  assign w23713 = w23469 ^ w23712 ;
  assign w23714 = ~w23551 & w23713 ;
  assign w23715 = ( w23449 & w23549 ) | ( w23449 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23716 = ~w23550 & w23715 ;
  assign w23717 = w23714 | w23716 ;
  assign w23718 = ~\pi068 & w23717 ;
  assign w23719 = ( \pi065 & w23462 ) | ( \pi065 & ~w23551 ) | ( w23462 & ~w23551 ) ;
  assign w23720 = ( \pi065 & w23464 ) | ( \pi065 & ~w23719 ) | ( w23464 & ~w23719 ) ;
  assign w23721 = w23465 ^ w23720 ;
  assign w23722 = ~w23551 & w23721 ;
  assign w23723 = ( w23457 & w23549 ) | ( w23457 & w23550 ) | ( w23549 & w23550 ) ;
  assign w23724 = ~w23550 & w23723 ;
  assign w23725 = w23722 | w23724 ;
  assign w23726 = ~\pi067 & w23725 ;
  assign w23727 = w3906 ^ w23462 ;
  assign w23728 = \pi065 ^ w23727 ;
  assign w23729 = w23551 ^ w23728 ;
  assign w23730 = ( w23462 & w23728 ) | ( w23462 & w23729 ) | ( w23728 & w23729 ) ;
  assign w23731 = ~\pi066 & w23730 ;
  assign w23732 = w23462 ^ w23551 ;
  assign w23733 = ( w23462 & w23728 ) | ( w23462 & ~w23732 ) | ( w23728 & ~w23732 ) ;
  assign w23734 = \pi066 ^ w23733 ;
  assign w23735 = ( \pi064 & ~w23551 ) | ( \pi064 & w23734 ) | ( ~w23551 & w23734 ) ;
  assign w23736 = \pi037 ^ w23735 ;
  assign w23737 = ( \pi065 & w4418 ) | ( \pi065 & ~w23736 ) | ( w4418 & ~w23736 ) ;
  assign w23738 = w23734 | w23737 ;
  assign w23739 = \pi067 ^ w23725 ;
  assign w23740 = ( ~w23731 & w23738 ) | ( ~w23731 & w23739 ) | ( w23738 & w23739 ) ;
  assign w23741 = w23739 | w23740 ;
  assign w23742 = \pi068 ^ w23717 ;
  assign w23743 = ( ~w23726 & w23741 ) | ( ~w23726 & w23742 ) | ( w23741 & w23742 ) ;
  assign w23744 = w23742 | w23743 ;
  assign w23745 = \pi069 ^ w23710 ;
  assign w23746 = ( ~w23718 & w23744 ) | ( ~w23718 & w23745 ) | ( w23744 & w23745 ) ;
  assign w23747 = w23745 | w23746 ;
  assign w23748 = \pi070 ^ w23703 ;
  assign w23749 = ( ~w23711 & w23747 ) | ( ~w23711 & w23748 ) | ( w23747 & w23748 ) ;
  assign w23750 = w23748 | w23749 ;
  assign w23751 = \pi071 ^ w23696 ;
  assign w23752 = ( ~w23704 & w23750 ) | ( ~w23704 & w23751 ) | ( w23750 & w23751 ) ;
  assign w23753 = w23751 | w23752 ;
  assign w23754 = \pi072 ^ w23689 ;
  assign w23755 = ( ~w23697 & w23753 ) | ( ~w23697 & w23754 ) | ( w23753 & w23754 ) ;
  assign w23756 = w23754 | w23755 ;
  assign w23757 = \pi073 ^ w23682 ;
  assign w23758 = ( ~w23690 & w23756 ) | ( ~w23690 & w23757 ) | ( w23756 & w23757 ) ;
  assign w23759 = w23757 | w23758 ;
  assign w23760 = \pi074 ^ w23675 ;
  assign w23761 = ( ~w23683 & w23759 ) | ( ~w23683 & w23760 ) | ( w23759 & w23760 ) ;
  assign w23762 = w23760 | w23761 ;
  assign w23763 = \pi075 ^ w23668 ;
  assign w23764 = ( ~w23676 & w23762 ) | ( ~w23676 & w23763 ) | ( w23762 & w23763 ) ;
  assign w23765 = w23763 | w23764 ;
  assign w23766 = \pi076 ^ w23661 ;
  assign w23767 = ( ~w23669 & w23765 ) | ( ~w23669 & w23766 ) | ( w23765 & w23766 ) ;
  assign w23768 = w23766 | w23767 ;
  assign w23769 = \pi077 ^ w23654 ;
  assign w23770 = ( ~w23662 & w23768 ) | ( ~w23662 & w23769 ) | ( w23768 & w23769 ) ;
  assign w23771 = w23769 | w23770 ;
  assign w23772 = \pi078 ^ w23647 ;
  assign w23773 = ( ~w23655 & w23771 ) | ( ~w23655 & w23772 ) | ( w23771 & w23772 ) ;
  assign w23774 = w23772 | w23773 ;
  assign w23775 = \pi079 ^ w23640 ;
  assign w23776 = ( ~w23648 & w23774 ) | ( ~w23648 & w23775 ) | ( w23774 & w23775 ) ;
  assign w23777 = w23775 | w23776 ;
  assign w23778 = \pi080 ^ w23633 ;
  assign w23779 = ( ~w23641 & w23777 ) | ( ~w23641 & w23778 ) | ( w23777 & w23778 ) ;
  assign w23780 = w23778 | w23779 ;
  assign w23781 = \pi081 ^ w23626 ;
  assign w23782 = ( ~w23634 & w23780 ) | ( ~w23634 & w23781 ) | ( w23780 & w23781 ) ;
  assign w23783 = w23781 | w23782 ;
  assign w23784 = \pi082 ^ w23619 ;
  assign w23785 = ( ~w23627 & w23783 ) | ( ~w23627 & w23784 ) | ( w23783 & w23784 ) ;
  assign w23786 = w23784 | w23785 ;
  assign w23787 = \pi083 ^ w23612 ;
  assign w23788 = ( ~w23620 & w23786 ) | ( ~w23620 & w23787 ) | ( w23786 & w23787 ) ;
  assign w23789 = w23787 | w23788 ;
  assign w23790 = \pi084 ^ w23605 ;
  assign w23791 = ( ~w23613 & w23789 ) | ( ~w23613 & w23790 ) | ( w23789 & w23790 ) ;
  assign w23792 = w23790 | w23791 ;
  assign w23793 = \pi085 ^ w23598 ;
  assign w23794 = ( ~w23606 & w23792 ) | ( ~w23606 & w23793 ) | ( w23792 & w23793 ) ;
  assign w23795 = w23793 | w23794 ;
  assign w23796 = \pi086 ^ w23591 ;
  assign w23797 = ( ~w23599 & w23795 ) | ( ~w23599 & w23796 ) | ( w23795 & w23796 ) ;
  assign w23798 = w23796 | w23797 ;
  assign w23799 = \pi087 ^ w23584 ;
  assign w23800 = ( ~w23592 & w23798 ) | ( ~w23592 & w23799 ) | ( w23798 & w23799 ) ;
  assign w23801 = w23799 | w23800 ;
  assign w23802 = \pi088 ^ w23577 ;
  assign w23803 = ( ~w23585 & w23801 ) | ( ~w23585 & w23802 ) | ( w23801 & w23802 ) ;
  assign w23804 = w23802 | w23803 ;
  assign w23805 = \pi089 ^ w23570 ;
  assign w23806 = ( ~w23578 & w23804 ) | ( ~w23578 & w23805 ) | ( w23804 & w23805 ) ;
  assign w23807 = w23805 | w23806 ;
  assign w23808 = \pi090 ^ w23557 ;
  assign w23809 = ( ~w23571 & w23807 ) | ( ~w23571 & w23808 ) | ( w23807 & w23808 ) ;
  assign w23810 = w23808 | w23809 ;
  assign w23811 = \pi091 ^ w23563 ;
  assign w23812 = w23564 & ~w23811 ;
  assign w23813 = ( w23810 & w23811 ) | ( w23810 & ~w23812 ) | ( w23811 & ~w23812 ) ;
  assign w23814 = ~\pi091 & w23563 ;
  assign w23815 = w23813 & ~w23814 ;
  assign w23816 = w4266 | w23815 ;
  assign w23817 = w23557 & w23816 ;
  assign w23818 = ~w23571 & w23807 ;
  assign w23819 = w23808 ^ w23818 ;
  assign w23820 = ~w23816 & w23819 ;
  assign w23821 = w23817 | w23820 ;
  assign w23822 = w23563 & w23816 ;
  assign w23823 = ~w23564 & w23810 ;
  assign w23824 = w23811 ^ w23823 ;
  assign w23825 = ~w23816 & w23824 ;
  assign w23826 = w23822 | w23825 ;
  assign w23827 = ~\pi091 & w23821 ;
  assign w23828 = w23570 & w23816 ;
  assign w23829 = ~w23578 & w23804 ;
  assign w23830 = w23805 ^ w23829 ;
  assign w23831 = ~w23816 & w23830 ;
  assign w23832 = w23828 | w23831 ;
  assign w23833 = ~\pi090 & w23832 ;
  assign w23834 = w23577 & w23816 ;
  assign w23835 = ~w23585 & w23801 ;
  assign w23836 = w23802 ^ w23835 ;
  assign w23837 = ~w23816 & w23836 ;
  assign w23838 = w23834 | w23837 ;
  assign w23839 = ~\pi089 & w23838 ;
  assign w23840 = w23584 & w23816 ;
  assign w23841 = ~w23592 & w23798 ;
  assign w23842 = w23799 ^ w23841 ;
  assign w23843 = ~w23816 & w23842 ;
  assign w23844 = w23840 | w23843 ;
  assign w23845 = ~\pi088 & w23844 ;
  assign w23846 = w23591 & w23816 ;
  assign w23847 = ~w23599 & w23795 ;
  assign w23848 = w23796 ^ w23847 ;
  assign w23849 = ~w23816 & w23848 ;
  assign w23850 = w23846 | w23849 ;
  assign w23851 = ~\pi087 & w23850 ;
  assign w23852 = w23598 & w23816 ;
  assign w23853 = ~w23606 & w23792 ;
  assign w23854 = w23793 ^ w23853 ;
  assign w23855 = ~w23816 & w23854 ;
  assign w23856 = w23852 | w23855 ;
  assign w23857 = ~\pi086 & w23856 ;
  assign w23858 = w23605 & w23816 ;
  assign w23859 = ~w23613 & w23789 ;
  assign w23860 = w23790 ^ w23859 ;
  assign w23861 = ~w23816 & w23860 ;
  assign w23862 = w23858 | w23861 ;
  assign w23863 = ~\pi085 & w23862 ;
  assign w23864 = w23612 & w23816 ;
  assign w23865 = ~w23620 & w23786 ;
  assign w23866 = w23787 ^ w23865 ;
  assign w23867 = ~w23816 & w23866 ;
  assign w23868 = w23864 | w23867 ;
  assign w23869 = ~\pi084 & w23868 ;
  assign w23870 = w23619 & w23816 ;
  assign w23871 = ~w23627 & w23783 ;
  assign w23872 = w23784 ^ w23871 ;
  assign w23873 = ~w23816 & w23872 ;
  assign w23874 = w23870 | w23873 ;
  assign w23875 = ~\pi083 & w23874 ;
  assign w23876 = w23626 & w23816 ;
  assign w23877 = ~w23634 & w23780 ;
  assign w23878 = w23781 ^ w23877 ;
  assign w23879 = ~w23816 & w23878 ;
  assign w23880 = w23876 | w23879 ;
  assign w23881 = ~\pi082 & w23880 ;
  assign w23882 = w23633 & w23816 ;
  assign w23883 = ~w23641 & w23777 ;
  assign w23884 = w23778 ^ w23883 ;
  assign w23885 = ~w23816 & w23884 ;
  assign w23886 = w23882 | w23885 ;
  assign w23887 = ~\pi081 & w23886 ;
  assign w23888 = w23640 & w23816 ;
  assign w23889 = ~w23648 & w23774 ;
  assign w23890 = w23775 ^ w23889 ;
  assign w23891 = ~w23816 & w23890 ;
  assign w23892 = w23888 | w23891 ;
  assign w23893 = ~\pi080 & w23892 ;
  assign w23894 = w23647 & w23816 ;
  assign w23895 = ~w23655 & w23771 ;
  assign w23896 = w23772 ^ w23895 ;
  assign w23897 = ~w23816 & w23896 ;
  assign w23898 = w23894 | w23897 ;
  assign w23899 = ~\pi079 & w23898 ;
  assign w23900 = w23654 & w23816 ;
  assign w23901 = ~w23662 & w23768 ;
  assign w23902 = w23769 ^ w23901 ;
  assign w23903 = ~w23816 & w23902 ;
  assign w23904 = w23900 | w23903 ;
  assign w23905 = ~\pi078 & w23904 ;
  assign w23906 = w23661 & w23816 ;
  assign w23907 = ~w23669 & w23765 ;
  assign w23908 = w23766 ^ w23907 ;
  assign w23909 = ~w23816 & w23908 ;
  assign w23910 = w23906 | w23909 ;
  assign w23911 = ~\pi077 & w23910 ;
  assign w23912 = w23668 & w23816 ;
  assign w23913 = ~w23676 & w23762 ;
  assign w23914 = w23763 ^ w23913 ;
  assign w23915 = ~w23816 & w23914 ;
  assign w23916 = w23912 | w23915 ;
  assign w23917 = ~\pi076 & w23916 ;
  assign w23918 = w23675 & w23816 ;
  assign w23919 = ~w23683 & w23759 ;
  assign w23920 = w23760 ^ w23919 ;
  assign w23921 = ~w23816 & w23920 ;
  assign w23922 = w23918 | w23921 ;
  assign w23923 = ~\pi075 & w23922 ;
  assign w23924 = w23682 & w23816 ;
  assign w23925 = ~w23690 & w23756 ;
  assign w23926 = w23757 ^ w23925 ;
  assign w23927 = ~w23816 & w23926 ;
  assign w23928 = w23924 | w23927 ;
  assign w23929 = ~\pi074 & w23928 ;
  assign w23930 = w23689 & w23816 ;
  assign w23931 = ~w23697 & w23753 ;
  assign w23932 = w23754 ^ w23931 ;
  assign w23933 = ~w23816 & w23932 ;
  assign w23934 = w23930 | w23933 ;
  assign w23935 = ~\pi073 & w23934 ;
  assign w23936 = w23696 & w23816 ;
  assign w23937 = ~w23704 & w23750 ;
  assign w23938 = w23751 ^ w23937 ;
  assign w23939 = ~w23816 & w23938 ;
  assign w23940 = w23936 | w23939 ;
  assign w23941 = ~\pi072 & w23940 ;
  assign w23942 = w23703 & w23816 ;
  assign w23943 = ~w23711 & w23747 ;
  assign w23944 = w23748 ^ w23943 ;
  assign w23945 = ~w23816 & w23944 ;
  assign w23946 = w23942 | w23945 ;
  assign w23947 = ~\pi071 & w23946 ;
  assign w23948 = w23710 & w23816 ;
  assign w23949 = ~w23718 & w23744 ;
  assign w23950 = w23745 ^ w23949 ;
  assign w23951 = ~w23816 & w23950 ;
  assign w23952 = w23948 | w23951 ;
  assign w23953 = ~\pi070 & w23952 ;
  assign w23954 = w23717 & w23816 ;
  assign w23955 = ~w23726 & w23741 ;
  assign w23956 = w23742 ^ w23955 ;
  assign w23957 = ~w23816 & w23956 ;
  assign w23958 = w23954 | w23957 ;
  assign w23959 = ~\pi069 & w23958 ;
  assign w23960 = w23725 & w23816 ;
  assign w23961 = ~w23731 & w23738 ;
  assign w23962 = w23739 ^ w23961 ;
  assign w23963 = ~w23816 & w23962 ;
  assign w23964 = w23960 | w23963 ;
  assign w23965 = ~\pi068 & w23964 ;
  assign w23966 = w23730 & w23816 ;
  assign w23967 = \pi064 & ~w23551 ;
  assign w23968 = \pi037 ^ w23967 ;
  assign w23969 = ( \pi065 & w4418 ) | ( \pi065 & ~w23968 ) | ( w4418 & ~w23968 ) ;
  assign w23970 = w23734 ^ w23969 ;
  assign w23971 = ( w4266 & w23815 ) | ( w4266 & w23970 ) | ( w23815 & w23970 ) ;
  assign w23972 = w23970 & ~w23971 ;
  assign w23973 = w23966 | w23972 ;
  assign w23974 = ~\pi067 & w23973 ;
  assign w23975 = \pi036 ^ w23551 ;
  assign w23976 = ( \pi064 & w4266 ) | ( \pi064 & w23975 ) | ( w4266 & w23975 ) ;
  assign w23977 = w4425 ^ w23976 ;
  assign w23978 = ~w4266 & w23977 ;
  assign w23979 = ~w23815 & w23978 ;
  assign w23980 = ( ~\pi064 & w23551 ) | ( ~\pi064 & w23816 ) | ( w23551 & w23816 ) ;
  assign w23981 = \pi037 ^ w23980 ;
  assign w23982 = w23816 & ~w23981 ;
  assign w23983 = w23979 | w23982 ;
  assign w23984 = ~\pi066 & w23983 ;
  assign w23985 = ( \pi036 & ~w4438 ) | ( \pi036 & w23815 ) | ( ~w4438 & w23815 ) ;
  assign w23986 = \pi036 & w23985 ;
  assign w23987 = w4442 & ~w23815 ;
  assign w23988 = w23986 | w23987 ;
  assign w23989 = \pi065 ^ w23988 ;
  assign w23990 = w4445 | w23989 ;
  assign w23991 = w23816 | w23979 ;
  assign w23992 = ( w23968 & w23979 ) | ( w23968 & w23991 ) | ( w23979 & w23991 ) ;
  assign w23993 = \pi066 ^ w23992 ;
  assign w23994 = ~\pi065 & w23988 ;
  assign w23995 = w23990 | w23994 ;
  assign w23996 = ( w23993 & ~w23994 ) | ( w23993 & w23995 ) | ( ~w23994 & w23995 ) ;
  assign w23997 = \pi067 ^ w23973 ;
  assign w23998 = ( ~w23984 & w23996 ) | ( ~w23984 & w23997 ) | ( w23996 & w23997 ) ;
  assign w23999 = w23997 | w23998 ;
  assign w24000 = \pi068 ^ w23964 ;
  assign w24001 = ( ~w23974 & w23999 ) | ( ~w23974 & w24000 ) | ( w23999 & w24000 ) ;
  assign w24002 = w24000 | w24001 ;
  assign w24003 = \pi069 ^ w23958 ;
  assign w24004 = ( ~w23965 & w24002 ) | ( ~w23965 & w24003 ) | ( w24002 & w24003 ) ;
  assign w24005 = w24003 | w24004 ;
  assign w24006 = \pi070 ^ w23952 ;
  assign w24007 = ( ~w23959 & w24005 ) | ( ~w23959 & w24006 ) | ( w24005 & w24006 ) ;
  assign w24008 = w24006 | w24007 ;
  assign w24009 = \pi071 ^ w23946 ;
  assign w24010 = ( ~w23953 & w24008 ) | ( ~w23953 & w24009 ) | ( w24008 & w24009 ) ;
  assign w24011 = w24009 | w24010 ;
  assign w24012 = \pi072 ^ w23940 ;
  assign w24013 = ( ~w23947 & w24011 ) | ( ~w23947 & w24012 ) | ( w24011 & w24012 ) ;
  assign w24014 = w24012 | w24013 ;
  assign w24015 = \pi073 ^ w23934 ;
  assign w24016 = ( ~w23941 & w24014 ) | ( ~w23941 & w24015 ) | ( w24014 & w24015 ) ;
  assign w24017 = w24015 | w24016 ;
  assign w24018 = \pi074 ^ w23928 ;
  assign w24019 = ( ~w23935 & w24017 ) | ( ~w23935 & w24018 ) | ( w24017 & w24018 ) ;
  assign w24020 = w24018 | w24019 ;
  assign w24021 = \pi075 ^ w23922 ;
  assign w24022 = ( ~w23929 & w24020 ) | ( ~w23929 & w24021 ) | ( w24020 & w24021 ) ;
  assign w24023 = w24021 | w24022 ;
  assign w24024 = \pi076 ^ w23916 ;
  assign w24025 = ( ~w23923 & w24023 ) | ( ~w23923 & w24024 ) | ( w24023 & w24024 ) ;
  assign w24026 = w24024 | w24025 ;
  assign w24027 = \pi077 ^ w23910 ;
  assign w24028 = ( ~w23917 & w24026 ) | ( ~w23917 & w24027 ) | ( w24026 & w24027 ) ;
  assign w24029 = w24027 | w24028 ;
  assign w24030 = \pi078 ^ w23904 ;
  assign w24031 = ( ~w23911 & w24029 ) | ( ~w23911 & w24030 ) | ( w24029 & w24030 ) ;
  assign w24032 = w24030 | w24031 ;
  assign w24033 = \pi079 ^ w23898 ;
  assign w24034 = ( ~w23905 & w24032 ) | ( ~w23905 & w24033 ) | ( w24032 & w24033 ) ;
  assign w24035 = w24033 | w24034 ;
  assign w24036 = \pi080 ^ w23892 ;
  assign w24037 = ( ~w23899 & w24035 ) | ( ~w23899 & w24036 ) | ( w24035 & w24036 ) ;
  assign w24038 = w24036 | w24037 ;
  assign w24039 = \pi081 ^ w23886 ;
  assign w24040 = ( ~w23893 & w24038 ) | ( ~w23893 & w24039 ) | ( w24038 & w24039 ) ;
  assign w24041 = w24039 | w24040 ;
  assign w24042 = \pi082 ^ w23880 ;
  assign w24043 = ( ~w23887 & w24041 ) | ( ~w23887 & w24042 ) | ( w24041 & w24042 ) ;
  assign w24044 = w24042 | w24043 ;
  assign w24045 = \pi083 ^ w23874 ;
  assign w24046 = ( ~w23881 & w24044 ) | ( ~w23881 & w24045 ) | ( w24044 & w24045 ) ;
  assign w24047 = w24045 | w24046 ;
  assign w24048 = \pi084 ^ w23868 ;
  assign w24049 = ( ~w23875 & w24047 ) | ( ~w23875 & w24048 ) | ( w24047 & w24048 ) ;
  assign w24050 = w24048 | w24049 ;
  assign w24051 = \pi085 ^ w23862 ;
  assign w24052 = ( ~w23869 & w24050 ) | ( ~w23869 & w24051 ) | ( w24050 & w24051 ) ;
  assign w24053 = w24051 | w24052 ;
  assign w24054 = \pi086 ^ w23856 ;
  assign w24055 = ( ~w23863 & w24053 ) | ( ~w23863 & w24054 ) | ( w24053 & w24054 ) ;
  assign w24056 = w24054 | w24055 ;
  assign w24057 = \pi087 ^ w23850 ;
  assign w24058 = ( ~w23857 & w24056 ) | ( ~w23857 & w24057 ) | ( w24056 & w24057 ) ;
  assign w24059 = w24057 | w24058 ;
  assign w24060 = \pi088 ^ w23844 ;
  assign w24061 = ( ~w23851 & w24059 ) | ( ~w23851 & w24060 ) | ( w24059 & w24060 ) ;
  assign w24062 = w24060 | w24061 ;
  assign w24063 = \pi089 ^ w23838 ;
  assign w24064 = ( ~w23845 & w24062 ) | ( ~w23845 & w24063 ) | ( w24062 & w24063 ) ;
  assign w24065 = w24063 | w24064 ;
  assign w24066 = \pi090 ^ w23832 ;
  assign w24067 = ( ~w23839 & w24065 ) | ( ~w23839 & w24066 ) | ( w24065 & w24066 ) ;
  assign w24068 = w24066 | w24067 ;
  assign w24069 = \pi091 ^ w23821 ;
  assign w24070 = ( ~w23833 & w24068 ) | ( ~w23833 & w24069 ) | ( w24068 & w24069 ) ;
  assign w24071 = w24069 | w24070 ;
  assign w24072 = \pi092 ^ w23826 ;
  assign w24073 = w23827 & ~w24072 ;
  assign w24074 = ( w24071 & w24072 ) | ( w24071 & ~w24073 ) | ( w24072 & ~w24073 ) ;
  assign w24075 = ~\pi092 & w23826 ;
  assign w24076 = w24074 & ~w24075 ;
  assign w24077 = w4535 | w24076 ;
  assign w24078 = w23821 & w24077 ;
  assign w24079 = ~w23833 & w24068 ;
  assign w24080 = w24069 ^ w24079 ;
  assign w24081 = ~w24077 & w24080 ;
  assign w24082 = w24078 | w24081 ;
  assign w24083 = ~\pi092 & w24082 ;
  assign w24084 = w23832 & w24077 ;
  assign w24085 = ~w23839 & w24065 ;
  assign w24086 = w24066 ^ w24085 ;
  assign w24087 = ~w24077 & w24086 ;
  assign w24088 = w24084 | w24087 ;
  assign w24089 = ~\pi091 & w24088 ;
  assign w24090 = w23838 & w24077 ;
  assign w24091 = ~w23845 & w24062 ;
  assign w24092 = w24063 ^ w24091 ;
  assign w24093 = ~w24077 & w24092 ;
  assign w24094 = w24090 | w24093 ;
  assign w24095 = ~\pi090 & w24094 ;
  assign w24096 = w23844 & w24077 ;
  assign w24097 = ~w23851 & w24059 ;
  assign w24098 = w24060 ^ w24097 ;
  assign w24099 = ~w24077 & w24098 ;
  assign w24100 = w24096 | w24099 ;
  assign w24101 = ~\pi089 & w24100 ;
  assign w24102 = w23850 & w24077 ;
  assign w24103 = ~w23857 & w24056 ;
  assign w24104 = w24057 ^ w24103 ;
  assign w24105 = ~w24077 & w24104 ;
  assign w24106 = w24102 | w24105 ;
  assign w24107 = ~\pi088 & w24106 ;
  assign w24108 = w23856 & w24077 ;
  assign w24109 = ~w23863 & w24053 ;
  assign w24110 = w24054 ^ w24109 ;
  assign w24111 = ~w24077 & w24110 ;
  assign w24112 = w24108 | w24111 ;
  assign w24113 = ~\pi087 & w24112 ;
  assign w24114 = w23862 & w24077 ;
  assign w24115 = ~w23869 & w24050 ;
  assign w24116 = w24051 ^ w24115 ;
  assign w24117 = ~w24077 & w24116 ;
  assign w24118 = w24114 | w24117 ;
  assign w24119 = ~\pi086 & w24118 ;
  assign w24120 = w23868 & w24077 ;
  assign w24121 = ~w23875 & w24047 ;
  assign w24122 = w24048 ^ w24121 ;
  assign w24123 = ~w24077 & w24122 ;
  assign w24124 = w24120 | w24123 ;
  assign w24125 = ~\pi085 & w24124 ;
  assign w24126 = w23874 & w24077 ;
  assign w24127 = ~w23881 & w24044 ;
  assign w24128 = w24045 ^ w24127 ;
  assign w24129 = ~w24077 & w24128 ;
  assign w24130 = w24126 | w24129 ;
  assign w24131 = ~\pi084 & w24130 ;
  assign w24132 = w23880 & w24077 ;
  assign w24133 = ~w23887 & w24041 ;
  assign w24134 = w24042 ^ w24133 ;
  assign w24135 = ~w24077 & w24134 ;
  assign w24136 = w24132 | w24135 ;
  assign w24137 = ~\pi083 & w24136 ;
  assign w24138 = w23886 & w24077 ;
  assign w24139 = ~w23893 & w24038 ;
  assign w24140 = w24039 ^ w24139 ;
  assign w24141 = ~w24077 & w24140 ;
  assign w24142 = w24138 | w24141 ;
  assign w24143 = ~\pi082 & w24142 ;
  assign w24144 = w23892 & w24077 ;
  assign w24145 = ~w23899 & w24035 ;
  assign w24146 = w24036 ^ w24145 ;
  assign w24147 = ~w24077 & w24146 ;
  assign w24148 = w24144 | w24147 ;
  assign w24149 = ~\pi081 & w24148 ;
  assign w24150 = w23898 & w24077 ;
  assign w24151 = ~w23905 & w24032 ;
  assign w24152 = w24033 ^ w24151 ;
  assign w24153 = ~w24077 & w24152 ;
  assign w24154 = w24150 | w24153 ;
  assign w24155 = ~\pi080 & w24154 ;
  assign w24156 = w23904 & w24077 ;
  assign w24157 = ~w23911 & w24029 ;
  assign w24158 = w24030 ^ w24157 ;
  assign w24159 = ~w24077 & w24158 ;
  assign w24160 = w24156 | w24159 ;
  assign w24161 = ~\pi079 & w24160 ;
  assign w24162 = w23910 & w24077 ;
  assign w24163 = ~w23917 & w24026 ;
  assign w24164 = w24027 ^ w24163 ;
  assign w24165 = ~w24077 & w24164 ;
  assign w24166 = w24162 | w24165 ;
  assign w24167 = ~\pi078 & w24166 ;
  assign w24168 = w23916 & w24077 ;
  assign w24169 = ~w23923 & w24023 ;
  assign w24170 = w24024 ^ w24169 ;
  assign w24171 = ~w24077 & w24170 ;
  assign w24172 = w24168 | w24171 ;
  assign w24173 = ~\pi077 & w24172 ;
  assign w24174 = w23922 & w24077 ;
  assign w24175 = ~w23929 & w24020 ;
  assign w24176 = w24021 ^ w24175 ;
  assign w24177 = ~w24077 & w24176 ;
  assign w24178 = w24174 | w24177 ;
  assign w24179 = ~\pi076 & w24178 ;
  assign w24180 = w23928 & w24077 ;
  assign w24181 = ~w23935 & w24017 ;
  assign w24182 = w24018 ^ w24181 ;
  assign w24183 = ~w24077 & w24182 ;
  assign w24184 = w24180 | w24183 ;
  assign w24185 = ~\pi075 & w24184 ;
  assign w24186 = w23934 & w24077 ;
  assign w24187 = ~w23941 & w24014 ;
  assign w24188 = w24015 ^ w24187 ;
  assign w24189 = ~w24077 & w24188 ;
  assign w24190 = w24186 | w24189 ;
  assign w24191 = ~\pi074 & w24190 ;
  assign w24192 = w23940 & w24077 ;
  assign w24193 = ~w23947 & w24011 ;
  assign w24194 = w24012 ^ w24193 ;
  assign w24195 = ~w24077 & w24194 ;
  assign w24196 = w24192 | w24195 ;
  assign w24197 = ~\pi073 & w24196 ;
  assign w24198 = w23946 & w24077 ;
  assign w24199 = ~w23953 & w24008 ;
  assign w24200 = w24009 ^ w24199 ;
  assign w24201 = ~w24077 & w24200 ;
  assign w24202 = w24198 | w24201 ;
  assign w24203 = ~\pi072 & w24202 ;
  assign w24204 = w23952 & w24077 ;
  assign w24205 = ~w23959 & w24005 ;
  assign w24206 = w24006 ^ w24205 ;
  assign w24207 = ~w24077 & w24206 ;
  assign w24208 = w24204 | w24207 ;
  assign w24209 = ~\pi071 & w24208 ;
  assign w24210 = w23958 & w24077 ;
  assign w24211 = ~w23965 & w24002 ;
  assign w24212 = w24003 ^ w24211 ;
  assign w24213 = ~w24077 & w24212 ;
  assign w24214 = w24210 | w24213 ;
  assign w24215 = ~\pi070 & w24214 ;
  assign w24216 = w23964 & w24077 ;
  assign w24217 = ~w23974 & w23999 ;
  assign w24218 = w24000 ^ w24217 ;
  assign w24219 = ~w24077 & w24218 ;
  assign w24220 = w24216 | w24219 ;
  assign w24221 = ~\pi069 & w24220 ;
  assign w24222 = w23973 & w24077 ;
  assign w24223 = ~w23984 & w23996 ;
  assign w24224 = w23997 ^ w24223 ;
  assign w24225 = ~w24077 & w24224 ;
  assign w24226 = w24222 | w24225 ;
  assign w24227 = ~\pi068 & w24226 ;
  assign w24228 = w23983 & w24077 ;
  assign w24229 = ~w23988 & w23990 ;
  assign w24230 = ( \pi065 & w23990 ) | ( \pi065 & w24229 ) | ( w23990 & w24229 ) ;
  assign w24231 = w23993 ^ w24230 ;
  assign w24232 = ~w24077 & w24231 ;
  assign w24233 = w24228 | w24232 ;
  assign w24234 = ~\pi067 & w24233 ;
  assign w24235 = ( ~w4535 & w23986 ) | ( ~w4535 & w23987 ) | ( w23986 & w23987 ) ;
  assign w24236 = \pi065 ^ w24235 ;
  assign w24237 = ( w4445 & ~w4535 ) | ( w4445 & w24236 ) | ( ~w4535 & w24236 ) ;
  assign w24238 = ( w4445 & w24076 ) | ( w4445 & w24236 ) | ( w24076 & w24236 ) ;
  assign w24239 = w24237 & ~w24238 ;
  assign w24240 = ( w23988 & w24077 ) | ( w23988 & w24239 ) | ( w24077 & w24239 ) ;
  assign w24241 = w24239 | w24240 ;
  assign w24242 = ~\pi066 & w24241 ;
  assign w24243 = ( \pi035 & ~w4707 ) | ( \pi035 & w24076 ) | ( ~w4707 & w24076 ) ;
  assign w24244 = \pi035 & w24243 ;
  assign w24245 = ( ~w275 & w290 ) | ( ~w275 & w24076 ) | ( w290 & w24076 ) ;
  assign w24246 = w4711 & ~w24245 ;
  assign w24247 = ~w23988 & w24077 ;
  assign w24248 = ( w24077 & w24239 ) | ( w24077 & ~w24247 ) | ( w24239 & ~w24247 ) ;
  assign w24249 = \pi066 ^ w24248 ;
  assign w24250 = w24244 | w24246 ;
  assign w24251 = ( \pi065 & w4714 ) | ( \pi065 & ~w24250 ) | ( w4714 & ~w24250 ) ;
  assign w24252 = w24249 | w24251 ;
  assign w24253 = \pi067 ^ w24233 ;
  assign w24254 = ( ~w24242 & w24252 ) | ( ~w24242 & w24253 ) | ( w24252 & w24253 ) ;
  assign w24255 = w24253 | w24254 ;
  assign w24256 = \pi068 ^ w24226 ;
  assign w24257 = ( ~w24234 & w24255 ) | ( ~w24234 & w24256 ) | ( w24255 & w24256 ) ;
  assign w24258 = w24256 | w24257 ;
  assign w24259 = \pi069 ^ w24220 ;
  assign w24260 = ( ~w24227 & w24258 ) | ( ~w24227 & w24259 ) | ( w24258 & w24259 ) ;
  assign w24261 = w24259 | w24260 ;
  assign w24262 = \pi070 ^ w24214 ;
  assign w24263 = ( ~w24221 & w24261 ) | ( ~w24221 & w24262 ) | ( w24261 & w24262 ) ;
  assign w24264 = w24262 | w24263 ;
  assign w24265 = \pi071 ^ w24208 ;
  assign w24266 = ( ~w24215 & w24264 ) | ( ~w24215 & w24265 ) | ( w24264 & w24265 ) ;
  assign w24267 = w24265 | w24266 ;
  assign w24268 = \pi072 ^ w24202 ;
  assign w24269 = ( ~w24209 & w24267 ) | ( ~w24209 & w24268 ) | ( w24267 & w24268 ) ;
  assign w24270 = w24268 | w24269 ;
  assign w24271 = \pi073 ^ w24196 ;
  assign w24272 = ( ~w24203 & w24270 ) | ( ~w24203 & w24271 ) | ( w24270 & w24271 ) ;
  assign w24273 = w24271 | w24272 ;
  assign w24274 = \pi074 ^ w24190 ;
  assign w24275 = ( ~w24197 & w24273 ) | ( ~w24197 & w24274 ) | ( w24273 & w24274 ) ;
  assign w24276 = w24274 | w24275 ;
  assign w24277 = \pi075 ^ w24184 ;
  assign w24278 = ( ~w24191 & w24276 ) | ( ~w24191 & w24277 ) | ( w24276 & w24277 ) ;
  assign w24279 = w24277 | w24278 ;
  assign w24280 = \pi076 ^ w24178 ;
  assign w24281 = ( ~w24185 & w24279 ) | ( ~w24185 & w24280 ) | ( w24279 & w24280 ) ;
  assign w24282 = w24280 | w24281 ;
  assign w24283 = \pi077 ^ w24172 ;
  assign w24284 = ( ~w24179 & w24282 ) | ( ~w24179 & w24283 ) | ( w24282 & w24283 ) ;
  assign w24285 = w24283 | w24284 ;
  assign w24286 = \pi078 ^ w24166 ;
  assign w24287 = ( ~w24173 & w24285 ) | ( ~w24173 & w24286 ) | ( w24285 & w24286 ) ;
  assign w24288 = w24286 | w24287 ;
  assign w24289 = \pi079 ^ w24160 ;
  assign w24290 = ( ~w24167 & w24288 ) | ( ~w24167 & w24289 ) | ( w24288 & w24289 ) ;
  assign w24291 = w24289 | w24290 ;
  assign w24292 = \pi080 ^ w24154 ;
  assign w24293 = ( ~w24161 & w24291 ) | ( ~w24161 & w24292 ) | ( w24291 & w24292 ) ;
  assign w24294 = w24292 | w24293 ;
  assign w24295 = \pi081 ^ w24148 ;
  assign w24296 = ( ~w24155 & w24294 ) | ( ~w24155 & w24295 ) | ( w24294 & w24295 ) ;
  assign w24297 = w24295 | w24296 ;
  assign w24298 = \pi082 ^ w24142 ;
  assign w24299 = ( ~w24149 & w24297 ) | ( ~w24149 & w24298 ) | ( w24297 & w24298 ) ;
  assign w24300 = w24298 | w24299 ;
  assign w24301 = \pi083 ^ w24136 ;
  assign w24302 = ( ~w24143 & w24300 ) | ( ~w24143 & w24301 ) | ( w24300 & w24301 ) ;
  assign w24303 = w24301 | w24302 ;
  assign w24304 = \pi084 ^ w24130 ;
  assign w24305 = ( ~w24137 & w24303 ) | ( ~w24137 & w24304 ) | ( w24303 & w24304 ) ;
  assign w24306 = w24304 | w24305 ;
  assign w24307 = \pi085 ^ w24124 ;
  assign w24308 = ( ~w24131 & w24306 ) | ( ~w24131 & w24307 ) | ( w24306 & w24307 ) ;
  assign w24309 = w24307 | w24308 ;
  assign w24310 = \pi086 ^ w24118 ;
  assign w24311 = ( ~w24125 & w24309 ) | ( ~w24125 & w24310 ) | ( w24309 & w24310 ) ;
  assign w24312 = w24310 | w24311 ;
  assign w24313 = \pi087 ^ w24112 ;
  assign w24314 = ( ~w24119 & w24312 ) | ( ~w24119 & w24313 ) | ( w24312 & w24313 ) ;
  assign w24315 = w24313 | w24314 ;
  assign w24316 = \pi088 ^ w24106 ;
  assign w24317 = ( ~w24113 & w24315 ) | ( ~w24113 & w24316 ) | ( w24315 & w24316 ) ;
  assign w24318 = w24316 | w24317 ;
  assign w24319 = \pi089 ^ w24100 ;
  assign w24320 = ( ~w24107 & w24318 ) | ( ~w24107 & w24319 ) | ( w24318 & w24319 ) ;
  assign w24321 = w24319 | w24320 ;
  assign w24322 = \pi090 ^ w24094 ;
  assign w24323 = ( ~w24101 & w24321 ) | ( ~w24101 & w24322 ) | ( w24321 & w24322 ) ;
  assign w24324 = w24322 | w24323 ;
  assign w24325 = \pi091 ^ w24088 ;
  assign w24326 = ( ~w24095 & w24324 ) | ( ~w24095 & w24325 ) | ( w24324 & w24325 ) ;
  assign w24327 = w24325 | w24326 ;
  assign w24328 = \pi092 ^ w24082 ;
  assign w24329 = ( ~w24089 & w24327 ) | ( ~w24089 & w24328 ) | ( w24327 & w24328 ) ;
  assign w24330 = w24328 | w24329 ;
  assign w24331 = w23826 & w24077 ;
  assign w24332 = ~w23827 & w24071 ;
  assign w24333 = w24072 ^ w24332 ;
  assign w24334 = ~w24077 & w24333 ;
  assign w24335 = w24331 | w24334 ;
  assign w24336 = ~\pi093 & w24335 ;
  assign w24337 = ( \pi093 & ~w24331 ) | ( \pi093 & w24334 ) | ( ~w24331 & w24334 ) ;
  assign w24338 = ~w24334 & w24337 ;
  assign w24339 = w24336 | w24338 ;
  assign w24340 = ( ~w24083 & w24330 ) | ( ~w24083 & w24339 ) | ( w24330 & w24339 ) ;
  assign w24341 = ( w4810 & ~w24339 ) | ( w4810 & w24340 ) | ( ~w24339 & w24340 ) ;
  assign w24342 = w24339 | w24341 ;
  assign w24343 = ~w4535 & w24335 ;
  assign w24344 = w24342 & ~w24343 ;
  assign w24345 = ~w24089 & w24327 ;
  assign w24346 = w24328 ^ w24345 ;
  assign w24347 = ~w24344 & w24346 ;
  assign w24348 = ( w24082 & w24342 ) | ( w24082 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24349 = ~w24343 & w24348 ;
  assign w24350 = w24347 | w24349 ;
  assign w24351 = ( ~w24083 & w24330 ) | ( ~w24083 & w24344 ) | ( w24330 & w24344 ) ;
  assign w24352 = w24339 ^ w24351 ;
  assign w24353 = ~w24344 & w24352 ;
  assign w24354 = ( w4535 & ~w24335 ) | ( w4535 & w24342 ) | ( ~w24335 & w24342 ) ;
  assign w24355 = w24335 & w24354 ;
  assign w24356 = w24353 | w24355 ;
  assign w24357 = ~\pi093 & w24350 ;
  assign w24358 = ~w24095 & w24324 ;
  assign w24359 = w24325 ^ w24358 ;
  assign w24360 = ~w24344 & w24359 ;
  assign w24361 = ( w24088 & w24342 ) | ( w24088 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24362 = ~w24343 & w24361 ;
  assign w24363 = w24360 | w24362 ;
  assign w24364 = ~\pi092 & w24363 ;
  assign w24365 = ~w24101 & w24321 ;
  assign w24366 = w24322 ^ w24365 ;
  assign w24367 = ~w24344 & w24366 ;
  assign w24368 = ( w24094 & w24342 ) | ( w24094 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24369 = ~w24343 & w24368 ;
  assign w24370 = w24367 | w24369 ;
  assign w24371 = ~\pi091 & w24370 ;
  assign w24372 = ~w24107 & w24318 ;
  assign w24373 = w24319 ^ w24372 ;
  assign w24374 = ~w24344 & w24373 ;
  assign w24375 = ( w24100 & w24342 ) | ( w24100 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24376 = ~w24343 & w24375 ;
  assign w24377 = w24374 | w24376 ;
  assign w24378 = ~\pi090 & w24377 ;
  assign w24379 = ~w24113 & w24315 ;
  assign w24380 = w24316 ^ w24379 ;
  assign w24381 = ~w24344 & w24380 ;
  assign w24382 = ( w24106 & w24342 ) | ( w24106 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24383 = ~w24343 & w24382 ;
  assign w24384 = w24381 | w24383 ;
  assign w24385 = ~\pi089 & w24384 ;
  assign w24386 = ~w24119 & w24312 ;
  assign w24387 = w24313 ^ w24386 ;
  assign w24388 = ~w24344 & w24387 ;
  assign w24389 = ( w24112 & w24342 ) | ( w24112 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24390 = ~w24343 & w24389 ;
  assign w24391 = w24388 | w24390 ;
  assign w24392 = ~\pi088 & w24391 ;
  assign w24393 = ~w24125 & w24309 ;
  assign w24394 = w24310 ^ w24393 ;
  assign w24395 = ~w24344 & w24394 ;
  assign w24396 = ( w24118 & w24342 ) | ( w24118 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24397 = ~w24343 & w24396 ;
  assign w24398 = w24395 | w24397 ;
  assign w24399 = ~\pi087 & w24398 ;
  assign w24400 = ~w24131 & w24306 ;
  assign w24401 = w24307 ^ w24400 ;
  assign w24402 = ~w24344 & w24401 ;
  assign w24403 = ( w24124 & w24342 ) | ( w24124 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24404 = ~w24343 & w24403 ;
  assign w24405 = w24402 | w24404 ;
  assign w24406 = ~\pi086 & w24405 ;
  assign w24407 = ~w24137 & w24303 ;
  assign w24408 = w24304 ^ w24407 ;
  assign w24409 = ~w24344 & w24408 ;
  assign w24410 = ( w24130 & w24342 ) | ( w24130 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24411 = ~w24343 & w24410 ;
  assign w24412 = w24409 | w24411 ;
  assign w24413 = ~\pi085 & w24412 ;
  assign w24414 = ~w24143 & w24300 ;
  assign w24415 = w24301 ^ w24414 ;
  assign w24416 = ~w24344 & w24415 ;
  assign w24417 = ( w24136 & w24342 ) | ( w24136 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24418 = ~w24343 & w24417 ;
  assign w24419 = w24416 | w24418 ;
  assign w24420 = ~\pi084 & w24419 ;
  assign w24421 = ~w24149 & w24297 ;
  assign w24422 = w24298 ^ w24421 ;
  assign w24423 = ~w24344 & w24422 ;
  assign w24424 = ( w24142 & w24342 ) | ( w24142 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24425 = ~w24343 & w24424 ;
  assign w24426 = w24423 | w24425 ;
  assign w24427 = ~\pi083 & w24426 ;
  assign w24428 = ~w24155 & w24294 ;
  assign w24429 = w24295 ^ w24428 ;
  assign w24430 = ~w24344 & w24429 ;
  assign w24431 = ( w24148 & w24342 ) | ( w24148 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24432 = ~w24343 & w24431 ;
  assign w24433 = w24430 | w24432 ;
  assign w24434 = ~\pi082 & w24433 ;
  assign w24435 = ~w24161 & w24291 ;
  assign w24436 = w24292 ^ w24435 ;
  assign w24437 = ~w24344 & w24436 ;
  assign w24438 = ( w24154 & w24342 ) | ( w24154 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24439 = ~w24343 & w24438 ;
  assign w24440 = w24437 | w24439 ;
  assign w24441 = ~\pi081 & w24440 ;
  assign w24442 = ~w24167 & w24288 ;
  assign w24443 = w24289 ^ w24442 ;
  assign w24444 = ~w24344 & w24443 ;
  assign w24445 = ( w24160 & w24342 ) | ( w24160 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24446 = ~w24343 & w24445 ;
  assign w24447 = w24444 | w24446 ;
  assign w24448 = ~\pi080 & w24447 ;
  assign w24449 = ~w24173 & w24285 ;
  assign w24450 = w24286 ^ w24449 ;
  assign w24451 = ~w24344 & w24450 ;
  assign w24452 = ( w24166 & w24342 ) | ( w24166 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24453 = ~w24343 & w24452 ;
  assign w24454 = w24451 | w24453 ;
  assign w24455 = ~\pi079 & w24454 ;
  assign w24456 = ~w24179 & w24282 ;
  assign w24457 = w24283 ^ w24456 ;
  assign w24458 = ~w24344 & w24457 ;
  assign w24459 = ( w24172 & w24342 ) | ( w24172 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24460 = ~w24343 & w24459 ;
  assign w24461 = w24458 | w24460 ;
  assign w24462 = ~\pi078 & w24461 ;
  assign w24463 = ~w24185 & w24279 ;
  assign w24464 = w24280 ^ w24463 ;
  assign w24465 = ~w24344 & w24464 ;
  assign w24466 = ( w24178 & w24342 ) | ( w24178 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24467 = ~w24343 & w24466 ;
  assign w24468 = w24465 | w24467 ;
  assign w24469 = ~\pi077 & w24468 ;
  assign w24470 = ~w24191 & w24276 ;
  assign w24471 = w24277 ^ w24470 ;
  assign w24472 = ~w24344 & w24471 ;
  assign w24473 = ( w24184 & w24342 ) | ( w24184 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24474 = ~w24343 & w24473 ;
  assign w24475 = w24472 | w24474 ;
  assign w24476 = ~\pi076 & w24475 ;
  assign w24477 = ~w24197 & w24273 ;
  assign w24478 = w24274 ^ w24477 ;
  assign w24479 = ~w24344 & w24478 ;
  assign w24480 = ( w24190 & w24342 ) | ( w24190 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24481 = ~w24343 & w24480 ;
  assign w24482 = w24479 | w24481 ;
  assign w24483 = ~\pi075 & w24482 ;
  assign w24484 = ~w24203 & w24270 ;
  assign w24485 = w24271 ^ w24484 ;
  assign w24486 = ~w24344 & w24485 ;
  assign w24487 = ( w24196 & w24342 ) | ( w24196 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24488 = ~w24343 & w24487 ;
  assign w24489 = w24486 | w24488 ;
  assign w24490 = ~\pi074 & w24489 ;
  assign w24491 = ~w24209 & w24267 ;
  assign w24492 = w24268 ^ w24491 ;
  assign w24493 = ~w24344 & w24492 ;
  assign w24494 = ( w24202 & w24342 ) | ( w24202 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24495 = ~w24343 & w24494 ;
  assign w24496 = w24493 | w24495 ;
  assign w24497 = ~\pi073 & w24496 ;
  assign w24498 = ~w24215 & w24264 ;
  assign w24499 = w24265 ^ w24498 ;
  assign w24500 = ~w24344 & w24499 ;
  assign w24501 = ( w24208 & w24342 ) | ( w24208 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24502 = ~w24343 & w24501 ;
  assign w24503 = w24500 | w24502 ;
  assign w24504 = ~\pi072 & w24503 ;
  assign w24505 = ~w24221 & w24261 ;
  assign w24506 = w24262 ^ w24505 ;
  assign w24507 = ~w24344 & w24506 ;
  assign w24508 = ( w24214 & w24342 ) | ( w24214 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24509 = ~w24343 & w24508 ;
  assign w24510 = w24507 | w24509 ;
  assign w24511 = ~\pi071 & w24510 ;
  assign w24512 = ~w24227 & w24258 ;
  assign w24513 = w24259 ^ w24512 ;
  assign w24514 = ~w24344 & w24513 ;
  assign w24515 = ( w24220 & w24342 ) | ( w24220 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24516 = ~w24343 & w24515 ;
  assign w24517 = w24514 | w24516 ;
  assign w24518 = ~\pi070 & w24517 ;
  assign w24519 = ~w24234 & w24255 ;
  assign w24520 = w24256 ^ w24519 ;
  assign w24521 = ~w24344 & w24520 ;
  assign w24522 = ( w24226 & w24342 ) | ( w24226 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24523 = ~w24343 & w24522 ;
  assign w24524 = w24521 | w24523 ;
  assign w24525 = ~\pi069 & w24524 ;
  assign w24526 = ~w24242 & w24252 ;
  assign w24527 = w24253 ^ w24526 ;
  assign w24528 = ~w24344 & w24527 ;
  assign w24529 = ( w24233 & w24342 ) | ( w24233 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24530 = ~w24343 & w24529 ;
  assign w24531 = w24528 | w24530 ;
  assign w24532 = ~\pi068 & w24531 ;
  assign w24533 = w24249 ^ w24251 ;
  assign w24534 = ~w24344 & w24533 ;
  assign w24535 = ( w24241 & w24342 ) | ( w24241 & w24343 ) | ( w24342 & w24343 ) ;
  assign w24536 = ~w24343 & w24535 ;
  assign w24537 = w24534 | w24536 ;
  assign w24538 = ~\pi067 & w24537 ;
  assign w24539 = w4714 ^ w24250 ;
  assign w24540 = \pi065 ^ w24539 ;
  assign w24541 = w24344 ^ w24540 ;
  assign w24542 = ( w24250 & w24540 ) | ( w24250 & w24541 ) | ( w24540 & w24541 ) ;
  assign w24543 = ~\pi066 & w24542 ;
  assign w24544 = w24250 ^ w24344 ;
  assign w24545 = ( w24250 & w24540 ) | ( w24250 & ~w24544 ) | ( w24540 & ~w24544 ) ;
  assign w24546 = \pi066 ^ w24545 ;
  assign w24547 = ( \pi064 & ~w24344 ) | ( \pi064 & w24546 ) | ( ~w24344 & w24546 ) ;
  assign w24548 = \pi034 ^ w24547 ;
  assign w24549 = ( \pi065 & w5287 ) | ( \pi065 & ~w24548 ) | ( w5287 & ~w24548 ) ;
  assign w24550 = w24546 | w24549 ;
  assign w24551 = \pi067 ^ w24537 ;
  assign w24552 = ( ~w24543 & w24550 ) | ( ~w24543 & w24551 ) | ( w24550 & w24551 ) ;
  assign w24553 = w24551 | w24552 ;
  assign w24554 = \pi068 ^ w24531 ;
  assign w24555 = ( ~w24538 & w24553 ) | ( ~w24538 & w24554 ) | ( w24553 & w24554 ) ;
  assign w24556 = w24554 | w24555 ;
  assign w24557 = \pi069 ^ w24524 ;
  assign w24558 = ( ~w24532 & w24556 ) | ( ~w24532 & w24557 ) | ( w24556 & w24557 ) ;
  assign w24559 = w24557 | w24558 ;
  assign w24560 = \pi070 ^ w24517 ;
  assign w24561 = ( ~w24525 & w24559 ) | ( ~w24525 & w24560 ) | ( w24559 & w24560 ) ;
  assign w24562 = w24560 | w24561 ;
  assign w24563 = \pi071 ^ w24510 ;
  assign w24564 = ( ~w24518 & w24562 ) | ( ~w24518 & w24563 ) | ( w24562 & w24563 ) ;
  assign w24565 = w24563 | w24564 ;
  assign w24566 = \pi072 ^ w24503 ;
  assign w24567 = ( ~w24511 & w24565 ) | ( ~w24511 & w24566 ) | ( w24565 & w24566 ) ;
  assign w24568 = w24566 | w24567 ;
  assign w24569 = \pi073 ^ w24496 ;
  assign w24570 = ( ~w24504 & w24568 ) | ( ~w24504 & w24569 ) | ( w24568 & w24569 ) ;
  assign w24571 = w24569 | w24570 ;
  assign w24572 = \pi074 ^ w24489 ;
  assign w24573 = ( ~w24497 & w24571 ) | ( ~w24497 & w24572 ) | ( w24571 & w24572 ) ;
  assign w24574 = w24572 | w24573 ;
  assign w24575 = \pi075 ^ w24482 ;
  assign w24576 = ( ~w24490 & w24574 ) | ( ~w24490 & w24575 ) | ( w24574 & w24575 ) ;
  assign w24577 = w24575 | w24576 ;
  assign w24578 = \pi076 ^ w24475 ;
  assign w24579 = ( ~w24483 & w24577 ) | ( ~w24483 & w24578 ) | ( w24577 & w24578 ) ;
  assign w24580 = w24578 | w24579 ;
  assign w24581 = \pi077 ^ w24468 ;
  assign w24582 = ( ~w24476 & w24580 ) | ( ~w24476 & w24581 ) | ( w24580 & w24581 ) ;
  assign w24583 = w24581 | w24582 ;
  assign w24584 = \pi078 ^ w24461 ;
  assign w24585 = ( ~w24469 & w24583 ) | ( ~w24469 & w24584 ) | ( w24583 & w24584 ) ;
  assign w24586 = w24584 | w24585 ;
  assign w24587 = \pi079 ^ w24454 ;
  assign w24588 = ( ~w24462 & w24586 ) | ( ~w24462 & w24587 ) | ( w24586 & w24587 ) ;
  assign w24589 = w24587 | w24588 ;
  assign w24590 = \pi080 ^ w24447 ;
  assign w24591 = ( ~w24455 & w24589 ) | ( ~w24455 & w24590 ) | ( w24589 & w24590 ) ;
  assign w24592 = w24590 | w24591 ;
  assign w24593 = \pi081 ^ w24440 ;
  assign w24594 = ( ~w24448 & w24592 ) | ( ~w24448 & w24593 ) | ( w24592 & w24593 ) ;
  assign w24595 = w24593 | w24594 ;
  assign w24596 = \pi082 ^ w24433 ;
  assign w24597 = ( ~w24441 & w24595 ) | ( ~w24441 & w24596 ) | ( w24595 & w24596 ) ;
  assign w24598 = w24596 | w24597 ;
  assign w24599 = \pi083 ^ w24426 ;
  assign w24600 = ( ~w24434 & w24598 ) | ( ~w24434 & w24599 ) | ( w24598 & w24599 ) ;
  assign w24601 = w24599 | w24600 ;
  assign w24602 = \pi084 ^ w24419 ;
  assign w24603 = ( ~w24427 & w24601 ) | ( ~w24427 & w24602 ) | ( w24601 & w24602 ) ;
  assign w24604 = w24602 | w24603 ;
  assign w24605 = \pi085 ^ w24412 ;
  assign w24606 = ( ~w24420 & w24604 ) | ( ~w24420 & w24605 ) | ( w24604 & w24605 ) ;
  assign w24607 = w24605 | w24606 ;
  assign w24608 = \pi086 ^ w24405 ;
  assign w24609 = ( ~w24413 & w24607 ) | ( ~w24413 & w24608 ) | ( w24607 & w24608 ) ;
  assign w24610 = w24608 | w24609 ;
  assign w24611 = \pi087 ^ w24398 ;
  assign w24612 = ( ~w24406 & w24610 ) | ( ~w24406 & w24611 ) | ( w24610 & w24611 ) ;
  assign w24613 = w24611 | w24612 ;
  assign w24614 = \pi088 ^ w24391 ;
  assign w24615 = ( ~w24399 & w24613 ) | ( ~w24399 & w24614 ) | ( w24613 & w24614 ) ;
  assign w24616 = w24614 | w24615 ;
  assign w24617 = \pi089 ^ w24384 ;
  assign w24618 = ( ~w24392 & w24616 ) | ( ~w24392 & w24617 ) | ( w24616 & w24617 ) ;
  assign w24619 = w24617 | w24618 ;
  assign w24620 = \pi090 ^ w24377 ;
  assign w24621 = ( ~w24385 & w24619 ) | ( ~w24385 & w24620 ) | ( w24619 & w24620 ) ;
  assign w24622 = w24620 | w24621 ;
  assign w24623 = \pi091 ^ w24370 ;
  assign w24624 = ( ~w24378 & w24622 ) | ( ~w24378 & w24623 ) | ( w24622 & w24623 ) ;
  assign w24625 = w24623 | w24624 ;
  assign w24626 = \pi092 ^ w24363 ;
  assign w24627 = ( ~w24371 & w24625 ) | ( ~w24371 & w24626 ) | ( w24625 & w24626 ) ;
  assign w24628 = w24626 | w24627 ;
  assign w24629 = \pi093 ^ w24350 ;
  assign w24630 = ( ~w24364 & w24628 ) | ( ~w24364 & w24629 ) | ( w24628 & w24629 ) ;
  assign w24631 = w24629 | w24630 ;
  assign w24632 = \pi094 ^ w24356 ;
  assign w24633 = w24357 & ~w24632 ;
  assign w24634 = ( w24631 & w24632 ) | ( w24631 & ~w24633 ) | ( w24632 & ~w24633 ) ;
  assign w24635 = ~\pi094 & w24356 ;
  assign w24636 = w24634 & ~w24635 ;
  assign w24637 = w5117 | w24636 ;
  assign w24638 = w24350 & w24637 ;
  assign w24639 = ~w24364 & w24628 ;
  assign w24640 = w24629 ^ w24639 ;
  assign w24641 = ~w24637 & w24640 ;
  assign w24642 = w24638 | w24641 ;
  assign w24643 = w24356 & w24637 ;
  assign w24644 = ~w24357 & w24631 ;
  assign w24645 = w24632 ^ w24644 ;
  assign w24646 = ~w24637 & w24645 ;
  assign w24647 = w24643 | w24646 ;
  assign w24648 = ~\pi094 & w24642 ;
  assign w24649 = w24363 & w24637 ;
  assign w24650 = ~w24371 & w24625 ;
  assign w24651 = w24626 ^ w24650 ;
  assign w24652 = ~w24637 & w24651 ;
  assign w24653 = w24649 | w24652 ;
  assign w24654 = ~\pi093 & w24653 ;
  assign w24655 = w24370 & w24637 ;
  assign w24656 = ~w24378 & w24622 ;
  assign w24657 = w24623 ^ w24656 ;
  assign w24658 = ~w24637 & w24657 ;
  assign w24659 = w24655 | w24658 ;
  assign w24660 = ~\pi092 & w24659 ;
  assign w24661 = w24377 & w24637 ;
  assign w24662 = ~w24385 & w24619 ;
  assign w24663 = w24620 ^ w24662 ;
  assign w24664 = ~w24637 & w24663 ;
  assign w24665 = w24661 | w24664 ;
  assign w24666 = ~\pi091 & w24665 ;
  assign w24667 = w24384 & w24637 ;
  assign w24668 = ~w24392 & w24616 ;
  assign w24669 = w24617 ^ w24668 ;
  assign w24670 = ~w24637 & w24669 ;
  assign w24671 = w24667 | w24670 ;
  assign w24672 = ~\pi090 & w24671 ;
  assign w24673 = w24391 & w24637 ;
  assign w24674 = ~w24399 & w24613 ;
  assign w24675 = w24614 ^ w24674 ;
  assign w24676 = ~w24637 & w24675 ;
  assign w24677 = w24673 | w24676 ;
  assign w24678 = ~\pi089 & w24677 ;
  assign w24679 = w24398 & w24637 ;
  assign w24680 = ~w24406 & w24610 ;
  assign w24681 = w24611 ^ w24680 ;
  assign w24682 = ~w24637 & w24681 ;
  assign w24683 = w24679 | w24682 ;
  assign w24684 = ~\pi088 & w24683 ;
  assign w24685 = w24405 & w24637 ;
  assign w24686 = ~w24413 & w24607 ;
  assign w24687 = w24608 ^ w24686 ;
  assign w24688 = ~w24637 & w24687 ;
  assign w24689 = w24685 | w24688 ;
  assign w24690 = ~\pi087 & w24689 ;
  assign w24691 = w24412 & w24637 ;
  assign w24692 = ~w24420 & w24604 ;
  assign w24693 = w24605 ^ w24692 ;
  assign w24694 = ~w24637 & w24693 ;
  assign w24695 = w24691 | w24694 ;
  assign w24696 = ~\pi086 & w24695 ;
  assign w24697 = w24419 & w24637 ;
  assign w24698 = ~w24427 & w24601 ;
  assign w24699 = w24602 ^ w24698 ;
  assign w24700 = ~w24637 & w24699 ;
  assign w24701 = w24697 | w24700 ;
  assign w24702 = ~\pi085 & w24701 ;
  assign w24703 = w24426 & w24637 ;
  assign w24704 = ~w24434 & w24598 ;
  assign w24705 = w24599 ^ w24704 ;
  assign w24706 = ~w24637 & w24705 ;
  assign w24707 = w24703 | w24706 ;
  assign w24708 = ~\pi084 & w24707 ;
  assign w24709 = w24433 & w24637 ;
  assign w24710 = ~w24441 & w24595 ;
  assign w24711 = w24596 ^ w24710 ;
  assign w24712 = ~w24637 & w24711 ;
  assign w24713 = w24709 | w24712 ;
  assign w24714 = ~\pi083 & w24713 ;
  assign w24715 = w24440 & w24637 ;
  assign w24716 = ~w24448 & w24592 ;
  assign w24717 = w24593 ^ w24716 ;
  assign w24718 = ~w24637 & w24717 ;
  assign w24719 = w24715 | w24718 ;
  assign w24720 = ~\pi082 & w24719 ;
  assign w24721 = w24447 & w24637 ;
  assign w24722 = ~w24455 & w24589 ;
  assign w24723 = w24590 ^ w24722 ;
  assign w24724 = ~w24637 & w24723 ;
  assign w24725 = w24721 | w24724 ;
  assign w24726 = ~\pi081 & w24725 ;
  assign w24727 = w24454 & w24637 ;
  assign w24728 = ~w24462 & w24586 ;
  assign w24729 = w24587 ^ w24728 ;
  assign w24730 = ~w24637 & w24729 ;
  assign w24731 = w24727 | w24730 ;
  assign w24732 = ~\pi080 & w24731 ;
  assign w24733 = w24461 & w24637 ;
  assign w24734 = ~w24469 & w24583 ;
  assign w24735 = w24584 ^ w24734 ;
  assign w24736 = ~w24637 & w24735 ;
  assign w24737 = w24733 | w24736 ;
  assign w24738 = ~\pi079 & w24737 ;
  assign w24739 = w24468 & w24637 ;
  assign w24740 = ~w24476 & w24580 ;
  assign w24741 = w24581 ^ w24740 ;
  assign w24742 = ~w24637 & w24741 ;
  assign w24743 = w24739 | w24742 ;
  assign w24744 = ~\pi078 & w24743 ;
  assign w24745 = w24475 & w24637 ;
  assign w24746 = ~w24483 & w24577 ;
  assign w24747 = w24578 ^ w24746 ;
  assign w24748 = ~w24637 & w24747 ;
  assign w24749 = w24745 | w24748 ;
  assign w24750 = ~\pi077 & w24749 ;
  assign w24751 = w24482 & w24637 ;
  assign w24752 = ~w24490 & w24574 ;
  assign w24753 = w24575 ^ w24752 ;
  assign w24754 = ~w24637 & w24753 ;
  assign w24755 = w24751 | w24754 ;
  assign w24756 = ~\pi076 & w24755 ;
  assign w24757 = w24489 & w24637 ;
  assign w24758 = ~w24497 & w24571 ;
  assign w24759 = w24572 ^ w24758 ;
  assign w24760 = ~w24637 & w24759 ;
  assign w24761 = w24757 | w24760 ;
  assign w24762 = ~\pi075 & w24761 ;
  assign w24763 = w24496 & w24637 ;
  assign w24764 = ~w24504 & w24568 ;
  assign w24765 = w24569 ^ w24764 ;
  assign w24766 = ~w24637 & w24765 ;
  assign w24767 = w24763 | w24766 ;
  assign w24768 = ~\pi074 & w24767 ;
  assign w24769 = w24503 & w24637 ;
  assign w24770 = ~w24511 & w24565 ;
  assign w24771 = w24566 ^ w24770 ;
  assign w24772 = ~w24637 & w24771 ;
  assign w24773 = w24769 | w24772 ;
  assign w24774 = ~\pi073 & w24773 ;
  assign w24775 = w24510 & w24637 ;
  assign w24776 = ~w24518 & w24562 ;
  assign w24777 = w24563 ^ w24776 ;
  assign w24778 = ~w24637 & w24777 ;
  assign w24779 = w24775 | w24778 ;
  assign w24780 = ~\pi072 & w24779 ;
  assign w24781 = w24517 & w24637 ;
  assign w24782 = ~w24525 & w24559 ;
  assign w24783 = w24560 ^ w24782 ;
  assign w24784 = ~w24637 & w24783 ;
  assign w24785 = w24781 | w24784 ;
  assign w24786 = ~\pi071 & w24785 ;
  assign w24787 = w24524 & w24637 ;
  assign w24788 = ~w24532 & w24556 ;
  assign w24789 = w24557 ^ w24788 ;
  assign w24790 = ~w24637 & w24789 ;
  assign w24791 = w24787 | w24790 ;
  assign w24792 = ~\pi070 & w24791 ;
  assign w24793 = w24531 & w24637 ;
  assign w24794 = ~w24538 & w24553 ;
  assign w24795 = w24554 ^ w24794 ;
  assign w24796 = ~w24637 & w24795 ;
  assign w24797 = w24793 | w24796 ;
  assign w24798 = ~\pi069 & w24797 ;
  assign w24799 = w24537 & w24637 ;
  assign w24800 = ~w24543 & w24550 ;
  assign w24801 = w24551 ^ w24800 ;
  assign w24802 = ~w24637 & w24801 ;
  assign w24803 = w24799 | w24802 ;
  assign w24804 = ~\pi068 & w24803 ;
  assign w24805 = w24542 & w24637 ;
  assign w24806 = \pi064 & ~w24344 ;
  assign w24807 = \pi034 ^ w24806 ;
  assign w24808 = ( \pi065 & w5287 ) | ( \pi065 & ~w24807 ) | ( w5287 & ~w24807 ) ;
  assign w24809 = w24546 ^ w24808 ;
  assign w24810 = ( w5117 & w24636 ) | ( w5117 & w24809 ) | ( w24636 & w24809 ) ;
  assign w24811 = w24809 & ~w24810 ;
  assign w24812 = w24805 | w24811 ;
  assign w24813 = ~\pi067 & w24812 ;
  assign w24814 = \pi033 ^ w24344 ;
  assign w24815 = ( \pi064 & w5117 ) | ( \pi064 & w24814 ) | ( w5117 & w24814 ) ;
  assign w24816 = w5294 ^ w24815 ;
  assign w24817 = ~w5117 & w24816 ;
  assign w24818 = ~w24636 & w24817 ;
  assign w24819 = ( ~\pi064 & w24344 ) | ( ~\pi064 & w24637 ) | ( w24344 & w24637 ) ;
  assign w24820 = \pi034 ^ w24819 ;
  assign w24821 = w24637 & ~w24820 ;
  assign w24822 = w24818 | w24821 ;
  assign w24823 = ~\pi066 & w24822 ;
  assign w24824 = ( \pi033 & ~w5307 ) | ( \pi033 & w24636 ) | ( ~w5307 & w24636 ) ;
  assign w24825 = \pi033 & w24824 ;
  assign w24826 = w5315 & ~w24636 ;
  assign w24827 = w24825 | w24826 ;
  assign w24828 = \pi065 ^ w24827 ;
  assign w24829 = w5318 | w24828 ;
  assign w24830 = w24637 | w24818 ;
  assign w24831 = ( w24807 & w24818 ) | ( w24807 & w24830 ) | ( w24818 & w24830 ) ;
  assign w24832 = \pi066 ^ w24831 ;
  assign w24833 = ~\pi065 & w24827 ;
  assign w24834 = w24829 | w24833 ;
  assign w24835 = ( w24832 & ~w24833 ) | ( w24832 & w24834 ) | ( ~w24833 & w24834 ) ;
  assign w24836 = \pi067 ^ w24812 ;
  assign w24837 = ( ~w24823 & w24835 ) | ( ~w24823 & w24836 ) | ( w24835 & w24836 ) ;
  assign w24838 = w24836 | w24837 ;
  assign w24839 = \pi068 ^ w24803 ;
  assign w24840 = ( ~w24813 & w24838 ) | ( ~w24813 & w24839 ) | ( w24838 & w24839 ) ;
  assign w24841 = w24839 | w24840 ;
  assign w24842 = \pi069 ^ w24797 ;
  assign w24843 = ( ~w24804 & w24841 ) | ( ~w24804 & w24842 ) | ( w24841 & w24842 ) ;
  assign w24844 = w24842 | w24843 ;
  assign w24845 = \pi070 ^ w24791 ;
  assign w24846 = ( ~w24798 & w24844 ) | ( ~w24798 & w24845 ) | ( w24844 & w24845 ) ;
  assign w24847 = w24845 | w24846 ;
  assign w24848 = \pi071 ^ w24785 ;
  assign w24849 = ( ~w24792 & w24847 ) | ( ~w24792 & w24848 ) | ( w24847 & w24848 ) ;
  assign w24850 = w24848 | w24849 ;
  assign w24851 = \pi072 ^ w24779 ;
  assign w24852 = ( ~w24786 & w24850 ) | ( ~w24786 & w24851 ) | ( w24850 & w24851 ) ;
  assign w24853 = w24851 | w24852 ;
  assign w24854 = \pi073 ^ w24773 ;
  assign w24855 = ( ~w24780 & w24853 ) | ( ~w24780 & w24854 ) | ( w24853 & w24854 ) ;
  assign w24856 = w24854 | w24855 ;
  assign w24857 = \pi074 ^ w24767 ;
  assign w24858 = ( ~w24774 & w24856 ) | ( ~w24774 & w24857 ) | ( w24856 & w24857 ) ;
  assign w24859 = w24857 | w24858 ;
  assign w24860 = \pi075 ^ w24761 ;
  assign w24861 = ( ~w24768 & w24859 ) | ( ~w24768 & w24860 ) | ( w24859 & w24860 ) ;
  assign w24862 = w24860 | w24861 ;
  assign w24863 = \pi076 ^ w24755 ;
  assign w24864 = ( ~w24762 & w24862 ) | ( ~w24762 & w24863 ) | ( w24862 & w24863 ) ;
  assign w24865 = w24863 | w24864 ;
  assign w24866 = \pi077 ^ w24749 ;
  assign w24867 = ( ~w24756 & w24865 ) | ( ~w24756 & w24866 ) | ( w24865 & w24866 ) ;
  assign w24868 = w24866 | w24867 ;
  assign w24869 = \pi078 ^ w24743 ;
  assign w24870 = ( ~w24750 & w24868 ) | ( ~w24750 & w24869 ) | ( w24868 & w24869 ) ;
  assign w24871 = w24869 | w24870 ;
  assign w24872 = \pi079 ^ w24737 ;
  assign w24873 = ( ~w24744 & w24871 ) | ( ~w24744 & w24872 ) | ( w24871 & w24872 ) ;
  assign w24874 = w24872 | w24873 ;
  assign w24875 = \pi080 ^ w24731 ;
  assign w24876 = ( ~w24738 & w24874 ) | ( ~w24738 & w24875 ) | ( w24874 & w24875 ) ;
  assign w24877 = w24875 | w24876 ;
  assign w24878 = \pi081 ^ w24725 ;
  assign w24879 = ( ~w24732 & w24877 ) | ( ~w24732 & w24878 ) | ( w24877 & w24878 ) ;
  assign w24880 = w24878 | w24879 ;
  assign w24881 = \pi082 ^ w24719 ;
  assign w24882 = ( ~w24726 & w24880 ) | ( ~w24726 & w24881 ) | ( w24880 & w24881 ) ;
  assign w24883 = w24881 | w24882 ;
  assign w24884 = \pi083 ^ w24713 ;
  assign w24885 = ( ~w24720 & w24883 ) | ( ~w24720 & w24884 ) | ( w24883 & w24884 ) ;
  assign w24886 = w24884 | w24885 ;
  assign w24887 = \pi084 ^ w24707 ;
  assign w24888 = ( ~w24714 & w24886 ) | ( ~w24714 & w24887 ) | ( w24886 & w24887 ) ;
  assign w24889 = w24887 | w24888 ;
  assign w24890 = \pi085 ^ w24701 ;
  assign w24891 = ( ~w24708 & w24889 ) | ( ~w24708 & w24890 ) | ( w24889 & w24890 ) ;
  assign w24892 = w24890 | w24891 ;
  assign w24893 = \pi086 ^ w24695 ;
  assign w24894 = ( ~w24702 & w24892 ) | ( ~w24702 & w24893 ) | ( w24892 & w24893 ) ;
  assign w24895 = w24893 | w24894 ;
  assign w24896 = \pi087 ^ w24689 ;
  assign w24897 = ( ~w24696 & w24895 ) | ( ~w24696 & w24896 ) | ( w24895 & w24896 ) ;
  assign w24898 = w24896 | w24897 ;
  assign w24899 = \pi088 ^ w24683 ;
  assign w24900 = ( ~w24690 & w24898 ) | ( ~w24690 & w24899 ) | ( w24898 & w24899 ) ;
  assign w24901 = w24899 | w24900 ;
  assign w24902 = \pi089 ^ w24677 ;
  assign w24903 = ( ~w24684 & w24901 ) | ( ~w24684 & w24902 ) | ( w24901 & w24902 ) ;
  assign w24904 = w24902 | w24903 ;
  assign w24905 = \pi090 ^ w24671 ;
  assign w24906 = ( ~w24678 & w24904 ) | ( ~w24678 & w24905 ) | ( w24904 & w24905 ) ;
  assign w24907 = w24905 | w24906 ;
  assign w24908 = \pi091 ^ w24665 ;
  assign w24909 = ( ~w24672 & w24907 ) | ( ~w24672 & w24908 ) | ( w24907 & w24908 ) ;
  assign w24910 = w24908 | w24909 ;
  assign w24911 = \pi092 ^ w24659 ;
  assign w24912 = ( ~w24666 & w24910 ) | ( ~w24666 & w24911 ) | ( w24910 & w24911 ) ;
  assign w24913 = w24911 | w24912 ;
  assign w24914 = \pi093 ^ w24653 ;
  assign w24915 = ( ~w24660 & w24913 ) | ( ~w24660 & w24914 ) | ( w24913 & w24914 ) ;
  assign w24916 = w24914 | w24915 ;
  assign w24917 = \pi094 ^ w24642 ;
  assign w24918 = ( ~w24654 & w24916 ) | ( ~w24654 & w24917 ) | ( w24916 & w24917 ) ;
  assign w24919 = w24917 | w24918 ;
  assign w24920 = \pi095 ^ w24647 ;
  assign w24921 = w24648 & ~w24920 ;
  assign w24922 = ( w24919 & w24920 ) | ( w24919 & ~w24921 ) | ( w24920 & ~w24921 ) ;
  assign w24923 = ~\pi095 & w24647 ;
  assign w24924 = w24922 & ~w24923 ;
  assign w24925 = w298 | w24924 ;
  assign w24926 = w24642 & w24925 ;
  assign w24927 = ~w24654 & w24916 ;
  assign w24928 = w24917 ^ w24927 ;
  assign w24929 = ~w24925 & w24928 ;
  assign w24930 = w24926 | w24929 ;
  assign w24931 = ~\pi095 & w24930 ;
  assign w24932 = w24653 & w24925 ;
  assign w24933 = ~w24660 & w24913 ;
  assign w24934 = w24914 ^ w24933 ;
  assign w24935 = ~w24925 & w24934 ;
  assign w24936 = w24932 | w24935 ;
  assign w24937 = ~\pi094 & w24936 ;
  assign w24938 = w24659 & w24925 ;
  assign w24939 = ~w24666 & w24910 ;
  assign w24940 = w24911 ^ w24939 ;
  assign w24941 = ~w24925 & w24940 ;
  assign w24942 = w24938 | w24941 ;
  assign w24943 = ~\pi093 & w24942 ;
  assign w24944 = w24665 & w24925 ;
  assign w24945 = ~w24672 & w24907 ;
  assign w24946 = w24908 ^ w24945 ;
  assign w24947 = ~w24925 & w24946 ;
  assign w24948 = w24944 | w24947 ;
  assign w24949 = ~\pi092 & w24948 ;
  assign w24950 = w24671 & w24925 ;
  assign w24951 = ~w24678 & w24904 ;
  assign w24952 = w24905 ^ w24951 ;
  assign w24953 = ~w24925 & w24952 ;
  assign w24954 = w24950 | w24953 ;
  assign w24955 = ~\pi091 & w24954 ;
  assign w24956 = w24677 & w24925 ;
  assign w24957 = ~w24684 & w24901 ;
  assign w24958 = w24902 ^ w24957 ;
  assign w24959 = ~w24925 & w24958 ;
  assign w24960 = w24956 | w24959 ;
  assign w24961 = ~\pi090 & w24960 ;
  assign w24962 = w24683 & w24925 ;
  assign w24963 = ~w24690 & w24898 ;
  assign w24964 = w24899 ^ w24963 ;
  assign w24965 = ~w24925 & w24964 ;
  assign w24966 = w24962 | w24965 ;
  assign w24967 = ~\pi089 & w24966 ;
  assign w24968 = w24689 & w24925 ;
  assign w24969 = ~w24696 & w24895 ;
  assign w24970 = w24896 ^ w24969 ;
  assign w24971 = ~w24925 & w24970 ;
  assign w24972 = w24968 | w24971 ;
  assign w24973 = ~\pi088 & w24972 ;
  assign w24974 = w24695 & w24925 ;
  assign w24975 = ~w24702 & w24892 ;
  assign w24976 = w24893 ^ w24975 ;
  assign w24977 = ~w24925 & w24976 ;
  assign w24978 = w24974 | w24977 ;
  assign w24979 = ~\pi087 & w24978 ;
  assign w24980 = w24701 & w24925 ;
  assign w24981 = ~w24708 & w24889 ;
  assign w24982 = w24890 ^ w24981 ;
  assign w24983 = ~w24925 & w24982 ;
  assign w24984 = w24980 | w24983 ;
  assign w24985 = ~\pi086 & w24984 ;
  assign w24986 = w24707 & w24925 ;
  assign w24987 = ~w24714 & w24886 ;
  assign w24988 = w24887 ^ w24987 ;
  assign w24989 = ~w24925 & w24988 ;
  assign w24990 = w24986 | w24989 ;
  assign w24991 = ~\pi085 & w24990 ;
  assign w24992 = w24713 & w24925 ;
  assign w24993 = ~w24720 & w24883 ;
  assign w24994 = w24884 ^ w24993 ;
  assign w24995 = ~w24925 & w24994 ;
  assign w24996 = w24992 | w24995 ;
  assign w24997 = ~\pi084 & w24996 ;
  assign w24998 = w24719 & w24925 ;
  assign w24999 = ~w24726 & w24880 ;
  assign w25000 = w24881 ^ w24999 ;
  assign w25001 = ~w24925 & w25000 ;
  assign w25002 = w24998 | w25001 ;
  assign w25003 = ~\pi083 & w25002 ;
  assign w25004 = w24725 & w24925 ;
  assign w25005 = ~w24732 & w24877 ;
  assign w25006 = w24878 ^ w25005 ;
  assign w25007 = ~w24925 & w25006 ;
  assign w25008 = w25004 | w25007 ;
  assign w25009 = ~\pi082 & w25008 ;
  assign w25010 = w24731 & w24925 ;
  assign w25011 = ~w24738 & w24874 ;
  assign w25012 = w24875 ^ w25011 ;
  assign w25013 = ~w24925 & w25012 ;
  assign w25014 = w25010 | w25013 ;
  assign w25015 = ~\pi081 & w25014 ;
  assign w25016 = w24737 & w24925 ;
  assign w25017 = ~w24744 & w24871 ;
  assign w25018 = w24872 ^ w25017 ;
  assign w25019 = ~w24925 & w25018 ;
  assign w25020 = w25016 | w25019 ;
  assign w25021 = ~\pi080 & w25020 ;
  assign w25022 = w24743 & w24925 ;
  assign w25023 = ~w24750 & w24868 ;
  assign w25024 = w24869 ^ w25023 ;
  assign w25025 = ~w24925 & w25024 ;
  assign w25026 = w25022 | w25025 ;
  assign w25027 = ~\pi079 & w25026 ;
  assign w25028 = w24749 & w24925 ;
  assign w25029 = ~w24756 & w24865 ;
  assign w25030 = w24866 ^ w25029 ;
  assign w25031 = ~w24925 & w25030 ;
  assign w25032 = w25028 | w25031 ;
  assign w25033 = ~\pi078 & w25032 ;
  assign w25034 = w24755 & w24925 ;
  assign w25035 = ~w24762 & w24862 ;
  assign w25036 = w24863 ^ w25035 ;
  assign w25037 = ~w24925 & w25036 ;
  assign w25038 = w25034 | w25037 ;
  assign w25039 = ~\pi077 & w25038 ;
  assign w25040 = w24761 & w24925 ;
  assign w25041 = ~w24768 & w24859 ;
  assign w25042 = w24860 ^ w25041 ;
  assign w25043 = ~w24925 & w25042 ;
  assign w25044 = w25040 | w25043 ;
  assign w25045 = ~\pi076 & w25044 ;
  assign w25046 = w24767 & w24925 ;
  assign w25047 = ~w24774 & w24856 ;
  assign w25048 = w24857 ^ w25047 ;
  assign w25049 = ~w24925 & w25048 ;
  assign w25050 = w25046 | w25049 ;
  assign w25051 = ~\pi075 & w25050 ;
  assign w25052 = w24773 & w24925 ;
  assign w25053 = ~w24780 & w24853 ;
  assign w25054 = w24854 ^ w25053 ;
  assign w25055 = ~w24925 & w25054 ;
  assign w25056 = w25052 | w25055 ;
  assign w25057 = ~\pi074 & w25056 ;
  assign w25058 = w24779 & w24925 ;
  assign w25059 = ~w24786 & w24850 ;
  assign w25060 = w24851 ^ w25059 ;
  assign w25061 = ~w24925 & w25060 ;
  assign w25062 = w25058 | w25061 ;
  assign w25063 = ~\pi073 & w25062 ;
  assign w25064 = w24785 & w24925 ;
  assign w25065 = ~w24792 & w24847 ;
  assign w25066 = w24848 ^ w25065 ;
  assign w25067 = ~w24925 & w25066 ;
  assign w25068 = w25064 | w25067 ;
  assign w25069 = ~\pi072 & w25068 ;
  assign w25070 = w24791 & w24925 ;
  assign w25071 = ~w24798 & w24844 ;
  assign w25072 = w24845 ^ w25071 ;
  assign w25073 = ~w24925 & w25072 ;
  assign w25074 = w25070 | w25073 ;
  assign w25075 = ~\pi071 & w25074 ;
  assign w25076 = w24797 & w24925 ;
  assign w25077 = ~w24804 & w24841 ;
  assign w25078 = w24842 ^ w25077 ;
  assign w25079 = ~w24925 & w25078 ;
  assign w25080 = w25076 | w25079 ;
  assign w25081 = ~\pi070 & w25080 ;
  assign w25082 = w24803 & w24925 ;
  assign w25083 = ~w24813 & w24838 ;
  assign w25084 = w24839 ^ w25083 ;
  assign w25085 = ~w24925 & w25084 ;
  assign w25086 = w25082 | w25085 ;
  assign w25087 = ~\pi069 & w25086 ;
  assign w25088 = w24812 & w24925 ;
  assign w25089 = ~w24823 & w24835 ;
  assign w25090 = w24836 ^ w25089 ;
  assign w25091 = ~w24925 & w25090 ;
  assign w25092 = w25088 | w25091 ;
  assign w25093 = ~\pi068 & w25092 ;
  assign w25094 = w24822 & w24925 ;
  assign w25095 = ~w24827 & w24829 ;
  assign w25096 = ( \pi065 & w24829 ) | ( \pi065 & w25095 ) | ( w24829 & w25095 ) ;
  assign w25097 = w24832 ^ w25096 ;
  assign w25098 = ~w24925 & w25097 ;
  assign w25099 = w25094 | w25098 ;
  assign w25100 = ~\pi067 & w25099 ;
  assign w25101 = ( ~w298 & w24825 ) | ( ~w298 & w24826 ) | ( w24825 & w24826 ) ;
  assign w25102 = \pi065 ^ w25101 ;
  assign w25103 = ( ~w298 & w5318 ) | ( ~w298 & w25102 ) | ( w5318 & w25102 ) ;
  assign w25104 = ( w5318 & w24924 ) | ( w5318 & w25102 ) | ( w24924 & w25102 ) ;
  assign w25105 = w25103 & ~w25104 ;
  assign w25106 = ( w24827 & w24925 ) | ( w24827 & w25105 ) | ( w24925 & w25105 ) ;
  assign w25107 = w25105 | w25106 ;
  assign w25108 = ~\pi066 & w25107 ;
  assign w25109 = ( \pi032 & ~w5602 ) | ( \pi032 & w24924 ) | ( ~w5602 & w24924 ) ;
  assign w25110 = \pi032 & w25109 ;
  assign w25111 = ( w155 & ~w170 ) | ( w155 & w24924 ) | ( ~w170 & w24924 ) ;
  assign w25112 = w5606 & ~w25111 ;
  assign w25113 = ~w24827 & w24925 ;
  assign w25114 = ( w24925 & w25105 ) | ( w24925 & ~w25113 ) | ( w25105 & ~w25113 ) ;
  assign w25115 = \pi066 ^ w25114 ;
  assign w25116 = w25110 | w25112 ;
  assign w25117 = ( \pi065 & w5609 ) | ( \pi065 & ~w25116 ) | ( w5609 & ~w25116 ) ;
  assign w25118 = w25115 | w25117 ;
  assign w25119 = \pi067 ^ w25099 ;
  assign w25120 = ( ~w25108 & w25118 ) | ( ~w25108 & w25119 ) | ( w25118 & w25119 ) ;
  assign w25121 = w25119 | w25120 ;
  assign w25122 = \pi068 ^ w25092 ;
  assign w25123 = ( ~w25100 & w25121 ) | ( ~w25100 & w25122 ) | ( w25121 & w25122 ) ;
  assign w25124 = w25122 | w25123 ;
  assign w25125 = \pi069 ^ w25086 ;
  assign w25126 = ( ~w25093 & w25124 ) | ( ~w25093 & w25125 ) | ( w25124 & w25125 ) ;
  assign w25127 = w25125 | w25126 ;
  assign w25128 = \pi070 ^ w25080 ;
  assign w25129 = ( ~w25087 & w25127 ) | ( ~w25087 & w25128 ) | ( w25127 & w25128 ) ;
  assign w25130 = w25128 | w25129 ;
  assign w25131 = \pi071 ^ w25074 ;
  assign w25132 = ( ~w25081 & w25130 ) | ( ~w25081 & w25131 ) | ( w25130 & w25131 ) ;
  assign w25133 = w25131 | w25132 ;
  assign w25134 = \pi072 ^ w25068 ;
  assign w25135 = ( ~w25075 & w25133 ) | ( ~w25075 & w25134 ) | ( w25133 & w25134 ) ;
  assign w25136 = w25134 | w25135 ;
  assign w25137 = \pi073 ^ w25062 ;
  assign w25138 = ( ~w25069 & w25136 ) | ( ~w25069 & w25137 ) | ( w25136 & w25137 ) ;
  assign w25139 = w25137 | w25138 ;
  assign w25140 = \pi074 ^ w25056 ;
  assign w25141 = ( ~w25063 & w25139 ) | ( ~w25063 & w25140 ) | ( w25139 & w25140 ) ;
  assign w25142 = w25140 | w25141 ;
  assign w25143 = \pi075 ^ w25050 ;
  assign w25144 = ( ~w25057 & w25142 ) | ( ~w25057 & w25143 ) | ( w25142 & w25143 ) ;
  assign w25145 = w25143 | w25144 ;
  assign w25146 = \pi076 ^ w25044 ;
  assign w25147 = ( ~w25051 & w25145 ) | ( ~w25051 & w25146 ) | ( w25145 & w25146 ) ;
  assign w25148 = w25146 | w25147 ;
  assign w25149 = \pi077 ^ w25038 ;
  assign w25150 = ( ~w25045 & w25148 ) | ( ~w25045 & w25149 ) | ( w25148 & w25149 ) ;
  assign w25151 = w25149 | w25150 ;
  assign w25152 = \pi078 ^ w25032 ;
  assign w25153 = ( ~w25039 & w25151 ) | ( ~w25039 & w25152 ) | ( w25151 & w25152 ) ;
  assign w25154 = w25152 | w25153 ;
  assign w25155 = \pi079 ^ w25026 ;
  assign w25156 = ( ~w25033 & w25154 ) | ( ~w25033 & w25155 ) | ( w25154 & w25155 ) ;
  assign w25157 = w25155 | w25156 ;
  assign w25158 = \pi080 ^ w25020 ;
  assign w25159 = ( ~w25027 & w25157 ) | ( ~w25027 & w25158 ) | ( w25157 & w25158 ) ;
  assign w25160 = w25158 | w25159 ;
  assign w25161 = \pi081 ^ w25014 ;
  assign w25162 = ( ~w25021 & w25160 ) | ( ~w25021 & w25161 ) | ( w25160 & w25161 ) ;
  assign w25163 = w25161 | w25162 ;
  assign w25164 = \pi082 ^ w25008 ;
  assign w25165 = ( ~w25015 & w25163 ) | ( ~w25015 & w25164 ) | ( w25163 & w25164 ) ;
  assign w25166 = w25164 | w25165 ;
  assign w25167 = \pi083 ^ w25002 ;
  assign w25168 = ( ~w25009 & w25166 ) | ( ~w25009 & w25167 ) | ( w25166 & w25167 ) ;
  assign w25169 = w25167 | w25168 ;
  assign w25170 = \pi084 ^ w24996 ;
  assign w25171 = ( ~w25003 & w25169 ) | ( ~w25003 & w25170 ) | ( w25169 & w25170 ) ;
  assign w25172 = w25170 | w25171 ;
  assign w25173 = \pi085 ^ w24990 ;
  assign w25174 = ( ~w24997 & w25172 ) | ( ~w24997 & w25173 ) | ( w25172 & w25173 ) ;
  assign w25175 = w25173 | w25174 ;
  assign w25176 = \pi086 ^ w24984 ;
  assign w25177 = ( ~w24991 & w25175 ) | ( ~w24991 & w25176 ) | ( w25175 & w25176 ) ;
  assign w25178 = w25176 | w25177 ;
  assign w25179 = \pi087 ^ w24978 ;
  assign w25180 = ( ~w24985 & w25178 ) | ( ~w24985 & w25179 ) | ( w25178 & w25179 ) ;
  assign w25181 = w25179 | w25180 ;
  assign w25182 = \pi088 ^ w24972 ;
  assign w25183 = ( ~w24979 & w25181 ) | ( ~w24979 & w25182 ) | ( w25181 & w25182 ) ;
  assign w25184 = w25182 | w25183 ;
  assign w25185 = \pi089 ^ w24966 ;
  assign w25186 = ( ~w24973 & w25184 ) | ( ~w24973 & w25185 ) | ( w25184 & w25185 ) ;
  assign w25187 = w25185 | w25186 ;
  assign w25188 = \pi090 ^ w24960 ;
  assign w25189 = ( ~w24967 & w25187 ) | ( ~w24967 & w25188 ) | ( w25187 & w25188 ) ;
  assign w25190 = w25188 | w25189 ;
  assign w25191 = \pi091 ^ w24954 ;
  assign w25192 = ( ~w24961 & w25190 ) | ( ~w24961 & w25191 ) | ( w25190 & w25191 ) ;
  assign w25193 = w25191 | w25192 ;
  assign w25194 = \pi092 ^ w24948 ;
  assign w25195 = ( ~w24955 & w25193 ) | ( ~w24955 & w25194 ) | ( w25193 & w25194 ) ;
  assign w25196 = w25194 | w25195 ;
  assign w25197 = \pi093 ^ w24942 ;
  assign w25198 = ( ~w24949 & w25196 ) | ( ~w24949 & w25197 ) | ( w25196 & w25197 ) ;
  assign w25199 = w25197 | w25198 ;
  assign w25200 = \pi094 ^ w24936 ;
  assign w25201 = ( ~w24943 & w25199 ) | ( ~w24943 & w25200 ) | ( w25199 & w25200 ) ;
  assign w25202 = w25200 | w25201 ;
  assign w25203 = \pi095 ^ w24930 ;
  assign w25204 = ( ~w24937 & w25202 ) | ( ~w24937 & w25203 ) | ( w25202 & w25203 ) ;
  assign w25205 = w25203 | w25204 ;
  assign w25206 = w24647 & w24925 ;
  assign w25207 = ~w24648 & w24919 ;
  assign w25208 = w24920 ^ w25207 ;
  assign w25209 = ~w24925 & w25208 ;
  assign w25210 = w25206 | w25209 ;
  assign w25211 = ~\pi096 & w25210 ;
  assign w25212 = ( \pi096 & ~w25206 ) | ( \pi096 & w25209 ) | ( ~w25206 & w25209 ) ;
  assign w25213 = ~w25209 & w25212 ;
  assign w25214 = w25211 | w25213 ;
  assign w25215 = ( ~w24931 & w25205 ) | ( ~w24931 & w25214 ) | ( w25205 & w25214 ) ;
  assign w25216 = ( w291 & ~w25214 ) | ( w291 & w25215 ) | ( ~w25214 & w25215 ) ;
  assign w25217 = w25214 | w25216 ;
  assign w25218 = ~w298 & w25210 ;
  assign w25219 = w25217 & ~w25218 ;
  assign w25220 = ~w24937 & w25202 ;
  assign w25221 = w25203 ^ w25220 ;
  assign w25222 = ~w25219 & w25221 ;
  assign w25223 = ( w24930 & w25217 ) | ( w24930 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25224 = ~w25218 & w25223 ;
  assign w25225 = w25222 | w25224 ;
  assign w25226 = ( ~w24931 & w25205 ) | ( ~w24931 & w25219 ) | ( w25205 & w25219 ) ;
  assign w25227 = w25214 ^ w25226 ;
  assign w25228 = ~w25219 & w25227 ;
  assign w25229 = ( w298 & ~w25210 ) | ( w298 & w25217 ) | ( ~w25210 & w25217 ) ;
  assign w25230 = w25210 & w25229 ;
  assign w25231 = w25228 | w25230 ;
  assign w25232 = ~\pi096 & w25225 ;
  assign w25233 = ~w24943 & w25199 ;
  assign w25234 = w25200 ^ w25233 ;
  assign w25235 = ~w25219 & w25234 ;
  assign w25236 = ( w24936 & w25217 ) | ( w24936 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25237 = ~w25218 & w25236 ;
  assign w25238 = w25235 | w25237 ;
  assign w25239 = ~\pi095 & w25238 ;
  assign w25240 = ~w24949 & w25196 ;
  assign w25241 = w25197 ^ w25240 ;
  assign w25242 = ~w25219 & w25241 ;
  assign w25243 = ( w24942 & w25217 ) | ( w24942 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25244 = ~w25218 & w25243 ;
  assign w25245 = w25242 | w25244 ;
  assign w25246 = ~\pi094 & w25245 ;
  assign w25247 = ~w24955 & w25193 ;
  assign w25248 = w25194 ^ w25247 ;
  assign w25249 = ~w25219 & w25248 ;
  assign w25250 = ( w24948 & w25217 ) | ( w24948 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25251 = ~w25218 & w25250 ;
  assign w25252 = w25249 | w25251 ;
  assign w25253 = ~\pi093 & w25252 ;
  assign w25254 = ~w24961 & w25190 ;
  assign w25255 = w25191 ^ w25254 ;
  assign w25256 = ~w25219 & w25255 ;
  assign w25257 = ( w24954 & w25217 ) | ( w24954 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25258 = ~w25218 & w25257 ;
  assign w25259 = w25256 | w25258 ;
  assign w25260 = ~\pi092 & w25259 ;
  assign w25261 = ~w24967 & w25187 ;
  assign w25262 = w25188 ^ w25261 ;
  assign w25263 = ~w25219 & w25262 ;
  assign w25264 = ( w24960 & w25217 ) | ( w24960 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25265 = ~w25218 & w25264 ;
  assign w25266 = w25263 | w25265 ;
  assign w25267 = ~\pi091 & w25266 ;
  assign w25268 = ~w24973 & w25184 ;
  assign w25269 = w25185 ^ w25268 ;
  assign w25270 = ~w25219 & w25269 ;
  assign w25271 = ( w24966 & w25217 ) | ( w24966 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25272 = ~w25218 & w25271 ;
  assign w25273 = w25270 | w25272 ;
  assign w25274 = ~\pi090 & w25273 ;
  assign w25275 = ~w24979 & w25181 ;
  assign w25276 = w25182 ^ w25275 ;
  assign w25277 = ~w25219 & w25276 ;
  assign w25278 = ( w24972 & w25217 ) | ( w24972 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25279 = ~w25218 & w25278 ;
  assign w25280 = w25277 | w25279 ;
  assign w25281 = ~\pi089 & w25280 ;
  assign w25282 = ~w24985 & w25178 ;
  assign w25283 = w25179 ^ w25282 ;
  assign w25284 = ~w25219 & w25283 ;
  assign w25285 = ( w24978 & w25217 ) | ( w24978 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25286 = ~w25218 & w25285 ;
  assign w25287 = w25284 | w25286 ;
  assign w25288 = ~\pi088 & w25287 ;
  assign w25289 = ~w24991 & w25175 ;
  assign w25290 = w25176 ^ w25289 ;
  assign w25291 = ~w25219 & w25290 ;
  assign w25292 = ( w24984 & w25217 ) | ( w24984 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25293 = ~w25218 & w25292 ;
  assign w25294 = w25291 | w25293 ;
  assign w25295 = ~\pi087 & w25294 ;
  assign w25296 = ~w24997 & w25172 ;
  assign w25297 = w25173 ^ w25296 ;
  assign w25298 = ~w25219 & w25297 ;
  assign w25299 = ( w24990 & w25217 ) | ( w24990 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25300 = ~w25218 & w25299 ;
  assign w25301 = w25298 | w25300 ;
  assign w25302 = ~\pi086 & w25301 ;
  assign w25303 = ~w25003 & w25169 ;
  assign w25304 = w25170 ^ w25303 ;
  assign w25305 = ~w25219 & w25304 ;
  assign w25306 = ( w24996 & w25217 ) | ( w24996 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25307 = ~w25218 & w25306 ;
  assign w25308 = w25305 | w25307 ;
  assign w25309 = ~\pi085 & w25308 ;
  assign w25310 = ~w25009 & w25166 ;
  assign w25311 = w25167 ^ w25310 ;
  assign w25312 = ~w25219 & w25311 ;
  assign w25313 = ( w25002 & w25217 ) | ( w25002 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25314 = ~w25218 & w25313 ;
  assign w25315 = w25312 | w25314 ;
  assign w25316 = ~\pi084 & w25315 ;
  assign w25317 = ~w25015 & w25163 ;
  assign w25318 = w25164 ^ w25317 ;
  assign w25319 = ~w25219 & w25318 ;
  assign w25320 = ( w25008 & w25217 ) | ( w25008 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25321 = ~w25218 & w25320 ;
  assign w25322 = w25319 | w25321 ;
  assign w25323 = ~\pi083 & w25322 ;
  assign w25324 = ~w25021 & w25160 ;
  assign w25325 = w25161 ^ w25324 ;
  assign w25326 = ~w25219 & w25325 ;
  assign w25327 = ( w25014 & w25217 ) | ( w25014 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25328 = ~w25218 & w25327 ;
  assign w25329 = w25326 | w25328 ;
  assign w25330 = ~\pi082 & w25329 ;
  assign w25331 = ~w25027 & w25157 ;
  assign w25332 = w25158 ^ w25331 ;
  assign w25333 = ~w25219 & w25332 ;
  assign w25334 = ( w25020 & w25217 ) | ( w25020 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25335 = ~w25218 & w25334 ;
  assign w25336 = w25333 | w25335 ;
  assign w25337 = ~\pi081 & w25336 ;
  assign w25338 = ~w25033 & w25154 ;
  assign w25339 = w25155 ^ w25338 ;
  assign w25340 = ~w25219 & w25339 ;
  assign w25341 = ( w25026 & w25217 ) | ( w25026 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25342 = ~w25218 & w25341 ;
  assign w25343 = w25340 | w25342 ;
  assign w25344 = ~\pi080 & w25343 ;
  assign w25345 = ~w25039 & w25151 ;
  assign w25346 = w25152 ^ w25345 ;
  assign w25347 = ~w25219 & w25346 ;
  assign w25348 = ( w25032 & w25217 ) | ( w25032 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25349 = ~w25218 & w25348 ;
  assign w25350 = w25347 | w25349 ;
  assign w25351 = ~\pi079 & w25350 ;
  assign w25352 = ~w25045 & w25148 ;
  assign w25353 = w25149 ^ w25352 ;
  assign w25354 = ~w25219 & w25353 ;
  assign w25355 = ( w25038 & w25217 ) | ( w25038 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25356 = ~w25218 & w25355 ;
  assign w25357 = w25354 | w25356 ;
  assign w25358 = ~\pi078 & w25357 ;
  assign w25359 = ~w25051 & w25145 ;
  assign w25360 = w25146 ^ w25359 ;
  assign w25361 = ~w25219 & w25360 ;
  assign w25362 = ( w25044 & w25217 ) | ( w25044 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25363 = ~w25218 & w25362 ;
  assign w25364 = w25361 | w25363 ;
  assign w25365 = ~\pi077 & w25364 ;
  assign w25366 = ~w25057 & w25142 ;
  assign w25367 = w25143 ^ w25366 ;
  assign w25368 = ~w25219 & w25367 ;
  assign w25369 = ( w25050 & w25217 ) | ( w25050 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25370 = ~w25218 & w25369 ;
  assign w25371 = w25368 | w25370 ;
  assign w25372 = ~\pi076 & w25371 ;
  assign w25373 = ~w25063 & w25139 ;
  assign w25374 = w25140 ^ w25373 ;
  assign w25375 = ~w25219 & w25374 ;
  assign w25376 = ( w25056 & w25217 ) | ( w25056 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25377 = ~w25218 & w25376 ;
  assign w25378 = w25375 | w25377 ;
  assign w25379 = ~\pi075 & w25378 ;
  assign w25380 = ~w25069 & w25136 ;
  assign w25381 = w25137 ^ w25380 ;
  assign w25382 = ~w25219 & w25381 ;
  assign w25383 = ( w25062 & w25217 ) | ( w25062 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25384 = ~w25218 & w25383 ;
  assign w25385 = w25382 | w25384 ;
  assign w25386 = ~\pi074 & w25385 ;
  assign w25387 = ~w25075 & w25133 ;
  assign w25388 = w25134 ^ w25387 ;
  assign w25389 = ~w25219 & w25388 ;
  assign w25390 = ( w25068 & w25217 ) | ( w25068 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25391 = ~w25218 & w25390 ;
  assign w25392 = w25389 | w25391 ;
  assign w25393 = ~\pi073 & w25392 ;
  assign w25394 = ~w25081 & w25130 ;
  assign w25395 = w25131 ^ w25394 ;
  assign w25396 = ~w25219 & w25395 ;
  assign w25397 = ( w25074 & w25217 ) | ( w25074 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25398 = ~w25218 & w25397 ;
  assign w25399 = w25396 | w25398 ;
  assign w25400 = ~\pi072 & w25399 ;
  assign w25401 = ~w25087 & w25127 ;
  assign w25402 = w25128 ^ w25401 ;
  assign w25403 = ~w25219 & w25402 ;
  assign w25404 = ( w25080 & w25217 ) | ( w25080 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25405 = ~w25218 & w25404 ;
  assign w25406 = w25403 | w25405 ;
  assign w25407 = ~\pi071 & w25406 ;
  assign w25408 = ~w25093 & w25124 ;
  assign w25409 = w25125 ^ w25408 ;
  assign w25410 = ~w25219 & w25409 ;
  assign w25411 = ( w25086 & w25217 ) | ( w25086 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25412 = ~w25218 & w25411 ;
  assign w25413 = w25410 | w25412 ;
  assign w25414 = ~\pi070 & w25413 ;
  assign w25415 = ~w25100 & w25121 ;
  assign w25416 = w25122 ^ w25415 ;
  assign w25417 = ~w25219 & w25416 ;
  assign w25418 = ( w25092 & w25217 ) | ( w25092 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25419 = ~w25218 & w25418 ;
  assign w25420 = w25417 | w25419 ;
  assign w25421 = ~\pi069 & w25420 ;
  assign w25422 = ~w25108 & w25118 ;
  assign w25423 = w25119 ^ w25422 ;
  assign w25424 = ~w25219 & w25423 ;
  assign w25425 = ( w25099 & w25217 ) | ( w25099 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25426 = ~w25218 & w25425 ;
  assign w25427 = w25424 | w25426 ;
  assign w25428 = ~\pi068 & w25427 ;
  assign w25429 = w25115 ^ w25117 ;
  assign w25430 = ~w25219 & w25429 ;
  assign w25431 = ( w25107 & w25217 ) | ( w25107 & w25218 ) | ( w25217 & w25218 ) ;
  assign w25432 = ~w25218 & w25431 ;
  assign w25433 = w25430 | w25432 ;
  assign w25434 = ~\pi067 & w25433 ;
  assign w25435 = w5609 ^ w25116 ;
  assign w25436 = \pi065 ^ w25435 ;
  assign w25437 = w25219 ^ w25436 ;
  assign w25438 = ( w25116 & w25436 ) | ( w25116 & w25437 ) | ( w25436 & w25437 ) ;
  assign w25439 = ~\pi066 & w25438 ;
  assign w25440 = w25116 ^ w25219 ;
  assign w25441 = ( w25116 & w25436 ) | ( w25116 & ~w25440 ) | ( w25436 & ~w25440 ) ;
  assign w25442 = \pi066 ^ w25441 ;
  assign w25443 = ( \pi064 & ~w25219 ) | ( \pi064 & w25442 ) | ( ~w25219 & w25442 ) ;
  assign w25444 = \pi031 ^ w25443 ;
  assign w25445 = ( \pi065 & w6235 ) | ( \pi065 & ~w25444 ) | ( w6235 & ~w25444 ) ;
  assign w25446 = w25442 | w25445 ;
  assign w25447 = \pi067 ^ w25433 ;
  assign w25448 = ( ~w25439 & w25446 ) | ( ~w25439 & w25447 ) | ( w25446 & w25447 ) ;
  assign w25449 = w25447 | w25448 ;
  assign w25450 = \pi068 ^ w25427 ;
  assign w25451 = ( ~w25434 & w25449 ) | ( ~w25434 & w25450 ) | ( w25449 & w25450 ) ;
  assign w25452 = w25450 | w25451 ;
  assign w25453 = \pi069 ^ w25420 ;
  assign w25454 = ( ~w25428 & w25452 ) | ( ~w25428 & w25453 ) | ( w25452 & w25453 ) ;
  assign w25455 = w25453 | w25454 ;
  assign w25456 = \pi070 ^ w25413 ;
  assign w25457 = ( ~w25421 & w25455 ) | ( ~w25421 & w25456 ) | ( w25455 & w25456 ) ;
  assign w25458 = w25456 | w25457 ;
  assign w25459 = \pi071 ^ w25406 ;
  assign w25460 = ( ~w25414 & w25458 ) | ( ~w25414 & w25459 ) | ( w25458 & w25459 ) ;
  assign w25461 = w25459 | w25460 ;
  assign w25462 = \pi072 ^ w25399 ;
  assign w25463 = ( ~w25407 & w25461 ) | ( ~w25407 & w25462 ) | ( w25461 & w25462 ) ;
  assign w25464 = w25462 | w25463 ;
  assign w25465 = \pi073 ^ w25392 ;
  assign w25466 = ( ~w25400 & w25464 ) | ( ~w25400 & w25465 ) | ( w25464 & w25465 ) ;
  assign w25467 = w25465 | w25466 ;
  assign w25468 = \pi074 ^ w25385 ;
  assign w25469 = ( ~w25393 & w25467 ) | ( ~w25393 & w25468 ) | ( w25467 & w25468 ) ;
  assign w25470 = w25468 | w25469 ;
  assign w25471 = \pi075 ^ w25378 ;
  assign w25472 = ( ~w25386 & w25470 ) | ( ~w25386 & w25471 ) | ( w25470 & w25471 ) ;
  assign w25473 = w25471 | w25472 ;
  assign w25474 = \pi076 ^ w25371 ;
  assign w25475 = ( ~w25379 & w25473 ) | ( ~w25379 & w25474 ) | ( w25473 & w25474 ) ;
  assign w25476 = w25474 | w25475 ;
  assign w25477 = \pi077 ^ w25364 ;
  assign w25478 = ( ~w25372 & w25476 ) | ( ~w25372 & w25477 ) | ( w25476 & w25477 ) ;
  assign w25479 = w25477 | w25478 ;
  assign w25480 = \pi078 ^ w25357 ;
  assign w25481 = ( ~w25365 & w25479 ) | ( ~w25365 & w25480 ) | ( w25479 & w25480 ) ;
  assign w25482 = w25480 | w25481 ;
  assign w25483 = \pi079 ^ w25350 ;
  assign w25484 = ( ~w25358 & w25482 ) | ( ~w25358 & w25483 ) | ( w25482 & w25483 ) ;
  assign w25485 = w25483 | w25484 ;
  assign w25486 = \pi080 ^ w25343 ;
  assign w25487 = ( ~w25351 & w25485 ) | ( ~w25351 & w25486 ) | ( w25485 & w25486 ) ;
  assign w25488 = w25486 | w25487 ;
  assign w25489 = \pi081 ^ w25336 ;
  assign w25490 = ( ~w25344 & w25488 ) | ( ~w25344 & w25489 ) | ( w25488 & w25489 ) ;
  assign w25491 = w25489 | w25490 ;
  assign w25492 = \pi082 ^ w25329 ;
  assign w25493 = ( ~w25337 & w25491 ) | ( ~w25337 & w25492 ) | ( w25491 & w25492 ) ;
  assign w25494 = w25492 | w25493 ;
  assign w25495 = \pi083 ^ w25322 ;
  assign w25496 = ( ~w25330 & w25494 ) | ( ~w25330 & w25495 ) | ( w25494 & w25495 ) ;
  assign w25497 = w25495 | w25496 ;
  assign w25498 = \pi084 ^ w25315 ;
  assign w25499 = ( ~w25323 & w25497 ) | ( ~w25323 & w25498 ) | ( w25497 & w25498 ) ;
  assign w25500 = w25498 | w25499 ;
  assign w25501 = \pi085 ^ w25308 ;
  assign w25502 = ( ~w25316 & w25500 ) | ( ~w25316 & w25501 ) | ( w25500 & w25501 ) ;
  assign w25503 = w25501 | w25502 ;
  assign w25504 = \pi086 ^ w25301 ;
  assign w25505 = ( ~w25309 & w25503 ) | ( ~w25309 & w25504 ) | ( w25503 & w25504 ) ;
  assign w25506 = w25504 | w25505 ;
  assign w25507 = \pi087 ^ w25294 ;
  assign w25508 = ( ~w25302 & w25506 ) | ( ~w25302 & w25507 ) | ( w25506 & w25507 ) ;
  assign w25509 = w25507 | w25508 ;
  assign w25510 = \pi088 ^ w25287 ;
  assign w25511 = ( ~w25295 & w25509 ) | ( ~w25295 & w25510 ) | ( w25509 & w25510 ) ;
  assign w25512 = w25510 | w25511 ;
  assign w25513 = \pi089 ^ w25280 ;
  assign w25514 = ( ~w25288 & w25512 ) | ( ~w25288 & w25513 ) | ( w25512 & w25513 ) ;
  assign w25515 = w25513 | w25514 ;
  assign w25516 = \pi090 ^ w25273 ;
  assign w25517 = ( ~w25281 & w25515 ) | ( ~w25281 & w25516 ) | ( w25515 & w25516 ) ;
  assign w25518 = w25516 | w25517 ;
  assign w25519 = \pi091 ^ w25266 ;
  assign w25520 = ( ~w25274 & w25518 ) | ( ~w25274 & w25519 ) | ( w25518 & w25519 ) ;
  assign w25521 = w25519 | w25520 ;
  assign w25522 = \pi092 ^ w25259 ;
  assign w25523 = ( ~w25267 & w25521 ) | ( ~w25267 & w25522 ) | ( w25521 & w25522 ) ;
  assign w25524 = w25522 | w25523 ;
  assign w25525 = \pi093 ^ w25252 ;
  assign w25526 = ( ~w25260 & w25524 ) | ( ~w25260 & w25525 ) | ( w25524 & w25525 ) ;
  assign w25527 = w25525 | w25526 ;
  assign w25528 = \pi094 ^ w25245 ;
  assign w25529 = ( ~w25253 & w25527 ) | ( ~w25253 & w25528 ) | ( w25527 & w25528 ) ;
  assign w25530 = w25528 | w25529 ;
  assign w25531 = \pi095 ^ w25238 ;
  assign w25532 = ( ~w25246 & w25530 ) | ( ~w25246 & w25531 ) | ( w25530 & w25531 ) ;
  assign w25533 = w25531 | w25532 ;
  assign w25534 = \pi096 ^ w25225 ;
  assign w25535 = ( ~w25239 & w25533 ) | ( ~w25239 & w25534 ) | ( w25533 & w25534 ) ;
  assign w25536 = w25534 | w25535 ;
  assign w25537 = \pi097 ^ w25231 ;
  assign w25538 = w25232 & ~w25537 ;
  assign w25539 = ( w25536 & w25537 ) | ( w25536 & ~w25538 ) | ( w25537 & ~w25538 ) ;
  assign w25540 = ~\pi097 & w25231 ;
  assign w25541 = w25539 & ~w25540 ;
  assign w25542 = w6047 | w25541 ;
  assign w25543 = w25225 & w25542 ;
  assign w25544 = ~w25239 & w25533 ;
  assign w25545 = w25534 ^ w25544 ;
  assign w25546 = ~w25542 & w25545 ;
  assign w25547 = w25543 | w25546 ;
  assign w25548 = w25231 & w25542 ;
  assign w25549 = ~w25232 & w25536 ;
  assign w25550 = w25537 ^ w25549 ;
  assign w25551 = ~w25542 & w25550 ;
  assign w25552 = w25548 | w25551 ;
  assign w25553 = ~\pi097 & w25547 ;
  assign w25554 = w25238 & w25542 ;
  assign w25555 = ~w25246 & w25530 ;
  assign w25556 = w25531 ^ w25555 ;
  assign w25557 = ~w25542 & w25556 ;
  assign w25558 = w25554 | w25557 ;
  assign w25559 = ~\pi096 & w25558 ;
  assign w25560 = w25245 & w25542 ;
  assign w25561 = ~w25253 & w25527 ;
  assign w25562 = w25528 ^ w25561 ;
  assign w25563 = ~w25542 & w25562 ;
  assign w25564 = w25560 | w25563 ;
  assign w25565 = ~\pi095 & w25564 ;
  assign w25566 = w25252 & w25542 ;
  assign w25567 = ~w25260 & w25524 ;
  assign w25568 = w25525 ^ w25567 ;
  assign w25569 = ~w25542 & w25568 ;
  assign w25570 = w25566 | w25569 ;
  assign w25571 = ~\pi094 & w25570 ;
  assign w25572 = w25259 & w25542 ;
  assign w25573 = ~w25267 & w25521 ;
  assign w25574 = w25522 ^ w25573 ;
  assign w25575 = ~w25542 & w25574 ;
  assign w25576 = w25572 | w25575 ;
  assign w25577 = ~\pi093 & w25576 ;
  assign w25578 = w25266 & w25542 ;
  assign w25579 = ~w25274 & w25518 ;
  assign w25580 = w25519 ^ w25579 ;
  assign w25581 = ~w25542 & w25580 ;
  assign w25582 = w25578 | w25581 ;
  assign w25583 = ~\pi092 & w25582 ;
  assign w25584 = w25273 & w25542 ;
  assign w25585 = ~w25281 & w25515 ;
  assign w25586 = w25516 ^ w25585 ;
  assign w25587 = ~w25542 & w25586 ;
  assign w25588 = w25584 | w25587 ;
  assign w25589 = ~\pi091 & w25588 ;
  assign w25590 = w25280 & w25542 ;
  assign w25591 = ~w25288 & w25512 ;
  assign w25592 = w25513 ^ w25591 ;
  assign w25593 = ~w25542 & w25592 ;
  assign w25594 = w25590 | w25593 ;
  assign w25595 = ~\pi090 & w25594 ;
  assign w25596 = w25287 & w25542 ;
  assign w25597 = ~w25295 & w25509 ;
  assign w25598 = w25510 ^ w25597 ;
  assign w25599 = ~w25542 & w25598 ;
  assign w25600 = w25596 | w25599 ;
  assign w25601 = ~\pi089 & w25600 ;
  assign w25602 = w25294 & w25542 ;
  assign w25603 = ~w25302 & w25506 ;
  assign w25604 = w25507 ^ w25603 ;
  assign w25605 = ~w25542 & w25604 ;
  assign w25606 = w25602 | w25605 ;
  assign w25607 = ~\pi088 & w25606 ;
  assign w25608 = w25301 & w25542 ;
  assign w25609 = ~w25309 & w25503 ;
  assign w25610 = w25504 ^ w25609 ;
  assign w25611 = ~w25542 & w25610 ;
  assign w25612 = w25608 | w25611 ;
  assign w25613 = ~\pi087 & w25612 ;
  assign w25614 = w25308 & w25542 ;
  assign w25615 = ~w25316 & w25500 ;
  assign w25616 = w25501 ^ w25615 ;
  assign w25617 = ~w25542 & w25616 ;
  assign w25618 = w25614 | w25617 ;
  assign w25619 = ~\pi086 & w25618 ;
  assign w25620 = w25315 & w25542 ;
  assign w25621 = ~w25323 & w25497 ;
  assign w25622 = w25498 ^ w25621 ;
  assign w25623 = ~w25542 & w25622 ;
  assign w25624 = w25620 | w25623 ;
  assign w25625 = ~\pi085 & w25624 ;
  assign w25626 = w25322 & w25542 ;
  assign w25627 = ~w25330 & w25494 ;
  assign w25628 = w25495 ^ w25627 ;
  assign w25629 = ~w25542 & w25628 ;
  assign w25630 = w25626 | w25629 ;
  assign w25631 = ~\pi084 & w25630 ;
  assign w25632 = w25329 & w25542 ;
  assign w25633 = ~w25337 & w25491 ;
  assign w25634 = w25492 ^ w25633 ;
  assign w25635 = ~w25542 & w25634 ;
  assign w25636 = w25632 | w25635 ;
  assign w25637 = ~\pi083 & w25636 ;
  assign w25638 = w25336 & w25542 ;
  assign w25639 = ~w25344 & w25488 ;
  assign w25640 = w25489 ^ w25639 ;
  assign w25641 = ~w25542 & w25640 ;
  assign w25642 = w25638 | w25641 ;
  assign w25643 = ~\pi082 & w25642 ;
  assign w25644 = w25343 & w25542 ;
  assign w25645 = ~w25351 & w25485 ;
  assign w25646 = w25486 ^ w25645 ;
  assign w25647 = ~w25542 & w25646 ;
  assign w25648 = w25644 | w25647 ;
  assign w25649 = ~\pi081 & w25648 ;
  assign w25650 = w25350 & w25542 ;
  assign w25651 = ~w25358 & w25482 ;
  assign w25652 = w25483 ^ w25651 ;
  assign w25653 = ~w25542 & w25652 ;
  assign w25654 = w25650 | w25653 ;
  assign w25655 = ~\pi080 & w25654 ;
  assign w25656 = w25357 & w25542 ;
  assign w25657 = ~w25365 & w25479 ;
  assign w25658 = w25480 ^ w25657 ;
  assign w25659 = ~w25542 & w25658 ;
  assign w25660 = w25656 | w25659 ;
  assign w25661 = ~\pi079 & w25660 ;
  assign w25662 = w25364 & w25542 ;
  assign w25663 = ~w25372 & w25476 ;
  assign w25664 = w25477 ^ w25663 ;
  assign w25665 = ~w25542 & w25664 ;
  assign w25666 = w25662 | w25665 ;
  assign w25667 = ~\pi078 & w25666 ;
  assign w25668 = w25371 & w25542 ;
  assign w25669 = ~w25379 & w25473 ;
  assign w25670 = w25474 ^ w25669 ;
  assign w25671 = ~w25542 & w25670 ;
  assign w25672 = w25668 | w25671 ;
  assign w25673 = ~\pi077 & w25672 ;
  assign w25674 = w25378 & w25542 ;
  assign w25675 = ~w25386 & w25470 ;
  assign w25676 = w25471 ^ w25675 ;
  assign w25677 = ~w25542 & w25676 ;
  assign w25678 = w25674 | w25677 ;
  assign w25679 = ~\pi076 & w25678 ;
  assign w25680 = w25385 & w25542 ;
  assign w25681 = ~w25393 & w25467 ;
  assign w25682 = w25468 ^ w25681 ;
  assign w25683 = ~w25542 & w25682 ;
  assign w25684 = w25680 | w25683 ;
  assign w25685 = ~\pi075 & w25684 ;
  assign w25686 = w25392 & w25542 ;
  assign w25687 = ~w25400 & w25464 ;
  assign w25688 = w25465 ^ w25687 ;
  assign w25689 = ~w25542 & w25688 ;
  assign w25690 = w25686 | w25689 ;
  assign w25691 = ~\pi074 & w25690 ;
  assign w25692 = w25399 & w25542 ;
  assign w25693 = ~w25407 & w25461 ;
  assign w25694 = w25462 ^ w25693 ;
  assign w25695 = ~w25542 & w25694 ;
  assign w25696 = w25692 | w25695 ;
  assign w25697 = ~\pi073 & w25696 ;
  assign w25698 = w25406 & w25542 ;
  assign w25699 = ~w25414 & w25458 ;
  assign w25700 = w25459 ^ w25699 ;
  assign w25701 = ~w25542 & w25700 ;
  assign w25702 = w25698 | w25701 ;
  assign w25703 = ~\pi072 & w25702 ;
  assign w25704 = w25413 & w25542 ;
  assign w25705 = ~w25421 & w25455 ;
  assign w25706 = w25456 ^ w25705 ;
  assign w25707 = ~w25542 & w25706 ;
  assign w25708 = w25704 | w25707 ;
  assign w25709 = ~\pi071 & w25708 ;
  assign w25710 = w25420 & w25542 ;
  assign w25711 = ~w25428 & w25452 ;
  assign w25712 = w25453 ^ w25711 ;
  assign w25713 = ~w25542 & w25712 ;
  assign w25714 = w25710 | w25713 ;
  assign w25715 = ~\pi070 & w25714 ;
  assign w25716 = w25427 & w25542 ;
  assign w25717 = ~w25434 & w25449 ;
  assign w25718 = w25450 ^ w25717 ;
  assign w25719 = ~w25542 & w25718 ;
  assign w25720 = w25716 | w25719 ;
  assign w25721 = ~\pi069 & w25720 ;
  assign w25722 = w25433 & w25542 ;
  assign w25723 = ~w25439 & w25446 ;
  assign w25724 = w25447 ^ w25723 ;
  assign w25725 = ~w25542 & w25724 ;
  assign w25726 = w25722 | w25725 ;
  assign w25727 = ~\pi068 & w25726 ;
  assign w25728 = w25438 & w25542 ;
  assign w25729 = \pi064 & ~w25219 ;
  assign w25730 = \pi031 ^ w25729 ;
  assign w25731 = ( \pi065 & w6235 ) | ( \pi065 & ~w25730 ) | ( w6235 & ~w25730 ) ;
  assign w25732 = w25442 ^ w25731 ;
  assign w25733 = ( w6047 & w25541 ) | ( w6047 & w25732 ) | ( w25541 & w25732 ) ;
  assign w25734 = w25732 & ~w25733 ;
  assign w25735 = w25728 | w25734 ;
  assign w25736 = ~\pi067 & w25735 ;
  assign w25737 = \pi030 ^ w25219 ;
  assign w25738 = ( \pi064 & w6047 ) | ( \pi064 & w25737 ) | ( w6047 & w25737 ) ;
  assign w25739 = w6242 ^ w25738 ;
  assign w25740 = ~w6047 & w25739 ;
  assign w25741 = ~w25541 & w25740 ;
  assign w25742 = ( ~\pi064 & w25219 ) | ( ~\pi064 & w25542 ) | ( w25219 & w25542 ) ;
  assign w25743 = \pi031 ^ w25742 ;
  assign w25744 = w25542 & ~w25743 ;
  assign w25745 = w25741 | w25744 ;
  assign w25746 = ~\pi066 & w25745 ;
  assign w25747 = ( \pi030 & ~w6258 ) | ( \pi030 & w25541 ) | ( ~w6258 & w25541 ) ;
  assign w25748 = \pi030 & w25747 ;
  assign w25749 = w6266 & ~w25541 ;
  assign w25750 = w25748 | w25749 ;
  assign w25751 = \pi065 ^ w25750 ;
  assign w25752 = w6269 | w25751 ;
  assign w25753 = w25542 | w25741 ;
  assign w25754 = ( w25730 & w25741 ) | ( w25730 & w25753 ) | ( w25741 & w25753 ) ;
  assign w25755 = \pi066 ^ w25754 ;
  assign w25756 = ~\pi065 & w25750 ;
  assign w25757 = w25752 | w25756 ;
  assign w25758 = ( w25755 & ~w25756 ) | ( w25755 & w25757 ) | ( ~w25756 & w25757 ) ;
  assign w25759 = \pi067 ^ w25735 ;
  assign w25760 = ( ~w25746 & w25758 ) | ( ~w25746 & w25759 ) | ( w25758 & w25759 ) ;
  assign w25761 = w25759 | w25760 ;
  assign w25762 = \pi068 ^ w25726 ;
  assign w25763 = ( ~w25736 & w25761 ) | ( ~w25736 & w25762 ) | ( w25761 & w25762 ) ;
  assign w25764 = w25762 | w25763 ;
  assign w25765 = \pi069 ^ w25720 ;
  assign w25766 = ( ~w25727 & w25764 ) | ( ~w25727 & w25765 ) | ( w25764 & w25765 ) ;
  assign w25767 = w25765 | w25766 ;
  assign w25768 = \pi070 ^ w25714 ;
  assign w25769 = ( ~w25721 & w25767 ) | ( ~w25721 & w25768 ) | ( w25767 & w25768 ) ;
  assign w25770 = w25768 | w25769 ;
  assign w25771 = \pi071 ^ w25708 ;
  assign w25772 = ( ~w25715 & w25770 ) | ( ~w25715 & w25771 ) | ( w25770 & w25771 ) ;
  assign w25773 = w25771 | w25772 ;
  assign w25774 = \pi072 ^ w25702 ;
  assign w25775 = ( ~w25709 & w25773 ) | ( ~w25709 & w25774 ) | ( w25773 & w25774 ) ;
  assign w25776 = w25774 | w25775 ;
  assign w25777 = \pi073 ^ w25696 ;
  assign w25778 = ( ~w25703 & w25776 ) | ( ~w25703 & w25777 ) | ( w25776 & w25777 ) ;
  assign w25779 = w25777 | w25778 ;
  assign w25780 = \pi074 ^ w25690 ;
  assign w25781 = ( ~w25697 & w25779 ) | ( ~w25697 & w25780 ) | ( w25779 & w25780 ) ;
  assign w25782 = w25780 | w25781 ;
  assign w25783 = \pi075 ^ w25684 ;
  assign w25784 = ( ~w25691 & w25782 ) | ( ~w25691 & w25783 ) | ( w25782 & w25783 ) ;
  assign w25785 = w25783 | w25784 ;
  assign w25786 = \pi076 ^ w25678 ;
  assign w25787 = ( ~w25685 & w25785 ) | ( ~w25685 & w25786 ) | ( w25785 & w25786 ) ;
  assign w25788 = w25786 | w25787 ;
  assign w25789 = \pi077 ^ w25672 ;
  assign w25790 = ( ~w25679 & w25788 ) | ( ~w25679 & w25789 ) | ( w25788 & w25789 ) ;
  assign w25791 = w25789 | w25790 ;
  assign w25792 = \pi078 ^ w25666 ;
  assign w25793 = ( ~w25673 & w25791 ) | ( ~w25673 & w25792 ) | ( w25791 & w25792 ) ;
  assign w25794 = w25792 | w25793 ;
  assign w25795 = \pi079 ^ w25660 ;
  assign w25796 = ( ~w25667 & w25794 ) | ( ~w25667 & w25795 ) | ( w25794 & w25795 ) ;
  assign w25797 = w25795 | w25796 ;
  assign w25798 = \pi080 ^ w25654 ;
  assign w25799 = ( ~w25661 & w25797 ) | ( ~w25661 & w25798 ) | ( w25797 & w25798 ) ;
  assign w25800 = w25798 | w25799 ;
  assign w25801 = \pi081 ^ w25648 ;
  assign w25802 = ( ~w25655 & w25800 ) | ( ~w25655 & w25801 ) | ( w25800 & w25801 ) ;
  assign w25803 = w25801 | w25802 ;
  assign w25804 = \pi082 ^ w25642 ;
  assign w25805 = ( ~w25649 & w25803 ) | ( ~w25649 & w25804 ) | ( w25803 & w25804 ) ;
  assign w25806 = w25804 | w25805 ;
  assign w25807 = \pi083 ^ w25636 ;
  assign w25808 = ( ~w25643 & w25806 ) | ( ~w25643 & w25807 ) | ( w25806 & w25807 ) ;
  assign w25809 = w25807 | w25808 ;
  assign w25810 = \pi084 ^ w25630 ;
  assign w25811 = ( ~w25637 & w25809 ) | ( ~w25637 & w25810 ) | ( w25809 & w25810 ) ;
  assign w25812 = w25810 | w25811 ;
  assign w25813 = \pi085 ^ w25624 ;
  assign w25814 = ( ~w25631 & w25812 ) | ( ~w25631 & w25813 ) | ( w25812 & w25813 ) ;
  assign w25815 = w25813 | w25814 ;
  assign w25816 = \pi086 ^ w25618 ;
  assign w25817 = ( ~w25625 & w25815 ) | ( ~w25625 & w25816 ) | ( w25815 & w25816 ) ;
  assign w25818 = w25816 | w25817 ;
  assign w25819 = \pi087 ^ w25612 ;
  assign w25820 = ( ~w25619 & w25818 ) | ( ~w25619 & w25819 ) | ( w25818 & w25819 ) ;
  assign w25821 = w25819 | w25820 ;
  assign w25822 = \pi088 ^ w25606 ;
  assign w25823 = ( ~w25613 & w25821 ) | ( ~w25613 & w25822 ) | ( w25821 & w25822 ) ;
  assign w25824 = w25822 | w25823 ;
  assign w25825 = \pi089 ^ w25600 ;
  assign w25826 = ( ~w25607 & w25824 ) | ( ~w25607 & w25825 ) | ( w25824 & w25825 ) ;
  assign w25827 = w25825 | w25826 ;
  assign w25828 = \pi090 ^ w25594 ;
  assign w25829 = ( ~w25601 & w25827 ) | ( ~w25601 & w25828 ) | ( w25827 & w25828 ) ;
  assign w25830 = w25828 | w25829 ;
  assign w25831 = \pi091 ^ w25588 ;
  assign w25832 = ( ~w25595 & w25830 ) | ( ~w25595 & w25831 ) | ( w25830 & w25831 ) ;
  assign w25833 = w25831 | w25832 ;
  assign w25834 = \pi092 ^ w25582 ;
  assign w25835 = ( ~w25589 & w25833 ) | ( ~w25589 & w25834 ) | ( w25833 & w25834 ) ;
  assign w25836 = w25834 | w25835 ;
  assign w25837 = \pi093 ^ w25576 ;
  assign w25838 = ( ~w25583 & w25836 ) | ( ~w25583 & w25837 ) | ( w25836 & w25837 ) ;
  assign w25839 = w25837 | w25838 ;
  assign w25840 = \pi094 ^ w25570 ;
  assign w25841 = ( ~w25577 & w25839 ) | ( ~w25577 & w25840 ) | ( w25839 & w25840 ) ;
  assign w25842 = w25840 | w25841 ;
  assign w25843 = \pi095 ^ w25564 ;
  assign w25844 = ( ~w25571 & w25842 ) | ( ~w25571 & w25843 ) | ( w25842 & w25843 ) ;
  assign w25845 = w25843 | w25844 ;
  assign w25846 = \pi096 ^ w25558 ;
  assign w25847 = ( ~w25565 & w25845 ) | ( ~w25565 & w25846 ) | ( w25845 & w25846 ) ;
  assign w25848 = w25846 | w25847 ;
  assign w25849 = \pi097 ^ w25547 ;
  assign w25850 = ( ~w25559 & w25848 ) | ( ~w25559 & w25849 ) | ( w25848 & w25849 ) ;
  assign w25851 = w25849 | w25850 ;
  assign w25852 = \pi098 ^ w25552 ;
  assign w25853 = w25553 & ~w25852 ;
  assign w25854 = ( w25851 & w25852 ) | ( w25851 & ~w25853 ) | ( w25852 & ~w25853 ) ;
  assign w25855 = ~\pi098 & w25552 ;
  assign w25856 = w25854 & ~w25855 ;
  assign w25857 = w6379 | w25856 ;
  assign w25858 = w25547 & w25857 ;
  assign w25859 = ~w25559 & w25848 ;
  assign w25860 = w25849 ^ w25859 ;
  assign w25861 = ~w25857 & w25860 ;
  assign w25862 = w25858 | w25861 ;
  assign w25863 = ~\pi098 & w25862 ;
  assign w25864 = w25558 & w25857 ;
  assign w25865 = ~w25565 & w25845 ;
  assign w25866 = w25846 ^ w25865 ;
  assign w25867 = ~w25857 & w25866 ;
  assign w25868 = w25864 | w25867 ;
  assign w25869 = ~\pi097 & w25868 ;
  assign w25870 = w25564 & w25857 ;
  assign w25871 = ~w25571 & w25842 ;
  assign w25872 = w25843 ^ w25871 ;
  assign w25873 = ~w25857 & w25872 ;
  assign w25874 = w25870 | w25873 ;
  assign w25875 = ~\pi096 & w25874 ;
  assign w25876 = w25570 & w25857 ;
  assign w25877 = ~w25577 & w25839 ;
  assign w25878 = w25840 ^ w25877 ;
  assign w25879 = ~w25857 & w25878 ;
  assign w25880 = w25876 | w25879 ;
  assign w25881 = ~\pi095 & w25880 ;
  assign w25882 = w25576 & w25857 ;
  assign w25883 = ~w25583 & w25836 ;
  assign w25884 = w25837 ^ w25883 ;
  assign w25885 = ~w25857 & w25884 ;
  assign w25886 = w25882 | w25885 ;
  assign w25887 = ~\pi094 & w25886 ;
  assign w25888 = w25582 & w25857 ;
  assign w25889 = ~w25589 & w25833 ;
  assign w25890 = w25834 ^ w25889 ;
  assign w25891 = ~w25857 & w25890 ;
  assign w25892 = w25888 | w25891 ;
  assign w25893 = ~\pi093 & w25892 ;
  assign w25894 = w25588 & w25857 ;
  assign w25895 = ~w25595 & w25830 ;
  assign w25896 = w25831 ^ w25895 ;
  assign w25897 = ~w25857 & w25896 ;
  assign w25898 = w25894 | w25897 ;
  assign w25899 = ~\pi092 & w25898 ;
  assign w25900 = w25594 & w25857 ;
  assign w25901 = ~w25601 & w25827 ;
  assign w25902 = w25828 ^ w25901 ;
  assign w25903 = ~w25857 & w25902 ;
  assign w25904 = w25900 | w25903 ;
  assign w25905 = ~\pi091 & w25904 ;
  assign w25906 = w25600 & w25857 ;
  assign w25907 = ~w25607 & w25824 ;
  assign w25908 = w25825 ^ w25907 ;
  assign w25909 = ~w25857 & w25908 ;
  assign w25910 = w25906 | w25909 ;
  assign w25911 = ~\pi090 & w25910 ;
  assign w25912 = w25606 & w25857 ;
  assign w25913 = ~w25613 & w25821 ;
  assign w25914 = w25822 ^ w25913 ;
  assign w25915 = ~w25857 & w25914 ;
  assign w25916 = w25912 | w25915 ;
  assign w25917 = ~\pi089 & w25916 ;
  assign w25918 = w25612 & w25857 ;
  assign w25919 = ~w25619 & w25818 ;
  assign w25920 = w25819 ^ w25919 ;
  assign w25921 = ~w25857 & w25920 ;
  assign w25922 = w25918 | w25921 ;
  assign w25923 = ~\pi088 & w25922 ;
  assign w25924 = w25618 & w25857 ;
  assign w25925 = ~w25625 & w25815 ;
  assign w25926 = w25816 ^ w25925 ;
  assign w25927 = ~w25857 & w25926 ;
  assign w25928 = w25924 | w25927 ;
  assign w25929 = ~\pi087 & w25928 ;
  assign w25930 = w25624 & w25857 ;
  assign w25931 = ~w25631 & w25812 ;
  assign w25932 = w25813 ^ w25931 ;
  assign w25933 = ~w25857 & w25932 ;
  assign w25934 = w25930 | w25933 ;
  assign w25935 = ~\pi086 & w25934 ;
  assign w25936 = w25630 & w25857 ;
  assign w25937 = ~w25637 & w25809 ;
  assign w25938 = w25810 ^ w25937 ;
  assign w25939 = ~w25857 & w25938 ;
  assign w25940 = w25936 | w25939 ;
  assign w25941 = ~\pi085 & w25940 ;
  assign w25942 = w25636 & w25857 ;
  assign w25943 = ~w25643 & w25806 ;
  assign w25944 = w25807 ^ w25943 ;
  assign w25945 = ~w25857 & w25944 ;
  assign w25946 = w25942 | w25945 ;
  assign w25947 = ~\pi084 & w25946 ;
  assign w25948 = w25642 & w25857 ;
  assign w25949 = ~w25649 & w25803 ;
  assign w25950 = w25804 ^ w25949 ;
  assign w25951 = ~w25857 & w25950 ;
  assign w25952 = w25948 | w25951 ;
  assign w25953 = ~\pi083 & w25952 ;
  assign w25954 = w25648 & w25857 ;
  assign w25955 = ~w25655 & w25800 ;
  assign w25956 = w25801 ^ w25955 ;
  assign w25957 = ~w25857 & w25956 ;
  assign w25958 = w25954 | w25957 ;
  assign w25959 = ~\pi082 & w25958 ;
  assign w25960 = w25654 & w25857 ;
  assign w25961 = ~w25661 & w25797 ;
  assign w25962 = w25798 ^ w25961 ;
  assign w25963 = ~w25857 & w25962 ;
  assign w25964 = w25960 | w25963 ;
  assign w25965 = ~\pi081 & w25964 ;
  assign w25966 = w25660 & w25857 ;
  assign w25967 = ~w25667 & w25794 ;
  assign w25968 = w25795 ^ w25967 ;
  assign w25969 = ~w25857 & w25968 ;
  assign w25970 = w25966 | w25969 ;
  assign w25971 = ~\pi080 & w25970 ;
  assign w25972 = w25666 & w25857 ;
  assign w25973 = ~w25673 & w25791 ;
  assign w25974 = w25792 ^ w25973 ;
  assign w25975 = ~w25857 & w25974 ;
  assign w25976 = w25972 | w25975 ;
  assign w25977 = ~\pi079 & w25976 ;
  assign w25978 = w25672 & w25857 ;
  assign w25979 = ~w25679 & w25788 ;
  assign w25980 = w25789 ^ w25979 ;
  assign w25981 = ~w25857 & w25980 ;
  assign w25982 = w25978 | w25981 ;
  assign w25983 = ~\pi078 & w25982 ;
  assign w25984 = w25678 & w25857 ;
  assign w25985 = ~w25685 & w25785 ;
  assign w25986 = w25786 ^ w25985 ;
  assign w25987 = ~w25857 & w25986 ;
  assign w25988 = w25984 | w25987 ;
  assign w25989 = ~\pi077 & w25988 ;
  assign w25990 = w25684 & w25857 ;
  assign w25991 = ~w25691 & w25782 ;
  assign w25992 = w25783 ^ w25991 ;
  assign w25993 = ~w25857 & w25992 ;
  assign w25994 = w25990 | w25993 ;
  assign w25995 = ~\pi076 & w25994 ;
  assign w25996 = w25690 & w25857 ;
  assign w25997 = ~w25697 & w25779 ;
  assign w25998 = w25780 ^ w25997 ;
  assign w25999 = ~w25857 & w25998 ;
  assign w26000 = w25996 | w25999 ;
  assign w26001 = ~\pi075 & w26000 ;
  assign w26002 = w25696 & w25857 ;
  assign w26003 = ~w25703 & w25776 ;
  assign w26004 = w25777 ^ w26003 ;
  assign w26005 = ~w25857 & w26004 ;
  assign w26006 = w26002 | w26005 ;
  assign w26007 = ~\pi074 & w26006 ;
  assign w26008 = w25702 & w25857 ;
  assign w26009 = ~w25709 & w25773 ;
  assign w26010 = w25774 ^ w26009 ;
  assign w26011 = ~w25857 & w26010 ;
  assign w26012 = w26008 | w26011 ;
  assign w26013 = ~\pi073 & w26012 ;
  assign w26014 = w25708 & w25857 ;
  assign w26015 = ~w25715 & w25770 ;
  assign w26016 = w25771 ^ w26015 ;
  assign w26017 = ~w25857 & w26016 ;
  assign w26018 = w26014 | w26017 ;
  assign w26019 = ~\pi072 & w26018 ;
  assign w26020 = w25714 & w25857 ;
  assign w26021 = ~w25721 & w25767 ;
  assign w26022 = w25768 ^ w26021 ;
  assign w26023 = ~w25857 & w26022 ;
  assign w26024 = w26020 | w26023 ;
  assign w26025 = ~\pi071 & w26024 ;
  assign w26026 = w25720 & w25857 ;
  assign w26027 = ~w25727 & w25764 ;
  assign w26028 = w25765 ^ w26027 ;
  assign w26029 = ~w25857 & w26028 ;
  assign w26030 = w26026 | w26029 ;
  assign w26031 = ~\pi070 & w26030 ;
  assign w26032 = w25726 & w25857 ;
  assign w26033 = ~w25736 & w25761 ;
  assign w26034 = w25762 ^ w26033 ;
  assign w26035 = ~w25857 & w26034 ;
  assign w26036 = w26032 | w26035 ;
  assign w26037 = ~\pi069 & w26036 ;
  assign w26038 = w25735 & w25857 ;
  assign w26039 = ~w25746 & w25758 ;
  assign w26040 = w25759 ^ w26039 ;
  assign w26041 = ~w25857 & w26040 ;
  assign w26042 = w26038 | w26041 ;
  assign w26043 = ~\pi068 & w26042 ;
  assign w26044 = w25745 & w25857 ;
  assign w26045 = ~w25750 & w25752 ;
  assign w26046 = ( \pi065 & w25752 ) | ( \pi065 & w26045 ) | ( w25752 & w26045 ) ;
  assign w26047 = w25755 ^ w26046 ;
  assign w26048 = ~w25857 & w26047 ;
  assign w26049 = w26044 | w26048 ;
  assign w26050 = ~\pi067 & w26049 ;
  assign w26051 = w25750 & w25857 ;
  assign w26052 = ( ~w6379 & w25748 ) | ( ~w6379 & w25749 ) | ( w25748 & w25749 ) ;
  assign w26053 = \pi065 ^ w26052 ;
  assign w26054 = ( w6269 & ~w6379 ) | ( w6269 & w26053 ) | ( ~w6379 & w26053 ) ;
  assign w26055 = ( w6269 & w25856 ) | ( w6269 & w26053 ) | ( w25856 & w26053 ) ;
  assign w26056 = w26054 & ~w26055 ;
  assign w26057 = w26051 | w26056 ;
  assign w26058 = ~\pi066 & w26057 ;
  assign w26059 = ( \pi029 & ~w6584 ) | ( \pi029 & w25856 ) | ( ~w6584 & w25856 ) ;
  assign w26060 = \pi029 & w26059 ;
  assign w26061 = w6591 & ~w25856 ;
  assign w26062 = w26060 | w26061 ;
  assign w26063 = \pi065 ^ w26062 ;
  assign w26064 = w6594 | w26063 ;
  assign w26065 = \pi066 ^ w26057 ;
  assign w26066 = ~\pi065 & w26062 ;
  assign w26067 = w26064 | w26066 ;
  assign w26068 = ( w26065 & ~w26066 ) | ( w26065 & w26067 ) | ( ~w26066 & w26067 ) ;
  assign w26069 = \pi067 ^ w26049 ;
  assign w26070 = ( ~w26058 & w26068 ) | ( ~w26058 & w26069 ) | ( w26068 & w26069 ) ;
  assign w26071 = w26069 | w26070 ;
  assign w26072 = \pi068 ^ w26042 ;
  assign w26073 = ( ~w26050 & w26071 ) | ( ~w26050 & w26072 ) | ( w26071 & w26072 ) ;
  assign w26074 = w26072 | w26073 ;
  assign w26075 = \pi069 ^ w26036 ;
  assign w26076 = ( ~w26043 & w26074 ) | ( ~w26043 & w26075 ) | ( w26074 & w26075 ) ;
  assign w26077 = w26075 | w26076 ;
  assign w26078 = \pi070 ^ w26030 ;
  assign w26079 = ( ~w26037 & w26077 ) | ( ~w26037 & w26078 ) | ( w26077 & w26078 ) ;
  assign w26080 = w26078 | w26079 ;
  assign w26081 = \pi071 ^ w26024 ;
  assign w26082 = ( ~w26031 & w26080 ) | ( ~w26031 & w26081 ) | ( w26080 & w26081 ) ;
  assign w26083 = w26081 | w26082 ;
  assign w26084 = \pi072 ^ w26018 ;
  assign w26085 = ( ~w26025 & w26083 ) | ( ~w26025 & w26084 ) | ( w26083 & w26084 ) ;
  assign w26086 = w26084 | w26085 ;
  assign w26087 = \pi073 ^ w26012 ;
  assign w26088 = ( ~w26019 & w26086 ) | ( ~w26019 & w26087 ) | ( w26086 & w26087 ) ;
  assign w26089 = w26087 | w26088 ;
  assign w26090 = \pi074 ^ w26006 ;
  assign w26091 = ( ~w26013 & w26089 ) | ( ~w26013 & w26090 ) | ( w26089 & w26090 ) ;
  assign w26092 = w26090 | w26091 ;
  assign w26093 = \pi075 ^ w26000 ;
  assign w26094 = ( ~w26007 & w26092 ) | ( ~w26007 & w26093 ) | ( w26092 & w26093 ) ;
  assign w26095 = w26093 | w26094 ;
  assign w26096 = \pi076 ^ w25994 ;
  assign w26097 = ( ~w26001 & w26095 ) | ( ~w26001 & w26096 ) | ( w26095 & w26096 ) ;
  assign w26098 = w26096 | w26097 ;
  assign w26099 = \pi077 ^ w25988 ;
  assign w26100 = ( ~w25995 & w26098 ) | ( ~w25995 & w26099 ) | ( w26098 & w26099 ) ;
  assign w26101 = w26099 | w26100 ;
  assign w26102 = \pi078 ^ w25982 ;
  assign w26103 = ( ~w25989 & w26101 ) | ( ~w25989 & w26102 ) | ( w26101 & w26102 ) ;
  assign w26104 = w26102 | w26103 ;
  assign w26105 = \pi079 ^ w25976 ;
  assign w26106 = ( ~w25983 & w26104 ) | ( ~w25983 & w26105 ) | ( w26104 & w26105 ) ;
  assign w26107 = w26105 | w26106 ;
  assign w26108 = \pi080 ^ w25970 ;
  assign w26109 = ( ~w25977 & w26107 ) | ( ~w25977 & w26108 ) | ( w26107 & w26108 ) ;
  assign w26110 = w26108 | w26109 ;
  assign w26111 = \pi081 ^ w25964 ;
  assign w26112 = ( ~w25971 & w26110 ) | ( ~w25971 & w26111 ) | ( w26110 & w26111 ) ;
  assign w26113 = w26111 | w26112 ;
  assign w26114 = \pi082 ^ w25958 ;
  assign w26115 = ( ~w25965 & w26113 ) | ( ~w25965 & w26114 ) | ( w26113 & w26114 ) ;
  assign w26116 = w26114 | w26115 ;
  assign w26117 = \pi083 ^ w25952 ;
  assign w26118 = ( ~w25959 & w26116 ) | ( ~w25959 & w26117 ) | ( w26116 & w26117 ) ;
  assign w26119 = w26117 | w26118 ;
  assign w26120 = \pi084 ^ w25946 ;
  assign w26121 = ( ~w25953 & w26119 ) | ( ~w25953 & w26120 ) | ( w26119 & w26120 ) ;
  assign w26122 = w26120 | w26121 ;
  assign w26123 = \pi085 ^ w25940 ;
  assign w26124 = ( ~w25947 & w26122 ) | ( ~w25947 & w26123 ) | ( w26122 & w26123 ) ;
  assign w26125 = w26123 | w26124 ;
  assign w26126 = \pi086 ^ w25934 ;
  assign w26127 = ( ~w25941 & w26125 ) | ( ~w25941 & w26126 ) | ( w26125 & w26126 ) ;
  assign w26128 = w26126 | w26127 ;
  assign w26129 = \pi087 ^ w25928 ;
  assign w26130 = ( ~w25935 & w26128 ) | ( ~w25935 & w26129 ) | ( w26128 & w26129 ) ;
  assign w26131 = w26129 | w26130 ;
  assign w26132 = \pi088 ^ w25922 ;
  assign w26133 = ( ~w25929 & w26131 ) | ( ~w25929 & w26132 ) | ( w26131 & w26132 ) ;
  assign w26134 = w26132 | w26133 ;
  assign w26135 = \pi089 ^ w25916 ;
  assign w26136 = ( ~w25923 & w26134 ) | ( ~w25923 & w26135 ) | ( w26134 & w26135 ) ;
  assign w26137 = w26135 | w26136 ;
  assign w26138 = \pi090 ^ w25910 ;
  assign w26139 = ( ~w25917 & w26137 ) | ( ~w25917 & w26138 ) | ( w26137 & w26138 ) ;
  assign w26140 = w26138 | w26139 ;
  assign w26141 = \pi091 ^ w25904 ;
  assign w26142 = ( ~w25911 & w26140 ) | ( ~w25911 & w26141 ) | ( w26140 & w26141 ) ;
  assign w26143 = w26141 | w26142 ;
  assign w26144 = \pi092 ^ w25898 ;
  assign w26145 = ( ~w25905 & w26143 ) | ( ~w25905 & w26144 ) | ( w26143 & w26144 ) ;
  assign w26146 = w26144 | w26145 ;
  assign w26147 = \pi093 ^ w25892 ;
  assign w26148 = ( ~w25899 & w26146 ) | ( ~w25899 & w26147 ) | ( w26146 & w26147 ) ;
  assign w26149 = w26147 | w26148 ;
  assign w26150 = \pi094 ^ w25886 ;
  assign w26151 = ( ~w25893 & w26149 ) | ( ~w25893 & w26150 ) | ( w26149 & w26150 ) ;
  assign w26152 = w26150 | w26151 ;
  assign w26153 = \pi095 ^ w25880 ;
  assign w26154 = ( ~w25887 & w26152 ) | ( ~w25887 & w26153 ) | ( w26152 & w26153 ) ;
  assign w26155 = w26153 | w26154 ;
  assign w26156 = \pi096 ^ w25874 ;
  assign w26157 = ( ~w25881 & w26155 ) | ( ~w25881 & w26156 ) | ( w26155 & w26156 ) ;
  assign w26158 = w26156 | w26157 ;
  assign w26159 = \pi097 ^ w25868 ;
  assign w26160 = ( ~w25875 & w26158 ) | ( ~w25875 & w26159 ) | ( w26158 & w26159 ) ;
  assign w26161 = w26159 | w26160 ;
  assign w26162 = \pi098 ^ w25862 ;
  assign w26163 = ( ~w25869 & w26161 ) | ( ~w25869 & w26162 ) | ( w26161 & w26162 ) ;
  assign w26164 = w26162 | w26163 ;
  assign w26165 = w25552 & w25857 ;
  assign w26166 = ~w25553 & w25851 ;
  assign w26167 = w25852 ^ w26166 ;
  assign w26168 = ~w25857 & w26167 ;
  assign w26169 = w26165 | w26168 ;
  assign w26170 = ~\pi099 & w26169 ;
  assign w26171 = ( \pi099 & ~w26165 ) | ( \pi099 & w26168 ) | ( ~w26165 & w26168 ) ;
  assign w26172 = ~w26168 & w26171 ;
  assign w26173 = w26170 | w26172 ;
  assign w26174 = ( ~w25863 & w26164 ) | ( ~w25863 & w26173 ) | ( w26164 & w26173 ) ;
  assign w26175 = ( w368 & ~w26173 ) | ( w368 & w26174 ) | ( ~w26173 & w26174 ) ;
  assign w26176 = w26173 | w26175 ;
  assign w26177 = ~w6379 & w26169 ;
  assign w26178 = w26176 & ~w26177 ;
  assign w26179 = ~w25869 & w26161 ;
  assign w26180 = w26162 ^ w26179 ;
  assign w26181 = ~w26178 & w26180 ;
  assign w26182 = ( w25862 & w26176 ) | ( w25862 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26183 = ~w26177 & w26182 ;
  assign w26184 = w26181 | w26183 ;
  assign w26185 = ( ~w25863 & w26164 ) | ( ~w25863 & w26178 ) | ( w26164 & w26178 ) ;
  assign w26186 = w26173 ^ w26185 ;
  assign w26187 = ~w26178 & w26186 ;
  assign w26188 = ( w6379 & ~w26169 ) | ( w6379 & w26176 ) | ( ~w26169 & w26176 ) ;
  assign w26189 = w26169 & w26188 ;
  assign w26190 = w26187 | w26189 ;
  assign w26191 = ~\pi099 & w26184 ;
  assign w26192 = ~w25875 & w26158 ;
  assign w26193 = w26159 ^ w26192 ;
  assign w26194 = ~w26178 & w26193 ;
  assign w26195 = ( w25868 & w26176 ) | ( w25868 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26196 = ~w26177 & w26195 ;
  assign w26197 = w26194 | w26196 ;
  assign w26198 = ~\pi098 & w26197 ;
  assign w26199 = ~w25881 & w26155 ;
  assign w26200 = w26156 ^ w26199 ;
  assign w26201 = ~w26178 & w26200 ;
  assign w26202 = ( w25874 & w26176 ) | ( w25874 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26203 = ~w26177 & w26202 ;
  assign w26204 = w26201 | w26203 ;
  assign w26205 = ~\pi097 & w26204 ;
  assign w26206 = ~w25887 & w26152 ;
  assign w26207 = w26153 ^ w26206 ;
  assign w26208 = ~w26178 & w26207 ;
  assign w26209 = ( w25880 & w26176 ) | ( w25880 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26210 = ~w26177 & w26209 ;
  assign w26211 = w26208 | w26210 ;
  assign w26212 = ~\pi096 & w26211 ;
  assign w26213 = ~w25893 & w26149 ;
  assign w26214 = w26150 ^ w26213 ;
  assign w26215 = ~w26178 & w26214 ;
  assign w26216 = ( w25886 & w26176 ) | ( w25886 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26217 = ~w26177 & w26216 ;
  assign w26218 = w26215 | w26217 ;
  assign w26219 = ~\pi095 & w26218 ;
  assign w26220 = ~w25899 & w26146 ;
  assign w26221 = w26147 ^ w26220 ;
  assign w26222 = ~w26178 & w26221 ;
  assign w26223 = ( w25892 & w26176 ) | ( w25892 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26224 = ~w26177 & w26223 ;
  assign w26225 = w26222 | w26224 ;
  assign w26226 = ~\pi094 & w26225 ;
  assign w26227 = ~w25905 & w26143 ;
  assign w26228 = w26144 ^ w26227 ;
  assign w26229 = ~w26178 & w26228 ;
  assign w26230 = ( w25898 & w26176 ) | ( w25898 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26231 = ~w26177 & w26230 ;
  assign w26232 = w26229 | w26231 ;
  assign w26233 = ~\pi093 & w26232 ;
  assign w26234 = ~w25911 & w26140 ;
  assign w26235 = w26141 ^ w26234 ;
  assign w26236 = ~w26178 & w26235 ;
  assign w26237 = ( w25904 & w26176 ) | ( w25904 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26238 = ~w26177 & w26237 ;
  assign w26239 = w26236 | w26238 ;
  assign w26240 = ~\pi092 & w26239 ;
  assign w26241 = ~w25917 & w26137 ;
  assign w26242 = w26138 ^ w26241 ;
  assign w26243 = ~w26178 & w26242 ;
  assign w26244 = ( w25910 & w26176 ) | ( w25910 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26245 = ~w26177 & w26244 ;
  assign w26246 = w26243 | w26245 ;
  assign w26247 = ~\pi091 & w26246 ;
  assign w26248 = ~w25923 & w26134 ;
  assign w26249 = w26135 ^ w26248 ;
  assign w26250 = ~w26178 & w26249 ;
  assign w26251 = ( w25916 & w26176 ) | ( w25916 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26252 = ~w26177 & w26251 ;
  assign w26253 = w26250 | w26252 ;
  assign w26254 = ~\pi090 & w26253 ;
  assign w26255 = ~w25929 & w26131 ;
  assign w26256 = w26132 ^ w26255 ;
  assign w26257 = ~w26178 & w26256 ;
  assign w26258 = ( w25922 & w26176 ) | ( w25922 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26259 = ~w26177 & w26258 ;
  assign w26260 = w26257 | w26259 ;
  assign w26261 = ~\pi089 & w26260 ;
  assign w26262 = ~w25935 & w26128 ;
  assign w26263 = w26129 ^ w26262 ;
  assign w26264 = ~w26178 & w26263 ;
  assign w26265 = ( w25928 & w26176 ) | ( w25928 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26266 = ~w26177 & w26265 ;
  assign w26267 = w26264 | w26266 ;
  assign w26268 = ~\pi088 & w26267 ;
  assign w26269 = ~w25941 & w26125 ;
  assign w26270 = w26126 ^ w26269 ;
  assign w26271 = ~w26178 & w26270 ;
  assign w26272 = ( w25934 & w26176 ) | ( w25934 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26273 = ~w26177 & w26272 ;
  assign w26274 = w26271 | w26273 ;
  assign w26275 = ~\pi087 & w26274 ;
  assign w26276 = ~w25947 & w26122 ;
  assign w26277 = w26123 ^ w26276 ;
  assign w26278 = ~w26178 & w26277 ;
  assign w26279 = ( w25940 & w26176 ) | ( w25940 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26280 = ~w26177 & w26279 ;
  assign w26281 = w26278 | w26280 ;
  assign w26282 = ~\pi086 & w26281 ;
  assign w26283 = ~w25953 & w26119 ;
  assign w26284 = w26120 ^ w26283 ;
  assign w26285 = ~w26178 & w26284 ;
  assign w26286 = ( w25946 & w26176 ) | ( w25946 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26287 = ~w26177 & w26286 ;
  assign w26288 = w26285 | w26287 ;
  assign w26289 = ~\pi085 & w26288 ;
  assign w26290 = ~w25959 & w26116 ;
  assign w26291 = w26117 ^ w26290 ;
  assign w26292 = ~w26178 & w26291 ;
  assign w26293 = ( w25952 & w26176 ) | ( w25952 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26294 = ~w26177 & w26293 ;
  assign w26295 = w26292 | w26294 ;
  assign w26296 = ~\pi084 & w26295 ;
  assign w26297 = ~w25965 & w26113 ;
  assign w26298 = w26114 ^ w26297 ;
  assign w26299 = ~w26178 & w26298 ;
  assign w26300 = ( w25958 & w26176 ) | ( w25958 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26301 = ~w26177 & w26300 ;
  assign w26302 = w26299 | w26301 ;
  assign w26303 = ~\pi083 & w26302 ;
  assign w26304 = ~w25971 & w26110 ;
  assign w26305 = w26111 ^ w26304 ;
  assign w26306 = ~w26178 & w26305 ;
  assign w26307 = ( w25964 & w26176 ) | ( w25964 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26308 = ~w26177 & w26307 ;
  assign w26309 = w26306 | w26308 ;
  assign w26310 = ~\pi082 & w26309 ;
  assign w26311 = ~w25977 & w26107 ;
  assign w26312 = w26108 ^ w26311 ;
  assign w26313 = ~w26178 & w26312 ;
  assign w26314 = ( w25970 & w26176 ) | ( w25970 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26315 = ~w26177 & w26314 ;
  assign w26316 = w26313 | w26315 ;
  assign w26317 = ~\pi081 & w26316 ;
  assign w26318 = ~w25983 & w26104 ;
  assign w26319 = w26105 ^ w26318 ;
  assign w26320 = ~w26178 & w26319 ;
  assign w26321 = ( w25976 & w26176 ) | ( w25976 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26322 = ~w26177 & w26321 ;
  assign w26323 = w26320 | w26322 ;
  assign w26324 = ~\pi080 & w26323 ;
  assign w26325 = ~w25989 & w26101 ;
  assign w26326 = w26102 ^ w26325 ;
  assign w26327 = ~w26178 & w26326 ;
  assign w26328 = ( w25982 & w26176 ) | ( w25982 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26329 = ~w26177 & w26328 ;
  assign w26330 = w26327 | w26329 ;
  assign w26331 = ~\pi079 & w26330 ;
  assign w26332 = ~w25995 & w26098 ;
  assign w26333 = w26099 ^ w26332 ;
  assign w26334 = ~w26178 & w26333 ;
  assign w26335 = ( w25988 & w26176 ) | ( w25988 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26336 = ~w26177 & w26335 ;
  assign w26337 = w26334 | w26336 ;
  assign w26338 = ~\pi078 & w26337 ;
  assign w26339 = ~w26001 & w26095 ;
  assign w26340 = w26096 ^ w26339 ;
  assign w26341 = ~w26178 & w26340 ;
  assign w26342 = ( w25994 & w26176 ) | ( w25994 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26343 = ~w26177 & w26342 ;
  assign w26344 = w26341 | w26343 ;
  assign w26345 = ~\pi077 & w26344 ;
  assign w26346 = ~w26007 & w26092 ;
  assign w26347 = w26093 ^ w26346 ;
  assign w26348 = ~w26178 & w26347 ;
  assign w26349 = ( w26000 & w26176 ) | ( w26000 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26350 = ~w26177 & w26349 ;
  assign w26351 = w26348 | w26350 ;
  assign w26352 = ~\pi076 & w26351 ;
  assign w26353 = ~w26013 & w26089 ;
  assign w26354 = w26090 ^ w26353 ;
  assign w26355 = ~w26178 & w26354 ;
  assign w26356 = ( w26006 & w26176 ) | ( w26006 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26357 = ~w26177 & w26356 ;
  assign w26358 = w26355 | w26357 ;
  assign w26359 = ~\pi075 & w26358 ;
  assign w26360 = ~w26019 & w26086 ;
  assign w26361 = w26087 ^ w26360 ;
  assign w26362 = ~w26178 & w26361 ;
  assign w26363 = ( w26012 & w26176 ) | ( w26012 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26364 = ~w26177 & w26363 ;
  assign w26365 = w26362 | w26364 ;
  assign w26366 = ~\pi074 & w26365 ;
  assign w26367 = ~w26025 & w26083 ;
  assign w26368 = w26084 ^ w26367 ;
  assign w26369 = ~w26178 & w26368 ;
  assign w26370 = ( w26018 & w26176 ) | ( w26018 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26371 = ~w26177 & w26370 ;
  assign w26372 = w26369 | w26371 ;
  assign w26373 = ~\pi073 & w26372 ;
  assign w26374 = ~w26031 & w26080 ;
  assign w26375 = w26081 ^ w26374 ;
  assign w26376 = ~w26178 & w26375 ;
  assign w26377 = ( w26024 & w26176 ) | ( w26024 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26378 = ~w26177 & w26377 ;
  assign w26379 = w26376 | w26378 ;
  assign w26380 = ~\pi072 & w26379 ;
  assign w26381 = ~w26037 & w26077 ;
  assign w26382 = w26078 ^ w26381 ;
  assign w26383 = ~w26178 & w26382 ;
  assign w26384 = ( w26030 & w26176 ) | ( w26030 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26385 = ~w26177 & w26384 ;
  assign w26386 = w26383 | w26385 ;
  assign w26387 = ~\pi071 & w26386 ;
  assign w26388 = ~w26043 & w26074 ;
  assign w26389 = w26075 ^ w26388 ;
  assign w26390 = ~w26178 & w26389 ;
  assign w26391 = ( w26036 & w26176 ) | ( w26036 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26392 = ~w26177 & w26391 ;
  assign w26393 = w26390 | w26392 ;
  assign w26394 = ~\pi070 & w26393 ;
  assign w26395 = ~w26050 & w26071 ;
  assign w26396 = w26072 ^ w26395 ;
  assign w26397 = ~w26178 & w26396 ;
  assign w26398 = ( w26042 & w26176 ) | ( w26042 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26399 = ~w26177 & w26398 ;
  assign w26400 = w26397 | w26399 ;
  assign w26401 = ~\pi069 & w26400 ;
  assign w26402 = ~w26058 & w26068 ;
  assign w26403 = w26069 ^ w26402 ;
  assign w26404 = ~w26178 & w26403 ;
  assign w26405 = ( w26049 & w26176 ) | ( w26049 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26406 = ~w26177 & w26405 ;
  assign w26407 = w26404 | w26406 ;
  assign w26408 = ~\pi068 & w26407 ;
  assign w26409 = ( \pi065 & w26062 ) | ( \pi065 & ~w26178 ) | ( w26062 & ~w26178 ) ;
  assign w26410 = ( \pi065 & w26064 ) | ( \pi065 & ~w26409 ) | ( w26064 & ~w26409 ) ;
  assign w26411 = w26065 ^ w26410 ;
  assign w26412 = ~w26178 & w26411 ;
  assign w26413 = ( w26057 & w26176 ) | ( w26057 & w26177 ) | ( w26176 & w26177 ) ;
  assign w26414 = ~w26177 & w26413 ;
  assign w26415 = w26412 | w26414 ;
  assign w26416 = ~\pi067 & w26415 ;
  assign w26417 = w6594 ^ w26062 ;
  assign w26418 = \pi065 ^ w26417 ;
  assign w26419 = w26178 ^ w26418 ;
  assign w26420 = ( w26062 & w26418 ) | ( w26062 & w26419 ) | ( w26418 & w26419 ) ;
  assign w26421 = ~\pi066 & w26420 ;
  assign w26422 = w26062 ^ w26178 ;
  assign w26423 = ( w26062 & w26418 ) | ( w26062 & ~w26422 ) | ( w26418 & ~w26422 ) ;
  assign w26424 = \pi066 ^ w26423 ;
  assign w26425 = ( \pi064 & ~w26178 ) | ( \pi064 & w26424 ) | ( ~w26178 & w26424 ) ;
  assign w26426 = \pi028 ^ w26425 ;
  assign w26427 = ( \pi065 & w7271 ) | ( \pi065 & ~w26426 ) | ( w7271 & ~w26426 ) ;
  assign w26428 = w26424 | w26427 ;
  assign w26429 = \pi067 ^ w26415 ;
  assign w26430 = ( ~w26421 & w26428 ) | ( ~w26421 & w26429 ) | ( w26428 & w26429 ) ;
  assign w26431 = w26429 | w26430 ;
  assign w26432 = \pi068 ^ w26407 ;
  assign w26433 = ( ~w26416 & w26431 ) | ( ~w26416 & w26432 ) | ( w26431 & w26432 ) ;
  assign w26434 = w26432 | w26433 ;
  assign w26435 = \pi069 ^ w26400 ;
  assign w26436 = ( ~w26408 & w26434 ) | ( ~w26408 & w26435 ) | ( w26434 & w26435 ) ;
  assign w26437 = w26435 | w26436 ;
  assign w26438 = \pi070 ^ w26393 ;
  assign w26439 = ( ~w26401 & w26437 ) | ( ~w26401 & w26438 ) | ( w26437 & w26438 ) ;
  assign w26440 = w26438 | w26439 ;
  assign w26441 = \pi071 ^ w26386 ;
  assign w26442 = ( ~w26394 & w26440 ) | ( ~w26394 & w26441 ) | ( w26440 & w26441 ) ;
  assign w26443 = w26441 | w26442 ;
  assign w26444 = \pi072 ^ w26379 ;
  assign w26445 = ( ~w26387 & w26443 ) | ( ~w26387 & w26444 ) | ( w26443 & w26444 ) ;
  assign w26446 = w26444 | w26445 ;
  assign w26447 = \pi073 ^ w26372 ;
  assign w26448 = ( ~w26380 & w26446 ) | ( ~w26380 & w26447 ) | ( w26446 & w26447 ) ;
  assign w26449 = w26447 | w26448 ;
  assign w26450 = \pi074 ^ w26365 ;
  assign w26451 = ( ~w26373 & w26449 ) | ( ~w26373 & w26450 ) | ( w26449 & w26450 ) ;
  assign w26452 = w26450 | w26451 ;
  assign w26453 = \pi075 ^ w26358 ;
  assign w26454 = ( ~w26366 & w26452 ) | ( ~w26366 & w26453 ) | ( w26452 & w26453 ) ;
  assign w26455 = w26453 | w26454 ;
  assign w26456 = \pi076 ^ w26351 ;
  assign w26457 = ( ~w26359 & w26455 ) | ( ~w26359 & w26456 ) | ( w26455 & w26456 ) ;
  assign w26458 = w26456 | w26457 ;
  assign w26459 = \pi077 ^ w26344 ;
  assign w26460 = ( ~w26352 & w26458 ) | ( ~w26352 & w26459 ) | ( w26458 & w26459 ) ;
  assign w26461 = w26459 | w26460 ;
  assign w26462 = \pi078 ^ w26337 ;
  assign w26463 = ( ~w26345 & w26461 ) | ( ~w26345 & w26462 ) | ( w26461 & w26462 ) ;
  assign w26464 = w26462 | w26463 ;
  assign w26465 = \pi079 ^ w26330 ;
  assign w26466 = ( ~w26338 & w26464 ) | ( ~w26338 & w26465 ) | ( w26464 & w26465 ) ;
  assign w26467 = w26465 | w26466 ;
  assign w26468 = \pi080 ^ w26323 ;
  assign w26469 = ( ~w26331 & w26467 ) | ( ~w26331 & w26468 ) | ( w26467 & w26468 ) ;
  assign w26470 = w26468 | w26469 ;
  assign w26471 = \pi081 ^ w26316 ;
  assign w26472 = ( ~w26324 & w26470 ) | ( ~w26324 & w26471 ) | ( w26470 & w26471 ) ;
  assign w26473 = w26471 | w26472 ;
  assign w26474 = \pi082 ^ w26309 ;
  assign w26475 = ( ~w26317 & w26473 ) | ( ~w26317 & w26474 ) | ( w26473 & w26474 ) ;
  assign w26476 = w26474 | w26475 ;
  assign w26477 = \pi083 ^ w26302 ;
  assign w26478 = ( ~w26310 & w26476 ) | ( ~w26310 & w26477 ) | ( w26476 & w26477 ) ;
  assign w26479 = w26477 | w26478 ;
  assign w26480 = \pi084 ^ w26295 ;
  assign w26481 = ( ~w26303 & w26479 ) | ( ~w26303 & w26480 ) | ( w26479 & w26480 ) ;
  assign w26482 = w26480 | w26481 ;
  assign w26483 = \pi085 ^ w26288 ;
  assign w26484 = ( ~w26296 & w26482 ) | ( ~w26296 & w26483 ) | ( w26482 & w26483 ) ;
  assign w26485 = w26483 | w26484 ;
  assign w26486 = \pi086 ^ w26281 ;
  assign w26487 = ( ~w26289 & w26485 ) | ( ~w26289 & w26486 ) | ( w26485 & w26486 ) ;
  assign w26488 = w26486 | w26487 ;
  assign w26489 = \pi087 ^ w26274 ;
  assign w26490 = ( ~w26282 & w26488 ) | ( ~w26282 & w26489 ) | ( w26488 & w26489 ) ;
  assign w26491 = w26489 | w26490 ;
  assign w26492 = \pi088 ^ w26267 ;
  assign w26493 = ( ~w26275 & w26491 ) | ( ~w26275 & w26492 ) | ( w26491 & w26492 ) ;
  assign w26494 = w26492 | w26493 ;
  assign w26495 = \pi089 ^ w26260 ;
  assign w26496 = ( ~w26268 & w26494 ) | ( ~w26268 & w26495 ) | ( w26494 & w26495 ) ;
  assign w26497 = w26495 | w26496 ;
  assign w26498 = \pi090 ^ w26253 ;
  assign w26499 = ( ~w26261 & w26497 ) | ( ~w26261 & w26498 ) | ( w26497 & w26498 ) ;
  assign w26500 = w26498 | w26499 ;
  assign w26501 = \pi091 ^ w26246 ;
  assign w26502 = ( ~w26254 & w26500 ) | ( ~w26254 & w26501 ) | ( w26500 & w26501 ) ;
  assign w26503 = w26501 | w26502 ;
  assign w26504 = \pi092 ^ w26239 ;
  assign w26505 = ( ~w26247 & w26503 ) | ( ~w26247 & w26504 ) | ( w26503 & w26504 ) ;
  assign w26506 = w26504 | w26505 ;
  assign w26507 = \pi093 ^ w26232 ;
  assign w26508 = ( ~w26240 & w26506 ) | ( ~w26240 & w26507 ) | ( w26506 & w26507 ) ;
  assign w26509 = w26507 | w26508 ;
  assign w26510 = \pi094 ^ w26225 ;
  assign w26511 = ( ~w26233 & w26509 ) | ( ~w26233 & w26510 ) | ( w26509 & w26510 ) ;
  assign w26512 = w26510 | w26511 ;
  assign w26513 = \pi095 ^ w26218 ;
  assign w26514 = ( ~w26226 & w26512 ) | ( ~w26226 & w26513 ) | ( w26512 & w26513 ) ;
  assign w26515 = w26513 | w26514 ;
  assign w26516 = \pi096 ^ w26211 ;
  assign w26517 = ( ~w26219 & w26515 ) | ( ~w26219 & w26516 ) | ( w26515 & w26516 ) ;
  assign w26518 = w26516 | w26517 ;
  assign w26519 = \pi097 ^ w26204 ;
  assign w26520 = ( ~w26212 & w26518 ) | ( ~w26212 & w26519 ) | ( w26518 & w26519 ) ;
  assign w26521 = w26519 | w26520 ;
  assign w26522 = \pi098 ^ w26197 ;
  assign w26523 = ( ~w26205 & w26521 ) | ( ~w26205 & w26522 ) | ( w26521 & w26522 ) ;
  assign w26524 = w26522 | w26523 ;
  assign w26525 = \pi099 ^ w26184 ;
  assign w26526 = ( ~w26198 & w26524 ) | ( ~w26198 & w26525 ) | ( w26524 & w26525 ) ;
  assign w26527 = w26525 | w26526 ;
  assign w26528 = \pi100 ^ w26190 ;
  assign w26529 = w26191 & ~w26528 ;
  assign w26530 = ( w26527 & w26528 ) | ( w26527 & ~w26529 ) | ( w26528 & ~w26529 ) ;
  assign w26531 = ~\pi100 & w26190 ;
  assign w26532 = w26530 & ~w26531 ;
  assign w26533 = w452 | w26532 ;
  assign w26534 = w26184 & w26533 ;
  assign w26535 = ~w26198 & w26524 ;
  assign w26536 = w26525 ^ w26535 ;
  assign w26537 = ~w26533 & w26536 ;
  assign w26538 = w26534 | w26537 ;
  assign w26539 = w26190 & w26533 ;
  assign w26540 = ~w26191 & w26527 ;
  assign w26541 = w26528 ^ w26540 ;
  assign w26542 = ~w26533 & w26541 ;
  assign w26543 = w26539 | w26542 ;
  assign w26544 = ~\pi100 & w26538 ;
  assign w26545 = w26197 & w26533 ;
  assign w26546 = ~w26205 & w26521 ;
  assign w26547 = w26522 ^ w26546 ;
  assign w26548 = ~w26533 & w26547 ;
  assign w26549 = w26545 | w26548 ;
  assign w26550 = ~\pi099 & w26549 ;
  assign w26551 = w26204 & w26533 ;
  assign w26552 = ~w26212 & w26518 ;
  assign w26553 = w26519 ^ w26552 ;
  assign w26554 = ~w26533 & w26553 ;
  assign w26555 = w26551 | w26554 ;
  assign w26556 = ~\pi098 & w26555 ;
  assign w26557 = w26211 & w26533 ;
  assign w26558 = ~w26219 & w26515 ;
  assign w26559 = w26516 ^ w26558 ;
  assign w26560 = ~w26533 & w26559 ;
  assign w26561 = w26557 | w26560 ;
  assign w26562 = ~\pi097 & w26561 ;
  assign w26563 = w26218 & w26533 ;
  assign w26564 = ~w26226 & w26512 ;
  assign w26565 = w26513 ^ w26564 ;
  assign w26566 = ~w26533 & w26565 ;
  assign w26567 = w26563 | w26566 ;
  assign w26568 = ~\pi096 & w26567 ;
  assign w26569 = w26225 & w26533 ;
  assign w26570 = ~w26233 & w26509 ;
  assign w26571 = w26510 ^ w26570 ;
  assign w26572 = ~w26533 & w26571 ;
  assign w26573 = w26569 | w26572 ;
  assign w26574 = ~\pi095 & w26573 ;
  assign w26575 = w26232 & w26533 ;
  assign w26576 = ~w26240 & w26506 ;
  assign w26577 = w26507 ^ w26576 ;
  assign w26578 = ~w26533 & w26577 ;
  assign w26579 = w26575 | w26578 ;
  assign w26580 = ~\pi094 & w26579 ;
  assign w26581 = w26239 & w26533 ;
  assign w26582 = ~w26247 & w26503 ;
  assign w26583 = w26504 ^ w26582 ;
  assign w26584 = ~w26533 & w26583 ;
  assign w26585 = w26581 | w26584 ;
  assign w26586 = ~\pi093 & w26585 ;
  assign w26587 = w26246 & w26533 ;
  assign w26588 = ~w26254 & w26500 ;
  assign w26589 = w26501 ^ w26588 ;
  assign w26590 = ~w26533 & w26589 ;
  assign w26591 = w26587 | w26590 ;
  assign w26592 = ~\pi092 & w26591 ;
  assign w26593 = w26253 & w26533 ;
  assign w26594 = ~w26261 & w26497 ;
  assign w26595 = w26498 ^ w26594 ;
  assign w26596 = ~w26533 & w26595 ;
  assign w26597 = w26593 | w26596 ;
  assign w26598 = ~\pi091 & w26597 ;
  assign w26599 = w26260 & w26533 ;
  assign w26600 = ~w26268 & w26494 ;
  assign w26601 = w26495 ^ w26600 ;
  assign w26602 = ~w26533 & w26601 ;
  assign w26603 = w26599 | w26602 ;
  assign w26604 = ~\pi090 & w26603 ;
  assign w26605 = w26267 & w26533 ;
  assign w26606 = ~w26275 & w26491 ;
  assign w26607 = w26492 ^ w26606 ;
  assign w26608 = ~w26533 & w26607 ;
  assign w26609 = w26605 | w26608 ;
  assign w26610 = ~\pi089 & w26609 ;
  assign w26611 = w26274 & w26533 ;
  assign w26612 = ~w26282 & w26488 ;
  assign w26613 = w26489 ^ w26612 ;
  assign w26614 = ~w26533 & w26613 ;
  assign w26615 = w26611 | w26614 ;
  assign w26616 = ~\pi088 & w26615 ;
  assign w26617 = w26281 & w26533 ;
  assign w26618 = ~w26289 & w26485 ;
  assign w26619 = w26486 ^ w26618 ;
  assign w26620 = ~w26533 & w26619 ;
  assign w26621 = w26617 | w26620 ;
  assign w26622 = ~\pi087 & w26621 ;
  assign w26623 = w26288 & w26533 ;
  assign w26624 = ~w26296 & w26482 ;
  assign w26625 = w26483 ^ w26624 ;
  assign w26626 = ~w26533 & w26625 ;
  assign w26627 = w26623 | w26626 ;
  assign w26628 = ~\pi086 & w26627 ;
  assign w26629 = w26295 & w26533 ;
  assign w26630 = ~w26303 & w26479 ;
  assign w26631 = w26480 ^ w26630 ;
  assign w26632 = ~w26533 & w26631 ;
  assign w26633 = w26629 | w26632 ;
  assign w26634 = ~\pi085 & w26633 ;
  assign w26635 = w26302 & w26533 ;
  assign w26636 = ~w26310 & w26476 ;
  assign w26637 = w26477 ^ w26636 ;
  assign w26638 = ~w26533 & w26637 ;
  assign w26639 = w26635 | w26638 ;
  assign w26640 = ~\pi084 & w26639 ;
  assign w26641 = w26309 & w26533 ;
  assign w26642 = ~w26317 & w26473 ;
  assign w26643 = w26474 ^ w26642 ;
  assign w26644 = ~w26533 & w26643 ;
  assign w26645 = w26641 | w26644 ;
  assign w26646 = ~\pi083 & w26645 ;
  assign w26647 = w26316 & w26533 ;
  assign w26648 = ~w26324 & w26470 ;
  assign w26649 = w26471 ^ w26648 ;
  assign w26650 = ~w26533 & w26649 ;
  assign w26651 = w26647 | w26650 ;
  assign w26652 = ~\pi082 & w26651 ;
  assign w26653 = w26323 & w26533 ;
  assign w26654 = ~w26331 & w26467 ;
  assign w26655 = w26468 ^ w26654 ;
  assign w26656 = ~w26533 & w26655 ;
  assign w26657 = w26653 | w26656 ;
  assign w26658 = ~\pi081 & w26657 ;
  assign w26659 = w26330 & w26533 ;
  assign w26660 = ~w26338 & w26464 ;
  assign w26661 = w26465 ^ w26660 ;
  assign w26662 = ~w26533 & w26661 ;
  assign w26663 = w26659 | w26662 ;
  assign w26664 = ~\pi080 & w26663 ;
  assign w26665 = w26337 & w26533 ;
  assign w26666 = ~w26345 & w26461 ;
  assign w26667 = w26462 ^ w26666 ;
  assign w26668 = ~w26533 & w26667 ;
  assign w26669 = w26665 | w26668 ;
  assign w26670 = ~\pi079 & w26669 ;
  assign w26671 = w26344 & w26533 ;
  assign w26672 = ~w26352 & w26458 ;
  assign w26673 = w26459 ^ w26672 ;
  assign w26674 = ~w26533 & w26673 ;
  assign w26675 = w26671 | w26674 ;
  assign w26676 = ~\pi078 & w26675 ;
  assign w26677 = w26351 & w26533 ;
  assign w26678 = ~w26359 & w26455 ;
  assign w26679 = w26456 ^ w26678 ;
  assign w26680 = ~w26533 & w26679 ;
  assign w26681 = w26677 | w26680 ;
  assign w26682 = ~\pi077 & w26681 ;
  assign w26683 = w26358 & w26533 ;
  assign w26684 = ~w26366 & w26452 ;
  assign w26685 = w26453 ^ w26684 ;
  assign w26686 = ~w26533 & w26685 ;
  assign w26687 = w26683 | w26686 ;
  assign w26688 = ~\pi076 & w26687 ;
  assign w26689 = w26365 & w26533 ;
  assign w26690 = ~w26373 & w26449 ;
  assign w26691 = w26450 ^ w26690 ;
  assign w26692 = ~w26533 & w26691 ;
  assign w26693 = w26689 | w26692 ;
  assign w26694 = ~\pi075 & w26693 ;
  assign w26695 = w26372 & w26533 ;
  assign w26696 = ~w26380 & w26446 ;
  assign w26697 = w26447 ^ w26696 ;
  assign w26698 = ~w26533 & w26697 ;
  assign w26699 = w26695 | w26698 ;
  assign w26700 = ~\pi074 & w26699 ;
  assign w26701 = w26379 & w26533 ;
  assign w26702 = ~w26387 & w26443 ;
  assign w26703 = w26444 ^ w26702 ;
  assign w26704 = ~w26533 & w26703 ;
  assign w26705 = w26701 | w26704 ;
  assign w26706 = ~\pi073 & w26705 ;
  assign w26707 = w26386 & w26533 ;
  assign w26708 = ~w26394 & w26440 ;
  assign w26709 = w26441 ^ w26708 ;
  assign w26710 = ~w26533 & w26709 ;
  assign w26711 = w26707 | w26710 ;
  assign w26712 = ~\pi072 & w26711 ;
  assign w26713 = w26393 & w26533 ;
  assign w26714 = ~w26401 & w26437 ;
  assign w26715 = w26438 ^ w26714 ;
  assign w26716 = ~w26533 & w26715 ;
  assign w26717 = w26713 | w26716 ;
  assign w26718 = ~\pi071 & w26717 ;
  assign w26719 = w26400 & w26533 ;
  assign w26720 = ~w26408 & w26434 ;
  assign w26721 = w26435 ^ w26720 ;
  assign w26722 = ~w26533 & w26721 ;
  assign w26723 = w26719 | w26722 ;
  assign w26724 = ~\pi070 & w26723 ;
  assign w26725 = w26407 & w26533 ;
  assign w26726 = ~w26416 & w26431 ;
  assign w26727 = w26432 ^ w26726 ;
  assign w26728 = ~w26533 & w26727 ;
  assign w26729 = w26725 | w26728 ;
  assign w26730 = ~\pi069 & w26729 ;
  assign w26731 = w26415 & w26533 ;
  assign w26732 = ~w26421 & w26428 ;
  assign w26733 = w26429 ^ w26732 ;
  assign w26734 = ~w26533 & w26733 ;
  assign w26735 = w26731 | w26734 ;
  assign w26736 = ~\pi068 & w26735 ;
  assign w26737 = w26420 & w26533 ;
  assign w26738 = \pi064 & ~w26178 ;
  assign w26739 = \pi028 ^ w26738 ;
  assign w26740 = ( \pi065 & w7271 ) | ( \pi065 & ~w26739 ) | ( w7271 & ~w26739 ) ;
  assign w26741 = w26424 ^ w26740 ;
  assign w26742 = ( w452 & w26532 ) | ( w452 & w26741 ) | ( w26532 & w26741 ) ;
  assign w26743 = w26741 & ~w26742 ;
  assign w26744 = w26737 | w26743 ;
  assign w26745 = ~\pi067 & w26744 ;
  assign w26746 = \pi027 ^ w26178 ;
  assign w26747 = ( \pi064 & w452 ) | ( \pi064 & w26746 ) | ( w452 & w26746 ) ;
  assign w26748 = w7278 ^ w26747 ;
  assign w26749 = ~w452 & w26748 ;
  assign w26750 = ~w26532 & w26749 ;
  assign w26751 = ( ~\pi064 & w26178 ) | ( ~\pi064 & w26533 ) | ( w26178 & w26533 ) ;
  assign w26752 = \pi028 ^ w26751 ;
  assign w26753 = w26533 & ~w26752 ;
  assign w26754 = w26750 | w26753 ;
  assign w26755 = ~\pi066 & w26754 ;
  assign w26756 = ( \pi027 & ~w7294 ) | ( \pi027 & w26532 ) | ( ~w7294 & w26532 ) ;
  assign w26757 = \pi027 & w26756 ;
  assign w26758 = w275 | w26532 ;
  assign w26759 = w7299 & ~w26758 ;
  assign w26760 = ~w7297 & w26759 ;
  assign w26761 = w26533 | w26750 ;
  assign w26762 = ( w26739 & w26750 ) | ( w26739 & w26761 ) | ( w26750 & w26761 ) ;
  assign w26763 = \pi066 ^ w26762 ;
  assign w26764 = w26757 | w26760 ;
  assign w26765 = ( \pi065 & w7302 ) | ( \pi065 & ~w26764 ) | ( w7302 & ~w26764 ) ;
  assign w26766 = w26763 | w26765 ;
  assign w26767 = \pi067 ^ w26744 ;
  assign w26768 = ( ~w26755 & w26766 ) | ( ~w26755 & w26767 ) | ( w26766 & w26767 ) ;
  assign w26769 = w26767 | w26768 ;
  assign w26770 = \pi068 ^ w26735 ;
  assign w26771 = ( ~w26745 & w26769 ) | ( ~w26745 & w26770 ) | ( w26769 & w26770 ) ;
  assign w26772 = w26770 | w26771 ;
  assign w26773 = \pi069 ^ w26729 ;
  assign w26774 = ( ~w26736 & w26772 ) | ( ~w26736 & w26773 ) | ( w26772 & w26773 ) ;
  assign w26775 = w26773 | w26774 ;
  assign w26776 = \pi070 ^ w26723 ;
  assign w26777 = ( ~w26730 & w26775 ) | ( ~w26730 & w26776 ) | ( w26775 & w26776 ) ;
  assign w26778 = w26776 | w26777 ;
  assign w26779 = \pi071 ^ w26717 ;
  assign w26780 = ( ~w26724 & w26778 ) | ( ~w26724 & w26779 ) | ( w26778 & w26779 ) ;
  assign w26781 = w26779 | w26780 ;
  assign w26782 = \pi072 ^ w26711 ;
  assign w26783 = ( ~w26718 & w26781 ) | ( ~w26718 & w26782 ) | ( w26781 & w26782 ) ;
  assign w26784 = w26782 | w26783 ;
  assign w26785 = \pi073 ^ w26705 ;
  assign w26786 = ( ~w26712 & w26784 ) | ( ~w26712 & w26785 ) | ( w26784 & w26785 ) ;
  assign w26787 = w26785 | w26786 ;
  assign w26788 = \pi074 ^ w26699 ;
  assign w26789 = ( ~w26706 & w26787 ) | ( ~w26706 & w26788 ) | ( w26787 & w26788 ) ;
  assign w26790 = w26788 | w26789 ;
  assign w26791 = \pi075 ^ w26693 ;
  assign w26792 = ( ~w26700 & w26790 ) | ( ~w26700 & w26791 ) | ( w26790 & w26791 ) ;
  assign w26793 = w26791 | w26792 ;
  assign w26794 = \pi076 ^ w26687 ;
  assign w26795 = ( ~w26694 & w26793 ) | ( ~w26694 & w26794 ) | ( w26793 & w26794 ) ;
  assign w26796 = w26794 | w26795 ;
  assign w26797 = \pi077 ^ w26681 ;
  assign w26798 = ( ~w26688 & w26796 ) | ( ~w26688 & w26797 ) | ( w26796 & w26797 ) ;
  assign w26799 = w26797 | w26798 ;
  assign w26800 = \pi078 ^ w26675 ;
  assign w26801 = ( ~w26682 & w26799 ) | ( ~w26682 & w26800 ) | ( w26799 & w26800 ) ;
  assign w26802 = w26800 | w26801 ;
  assign w26803 = \pi079 ^ w26669 ;
  assign w26804 = ( ~w26676 & w26802 ) | ( ~w26676 & w26803 ) | ( w26802 & w26803 ) ;
  assign w26805 = w26803 | w26804 ;
  assign w26806 = \pi080 ^ w26663 ;
  assign w26807 = ( ~w26670 & w26805 ) | ( ~w26670 & w26806 ) | ( w26805 & w26806 ) ;
  assign w26808 = w26806 | w26807 ;
  assign w26809 = \pi081 ^ w26657 ;
  assign w26810 = ( ~w26664 & w26808 ) | ( ~w26664 & w26809 ) | ( w26808 & w26809 ) ;
  assign w26811 = w26809 | w26810 ;
  assign w26812 = \pi082 ^ w26651 ;
  assign w26813 = ( ~w26658 & w26811 ) | ( ~w26658 & w26812 ) | ( w26811 & w26812 ) ;
  assign w26814 = w26812 | w26813 ;
  assign w26815 = \pi083 ^ w26645 ;
  assign w26816 = ( ~w26652 & w26814 ) | ( ~w26652 & w26815 ) | ( w26814 & w26815 ) ;
  assign w26817 = w26815 | w26816 ;
  assign w26818 = \pi084 ^ w26639 ;
  assign w26819 = ( ~w26646 & w26817 ) | ( ~w26646 & w26818 ) | ( w26817 & w26818 ) ;
  assign w26820 = w26818 | w26819 ;
  assign w26821 = \pi085 ^ w26633 ;
  assign w26822 = ( ~w26640 & w26820 ) | ( ~w26640 & w26821 ) | ( w26820 & w26821 ) ;
  assign w26823 = w26821 | w26822 ;
  assign w26824 = \pi086 ^ w26627 ;
  assign w26825 = ( ~w26634 & w26823 ) | ( ~w26634 & w26824 ) | ( w26823 & w26824 ) ;
  assign w26826 = w26824 | w26825 ;
  assign w26827 = \pi087 ^ w26621 ;
  assign w26828 = ( ~w26628 & w26826 ) | ( ~w26628 & w26827 ) | ( w26826 & w26827 ) ;
  assign w26829 = w26827 | w26828 ;
  assign w26830 = \pi088 ^ w26615 ;
  assign w26831 = ( ~w26622 & w26829 ) | ( ~w26622 & w26830 ) | ( w26829 & w26830 ) ;
  assign w26832 = w26830 | w26831 ;
  assign w26833 = \pi089 ^ w26609 ;
  assign w26834 = ( ~w26616 & w26832 ) | ( ~w26616 & w26833 ) | ( w26832 & w26833 ) ;
  assign w26835 = w26833 | w26834 ;
  assign w26836 = \pi090 ^ w26603 ;
  assign w26837 = ( ~w26610 & w26835 ) | ( ~w26610 & w26836 ) | ( w26835 & w26836 ) ;
  assign w26838 = w26836 | w26837 ;
  assign w26839 = \pi091 ^ w26597 ;
  assign w26840 = ( ~w26604 & w26838 ) | ( ~w26604 & w26839 ) | ( w26838 & w26839 ) ;
  assign w26841 = w26839 | w26840 ;
  assign w26842 = \pi092 ^ w26591 ;
  assign w26843 = ( ~w26598 & w26841 ) | ( ~w26598 & w26842 ) | ( w26841 & w26842 ) ;
  assign w26844 = w26842 | w26843 ;
  assign w26845 = \pi093 ^ w26585 ;
  assign w26846 = ( ~w26592 & w26844 ) | ( ~w26592 & w26845 ) | ( w26844 & w26845 ) ;
  assign w26847 = w26845 | w26846 ;
  assign w26848 = \pi094 ^ w26579 ;
  assign w26849 = ( ~w26586 & w26847 ) | ( ~w26586 & w26848 ) | ( w26847 & w26848 ) ;
  assign w26850 = w26848 | w26849 ;
  assign w26851 = \pi095 ^ w26573 ;
  assign w26852 = ( ~w26580 & w26850 ) | ( ~w26580 & w26851 ) | ( w26850 & w26851 ) ;
  assign w26853 = w26851 | w26852 ;
  assign w26854 = \pi096 ^ w26567 ;
  assign w26855 = ( ~w26574 & w26853 ) | ( ~w26574 & w26854 ) | ( w26853 & w26854 ) ;
  assign w26856 = w26854 | w26855 ;
  assign w26857 = \pi097 ^ w26561 ;
  assign w26858 = ( ~w26568 & w26856 ) | ( ~w26568 & w26857 ) | ( w26856 & w26857 ) ;
  assign w26859 = w26857 | w26858 ;
  assign w26860 = \pi098 ^ w26555 ;
  assign w26861 = ( ~w26562 & w26859 ) | ( ~w26562 & w26860 ) | ( w26859 & w26860 ) ;
  assign w26862 = w26860 | w26861 ;
  assign w26863 = \pi099 ^ w26549 ;
  assign w26864 = ( ~w26556 & w26862 ) | ( ~w26556 & w26863 ) | ( w26862 & w26863 ) ;
  assign w26865 = w26863 | w26864 ;
  assign w26866 = \pi100 ^ w26538 ;
  assign w26867 = ( ~w26550 & w26865 ) | ( ~w26550 & w26866 ) | ( w26865 & w26866 ) ;
  assign w26868 = w26866 | w26867 ;
  assign w26869 = \pi101 ^ w26543 ;
  assign w26870 = w26544 & ~w26869 ;
  assign w26871 = ( w26868 & w26869 ) | ( w26868 & ~w26870 ) | ( w26869 & ~w26870 ) ;
  assign w26872 = ~\pi101 & w26543 ;
  assign w26873 = w26871 & ~w26872 ;
  assign w26874 = w7419 | w26873 ;
  assign w26875 = w26538 & w26874 ;
  assign w26876 = ~w26550 & w26865 ;
  assign w26877 = w26866 ^ w26876 ;
  assign w26878 = ~w26874 & w26877 ;
  assign w26879 = w26875 | w26878 ;
  assign w26880 = ~\pi101 & w26879 ;
  assign w26881 = w26549 & w26874 ;
  assign w26882 = ~w26556 & w26862 ;
  assign w26883 = w26863 ^ w26882 ;
  assign w26884 = ~w26874 & w26883 ;
  assign w26885 = w26881 | w26884 ;
  assign w26886 = ~\pi100 & w26885 ;
  assign w26887 = w26555 & w26874 ;
  assign w26888 = ~w26562 & w26859 ;
  assign w26889 = w26860 ^ w26888 ;
  assign w26890 = ~w26874 & w26889 ;
  assign w26891 = w26887 | w26890 ;
  assign w26892 = ~\pi099 & w26891 ;
  assign w26893 = w26561 & w26874 ;
  assign w26894 = ~w26568 & w26856 ;
  assign w26895 = w26857 ^ w26894 ;
  assign w26896 = ~w26874 & w26895 ;
  assign w26897 = w26893 | w26896 ;
  assign w26898 = ~\pi098 & w26897 ;
  assign w26899 = w26567 & w26874 ;
  assign w26900 = ~w26574 & w26853 ;
  assign w26901 = w26854 ^ w26900 ;
  assign w26902 = ~w26874 & w26901 ;
  assign w26903 = w26899 | w26902 ;
  assign w26904 = ~\pi097 & w26903 ;
  assign w26905 = w26573 & w26874 ;
  assign w26906 = ~w26580 & w26850 ;
  assign w26907 = w26851 ^ w26906 ;
  assign w26908 = ~w26874 & w26907 ;
  assign w26909 = w26905 | w26908 ;
  assign w26910 = ~\pi096 & w26909 ;
  assign w26911 = w26579 & w26874 ;
  assign w26912 = ~w26586 & w26847 ;
  assign w26913 = w26848 ^ w26912 ;
  assign w26914 = ~w26874 & w26913 ;
  assign w26915 = w26911 | w26914 ;
  assign w26916 = ~\pi095 & w26915 ;
  assign w26917 = w26585 & w26874 ;
  assign w26918 = ~w26592 & w26844 ;
  assign w26919 = w26845 ^ w26918 ;
  assign w26920 = ~w26874 & w26919 ;
  assign w26921 = w26917 | w26920 ;
  assign w26922 = ~\pi094 & w26921 ;
  assign w26923 = w26591 & w26874 ;
  assign w26924 = ~w26598 & w26841 ;
  assign w26925 = w26842 ^ w26924 ;
  assign w26926 = ~w26874 & w26925 ;
  assign w26927 = w26923 | w26926 ;
  assign w26928 = ~\pi093 & w26927 ;
  assign w26929 = w26597 & w26874 ;
  assign w26930 = ~w26604 & w26838 ;
  assign w26931 = w26839 ^ w26930 ;
  assign w26932 = ~w26874 & w26931 ;
  assign w26933 = w26929 | w26932 ;
  assign w26934 = ~\pi092 & w26933 ;
  assign w26935 = w26603 & w26874 ;
  assign w26936 = ~w26610 & w26835 ;
  assign w26937 = w26836 ^ w26936 ;
  assign w26938 = ~w26874 & w26937 ;
  assign w26939 = w26935 | w26938 ;
  assign w26940 = ~\pi091 & w26939 ;
  assign w26941 = w26609 & w26874 ;
  assign w26942 = ~w26616 & w26832 ;
  assign w26943 = w26833 ^ w26942 ;
  assign w26944 = ~w26874 & w26943 ;
  assign w26945 = w26941 | w26944 ;
  assign w26946 = ~\pi090 & w26945 ;
  assign w26947 = w26615 & w26874 ;
  assign w26948 = ~w26622 & w26829 ;
  assign w26949 = w26830 ^ w26948 ;
  assign w26950 = ~w26874 & w26949 ;
  assign w26951 = w26947 | w26950 ;
  assign w26952 = ~\pi089 & w26951 ;
  assign w26953 = w26621 & w26874 ;
  assign w26954 = ~w26628 & w26826 ;
  assign w26955 = w26827 ^ w26954 ;
  assign w26956 = ~w26874 & w26955 ;
  assign w26957 = w26953 | w26956 ;
  assign w26958 = ~\pi088 & w26957 ;
  assign w26959 = w26627 & w26874 ;
  assign w26960 = ~w26634 & w26823 ;
  assign w26961 = w26824 ^ w26960 ;
  assign w26962 = ~w26874 & w26961 ;
  assign w26963 = w26959 | w26962 ;
  assign w26964 = ~\pi087 & w26963 ;
  assign w26965 = w26633 & w26874 ;
  assign w26966 = ~w26640 & w26820 ;
  assign w26967 = w26821 ^ w26966 ;
  assign w26968 = ~w26874 & w26967 ;
  assign w26969 = w26965 | w26968 ;
  assign w26970 = ~\pi086 & w26969 ;
  assign w26971 = w26639 & w26874 ;
  assign w26972 = ~w26646 & w26817 ;
  assign w26973 = w26818 ^ w26972 ;
  assign w26974 = ~w26874 & w26973 ;
  assign w26975 = w26971 | w26974 ;
  assign w26976 = ~\pi085 & w26975 ;
  assign w26977 = w26645 & w26874 ;
  assign w26978 = ~w26652 & w26814 ;
  assign w26979 = w26815 ^ w26978 ;
  assign w26980 = ~w26874 & w26979 ;
  assign w26981 = w26977 | w26980 ;
  assign w26982 = ~\pi084 & w26981 ;
  assign w26983 = w26651 & w26874 ;
  assign w26984 = ~w26658 & w26811 ;
  assign w26985 = w26812 ^ w26984 ;
  assign w26986 = ~w26874 & w26985 ;
  assign w26987 = w26983 | w26986 ;
  assign w26988 = ~\pi083 & w26987 ;
  assign w26989 = w26657 & w26874 ;
  assign w26990 = ~w26664 & w26808 ;
  assign w26991 = w26809 ^ w26990 ;
  assign w26992 = ~w26874 & w26991 ;
  assign w26993 = w26989 | w26992 ;
  assign w26994 = ~\pi082 & w26993 ;
  assign w26995 = w26663 & w26874 ;
  assign w26996 = ~w26670 & w26805 ;
  assign w26997 = w26806 ^ w26996 ;
  assign w26998 = ~w26874 & w26997 ;
  assign w26999 = w26995 | w26998 ;
  assign w27000 = ~\pi081 & w26999 ;
  assign w27001 = w26669 & w26874 ;
  assign w27002 = ~w26676 & w26802 ;
  assign w27003 = w26803 ^ w27002 ;
  assign w27004 = ~w26874 & w27003 ;
  assign w27005 = w27001 | w27004 ;
  assign w27006 = ~\pi080 & w27005 ;
  assign w27007 = w26675 & w26874 ;
  assign w27008 = ~w26682 & w26799 ;
  assign w27009 = w26800 ^ w27008 ;
  assign w27010 = ~w26874 & w27009 ;
  assign w27011 = w27007 | w27010 ;
  assign w27012 = ~\pi079 & w27011 ;
  assign w27013 = w26681 & w26874 ;
  assign w27014 = ~w26688 & w26796 ;
  assign w27015 = w26797 ^ w27014 ;
  assign w27016 = ~w26874 & w27015 ;
  assign w27017 = w27013 | w27016 ;
  assign w27018 = ~\pi078 & w27017 ;
  assign w27019 = w26687 & w26874 ;
  assign w27020 = ~w26694 & w26793 ;
  assign w27021 = w26794 ^ w27020 ;
  assign w27022 = ~w26874 & w27021 ;
  assign w27023 = w27019 | w27022 ;
  assign w27024 = ~\pi077 & w27023 ;
  assign w27025 = w26693 & w26874 ;
  assign w27026 = ~w26700 & w26790 ;
  assign w27027 = w26791 ^ w27026 ;
  assign w27028 = ~w26874 & w27027 ;
  assign w27029 = w27025 | w27028 ;
  assign w27030 = ~\pi076 & w27029 ;
  assign w27031 = w26699 & w26874 ;
  assign w27032 = ~w26706 & w26787 ;
  assign w27033 = w26788 ^ w27032 ;
  assign w27034 = ~w26874 & w27033 ;
  assign w27035 = w27031 | w27034 ;
  assign w27036 = ~\pi075 & w27035 ;
  assign w27037 = w26705 & w26874 ;
  assign w27038 = ~w26712 & w26784 ;
  assign w27039 = w26785 ^ w27038 ;
  assign w27040 = ~w26874 & w27039 ;
  assign w27041 = w27037 | w27040 ;
  assign w27042 = ~\pi074 & w27041 ;
  assign w27043 = w26711 & w26874 ;
  assign w27044 = ~w26718 & w26781 ;
  assign w27045 = w26782 ^ w27044 ;
  assign w27046 = ~w26874 & w27045 ;
  assign w27047 = w27043 | w27046 ;
  assign w27048 = ~\pi073 & w27047 ;
  assign w27049 = w26717 & w26874 ;
  assign w27050 = ~w26724 & w26778 ;
  assign w27051 = w26779 ^ w27050 ;
  assign w27052 = ~w26874 & w27051 ;
  assign w27053 = w27049 | w27052 ;
  assign w27054 = ~\pi072 & w27053 ;
  assign w27055 = w26723 & w26874 ;
  assign w27056 = ~w26730 & w26775 ;
  assign w27057 = w26776 ^ w27056 ;
  assign w27058 = ~w26874 & w27057 ;
  assign w27059 = w27055 | w27058 ;
  assign w27060 = ~\pi071 & w27059 ;
  assign w27061 = w26729 & w26874 ;
  assign w27062 = ~w26736 & w26772 ;
  assign w27063 = w26773 ^ w27062 ;
  assign w27064 = ~w26874 & w27063 ;
  assign w27065 = w27061 | w27064 ;
  assign w27066 = ~\pi070 & w27065 ;
  assign w27067 = w26735 & w26874 ;
  assign w27068 = ~w26745 & w26769 ;
  assign w27069 = w26770 ^ w27068 ;
  assign w27070 = ~w26874 & w27069 ;
  assign w27071 = w27067 | w27070 ;
  assign w27072 = ~\pi069 & w27071 ;
  assign w27073 = w26744 & w26874 ;
  assign w27074 = ~w26755 & w26766 ;
  assign w27075 = w26767 ^ w27074 ;
  assign w27076 = ~w26874 & w27075 ;
  assign w27077 = w27073 | w27076 ;
  assign w27078 = ~\pi068 & w27077 ;
  assign w27079 = w26754 & w26874 ;
  assign w27080 = w26763 ^ w26765 ;
  assign w27081 = ( w7419 & w26873 ) | ( w7419 & w27080 ) | ( w26873 & w27080 ) ;
  assign w27082 = w27080 & ~w27081 ;
  assign w27083 = w27079 | w27082 ;
  assign w27084 = ~\pi067 & w27083 ;
  assign w27085 = ( ~w7419 & w26757 ) | ( ~w7419 & w26760 ) | ( w26757 & w26760 ) ;
  assign w27086 = \pi065 ^ w27085 ;
  assign w27087 = ( w7302 & ~w7419 ) | ( w7302 & w27086 ) | ( ~w7419 & w27086 ) ;
  assign w27088 = ( w7302 & w26873 ) | ( w7302 & w27086 ) | ( w26873 & w27086 ) ;
  assign w27089 = w27087 & ~w27088 ;
  assign w27090 = w26764 & ~w26874 ;
  assign w27091 = ( w26764 & w27089 ) | ( w26764 & ~w27090 ) | ( w27089 & ~w27090 ) ;
  assign w27092 = ~\pi066 & w27091 ;
  assign w27093 = ( \pi026 & ~w7644 ) | ( \pi026 & w26873 ) | ( ~w7644 & w26873 ) ;
  assign w27094 = \pi026 & w27093 ;
  assign w27095 = w7651 & ~w26873 ;
  assign w27096 = w27094 | w27095 ;
  assign w27097 = \pi065 ^ w27096 ;
  assign w27098 = w7654 | w27097 ;
  assign w27099 = \pi066 ^ w27091 ;
  assign w27100 = ~\pi065 & w27096 ;
  assign w27101 = w27098 | w27100 ;
  assign w27102 = ( w27099 & ~w27100 ) | ( w27099 & w27101 ) | ( ~w27100 & w27101 ) ;
  assign w27103 = \pi067 ^ w27083 ;
  assign w27104 = ( ~w27092 & w27102 ) | ( ~w27092 & w27103 ) | ( w27102 & w27103 ) ;
  assign w27105 = w27103 | w27104 ;
  assign w27106 = \pi068 ^ w27077 ;
  assign w27107 = ( ~w27084 & w27105 ) | ( ~w27084 & w27106 ) | ( w27105 & w27106 ) ;
  assign w27108 = w27106 | w27107 ;
  assign w27109 = \pi069 ^ w27071 ;
  assign w27110 = ( ~w27078 & w27108 ) | ( ~w27078 & w27109 ) | ( w27108 & w27109 ) ;
  assign w27111 = w27109 | w27110 ;
  assign w27112 = \pi070 ^ w27065 ;
  assign w27113 = ( ~w27072 & w27111 ) | ( ~w27072 & w27112 ) | ( w27111 & w27112 ) ;
  assign w27114 = w27112 | w27113 ;
  assign w27115 = \pi071 ^ w27059 ;
  assign w27116 = ( ~w27066 & w27114 ) | ( ~w27066 & w27115 ) | ( w27114 & w27115 ) ;
  assign w27117 = w27115 | w27116 ;
  assign w27118 = \pi072 ^ w27053 ;
  assign w27119 = ( ~w27060 & w27117 ) | ( ~w27060 & w27118 ) | ( w27117 & w27118 ) ;
  assign w27120 = w27118 | w27119 ;
  assign w27121 = \pi073 ^ w27047 ;
  assign w27122 = ( ~w27054 & w27120 ) | ( ~w27054 & w27121 ) | ( w27120 & w27121 ) ;
  assign w27123 = w27121 | w27122 ;
  assign w27124 = \pi074 ^ w27041 ;
  assign w27125 = ( ~w27048 & w27123 ) | ( ~w27048 & w27124 ) | ( w27123 & w27124 ) ;
  assign w27126 = w27124 | w27125 ;
  assign w27127 = \pi075 ^ w27035 ;
  assign w27128 = ( ~w27042 & w27126 ) | ( ~w27042 & w27127 ) | ( w27126 & w27127 ) ;
  assign w27129 = w27127 | w27128 ;
  assign w27130 = \pi076 ^ w27029 ;
  assign w27131 = ( ~w27036 & w27129 ) | ( ~w27036 & w27130 ) | ( w27129 & w27130 ) ;
  assign w27132 = w27130 | w27131 ;
  assign w27133 = \pi077 ^ w27023 ;
  assign w27134 = ( ~w27030 & w27132 ) | ( ~w27030 & w27133 ) | ( w27132 & w27133 ) ;
  assign w27135 = w27133 | w27134 ;
  assign w27136 = \pi078 ^ w27017 ;
  assign w27137 = ( ~w27024 & w27135 ) | ( ~w27024 & w27136 ) | ( w27135 & w27136 ) ;
  assign w27138 = w27136 | w27137 ;
  assign w27139 = \pi079 ^ w27011 ;
  assign w27140 = ( ~w27018 & w27138 ) | ( ~w27018 & w27139 ) | ( w27138 & w27139 ) ;
  assign w27141 = w27139 | w27140 ;
  assign w27142 = \pi080 ^ w27005 ;
  assign w27143 = ( ~w27012 & w27141 ) | ( ~w27012 & w27142 ) | ( w27141 & w27142 ) ;
  assign w27144 = w27142 | w27143 ;
  assign w27145 = \pi081 ^ w26999 ;
  assign w27146 = ( ~w27006 & w27144 ) | ( ~w27006 & w27145 ) | ( w27144 & w27145 ) ;
  assign w27147 = w27145 | w27146 ;
  assign w27148 = \pi082 ^ w26993 ;
  assign w27149 = ( ~w27000 & w27147 ) | ( ~w27000 & w27148 ) | ( w27147 & w27148 ) ;
  assign w27150 = w27148 | w27149 ;
  assign w27151 = \pi083 ^ w26987 ;
  assign w27152 = ( ~w26994 & w27150 ) | ( ~w26994 & w27151 ) | ( w27150 & w27151 ) ;
  assign w27153 = w27151 | w27152 ;
  assign w27154 = \pi084 ^ w26981 ;
  assign w27155 = ( ~w26988 & w27153 ) | ( ~w26988 & w27154 ) | ( w27153 & w27154 ) ;
  assign w27156 = w27154 | w27155 ;
  assign w27157 = \pi085 ^ w26975 ;
  assign w27158 = ( ~w26982 & w27156 ) | ( ~w26982 & w27157 ) | ( w27156 & w27157 ) ;
  assign w27159 = w27157 | w27158 ;
  assign w27160 = \pi086 ^ w26969 ;
  assign w27161 = ( ~w26976 & w27159 ) | ( ~w26976 & w27160 ) | ( w27159 & w27160 ) ;
  assign w27162 = w27160 | w27161 ;
  assign w27163 = \pi087 ^ w26963 ;
  assign w27164 = ( ~w26970 & w27162 ) | ( ~w26970 & w27163 ) | ( w27162 & w27163 ) ;
  assign w27165 = w27163 | w27164 ;
  assign w27166 = \pi088 ^ w26957 ;
  assign w27167 = ( ~w26964 & w27165 ) | ( ~w26964 & w27166 ) | ( w27165 & w27166 ) ;
  assign w27168 = w27166 | w27167 ;
  assign w27169 = \pi089 ^ w26951 ;
  assign w27170 = ( ~w26958 & w27168 ) | ( ~w26958 & w27169 ) | ( w27168 & w27169 ) ;
  assign w27171 = w27169 | w27170 ;
  assign w27172 = \pi090 ^ w26945 ;
  assign w27173 = ( ~w26952 & w27171 ) | ( ~w26952 & w27172 ) | ( w27171 & w27172 ) ;
  assign w27174 = w27172 | w27173 ;
  assign w27175 = \pi091 ^ w26939 ;
  assign w27176 = ( ~w26946 & w27174 ) | ( ~w26946 & w27175 ) | ( w27174 & w27175 ) ;
  assign w27177 = w27175 | w27176 ;
  assign w27178 = \pi092 ^ w26933 ;
  assign w27179 = ( ~w26940 & w27177 ) | ( ~w26940 & w27178 ) | ( w27177 & w27178 ) ;
  assign w27180 = w27178 | w27179 ;
  assign w27181 = \pi093 ^ w26927 ;
  assign w27182 = ( ~w26934 & w27180 ) | ( ~w26934 & w27181 ) | ( w27180 & w27181 ) ;
  assign w27183 = w27181 | w27182 ;
  assign w27184 = \pi094 ^ w26921 ;
  assign w27185 = ( ~w26928 & w27183 ) | ( ~w26928 & w27184 ) | ( w27183 & w27184 ) ;
  assign w27186 = w27184 | w27185 ;
  assign w27187 = \pi095 ^ w26915 ;
  assign w27188 = ( ~w26922 & w27186 ) | ( ~w26922 & w27187 ) | ( w27186 & w27187 ) ;
  assign w27189 = w27187 | w27188 ;
  assign w27190 = \pi096 ^ w26909 ;
  assign w27191 = ( ~w26916 & w27189 ) | ( ~w26916 & w27190 ) | ( w27189 & w27190 ) ;
  assign w27192 = w27190 | w27191 ;
  assign w27193 = \pi097 ^ w26903 ;
  assign w27194 = ( ~w26910 & w27192 ) | ( ~w26910 & w27193 ) | ( w27192 & w27193 ) ;
  assign w27195 = w27193 | w27194 ;
  assign w27196 = \pi098 ^ w26897 ;
  assign w27197 = ( ~w26904 & w27195 ) | ( ~w26904 & w27196 ) | ( w27195 & w27196 ) ;
  assign w27198 = w27196 | w27197 ;
  assign w27199 = \pi099 ^ w26891 ;
  assign w27200 = ( ~w26898 & w27198 ) | ( ~w26898 & w27199 ) | ( w27198 & w27199 ) ;
  assign w27201 = w27199 | w27200 ;
  assign w27202 = \pi100 ^ w26885 ;
  assign w27203 = ( ~w26892 & w27201 ) | ( ~w26892 & w27202 ) | ( w27201 & w27202 ) ;
  assign w27204 = w27202 | w27203 ;
  assign w27205 = \pi101 ^ w26879 ;
  assign w27206 = ( ~w26886 & w27204 ) | ( ~w26886 & w27205 ) | ( w27204 & w27205 ) ;
  assign w27207 = w27205 | w27206 ;
  assign w27208 = w26543 & w26874 ;
  assign w27209 = ~w26544 & w26868 ;
  assign w27210 = w26869 ^ w27209 ;
  assign w27211 = ~w26874 & w27210 ;
  assign w27212 = w27208 | w27211 ;
  assign w27213 = ~\pi102 & w27212 ;
  assign w27214 = ( \pi102 & ~w27208 ) | ( \pi102 & w27211 ) | ( ~w27208 & w27211 ) ;
  assign w27215 = ~w27211 & w27214 ;
  assign w27216 = w27213 | w27215 ;
  assign w27217 = ( ~w26880 & w27207 ) | ( ~w26880 & w27216 ) | ( w27207 & w27216 ) ;
  assign w27218 = ( w7777 & ~w27216 ) | ( w7777 & w27217 ) | ( ~w27216 & w27217 ) ;
  assign w27219 = w27216 | w27218 ;
  assign w27220 = ~w7419 & w27212 ;
  assign w27221 = w27219 & ~w27220 ;
  assign w27222 = ~w26886 & w27204 ;
  assign w27223 = w27205 ^ w27222 ;
  assign w27224 = ~w27221 & w27223 ;
  assign w27225 = ( w26879 & w27219 ) | ( w26879 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27226 = ~w27220 & w27225 ;
  assign w27227 = w27224 | w27226 ;
  assign w27228 = ( ~w26880 & w27207 ) | ( ~w26880 & w27221 ) | ( w27207 & w27221 ) ;
  assign w27229 = w27216 ^ w27228 ;
  assign w27230 = ~w27221 & w27229 ;
  assign w27231 = ( w7419 & ~w27212 ) | ( w7419 & w27219 ) | ( ~w27212 & w27219 ) ;
  assign w27232 = w27212 & w27231 ;
  assign w27233 = w27230 | w27232 ;
  assign w27234 = ~\pi102 & w27227 ;
  assign w27235 = ~w26892 & w27201 ;
  assign w27236 = w27202 ^ w27235 ;
  assign w27237 = ~w27221 & w27236 ;
  assign w27238 = ( w26885 & w27219 ) | ( w26885 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27239 = ~w27220 & w27238 ;
  assign w27240 = w27237 | w27239 ;
  assign w27241 = ~\pi101 & w27240 ;
  assign w27242 = ~w26898 & w27198 ;
  assign w27243 = w27199 ^ w27242 ;
  assign w27244 = ~w27221 & w27243 ;
  assign w27245 = ( w26891 & w27219 ) | ( w26891 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27246 = ~w27220 & w27245 ;
  assign w27247 = w27244 | w27246 ;
  assign w27248 = ~\pi100 & w27247 ;
  assign w27249 = ~w26904 & w27195 ;
  assign w27250 = w27196 ^ w27249 ;
  assign w27251 = ~w27221 & w27250 ;
  assign w27252 = ( w26897 & w27219 ) | ( w26897 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27253 = ~w27220 & w27252 ;
  assign w27254 = w27251 | w27253 ;
  assign w27255 = ~\pi099 & w27254 ;
  assign w27256 = ~w26910 & w27192 ;
  assign w27257 = w27193 ^ w27256 ;
  assign w27258 = ~w27221 & w27257 ;
  assign w27259 = ( w26903 & w27219 ) | ( w26903 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27260 = ~w27220 & w27259 ;
  assign w27261 = w27258 | w27260 ;
  assign w27262 = ~\pi098 & w27261 ;
  assign w27263 = ~w26916 & w27189 ;
  assign w27264 = w27190 ^ w27263 ;
  assign w27265 = ~w27221 & w27264 ;
  assign w27266 = ( w26909 & w27219 ) | ( w26909 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27267 = ~w27220 & w27266 ;
  assign w27268 = w27265 | w27267 ;
  assign w27269 = ~\pi097 & w27268 ;
  assign w27270 = ~w26922 & w27186 ;
  assign w27271 = w27187 ^ w27270 ;
  assign w27272 = ~w27221 & w27271 ;
  assign w27273 = ( w26915 & w27219 ) | ( w26915 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27274 = ~w27220 & w27273 ;
  assign w27275 = w27272 | w27274 ;
  assign w27276 = ~\pi096 & w27275 ;
  assign w27277 = ~w26928 & w27183 ;
  assign w27278 = w27184 ^ w27277 ;
  assign w27279 = ~w27221 & w27278 ;
  assign w27280 = ( w26921 & w27219 ) | ( w26921 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27281 = ~w27220 & w27280 ;
  assign w27282 = w27279 | w27281 ;
  assign w27283 = ~\pi095 & w27282 ;
  assign w27284 = ~w26934 & w27180 ;
  assign w27285 = w27181 ^ w27284 ;
  assign w27286 = ~w27221 & w27285 ;
  assign w27287 = ( w26927 & w27219 ) | ( w26927 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27288 = ~w27220 & w27287 ;
  assign w27289 = w27286 | w27288 ;
  assign w27290 = ~\pi094 & w27289 ;
  assign w27291 = ~w26940 & w27177 ;
  assign w27292 = w27178 ^ w27291 ;
  assign w27293 = ~w27221 & w27292 ;
  assign w27294 = ( w26933 & w27219 ) | ( w26933 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27295 = ~w27220 & w27294 ;
  assign w27296 = w27293 | w27295 ;
  assign w27297 = ~\pi093 & w27296 ;
  assign w27298 = ~w26946 & w27174 ;
  assign w27299 = w27175 ^ w27298 ;
  assign w27300 = ~w27221 & w27299 ;
  assign w27301 = ( w26939 & w27219 ) | ( w26939 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27302 = ~w27220 & w27301 ;
  assign w27303 = w27300 | w27302 ;
  assign w27304 = ~\pi092 & w27303 ;
  assign w27305 = ~w26952 & w27171 ;
  assign w27306 = w27172 ^ w27305 ;
  assign w27307 = ~w27221 & w27306 ;
  assign w27308 = ( w26945 & w27219 ) | ( w26945 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27309 = ~w27220 & w27308 ;
  assign w27310 = w27307 | w27309 ;
  assign w27311 = ~\pi091 & w27310 ;
  assign w27312 = ~w26958 & w27168 ;
  assign w27313 = w27169 ^ w27312 ;
  assign w27314 = ~w27221 & w27313 ;
  assign w27315 = ( w26951 & w27219 ) | ( w26951 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27316 = ~w27220 & w27315 ;
  assign w27317 = w27314 | w27316 ;
  assign w27318 = ~\pi090 & w27317 ;
  assign w27319 = ~w26964 & w27165 ;
  assign w27320 = w27166 ^ w27319 ;
  assign w27321 = ~w27221 & w27320 ;
  assign w27322 = ( w26957 & w27219 ) | ( w26957 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27323 = ~w27220 & w27322 ;
  assign w27324 = w27321 | w27323 ;
  assign w27325 = ~\pi089 & w27324 ;
  assign w27326 = ~w26970 & w27162 ;
  assign w27327 = w27163 ^ w27326 ;
  assign w27328 = ~w27221 & w27327 ;
  assign w27329 = ( w26963 & w27219 ) | ( w26963 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27330 = ~w27220 & w27329 ;
  assign w27331 = w27328 | w27330 ;
  assign w27332 = ~\pi088 & w27331 ;
  assign w27333 = ~w26976 & w27159 ;
  assign w27334 = w27160 ^ w27333 ;
  assign w27335 = ~w27221 & w27334 ;
  assign w27336 = ( w26969 & w27219 ) | ( w26969 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27337 = ~w27220 & w27336 ;
  assign w27338 = w27335 | w27337 ;
  assign w27339 = ~\pi087 & w27338 ;
  assign w27340 = ~w26982 & w27156 ;
  assign w27341 = w27157 ^ w27340 ;
  assign w27342 = ~w27221 & w27341 ;
  assign w27343 = ( w26975 & w27219 ) | ( w26975 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27344 = ~w27220 & w27343 ;
  assign w27345 = w27342 | w27344 ;
  assign w27346 = ~\pi086 & w27345 ;
  assign w27347 = ~w26988 & w27153 ;
  assign w27348 = w27154 ^ w27347 ;
  assign w27349 = ~w27221 & w27348 ;
  assign w27350 = ( w26981 & w27219 ) | ( w26981 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27351 = ~w27220 & w27350 ;
  assign w27352 = w27349 | w27351 ;
  assign w27353 = ~\pi085 & w27352 ;
  assign w27354 = ~w26994 & w27150 ;
  assign w27355 = w27151 ^ w27354 ;
  assign w27356 = ~w27221 & w27355 ;
  assign w27357 = ( w26987 & w27219 ) | ( w26987 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27358 = ~w27220 & w27357 ;
  assign w27359 = w27356 | w27358 ;
  assign w27360 = ~\pi084 & w27359 ;
  assign w27361 = ~w27000 & w27147 ;
  assign w27362 = w27148 ^ w27361 ;
  assign w27363 = ~w27221 & w27362 ;
  assign w27364 = ( w26993 & w27219 ) | ( w26993 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27365 = ~w27220 & w27364 ;
  assign w27366 = w27363 | w27365 ;
  assign w27367 = ~\pi083 & w27366 ;
  assign w27368 = ~w27006 & w27144 ;
  assign w27369 = w27145 ^ w27368 ;
  assign w27370 = ~w27221 & w27369 ;
  assign w27371 = ( w26999 & w27219 ) | ( w26999 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27372 = ~w27220 & w27371 ;
  assign w27373 = w27370 | w27372 ;
  assign w27374 = ~\pi082 & w27373 ;
  assign w27375 = ~w27012 & w27141 ;
  assign w27376 = w27142 ^ w27375 ;
  assign w27377 = ~w27221 & w27376 ;
  assign w27378 = ( w27005 & w27219 ) | ( w27005 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27379 = ~w27220 & w27378 ;
  assign w27380 = w27377 | w27379 ;
  assign w27381 = ~\pi081 & w27380 ;
  assign w27382 = ~w27018 & w27138 ;
  assign w27383 = w27139 ^ w27382 ;
  assign w27384 = ~w27221 & w27383 ;
  assign w27385 = ( w27011 & w27219 ) | ( w27011 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27386 = ~w27220 & w27385 ;
  assign w27387 = w27384 | w27386 ;
  assign w27388 = ~\pi080 & w27387 ;
  assign w27389 = ~w27024 & w27135 ;
  assign w27390 = w27136 ^ w27389 ;
  assign w27391 = ~w27221 & w27390 ;
  assign w27392 = ( w27017 & w27219 ) | ( w27017 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27393 = ~w27220 & w27392 ;
  assign w27394 = w27391 | w27393 ;
  assign w27395 = ~\pi079 & w27394 ;
  assign w27396 = ~w27030 & w27132 ;
  assign w27397 = w27133 ^ w27396 ;
  assign w27398 = ~w27221 & w27397 ;
  assign w27399 = ( w27023 & w27219 ) | ( w27023 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27400 = ~w27220 & w27399 ;
  assign w27401 = w27398 | w27400 ;
  assign w27402 = ~\pi078 & w27401 ;
  assign w27403 = ~w27036 & w27129 ;
  assign w27404 = w27130 ^ w27403 ;
  assign w27405 = ~w27221 & w27404 ;
  assign w27406 = ( w27029 & w27219 ) | ( w27029 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27407 = ~w27220 & w27406 ;
  assign w27408 = w27405 | w27407 ;
  assign w27409 = ~\pi077 & w27408 ;
  assign w27410 = ~w27042 & w27126 ;
  assign w27411 = w27127 ^ w27410 ;
  assign w27412 = ~w27221 & w27411 ;
  assign w27413 = ( w27035 & w27219 ) | ( w27035 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27414 = ~w27220 & w27413 ;
  assign w27415 = w27412 | w27414 ;
  assign w27416 = ~\pi076 & w27415 ;
  assign w27417 = ~w27048 & w27123 ;
  assign w27418 = w27124 ^ w27417 ;
  assign w27419 = ~w27221 & w27418 ;
  assign w27420 = ( w27041 & w27219 ) | ( w27041 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27421 = ~w27220 & w27420 ;
  assign w27422 = w27419 | w27421 ;
  assign w27423 = ~\pi075 & w27422 ;
  assign w27424 = ~w27054 & w27120 ;
  assign w27425 = w27121 ^ w27424 ;
  assign w27426 = ~w27221 & w27425 ;
  assign w27427 = ( w27047 & w27219 ) | ( w27047 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27428 = ~w27220 & w27427 ;
  assign w27429 = w27426 | w27428 ;
  assign w27430 = ~\pi074 & w27429 ;
  assign w27431 = ~w27060 & w27117 ;
  assign w27432 = w27118 ^ w27431 ;
  assign w27433 = ~w27221 & w27432 ;
  assign w27434 = ( w27053 & w27219 ) | ( w27053 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27435 = ~w27220 & w27434 ;
  assign w27436 = w27433 | w27435 ;
  assign w27437 = ~\pi073 & w27436 ;
  assign w27438 = ~w27066 & w27114 ;
  assign w27439 = w27115 ^ w27438 ;
  assign w27440 = ~w27221 & w27439 ;
  assign w27441 = ( w27059 & w27219 ) | ( w27059 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27442 = ~w27220 & w27441 ;
  assign w27443 = w27440 | w27442 ;
  assign w27444 = ~\pi072 & w27443 ;
  assign w27445 = ~w27072 & w27111 ;
  assign w27446 = w27112 ^ w27445 ;
  assign w27447 = ~w27221 & w27446 ;
  assign w27448 = ( w27065 & w27219 ) | ( w27065 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27449 = ~w27220 & w27448 ;
  assign w27450 = w27447 | w27449 ;
  assign w27451 = ~\pi071 & w27450 ;
  assign w27452 = ~w27078 & w27108 ;
  assign w27453 = w27109 ^ w27452 ;
  assign w27454 = ~w27221 & w27453 ;
  assign w27455 = ( w27071 & w27219 ) | ( w27071 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27456 = ~w27220 & w27455 ;
  assign w27457 = w27454 | w27456 ;
  assign w27458 = ~\pi070 & w27457 ;
  assign w27459 = ~w27084 & w27105 ;
  assign w27460 = w27106 ^ w27459 ;
  assign w27461 = ~w27221 & w27460 ;
  assign w27462 = ( w27077 & w27219 ) | ( w27077 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27463 = ~w27220 & w27462 ;
  assign w27464 = w27461 | w27463 ;
  assign w27465 = ~\pi069 & w27464 ;
  assign w27466 = ~w27092 & w27102 ;
  assign w27467 = w27103 ^ w27466 ;
  assign w27468 = ~w27221 & w27467 ;
  assign w27469 = ( w27083 & w27219 ) | ( w27083 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27470 = ~w27220 & w27469 ;
  assign w27471 = w27468 | w27470 ;
  assign w27472 = ~\pi068 & w27471 ;
  assign w27473 = ( \pi065 & w27096 ) | ( \pi065 & ~w27221 ) | ( w27096 & ~w27221 ) ;
  assign w27474 = ( \pi065 & w27098 ) | ( \pi065 & ~w27473 ) | ( w27098 & ~w27473 ) ;
  assign w27475 = w27099 ^ w27474 ;
  assign w27476 = ~w27221 & w27475 ;
  assign w27477 = ( w27091 & w27219 ) | ( w27091 & w27220 ) | ( w27219 & w27220 ) ;
  assign w27478 = ~w27220 & w27477 ;
  assign w27479 = w27476 | w27478 ;
  assign w27480 = ~\pi067 & w27479 ;
  assign w27481 = w7654 ^ w27096 ;
  assign w27482 = \pi065 ^ w27481 ;
  assign w27483 = w27221 ^ w27482 ;
  assign w27484 = ( w27096 & w27482 ) | ( w27096 & w27483 ) | ( w27482 & w27483 ) ;
  assign w27485 = ~\pi066 & w27484 ;
  assign w27486 = w27096 ^ w27221 ;
  assign w27487 = ( w27096 & w27482 ) | ( w27096 & ~w27486 ) | ( w27482 & ~w27486 ) ;
  assign w27488 = \pi066 ^ w27487 ;
  assign w27489 = ( \pi064 & ~w27221 ) | ( \pi064 & w27488 ) | ( ~w27221 & w27488 ) ;
  assign w27490 = \pi025 ^ w27489 ;
  assign w27491 = ( \pi065 & w8393 ) | ( \pi065 & ~w27490 ) | ( w8393 & ~w27490 ) ;
  assign w27492 = w27488 | w27491 ;
  assign w27493 = \pi067 ^ w27479 ;
  assign w27494 = ( ~w27485 & w27492 ) | ( ~w27485 & w27493 ) | ( w27492 & w27493 ) ;
  assign w27495 = w27493 | w27494 ;
  assign w27496 = \pi068 ^ w27471 ;
  assign w27497 = ( ~w27480 & w27495 ) | ( ~w27480 & w27496 ) | ( w27495 & w27496 ) ;
  assign w27498 = w27496 | w27497 ;
  assign w27499 = \pi069 ^ w27464 ;
  assign w27500 = ( ~w27472 & w27498 ) | ( ~w27472 & w27499 ) | ( w27498 & w27499 ) ;
  assign w27501 = w27499 | w27500 ;
  assign w27502 = \pi070 ^ w27457 ;
  assign w27503 = ( ~w27465 & w27501 ) | ( ~w27465 & w27502 ) | ( w27501 & w27502 ) ;
  assign w27504 = w27502 | w27503 ;
  assign w27505 = \pi071 ^ w27450 ;
  assign w27506 = ( ~w27458 & w27504 ) | ( ~w27458 & w27505 ) | ( w27504 & w27505 ) ;
  assign w27507 = w27505 | w27506 ;
  assign w27508 = \pi072 ^ w27443 ;
  assign w27509 = ( ~w27451 & w27507 ) | ( ~w27451 & w27508 ) | ( w27507 & w27508 ) ;
  assign w27510 = w27508 | w27509 ;
  assign w27511 = \pi073 ^ w27436 ;
  assign w27512 = ( ~w27444 & w27510 ) | ( ~w27444 & w27511 ) | ( w27510 & w27511 ) ;
  assign w27513 = w27511 | w27512 ;
  assign w27514 = \pi074 ^ w27429 ;
  assign w27515 = ( ~w27437 & w27513 ) | ( ~w27437 & w27514 ) | ( w27513 & w27514 ) ;
  assign w27516 = w27514 | w27515 ;
  assign w27517 = \pi075 ^ w27422 ;
  assign w27518 = ( ~w27430 & w27516 ) | ( ~w27430 & w27517 ) | ( w27516 & w27517 ) ;
  assign w27519 = w27517 | w27518 ;
  assign w27520 = \pi076 ^ w27415 ;
  assign w27521 = ( ~w27423 & w27519 ) | ( ~w27423 & w27520 ) | ( w27519 & w27520 ) ;
  assign w27522 = w27520 | w27521 ;
  assign w27523 = \pi077 ^ w27408 ;
  assign w27524 = ( ~w27416 & w27522 ) | ( ~w27416 & w27523 ) | ( w27522 & w27523 ) ;
  assign w27525 = w27523 | w27524 ;
  assign w27526 = \pi078 ^ w27401 ;
  assign w27527 = ( ~w27409 & w27525 ) | ( ~w27409 & w27526 ) | ( w27525 & w27526 ) ;
  assign w27528 = w27526 | w27527 ;
  assign w27529 = \pi079 ^ w27394 ;
  assign w27530 = ( ~w27402 & w27528 ) | ( ~w27402 & w27529 ) | ( w27528 & w27529 ) ;
  assign w27531 = w27529 | w27530 ;
  assign w27532 = \pi080 ^ w27387 ;
  assign w27533 = ( ~w27395 & w27531 ) | ( ~w27395 & w27532 ) | ( w27531 & w27532 ) ;
  assign w27534 = w27532 | w27533 ;
  assign w27535 = \pi081 ^ w27380 ;
  assign w27536 = ( ~w27388 & w27534 ) | ( ~w27388 & w27535 ) | ( w27534 & w27535 ) ;
  assign w27537 = w27535 | w27536 ;
  assign w27538 = \pi082 ^ w27373 ;
  assign w27539 = ( ~w27381 & w27537 ) | ( ~w27381 & w27538 ) | ( w27537 & w27538 ) ;
  assign w27540 = w27538 | w27539 ;
  assign w27541 = \pi083 ^ w27366 ;
  assign w27542 = ( ~w27374 & w27540 ) | ( ~w27374 & w27541 ) | ( w27540 & w27541 ) ;
  assign w27543 = w27541 | w27542 ;
  assign w27544 = \pi084 ^ w27359 ;
  assign w27545 = ( ~w27367 & w27543 ) | ( ~w27367 & w27544 ) | ( w27543 & w27544 ) ;
  assign w27546 = w27544 | w27545 ;
  assign w27547 = \pi085 ^ w27352 ;
  assign w27548 = ( ~w27360 & w27546 ) | ( ~w27360 & w27547 ) | ( w27546 & w27547 ) ;
  assign w27549 = w27547 | w27548 ;
  assign w27550 = \pi086 ^ w27345 ;
  assign w27551 = ( ~w27353 & w27549 ) | ( ~w27353 & w27550 ) | ( w27549 & w27550 ) ;
  assign w27552 = w27550 | w27551 ;
  assign w27553 = \pi087 ^ w27338 ;
  assign w27554 = ( ~w27346 & w27552 ) | ( ~w27346 & w27553 ) | ( w27552 & w27553 ) ;
  assign w27555 = w27553 | w27554 ;
  assign w27556 = \pi088 ^ w27331 ;
  assign w27557 = ( ~w27339 & w27555 ) | ( ~w27339 & w27556 ) | ( w27555 & w27556 ) ;
  assign w27558 = w27556 | w27557 ;
  assign w27559 = \pi089 ^ w27324 ;
  assign w27560 = ( ~w27332 & w27558 ) | ( ~w27332 & w27559 ) | ( w27558 & w27559 ) ;
  assign w27561 = w27559 | w27560 ;
  assign w27562 = \pi090 ^ w27317 ;
  assign w27563 = ( ~w27325 & w27561 ) | ( ~w27325 & w27562 ) | ( w27561 & w27562 ) ;
  assign w27564 = w27562 | w27563 ;
  assign w27565 = \pi091 ^ w27310 ;
  assign w27566 = ( ~w27318 & w27564 ) | ( ~w27318 & w27565 ) | ( w27564 & w27565 ) ;
  assign w27567 = w27565 | w27566 ;
  assign w27568 = \pi092 ^ w27303 ;
  assign w27569 = ( ~w27311 & w27567 ) | ( ~w27311 & w27568 ) | ( w27567 & w27568 ) ;
  assign w27570 = w27568 | w27569 ;
  assign w27571 = \pi093 ^ w27296 ;
  assign w27572 = ( ~w27304 & w27570 ) | ( ~w27304 & w27571 ) | ( w27570 & w27571 ) ;
  assign w27573 = w27571 | w27572 ;
  assign w27574 = \pi094 ^ w27289 ;
  assign w27575 = ( ~w27297 & w27573 ) | ( ~w27297 & w27574 ) | ( w27573 & w27574 ) ;
  assign w27576 = w27574 | w27575 ;
  assign w27577 = \pi095 ^ w27282 ;
  assign w27578 = ( ~w27290 & w27576 ) | ( ~w27290 & w27577 ) | ( w27576 & w27577 ) ;
  assign w27579 = w27577 | w27578 ;
  assign w27580 = \pi096 ^ w27275 ;
  assign w27581 = ( ~w27283 & w27579 ) | ( ~w27283 & w27580 ) | ( w27579 & w27580 ) ;
  assign w27582 = w27580 | w27581 ;
  assign w27583 = \pi097 ^ w27268 ;
  assign w27584 = ( ~w27276 & w27582 ) | ( ~w27276 & w27583 ) | ( w27582 & w27583 ) ;
  assign w27585 = w27583 | w27584 ;
  assign w27586 = \pi098 ^ w27261 ;
  assign w27587 = ( ~w27269 & w27585 ) | ( ~w27269 & w27586 ) | ( w27585 & w27586 ) ;
  assign w27588 = w27586 | w27587 ;
  assign w27589 = \pi099 ^ w27254 ;
  assign w27590 = ( ~w27262 & w27588 ) | ( ~w27262 & w27589 ) | ( w27588 & w27589 ) ;
  assign w27591 = w27589 | w27590 ;
  assign w27592 = \pi100 ^ w27247 ;
  assign w27593 = ( ~w27255 & w27591 ) | ( ~w27255 & w27592 ) | ( w27591 & w27592 ) ;
  assign w27594 = w27592 | w27593 ;
  assign w27595 = \pi101 ^ w27240 ;
  assign w27596 = ( ~w27248 & w27594 ) | ( ~w27248 & w27595 ) | ( w27594 & w27595 ) ;
  assign w27597 = w27595 | w27596 ;
  assign w27598 = \pi102 ^ w27227 ;
  assign w27599 = ( ~w27241 & w27597 ) | ( ~w27241 & w27598 ) | ( w27597 & w27598 ) ;
  assign w27600 = w27598 | w27599 ;
  assign w27601 = \pi103 ^ w27233 ;
  assign w27602 = w27234 & ~w27601 ;
  assign w27603 = ( w27600 & w27601 ) | ( w27600 & ~w27602 ) | ( w27601 & ~w27602 ) ;
  assign w27604 = ~\pi103 & w27233 ;
  assign w27605 = w27603 & ~w27604 ;
  assign w27606 = w8169 | w27605 ;
  assign w27607 = w27227 & w27606 ;
  assign w27608 = ~w27241 & w27597 ;
  assign w27609 = w27598 ^ w27608 ;
  assign w27610 = ~w27606 & w27609 ;
  assign w27611 = w27607 | w27610 ;
  assign w27612 = w27233 & w27606 ;
  assign w27613 = ~w27234 & w27600 ;
  assign w27614 = w27601 ^ w27613 ;
  assign w27615 = ~w27606 & w27614 ;
  assign w27616 = w27612 | w27615 ;
  assign w27617 = ~\pi103 & w27611 ;
  assign w27618 = w27240 & w27606 ;
  assign w27619 = ~w27248 & w27594 ;
  assign w27620 = w27595 ^ w27619 ;
  assign w27621 = ~w27606 & w27620 ;
  assign w27622 = w27618 | w27621 ;
  assign w27623 = ~\pi102 & w27622 ;
  assign w27624 = w27247 & w27606 ;
  assign w27625 = ~w27255 & w27591 ;
  assign w27626 = w27592 ^ w27625 ;
  assign w27627 = ~w27606 & w27626 ;
  assign w27628 = w27624 | w27627 ;
  assign w27629 = ~\pi101 & w27628 ;
  assign w27630 = w27254 & w27606 ;
  assign w27631 = ~w27262 & w27588 ;
  assign w27632 = w27589 ^ w27631 ;
  assign w27633 = ~w27606 & w27632 ;
  assign w27634 = w27630 | w27633 ;
  assign w27635 = ~\pi100 & w27634 ;
  assign w27636 = w27261 & w27606 ;
  assign w27637 = ~w27269 & w27585 ;
  assign w27638 = w27586 ^ w27637 ;
  assign w27639 = ~w27606 & w27638 ;
  assign w27640 = w27636 | w27639 ;
  assign w27641 = ~\pi099 & w27640 ;
  assign w27642 = w27268 & w27606 ;
  assign w27643 = ~w27276 & w27582 ;
  assign w27644 = w27583 ^ w27643 ;
  assign w27645 = ~w27606 & w27644 ;
  assign w27646 = w27642 | w27645 ;
  assign w27647 = ~\pi098 & w27646 ;
  assign w27648 = w27275 & w27606 ;
  assign w27649 = ~w27283 & w27579 ;
  assign w27650 = w27580 ^ w27649 ;
  assign w27651 = ~w27606 & w27650 ;
  assign w27652 = w27648 | w27651 ;
  assign w27653 = ~\pi097 & w27652 ;
  assign w27654 = w27282 & w27606 ;
  assign w27655 = ~w27290 & w27576 ;
  assign w27656 = w27577 ^ w27655 ;
  assign w27657 = ~w27606 & w27656 ;
  assign w27658 = w27654 | w27657 ;
  assign w27659 = ~\pi096 & w27658 ;
  assign w27660 = w27289 & w27606 ;
  assign w27661 = ~w27297 & w27573 ;
  assign w27662 = w27574 ^ w27661 ;
  assign w27663 = ~w27606 & w27662 ;
  assign w27664 = w27660 | w27663 ;
  assign w27665 = ~\pi095 & w27664 ;
  assign w27666 = w27296 & w27606 ;
  assign w27667 = ~w27304 & w27570 ;
  assign w27668 = w27571 ^ w27667 ;
  assign w27669 = ~w27606 & w27668 ;
  assign w27670 = w27666 | w27669 ;
  assign w27671 = ~\pi094 & w27670 ;
  assign w27672 = w27303 & w27606 ;
  assign w27673 = ~w27311 & w27567 ;
  assign w27674 = w27568 ^ w27673 ;
  assign w27675 = ~w27606 & w27674 ;
  assign w27676 = w27672 | w27675 ;
  assign w27677 = ~\pi093 & w27676 ;
  assign w27678 = w27310 & w27606 ;
  assign w27679 = ~w27318 & w27564 ;
  assign w27680 = w27565 ^ w27679 ;
  assign w27681 = ~w27606 & w27680 ;
  assign w27682 = w27678 | w27681 ;
  assign w27683 = ~\pi092 & w27682 ;
  assign w27684 = w27317 & w27606 ;
  assign w27685 = ~w27325 & w27561 ;
  assign w27686 = w27562 ^ w27685 ;
  assign w27687 = ~w27606 & w27686 ;
  assign w27688 = w27684 | w27687 ;
  assign w27689 = ~\pi091 & w27688 ;
  assign w27690 = w27324 & w27606 ;
  assign w27691 = ~w27332 & w27558 ;
  assign w27692 = w27559 ^ w27691 ;
  assign w27693 = ~w27606 & w27692 ;
  assign w27694 = w27690 | w27693 ;
  assign w27695 = ~\pi090 & w27694 ;
  assign w27696 = w27331 & w27606 ;
  assign w27697 = ~w27339 & w27555 ;
  assign w27698 = w27556 ^ w27697 ;
  assign w27699 = ~w27606 & w27698 ;
  assign w27700 = w27696 | w27699 ;
  assign w27701 = ~\pi089 & w27700 ;
  assign w27702 = w27338 & w27606 ;
  assign w27703 = ~w27346 & w27552 ;
  assign w27704 = w27553 ^ w27703 ;
  assign w27705 = ~w27606 & w27704 ;
  assign w27706 = w27702 | w27705 ;
  assign w27707 = ~\pi088 & w27706 ;
  assign w27708 = w27345 & w27606 ;
  assign w27709 = ~w27353 & w27549 ;
  assign w27710 = w27550 ^ w27709 ;
  assign w27711 = ~w27606 & w27710 ;
  assign w27712 = w27708 | w27711 ;
  assign w27713 = ~\pi087 & w27712 ;
  assign w27714 = w27352 & w27606 ;
  assign w27715 = ~w27360 & w27546 ;
  assign w27716 = w27547 ^ w27715 ;
  assign w27717 = ~w27606 & w27716 ;
  assign w27718 = w27714 | w27717 ;
  assign w27719 = ~\pi086 & w27718 ;
  assign w27720 = w27359 & w27606 ;
  assign w27721 = ~w27367 & w27543 ;
  assign w27722 = w27544 ^ w27721 ;
  assign w27723 = ~w27606 & w27722 ;
  assign w27724 = w27720 | w27723 ;
  assign w27725 = ~\pi085 & w27724 ;
  assign w27726 = w27366 & w27606 ;
  assign w27727 = ~w27374 & w27540 ;
  assign w27728 = w27541 ^ w27727 ;
  assign w27729 = ~w27606 & w27728 ;
  assign w27730 = w27726 | w27729 ;
  assign w27731 = ~\pi084 & w27730 ;
  assign w27732 = w27373 & w27606 ;
  assign w27733 = ~w27381 & w27537 ;
  assign w27734 = w27538 ^ w27733 ;
  assign w27735 = ~w27606 & w27734 ;
  assign w27736 = w27732 | w27735 ;
  assign w27737 = ~\pi083 & w27736 ;
  assign w27738 = w27380 & w27606 ;
  assign w27739 = ~w27388 & w27534 ;
  assign w27740 = w27535 ^ w27739 ;
  assign w27741 = ~w27606 & w27740 ;
  assign w27742 = w27738 | w27741 ;
  assign w27743 = ~\pi082 & w27742 ;
  assign w27744 = w27387 & w27606 ;
  assign w27745 = ~w27395 & w27531 ;
  assign w27746 = w27532 ^ w27745 ;
  assign w27747 = ~w27606 & w27746 ;
  assign w27748 = w27744 | w27747 ;
  assign w27749 = ~\pi081 & w27748 ;
  assign w27750 = w27394 & w27606 ;
  assign w27751 = ~w27402 & w27528 ;
  assign w27752 = w27529 ^ w27751 ;
  assign w27753 = ~w27606 & w27752 ;
  assign w27754 = w27750 | w27753 ;
  assign w27755 = ~\pi080 & w27754 ;
  assign w27756 = w27401 & w27606 ;
  assign w27757 = ~w27409 & w27525 ;
  assign w27758 = w27526 ^ w27757 ;
  assign w27759 = ~w27606 & w27758 ;
  assign w27760 = w27756 | w27759 ;
  assign w27761 = ~\pi079 & w27760 ;
  assign w27762 = w27408 & w27606 ;
  assign w27763 = ~w27416 & w27522 ;
  assign w27764 = w27523 ^ w27763 ;
  assign w27765 = ~w27606 & w27764 ;
  assign w27766 = w27762 | w27765 ;
  assign w27767 = ~\pi078 & w27766 ;
  assign w27768 = w27415 & w27606 ;
  assign w27769 = ~w27423 & w27519 ;
  assign w27770 = w27520 ^ w27769 ;
  assign w27771 = ~w27606 & w27770 ;
  assign w27772 = w27768 | w27771 ;
  assign w27773 = ~\pi077 & w27772 ;
  assign w27774 = w27422 & w27606 ;
  assign w27775 = ~w27430 & w27516 ;
  assign w27776 = w27517 ^ w27775 ;
  assign w27777 = ~w27606 & w27776 ;
  assign w27778 = w27774 | w27777 ;
  assign w27779 = ~\pi076 & w27778 ;
  assign w27780 = w27429 & w27606 ;
  assign w27781 = ~w27437 & w27513 ;
  assign w27782 = w27514 ^ w27781 ;
  assign w27783 = ~w27606 & w27782 ;
  assign w27784 = w27780 | w27783 ;
  assign w27785 = ~\pi075 & w27784 ;
  assign w27786 = w27436 & w27606 ;
  assign w27787 = ~w27444 & w27510 ;
  assign w27788 = w27511 ^ w27787 ;
  assign w27789 = ~w27606 & w27788 ;
  assign w27790 = w27786 | w27789 ;
  assign w27791 = ~\pi074 & w27790 ;
  assign w27792 = w27443 & w27606 ;
  assign w27793 = ~w27451 & w27507 ;
  assign w27794 = w27508 ^ w27793 ;
  assign w27795 = ~w27606 & w27794 ;
  assign w27796 = w27792 | w27795 ;
  assign w27797 = ~\pi073 & w27796 ;
  assign w27798 = w27450 & w27606 ;
  assign w27799 = ~w27458 & w27504 ;
  assign w27800 = w27505 ^ w27799 ;
  assign w27801 = ~w27606 & w27800 ;
  assign w27802 = w27798 | w27801 ;
  assign w27803 = ~\pi072 & w27802 ;
  assign w27804 = w27457 & w27606 ;
  assign w27805 = ~w27465 & w27501 ;
  assign w27806 = w27502 ^ w27805 ;
  assign w27807 = ~w27606 & w27806 ;
  assign w27808 = w27804 | w27807 ;
  assign w27809 = ~\pi071 & w27808 ;
  assign w27810 = w27464 & w27606 ;
  assign w27811 = ~w27472 & w27498 ;
  assign w27812 = w27499 ^ w27811 ;
  assign w27813 = ~w27606 & w27812 ;
  assign w27814 = w27810 | w27813 ;
  assign w27815 = ~\pi070 & w27814 ;
  assign w27816 = w27471 & w27606 ;
  assign w27817 = ~w27480 & w27495 ;
  assign w27818 = w27496 ^ w27817 ;
  assign w27819 = ~w27606 & w27818 ;
  assign w27820 = w27816 | w27819 ;
  assign w27821 = ~\pi069 & w27820 ;
  assign w27822 = w27479 & w27606 ;
  assign w27823 = ~w27485 & w27492 ;
  assign w27824 = w27493 ^ w27823 ;
  assign w27825 = ~w27606 & w27824 ;
  assign w27826 = w27822 | w27825 ;
  assign w27827 = ~\pi068 & w27826 ;
  assign w27828 = w27484 & w27606 ;
  assign w27829 = \pi064 & ~w27221 ;
  assign w27830 = \pi025 ^ w27829 ;
  assign w27831 = ( \pi065 & w8393 ) | ( \pi065 & ~w27830 ) | ( w8393 & ~w27830 ) ;
  assign w27832 = w27488 ^ w27831 ;
  assign w27833 = ( w8169 & w27605 ) | ( w8169 & w27832 ) | ( w27605 & w27832 ) ;
  assign w27834 = w27832 & ~w27833 ;
  assign w27835 = w27828 | w27834 ;
  assign w27836 = ~\pi067 & w27835 ;
  assign w27837 = \pi024 ^ w27221 ;
  assign w27838 = ( \pi064 & w8169 ) | ( \pi064 & w27837 ) | ( w8169 & w27837 ) ;
  assign w27839 = w8400 ^ w27838 ;
  assign w27840 = ~w8169 & w27839 ;
  assign w27841 = ~w27605 & w27840 ;
  assign w27842 = ( ~\pi064 & w27221 ) | ( ~\pi064 & w27606 ) | ( w27221 & w27606 ) ;
  assign w27843 = \pi025 ^ w27842 ;
  assign w27844 = w27606 & ~w27843 ;
  assign w27845 = w27841 | w27844 ;
  assign w27846 = ~\pi066 & w27845 ;
  assign w27847 = ( \pi024 & ~w8413 ) | ( \pi024 & w27605 ) | ( ~w8413 & w27605 ) ;
  assign w27848 = \pi024 & w27847 ;
  assign w27849 = w155 | w27605 ;
  assign w27850 = w8418 & ~w27849 ;
  assign w27851 = ~w8416 & w27850 ;
  assign w27852 = w27606 | w27841 ;
  assign w27853 = ( w27830 & w27841 ) | ( w27830 & w27852 ) | ( w27841 & w27852 ) ;
  assign w27854 = \pi066 ^ w27853 ;
  assign w27855 = w27848 | w27851 ;
  assign w27856 = ( \pi065 & w8422 ) | ( \pi065 & ~w27855 ) | ( w8422 & ~w27855 ) ;
  assign w27857 = w27854 | w27856 ;
  assign w27858 = \pi067 ^ w27835 ;
  assign w27859 = ( ~w27846 & w27857 ) | ( ~w27846 & w27858 ) | ( w27857 & w27858 ) ;
  assign w27860 = w27858 | w27859 ;
  assign w27861 = \pi068 ^ w27826 ;
  assign w27862 = ( ~w27836 & w27860 ) | ( ~w27836 & w27861 ) | ( w27860 & w27861 ) ;
  assign w27863 = w27861 | w27862 ;
  assign w27864 = \pi069 ^ w27820 ;
  assign w27865 = ( ~w27827 & w27863 ) | ( ~w27827 & w27864 ) | ( w27863 & w27864 ) ;
  assign w27866 = w27864 | w27865 ;
  assign w27867 = \pi070 ^ w27814 ;
  assign w27868 = ( ~w27821 & w27866 ) | ( ~w27821 & w27867 ) | ( w27866 & w27867 ) ;
  assign w27869 = w27867 | w27868 ;
  assign w27870 = \pi071 ^ w27808 ;
  assign w27871 = ( ~w27815 & w27869 ) | ( ~w27815 & w27870 ) | ( w27869 & w27870 ) ;
  assign w27872 = w27870 | w27871 ;
  assign w27873 = \pi072 ^ w27802 ;
  assign w27874 = ( ~w27809 & w27872 ) | ( ~w27809 & w27873 ) | ( w27872 & w27873 ) ;
  assign w27875 = w27873 | w27874 ;
  assign w27876 = \pi073 ^ w27796 ;
  assign w27877 = ( ~w27803 & w27875 ) | ( ~w27803 & w27876 ) | ( w27875 & w27876 ) ;
  assign w27878 = w27876 | w27877 ;
  assign w27879 = \pi074 ^ w27790 ;
  assign w27880 = ( ~w27797 & w27878 ) | ( ~w27797 & w27879 ) | ( w27878 & w27879 ) ;
  assign w27881 = w27879 | w27880 ;
  assign w27882 = \pi075 ^ w27784 ;
  assign w27883 = ( ~w27791 & w27881 ) | ( ~w27791 & w27882 ) | ( w27881 & w27882 ) ;
  assign w27884 = w27882 | w27883 ;
  assign w27885 = \pi076 ^ w27778 ;
  assign w27886 = ( ~w27785 & w27884 ) | ( ~w27785 & w27885 ) | ( w27884 & w27885 ) ;
  assign w27887 = w27885 | w27886 ;
  assign w27888 = \pi077 ^ w27772 ;
  assign w27889 = ( ~w27779 & w27887 ) | ( ~w27779 & w27888 ) | ( w27887 & w27888 ) ;
  assign w27890 = w27888 | w27889 ;
  assign w27891 = \pi078 ^ w27766 ;
  assign w27892 = ( ~w27773 & w27890 ) | ( ~w27773 & w27891 ) | ( w27890 & w27891 ) ;
  assign w27893 = w27891 | w27892 ;
  assign w27894 = \pi079 ^ w27760 ;
  assign w27895 = ( ~w27767 & w27893 ) | ( ~w27767 & w27894 ) | ( w27893 & w27894 ) ;
  assign w27896 = w27894 | w27895 ;
  assign w27897 = \pi080 ^ w27754 ;
  assign w27898 = ( ~w27761 & w27896 ) | ( ~w27761 & w27897 ) | ( w27896 & w27897 ) ;
  assign w27899 = w27897 | w27898 ;
  assign w27900 = \pi081 ^ w27748 ;
  assign w27901 = ( ~w27755 & w27899 ) | ( ~w27755 & w27900 ) | ( w27899 & w27900 ) ;
  assign w27902 = w27900 | w27901 ;
  assign w27903 = \pi082 ^ w27742 ;
  assign w27904 = ( ~w27749 & w27902 ) | ( ~w27749 & w27903 ) | ( w27902 & w27903 ) ;
  assign w27905 = w27903 | w27904 ;
  assign w27906 = \pi083 ^ w27736 ;
  assign w27907 = ( ~w27743 & w27905 ) | ( ~w27743 & w27906 ) | ( w27905 & w27906 ) ;
  assign w27908 = w27906 | w27907 ;
  assign w27909 = \pi084 ^ w27730 ;
  assign w27910 = ( ~w27737 & w27908 ) | ( ~w27737 & w27909 ) | ( w27908 & w27909 ) ;
  assign w27911 = w27909 | w27910 ;
  assign w27912 = \pi085 ^ w27724 ;
  assign w27913 = ( ~w27731 & w27911 ) | ( ~w27731 & w27912 ) | ( w27911 & w27912 ) ;
  assign w27914 = w27912 | w27913 ;
  assign w27915 = \pi086 ^ w27718 ;
  assign w27916 = ( ~w27725 & w27914 ) | ( ~w27725 & w27915 ) | ( w27914 & w27915 ) ;
  assign w27917 = w27915 | w27916 ;
  assign w27918 = \pi087 ^ w27712 ;
  assign w27919 = ( ~w27719 & w27917 ) | ( ~w27719 & w27918 ) | ( w27917 & w27918 ) ;
  assign w27920 = w27918 | w27919 ;
  assign w27921 = \pi088 ^ w27706 ;
  assign w27922 = ( ~w27713 & w27920 ) | ( ~w27713 & w27921 ) | ( w27920 & w27921 ) ;
  assign w27923 = w27921 | w27922 ;
  assign w27924 = \pi089 ^ w27700 ;
  assign w27925 = ( ~w27707 & w27923 ) | ( ~w27707 & w27924 ) | ( w27923 & w27924 ) ;
  assign w27926 = w27924 | w27925 ;
  assign w27927 = \pi090 ^ w27694 ;
  assign w27928 = ( ~w27701 & w27926 ) | ( ~w27701 & w27927 ) | ( w27926 & w27927 ) ;
  assign w27929 = w27927 | w27928 ;
  assign w27930 = \pi091 ^ w27688 ;
  assign w27931 = ( ~w27695 & w27929 ) | ( ~w27695 & w27930 ) | ( w27929 & w27930 ) ;
  assign w27932 = w27930 | w27931 ;
  assign w27933 = \pi092 ^ w27682 ;
  assign w27934 = ( ~w27689 & w27932 ) | ( ~w27689 & w27933 ) | ( w27932 & w27933 ) ;
  assign w27935 = w27933 | w27934 ;
  assign w27936 = \pi093 ^ w27676 ;
  assign w27937 = ( ~w27683 & w27935 ) | ( ~w27683 & w27936 ) | ( w27935 & w27936 ) ;
  assign w27938 = w27936 | w27937 ;
  assign w27939 = \pi094 ^ w27670 ;
  assign w27940 = ( ~w27677 & w27938 ) | ( ~w27677 & w27939 ) | ( w27938 & w27939 ) ;
  assign w27941 = w27939 | w27940 ;
  assign w27942 = \pi095 ^ w27664 ;
  assign w27943 = ( ~w27671 & w27941 ) | ( ~w27671 & w27942 ) | ( w27941 & w27942 ) ;
  assign w27944 = w27942 | w27943 ;
  assign w27945 = \pi096 ^ w27658 ;
  assign w27946 = ( ~w27665 & w27944 ) | ( ~w27665 & w27945 ) | ( w27944 & w27945 ) ;
  assign w27947 = w27945 | w27946 ;
  assign w27948 = \pi097 ^ w27652 ;
  assign w27949 = ( ~w27659 & w27947 ) | ( ~w27659 & w27948 ) | ( w27947 & w27948 ) ;
  assign w27950 = w27948 | w27949 ;
  assign w27951 = \pi098 ^ w27646 ;
  assign w27952 = ( ~w27653 & w27950 ) | ( ~w27653 & w27951 ) | ( w27950 & w27951 ) ;
  assign w27953 = w27951 | w27952 ;
  assign w27954 = \pi099 ^ w27640 ;
  assign w27955 = ( ~w27647 & w27953 ) | ( ~w27647 & w27954 ) | ( w27953 & w27954 ) ;
  assign w27956 = w27954 | w27955 ;
  assign w27957 = \pi100 ^ w27634 ;
  assign w27958 = ( ~w27641 & w27956 ) | ( ~w27641 & w27957 ) | ( w27956 & w27957 ) ;
  assign w27959 = w27957 | w27958 ;
  assign w27960 = \pi101 ^ w27628 ;
  assign w27961 = ( ~w27635 & w27959 ) | ( ~w27635 & w27960 ) | ( w27959 & w27960 ) ;
  assign w27962 = w27960 | w27961 ;
  assign w27963 = \pi102 ^ w27622 ;
  assign w27964 = ( ~w27629 & w27962 ) | ( ~w27629 & w27963 ) | ( w27962 & w27963 ) ;
  assign w27965 = w27963 | w27964 ;
  assign w27966 = \pi103 ^ w27611 ;
  assign w27967 = ( ~w27623 & w27965 ) | ( ~w27623 & w27966 ) | ( w27965 & w27966 ) ;
  assign w27968 = w27966 | w27967 ;
  assign w27969 = \pi104 ^ w27616 ;
  assign w27970 = w27617 & ~w27969 ;
  assign w27971 = ( w27968 & w27969 ) | ( w27968 & ~w27970 ) | ( w27969 & ~w27970 ) ;
  assign w27972 = ~\pi104 & w27616 ;
  assign w27973 = w27971 & ~w27972 ;
  assign w27974 = w6588 | w27973 ;
  assign w27975 = w27611 & w27974 ;
  assign w27976 = ~w27623 & w27965 ;
  assign w27977 = w27966 ^ w27976 ;
  assign w27978 = ~w27974 & w27977 ;
  assign w27979 = w27975 | w27978 ;
  assign w27980 = ~\pi104 & w27979 ;
  assign w27981 = w27622 & w27974 ;
  assign w27982 = ~w27629 & w27962 ;
  assign w27983 = w27963 ^ w27982 ;
  assign w27984 = ~w27974 & w27983 ;
  assign w27985 = w27981 | w27984 ;
  assign w27986 = ~\pi103 & w27985 ;
  assign w27987 = w27628 & w27974 ;
  assign w27988 = ~w27635 & w27959 ;
  assign w27989 = w27960 ^ w27988 ;
  assign w27990 = ~w27974 & w27989 ;
  assign w27991 = w27987 | w27990 ;
  assign w27992 = ~\pi102 & w27991 ;
  assign w27993 = w27634 & w27974 ;
  assign w27994 = ~w27641 & w27956 ;
  assign w27995 = w27957 ^ w27994 ;
  assign w27996 = ~w27974 & w27995 ;
  assign w27997 = w27993 | w27996 ;
  assign w27998 = ~\pi101 & w27997 ;
  assign w27999 = w27640 & w27974 ;
  assign w28000 = ~w27647 & w27953 ;
  assign w28001 = w27954 ^ w28000 ;
  assign w28002 = ~w27974 & w28001 ;
  assign w28003 = w27999 | w28002 ;
  assign w28004 = ~\pi100 & w28003 ;
  assign w28005 = w27646 & w27974 ;
  assign w28006 = ~w27653 & w27950 ;
  assign w28007 = w27951 ^ w28006 ;
  assign w28008 = ~w27974 & w28007 ;
  assign w28009 = w28005 | w28008 ;
  assign w28010 = ~\pi099 & w28009 ;
  assign w28011 = w27652 & w27974 ;
  assign w28012 = ~w27659 & w27947 ;
  assign w28013 = w27948 ^ w28012 ;
  assign w28014 = ~w27974 & w28013 ;
  assign w28015 = w28011 | w28014 ;
  assign w28016 = ~\pi098 & w28015 ;
  assign w28017 = w27658 & w27974 ;
  assign w28018 = ~w27665 & w27944 ;
  assign w28019 = w27945 ^ w28018 ;
  assign w28020 = ~w27974 & w28019 ;
  assign w28021 = w28017 | w28020 ;
  assign w28022 = ~\pi097 & w28021 ;
  assign w28023 = w27664 & w27974 ;
  assign w28024 = ~w27671 & w27941 ;
  assign w28025 = w27942 ^ w28024 ;
  assign w28026 = ~w27974 & w28025 ;
  assign w28027 = w28023 | w28026 ;
  assign w28028 = ~\pi096 & w28027 ;
  assign w28029 = w27670 & w27974 ;
  assign w28030 = ~w27677 & w27938 ;
  assign w28031 = w27939 ^ w28030 ;
  assign w28032 = ~w27974 & w28031 ;
  assign w28033 = w28029 | w28032 ;
  assign w28034 = ~\pi095 & w28033 ;
  assign w28035 = w27676 & w27974 ;
  assign w28036 = ~w27683 & w27935 ;
  assign w28037 = w27936 ^ w28036 ;
  assign w28038 = ~w27974 & w28037 ;
  assign w28039 = w28035 | w28038 ;
  assign w28040 = ~\pi094 & w28039 ;
  assign w28041 = w27682 & w27974 ;
  assign w28042 = ~w27689 & w27932 ;
  assign w28043 = w27933 ^ w28042 ;
  assign w28044 = ~w27974 & w28043 ;
  assign w28045 = w28041 | w28044 ;
  assign w28046 = ~\pi093 & w28045 ;
  assign w28047 = w27688 & w27974 ;
  assign w28048 = ~w27695 & w27929 ;
  assign w28049 = w27930 ^ w28048 ;
  assign w28050 = ~w27974 & w28049 ;
  assign w28051 = w28047 | w28050 ;
  assign w28052 = ~\pi092 & w28051 ;
  assign w28053 = w27694 & w27974 ;
  assign w28054 = ~w27701 & w27926 ;
  assign w28055 = w27927 ^ w28054 ;
  assign w28056 = ~w27974 & w28055 ;
  assign w28057 = w28053 | w28056 ;
  assign w28058 = ~\pi091 & w28057 ;
  assign w28059 = w27700 & w27974 ;
  assign w28060 = ~w27707 & w27923 ;
  assign w28061 = w27924 ^ w28060 ;
  assign w28062 = ~w27974 & w28061 ;
  assign w28063 = w28059 | w28062 ;
  assign w28064 = ~\pi090 & w28063 ;
  assign w28065 = w27706 & w27974 ;
  assign w28066 = ~w27713 & w27920 ;
  assign w28067 = w27921 ^ w28066 ;
  assign w28068 = ~w27974 & w28067 ;
  assign w28069 = w28065 | w28068 ;
  assign w28070 = ~\pi089 & w28069 ;
  assign w28071 = w27712 & w27974 ;
  assign w28072 = ~w27719 & w27917 ;
  assign w28073 = w27918 ^ w28072 ;
  assign w28074 = ~w27974 & w28073 ;
  assign w28075 = w28071 | w28074 ;
  assign w28076 = ~\pi088 & w28075 ;
  assign w28077 = w27718 & w27974 ;
  assign w28078 = ~w27725 & w27914 ;
  assign w28079 = w27915 ^ w28078 ;
  assign w28080 = ~w27974 & w28079 ;
  assign w28081 = w28077 | w28080 ;
  assign w28082 = ~\pi087 & w28081 ;
  assign w28083 = w27724 & w27974 ;
  assign w28084 = ~w27731 & w27911 ;
  assign w28085 = w27912 ^ w28084 ;
  assign w28086 = ~w27974 & w28085 ;
  assign w28087 = w28083 | w28086 ;
  assign w28088 = ~\pi086 & w28087 ;
  assign w28089 = w27730 & w27974 ;
  assign w28090 = ~w27737 & w27908 ;
  assign w28091 = w27909 ^ w28090 ;
  assign w28092 = ~w27974 & w28091 ;
  assign w28093 = w28089 | w28092 ;
  assign w28094 = ~\pi085 & w28093 ;
  assign w28095 = w27736 & w27974 ;
  assign w28096 = ~w27743 & w27905 ;
  assign w28097 = w27906 ^ w28096 ;
  assign w28098 = ~w27974 & w28097 ;
  assign w28099 = w28095 | w28098 ;
  assign w28100 = ~\pi084 & w28099 ;
  assign w28101 = w27742 & w27974 ;
  assign w28102 = ~w27749 & w27902 ;
  assign w28103 = w27903 ^ w28102 ;
  assign w28104 = ~w27974 & w28103 ;
  assign w28105 = w28101 | w28104 ;
  assign w28106 = ~\pi083 & w28105 ;
  assign w28107 = w27748 & w27974 ;
  assign w28108 = ~w27755 & w27899 ;
  assign w28109 = w27900 ^ w28108 ;
  assign w28110 = ~w27974 & w28109 ;
  assign w28111 = w28107 | w28110 ;
  assign w28112 = ~\pi082 & w28111 ;
  assign w28113 = w27754 & w27974 ;
  assign w28114 = ~w27761 & w27896 ;
  assign w28115 = w27897 ^ w28114 ;
  assign w28116 = ~w27974 & w28115 ;
  assign w28117 = w28113 | w28116 ;
  assign w28118 = ~\pi081 & w28117 ;
  assign w28119 = w27760 & w27974 ;
  assign w28120 = ~w27767 & w27893 ;
  assign w28121 = w27894 ^ w28120 ;
  assign w28122 = ~w27974 & w28121 ;
  assign w28123 = w28119 | w28122 ;
  assign w28124 = ~\pi080 & w28123 ;
  assign w28125 = w27766 & w27974 ;
  assign w28126 = ~w27773 & w27890 ;
  assign w28127 = w27891 ^ w28126 ;
  assign w28128 = ~w27974 & w28127 ;
  assign w28129 = w28125 | w28128 ;
  assign w28130 = ~\pi079 & w28129 ;
  assign w28131 = w27772 & w27974 ;
  assign w28132 = ~w27779 & w27887 ;
  assign w28133 = w27888 ^ w28132 ;
  assign w28134 = ~w27974 & w28133 ;
  assign w28135 = w28131 | w28134 ;
  assign w28136 = ~\pi078 & w28135 ;
  assign w28137 = w27778 & w27974 ;
  assign w28138 = ~w27785 & w27884 ;
  assign w28139 = w27885 ^ w28138 ;
  assign w28140 = ~w27974 & w28139 ;
  assign w28141 = w28137 | w28140 ;
  assign w28142 = ~\pi077 & w28141 ;
  assign w28143 = w27784 & w27974 ;
  assign w28144 = ~w27791 & w27881 ;
  assign w28145 = w27882 ^ w28144 ;
  assign w28146 = ~w27974 & w28145 ;
  assign w28147 = w28143 | w28146 ;
  assign w28148 = ~\pi076 & w28147 ;
  assign w28149 = w27790 & w27974 ;
  assign w28150 = ~w27797 & w27878 ;
  assign w28151 = w27879 ^ w28150 ;
  assign w28152 = ~w27974 & w28151 ;
  assign w28153 = w28149 | w28152 ;
  assign w28154 = ~\pi075 & w28153 ;
  assign w28155 = w27796 & w27974 ;
  assign w28156 = ~w27803 & w27875 ;
  assign w28157 = w27876 ^ w28156 ;
  assign w28158 = ~w27974 & w28157 ;
  assign w28159 = w28155 | w28158 ;
  assign w28160 = ~\pi074 & w28159 ;
  assign w28161 = w27802 & w27974 ;
  assign w28162 = ~w27809 & w27872 ;
  assign w28163 = w27873 ^ w28162 ;
  assign w28164 = ~w27974 & w28163 ;
  assign w28165 = w28161 | w28164 ;
  assign w28166 = ~\pi073 & w28165 ;
  assign w28167 = w27808 & w27974 ;
  assign w28168 = ~w27815 & w27869 ;
  assign w28169 = w27870 ^ w28168 ;
  assign w28170 = ~w27974 & w28169 ;
  assign w28171 = w28167 | w28170 ;
  assign w28172 = ~\pi072 & w28171 ;
  assign w28173 = w27814 & w27974 ;
  assign w28174 = ~w27821 & w27866 ;
  assign w28175 = w27867 ^ w28174 ;
  assign w28176 = ~w27974 & w28175 ;
  assign w28177 = w28173 | w28176 ;
  assign w28178 = ~\pi071 & w28177 ;
  assign w28179 = w27820 & w27974 ;
  assign w28180 = ~w27827 & w27863 ;
  assign w28181 = w27864 ^ w28180 ;
  assign w28182 = ~w27974 & w28181 ;
  assign w28183 = w28179 | w28182 ;
  assign w28184 = ~\pi070 & w28183 ;
  assign w28185 = w27826 & w27974 ;
  assign w28186 = ~w27836 & w27860 ;
  assign w28187 = w27861 ^ w28186 ;
  assign w28188 = ~w27974 & w28187 ;
  assign w28189 = w28185 | w28188 ;
  assign w28190 = ~\pi069 & w28189 ;
  assign w28191 = w27835 & w27974 ;
  assign w28192 = ~w27846 & w27857 ;
  assign w28193 = w27858 ^ w28192 ;
  assign w28194 = ~w27974 & w28193 ;
  assign w28195 = w28191 | w28194 ;
  assign w28196 = ~\pi068 & w28195 ;
  assign w28197 = w27845 & w27974 ;
  assign w28198 = w27854 ^ w27856 ;
  assign w28199 = ( w6588 & w27973 ) | ( w6588 & w28198 ) | ( w27973 & w28198 ) ;
  assign w28200 = w28198 & ~w28199 ;
  assign w28201 = w28197 | w28200 ;
  assign w28202 = ~\pi067 & w28201 ;
  assign w28203 = ( ~w6588 & w27848 ) | ( ~w6588 & w27851 ) | ( w27848 & w27851 ) ;
  assign w28204 = \pi065 ^ w28203 ;
  assign w28205 = ( ~w6588 & w8422 ) | ( ~w6588 & w28204 ) | ( w8422 & w28204 ) ;
  assign w28206 = ( w8422 & w27973 ) | ( w8422 & w28204 ) | ( w27973 & w28204 ) ;
  assign w28207 = w28205 & ~w28206 ;
  assign w28208 = w27855 & ~w27974 ;
  assign w28209 = ( w27855 & w28207 ) | ( w27855 & ~w28208 ) | ( w28207 & ~w28208 ) ;
  assign w28210 = ~\pi066 & w28209 ;
  assign w28211 = ( \pi023 & ~w8785 ) | ( \pi023 & w27973 ) | ( ~w8785 & w27973 ) ;
  assign w28212 = \pi023 & w28211 ;
  assign w28213 = w8789 & ~w27973 ;
  assign w28214 = w28212 | w28213 ;
  assign w28215 = \pi065 ^ w28214 ;
  assign w28216 = w8792 | w28215 ;
  assign w28217 = \pi066 ^ w28209 ;
  assign w28218 = ~\pi065 & w28214 ;
  assign w28219 = w28216 | w28218 ;
  assign w28220 = ( w28217 & ~w28218 ) | ( w28217 & w28219 ) | ( ~w28218 & w28219 ) ;
  assign w28221 = \pi067 ^ w28201 ;
  assign w28222 = ( ~w28210 & w28220 ) | ( ~w28210 & w28221 ) | ( w28220 & w28221 ) ;
  assign w28223 = w28221 | w28222 ;
  assign w28224 = \pi068 ^ w28195 ;
  assign w28225 = ( ~w28202 & w28223 ) | ( ~w28202 & w28224 ) | ( w28223 & w28224 ) ;
  assign w28226 = w28224 | w28225 ;
  assign w28227 = \pi069 ^ w28189 ;
  assign w28228 = ( ~w28196 & w28226 ) | ( ~w28196 & w28227 ) | ( w28226 & w28227 ) ;
  assign w28229 = w28227 | w28228 ;
  assign w28230 = \pi070 ^ w28183 ;
  assign w28231 = ( ~w28190 & w28229 ) | ( ~w28190 & w28230 ) | ( w28229 & w28230 ) ;
  assign w28232 = w28230 | w28231 ;
  assign w28233 = \pi071 ^ w28177 ;
  assign w28234 = ( ~w28184 & w28232 ) | ( ~w28184 & w28233 ) | ( w28232 & w28233 ) ;
  assign w28235 = w28233 | w28234 ;
  assign w28236 = \pi072 ^ w28171 ;
  assign w28237 = ( ~w28178 & w28235 ) | ( ~w28178 & w28236 ) | ( w28235 & w28236 ) ;
  assign w28238 = w28236 | w28237 ;
  assign w28239 = \pi073 ^ w28165 ;
  assign w28240 = ( ~w28172 & w28238 ) | ( ~w28172 & w28239 ) | ( w28238 & w28239 ) ;
  assign w28241 = w28239 | w28240 ;
  assign w28242 = \pi074 ^ w28159 ;
  assign w28243 = ( ~w28166 & w28241 ) | ( ~w28166 & w28242 ) | ( w28241 & w28242 ) ;
  assign w28244 = w28242 | w28243 ;
  assign w28245 = \pi075 ^ w28153 ;
  assign w28246 = ( ~w28160 & w28244 ) | ( ~w28160 & w28245 ) | ( w28244 & w28245 ) ;
  assign w28247 = w28245 | w28246 ;
  assign w28248 = \pi076 ^ w28147 ;
  assign w28249 = ( ~w28154 & w28247 ) | ( ~w28154 & w28248 ) | ( w28247 & w28248 ) ;
  assign w28250 = w28248 | w28249 ;
  assign w28251 = \pi077 ^ w28141 ;
  assign w28252 = ( ~w28148 & w28250 ) | ( ~w28148 & w28251 ) | ( w28250 & w28251 ) ;
  assign w28253 = w28251 | w28252 ;
  assign w28254 = \pi078 ^ w28135 ;
  assign w28255 = ( ~w28142 & w28253 ) | ( ~w28142 & w28254 ) | ( w28253 & w28254 ) ;
  assign w28256 = w28254 | w28255 ;
  assign w28257 = \pi079 ^ w28129 ;
  assign w28258 = ( ~w28136 & w28256 ) | ( ~w28136 & w28257 ) | ( w28256 & w28257 ) ;
  assign w28259 = w28257 | w28258 ;
  assign w28260 = \pi080 ^ w28123 ;
  assign w28261 = ( ~w28130 & w28259 ) | ( ~w28130 & w28260 ) | ( w28259 & w28260 ) ;
  assign w28262 = w28260 | w28261 ;
  assign w28263 = \pi081 ^ w28117 ;
  assign w28264 = ( ~w28124 & w28262 ) | ( ~w28124 & w28263 ) | ( w28262 & w28263 ) ;
  assign w28265 = w28263 | w28264 ;
  assign w28266 = \pi082 ^ w28111 ;
  assign w28267 = ( ~w28118 & w28265 ) | ( ~w28118 & w28266 ) | ( w28265 & w28266 ) ;
  assign w28268 = w28266 | w28267 ;
  assign w28269 = \pi083 ^ w28105 ;
  assign w28270 = ( ~w28112 & w28268 ) | ( ~w28112 & w28269 ) | ( w28268 & w28269 ) ;
  assign w28271 = w28269 | w28270 ;
  assign w28272 = \pi084 ^ w28099 ;
  assign w28273 = ( ~w28106 & w28271 ) | ( ~w28106 & w28272 ) | ( w28271 & w28272 ) ;
  assign w28274 = w28272 | w28273 ;
  assign w28275 = \pi085 ^ w28093 ;
  assign w28276 = ( ~w28100 & w28274 ) | ( ~w28100 & w28275 ) | ( w28274 & w28275 ) ;
  assign w28277 = w28275 | w28276 ;
  assign w28278 = \pi086 ^ w28087 ;
  assign w28279 = ( ~w28094 & w28277 ) | ( ~w28094 & w28278 ) | ( w28277 & w28278 ) ;
  assign w28280 = w28278 | w28279 ;
  assign w28281 = \pi087 ^ w28081 ;
  assign w28282 = ( ~w28088 & w28280 ) | ( ~w28088 & w28281 ) | ( w28280 & w28281 ) ;
  assign w28283 = w28281 | w28282 ;
  assign w28284 = \pi088 ^ w28075 ;
  assign w28285 = ( ~w28082 & w28283 ) | ( ~w28082 & w28284 ) | ( w28283 & w28284 ) ;
  assign w28286 = w28284 | w28285 ;
  assign w28287 = \pi089 ^ w28069 ;
  assign w28288 = ( ~w28076 & w28286 ) | ( ~w28076 & w28287 ) | ( w28286 & w28287 ) ;
  assign w28289 = w28287 | w28288 ;
  assign w28290 = \pi090 ^ w28063 ;
  assign w28291 = ( ~w28070 & w28289 ) | ( ~w28070 & w28290 ) | ( w28289 & w28290 ) ;
  assign w28292 = w28290 | w28291 ;
  assign w28293 = \pi091 ^ w28057 ;
  assign w28294 = ( ~w28064 & w28292 ) | ( ~w28064 & w28293 ) | ( w28292 & w28293 ) ;
  assign w28295 = w28293 | w28294 ;
  assign w28296 = \pi092 ^ w28051 ;
  assign w28297 = ( ~w28058 & w28295 ) | ( ~w28058 & w28296 ) | ( w28295 & w28296 ) ;
  assign w28298 = w28296 | w28297 ;
  assign w28299 = \pi093 ^ w28045 ;
  assign w28300 = ( ~w28052 & w28298 ) | ( ~w28052 & w28299 ) | ( w28298 & w28299 ) ;
  assign w28301 = w28299 | w28300 ;
  assign w28302 = \pi094 ^ w28039 ;
  assign w28303 = ( ~w28046 & w28301 ) | ( ~w28046 & w28302 ) | ( w28301 & w28302 ) ;
  assign w28304 = w28302 | w28303 ;
  assign w28305 = \pi095 ^ w28033 ;
  assign w28306 = ( ~w28040 & w28304 ) | ( ~w28040 & w28305 ) | ( w28304 & w28305 ) ;
  assign w28307 = w28305 | w28306 ;
  assign w28308 = \pi096 ^ w28027 ;
  assign w28309 = ( ~w28034 & w28307 ) | ( ~w28034 & w28308 ) | ( w28307 & w28308 ) ;
  assign w28310 = w28308 | w28309 ;
  assign w28311 = \pi097 ^ w28021 ;
  assign w28312 = ( ~w28028 & w28310 ) | ( ~w28028 & w28311 ) | ( w28310 & w28311 ) ;
  assign w28313 = w28311 | w28312 ;
  assign w28314 = \pi098 ^ w28015 ;
  assign w28315 = ( ~w28022 & w28313 ) | ( ~w28022 & w28314 ) | ( w28313 & w28314 ) ;
  assign w28316 = w28314 | w28315 ;
  assign w28317 = \pi099 ^ w28009 ;
  assign w28318 = ( ~w28016 & w28316 ) | ( ~w28016 & w28317 ) | ( w28316 & w28317 ) ;
  assign w28319 = w28317 | w28318 ;
  assign w28320 = \pi100 ^ w28003 ;
  assign w28321 = ( ~w28010 & w28319 ) | ( ~w28010 & w28320 ) | ( w28319 & w28320 ) ;
  assign w28322 = w28320 | w28321 ;
  assign w28323 = \pi101 ^ w27997 ;
  assign w28324 = ( ~w28004 & w28322 ) | ( ~w28004 & w28323 ) | ( w28322 & w28323 ) ;
  assign w28325 = w28323 | w28324 ;
  assign w28326 = \pi102 ^ w27991 ;
  assign w28327 = ( ~w27998 & w28325 ) | ( ~w27998 & w28326 ) | ( w28325 & w28326 ) ;
  assign w28328 = w28326 | w28327 ;
  assign w28329 = \pi103 ^ w27985 ;
  assign w28330 = ( ~w27992 & w28328 ) | ( ~w27992 & w28329 ) | ( w28328 & w28329 ) ;
  assign w28331 = w28329 | w28330 ;
  assign w28332 = \pi104 ^ w27979 ;
  assign w28333 = ( ~w27986 & w28331 ) | ( ~w27986 & w28332 ) | ( w28331 & w28332 ) ;
  assign w28334 = w28332 | w28333 ;
  assign w28335 = w27616 & w27974 ;
  assign w28336 = ~w27617 & w27968 ;
  assign w28337 = w27969 ^ w28336 ;
  assign w28338 = ~w27974 & w28337 ;
  assign w28339 = w28335 | w28338 ;
  assign w28340 = ~\pi105 & w28339 ;
  assign w28341 = ( \pi105 & ~w28335 ) | ( \pi105 & w28338 ) | ( ~w28335 & w28338 ) ;
  assign w28342 = ~w28338 & w28341 ;
  assign w28343 = ( ~w27980 & w28334 ) | ( ~w27980 & w28340 ) | ( w28334 & w28340 ) ;
  assign w28344 = ( w8924 & w28340 ) | ( w8924 & ~w28343 ) | ( w28340 & ~w28343 ) ;
  assign w28345 = ( w201 & w28342 ) | ( w201 & ~w28343 ) | ( w28342 & ~w28343 ) ;
  assign w28346 = ( w28343 & ~w28344 ) | ( w28343 & w28345 ) | ( ~w28344 & w28345 ) ;
  assign w28347 = w28344 | w28346 ;
  assign w28348 = ~w6588 & w28339 ;
  assign w28349 = w28347 & ~w28348 ;
  assign w28350 = ~w27986 & w28331 ;
  assign w28351 = w28332 ^ w28350 ;
  assign w28352 = ~w28349 & w28351 ;
  assign w28353 = ( w27979 & w28347 ) | ( w27979 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28354 = ~w28348 & w28353 ;
  assign w28355 = w28352 | w28354 ;
  assign w28356 = w28340 | w28342 ;
  assign w28357 = ( ~w27980 & w28334 ) | ( ~w27980 & w28349 ) | ( w28334 & w28349 ) ;
  assign w28358 = w28356 ^ w28357 ;
  assign w28359 = ~w28349 & w28358 ;
  assign w28360 = ( w6588 & ~w28339 ) | ( w6588 & w28347 ) | ( ~w28339 & w28347 ) ;
  assign w28361 = w28339 & w28360 ;
  assign w28362 = w28359 | w28361 ;
  assign w28363 = ~\pi105 & w28355 ;
  assign w28364 = ~w27992 & w28328 ;
  assign w28365 = w28329 ^ w28364 ;
  assign w28366 = ~w28349 & w28365 ;
  assign w28367 = ( w27985 & w28347 ) | ( w27985 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28368 = ~w28348 & w28367 ;
  assign w28369 = w28366 | w28368 ;
  assign w28370 = ~\pi104 & w28369 ;
  assign w28371 = ~w27998 & w28325 ;
  assign w28372 = w28326 ^ w28371 ;
  assign w28373 = ~w28349 & w28372 ;
  assign w28374 = ( w27991 & w28347 ) | ( w27991 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28375 = ~w28348 & w28374 ;
  assign w28376 = w28373 | w28375 ;
  assign w28377 = ~\pi103 & w28376 ;
  assign w28378 = ~w28004 & w28322 ;
  assign w28379 = w28323 ^ w28378 ;
  assign w28380 = ~w28349 & w28379 ;
  assign w28381 = ( w27997 & w28347 ) | ( w27997 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28382 = ~w28348 & w28381 ;
  assign w28383 = w28380 | w28382 ;
  assign w28384 = ~\pi102 & w28383 ;
  assign w28385 = ~w28010 & w28319 ;
  assign w28386 = w28320 ^ w28385 ;
  assign w28387 = ~w28349 & w28386 ;
  assign w28388 = ( w28003 & w28347 ) | ( w28003 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28389 = ~w28348 & w28388 ;
  assign w28390 = w28387 | w28389 ;
  assign w28391 = ~\pi101 & w28390 ;
  assign w28392 = ~w28016 & w28316 ;
  assign w28393 = w28317 ^ w28392 ;
  assign w28394 = ~w28349 & w28393 ;
  assign w28395 = ( w28009 & w28347 ) | ( w28009 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28396 = ~w28348 & w28395 ;
  assign w28397 = w28394 | w28396 ;
  assign w28398 = ~\pi100 & w28397 ;
  assign w28399 = ~w28022 & w28313 ;
  assign w28400 = w28314 ^ w28399 ;
  assign w28401 = ~w28349 & w28400 ;
  assign w28402 = ( w28015 & w28347 ) | ( w28015 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28403 = ~w28348 & w28402 ;
  assign w28404 = w28401 | w28403 ;
  assign w28405 = ~\pi099 & w28404 ;
  assign w28406 = ~w28028 & w28310 ;
  assign w28407 = w28311 ^ w28406 ;
  assign w28408 = ~w28349 & w28407 ;
  assign w28409 = ( w28021 & w28347 ) | ( w28021 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28410 = ~w28348 & w28409 ;
  assign w28411 = w28408 | w28410 ;
  assign w28412 = ~\pi098 & w28411 ;
  assign w28413 = ~w28034 & w28307 ;
  assign w28414 = w28308 ^ w28413 ;
  assign w28415 = ~w28349 & w28414 ;
  assign w28416 = ( w28027 & w28347 ) | ( w28027 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28417 = ~w28348 & w28416 ;
  assign w28418 = w28415 | w28417 ;
  assign w28419 = ~\pi097 & w28418 ;
  assign w28420 = ~w28040 & w28304 ;
  assign w28421 = w28305 ^ w28420 ;
  assign w28422 = ~w28349 & w28421 ;
  assign w28423 = ( w28033 & w28347 ) | ( w28033 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28424 = ~w28348 & w28423 ;
  assign w28425 = w28422 | w28424 ;
  assign w28426 = ~\pi096 & w28425 ;
  assign w28427 = ~w28046 & w28301 ;
  assign w28428 = w28302 ^ w28427 ;
  assign w28429 = ~w28349 & w28428 ;
  assign w28430 = ( w28039 & w28347 ) | ( w28039 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28431 = ~w28348 & w28430 ;
  assign w28432 = w28429 | w28431 ;
  assign w28433 = ~\pi095 & w28432 ;
  assign w28434 = ~w28052 & w28298 ;
  assign w28435 = w28299 ^ w28434 ;
  assign w28436 = ~w28349 & w28435 ;
  assign w28437 = ( w28045 & w28347 ) | ( w28045 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28438 = ~w28348 & w28437 ;
  assign w28439 = w28436 | w28438 ;
  assign w28440 = ~\pi094 & w28439 ;
  assign w28441 = ~w28058 & w28295 ;
  assign w28442 = w28296 ^ w28441 ;
  assign w28443 = ~w28349 & w28442 ;
  assign w28444 = ( w28051 & w28347 ) | ( w28051 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28445 = ~w28348 & w28444 ;
  assign w28446 = w28443 | w28445 ;
  assign w28447 = ~\pi093 & w28446 ;
  assign w28448 = ~w28064 & w28292 ;
  assign w28449 = w28293 ^ w28448 ;
  assign w28450 = ~w28349 & w28449 ;
  assign w28451 = ( w28057 & w28347 ) | ( w28057 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28452 = ~w28348 & w28451 ;
  assign w28453 = w28450 | w28452 ;
  assign w28454 = ~\pi092 & w28453 ;
  assign w28455 = ~w28070 & w28289 ;
  assign w28456 = w28290 ^ w28455 ;
  assign w28457 = ~w28349 & w28456 ;
  assign w28458 = ( w28063 & w28347 ) | ( w28063 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28459 = ~w28348 & w28458 ;
  assign w28460 = w28457 | w28459 ;
  assign w28461 = ~\pi091 & w28460 ;
  assign w28462 = ~w28076 & w28286 ;
  assign w28463 = w28287 ^ w28462 ;
  assign w28464 = ~w28349 & w28463 ;
  assign w28465 = ( w28069 & w28347 ) | ( w28069 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28466 = ~w28348 & w28465 ;
  assign w28467 = w28464 | w28466 ;
  assign w28468 = ~\pi090 & w28467 ;
  assign w28469 = ~w28082 & w28283 ;
  assign w28470 = w28284 ^ w28469 ;
  assign w28471 = ~w28349 & w28470 ;
  assign w28472 = ( w28075 & w28347 ) | ( w28075 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28473 = ~w28348 & w28472 ;
  assign w28474 = w28471 | w28473 ;
  assign w28475 = ~\pi089 & w28474 ;
  assign w28476 = ~w28088 & w28280 ;
  assign w28477 = w28281 ^ w28476 ;
  assign w28478 = ~w28349 & w28477 ;
  assign w28479 = ( w28081 & w28347 ) | ( w28081 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28480 = ~w28348 & w28479 ;
  assign w28481 = w28478 | w28480 ;
  assign w28482 = ~\pi088 & w28481 ;
  assign w28483 = ~w28094 & w28277 ;
  assign w28484 = w28278 ^ w28483 ;
  assign w28485 = ~w28349 & w28484 ;
  assign w28486 = ( w28087 & w28347 ) | ( w28087 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28487 = ~w28348 & w28486 ;
  assign w28488 = w28485 | w28487 ;
  assign w28489 = ~\pi087 & w28488 ;
  assign w28490 = ~w28100 & w28274 ;
  assign w28491 = w28275 ^ w28490 ;
  assign w28492 = ~w28349 & w28491 ;
  assign w28493 = ( w28093 & w28347 ) | ( w28093 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28494 = ~w28348 & w28493 ;
  assign w28495 = w28492 | w28494 ;
  assign w28496 = ~\pi086 & w28495 ;
  assign w28497 = ~w28106 & w28271 ;
  assign w28498 = w28272 ^ w28497 ;
  assign w28499 = ~w28349 & w28498 ;
  assign w28500 = ( w28099 & w28347 ) | ( w28099 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28501 = ~w28348 & w28500 ;
  assign w28502 = w28499 | w28501 ;
  assign w28503 = ~\pi085 & w28502 ;
  assign w28504 = ~w28112 & w28268 ;
  assign w28505 = w28269 ^ w28504 ;
  assign w28506 = ~w28349 & w28505 ;
  assign w28507 = ( w28105 & w28347 ) | ( w28105 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28508 = ~w28348 & w28507 ;
  assign w28509 = w28506 | w28508 ;
  assign w28510 = ~\pi084 & w28509 ;
  assign w28511 = ~w28118 & w28265 ;
  assign w28512 = w28266 ^ w28511 ;
  assign w28513 = ~w28349 & w28512 ;
  assign w28514 = ( w28111 & w28347 ) | ( w28111 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28515 = ~w28348 & w28514 ;
  assign w28516 = w28513 | w28515 ;
  assign w28517 = ~\pi083 & w28516 ;
  assign w28518 = ~w28124 & w28262 ;
  assign w28519 = w28263 ^ w28518 ;
  assign w28520 = ~w28349 & w28519 ;
  assign w28521 = ( w28117 & w28347 ) | ( w28117 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28522 = ~w28348 & w28521 ;
  assign w28523 = w28520 | w28522 ;
  assign w28524 = ~\pi082 & w28523 ;
  assign w28525 = ~w28130 & w28259 ;
  assign w28526 = w28260 ^ w28525 ;
  assign w28527 = ~w28349 & w28526 ;
  assign w28528 = ( w28123 & w28347 ) | ( w28123 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28529 = ~w28348 & w28528 ;
  assign w28530 = w28527 | w28529 ;
  assign w28531 = ~\pi081 & w28530 ;
  assign w28532 = ~w28136 & w28256 ;
  assign w28533 = w28257 ^ w28532 ;
  assign w28534 = ~w28349 & w28533 ;
  assign w28535 = ( w28129 & w28347 ) | ( w28129 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28536 = ~w28348 & w28535 ;
  assign w28537 = w28534 | w28536 ;
  assign w28538 = ~\pi080 & w28537 ;
  assign w28539 = ~w28142 & w28253 ;
  assign w28540 = w28254 ^ w28539 ;
  assign w28541 = ~w28349 & w28540 ;
  assign w28542 = ( w28135 & w28347 ) | ( w28135 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28543 = ~w28348 & w28542 ;
  assign w28544 = w28541 | w28543 ;
  assign w28545 = ~\pi079 & w28544 ;
  assign w28546 = ~w28148 & w28250 ;
  assign w28547 = w28251 ^ w28546 ;
  assign w28548 = ~w28349 & w28547 ;
  assign w28549 = ( w28141 & w28347 ) | ( w28141 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28550 = ~w28348 & w28549 ;
  assign w28551 = w28548 | w28550 ;
  assign w28552 = ~\pi078 & w28551 ;
  assign w28553 = ~w28154 & w28247 ;
  assign w28554 = w28248 ^ w28553 ;
  assign w28555 = ~w28349 & w28554 ;
  assign w28556 = ( w28147 & w28347 ) | ( w28147 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28557 = ~w28348 & w28556 ;
  assign w28558 = w28555 | w28557 ;
  assign w28559 = ~\pi077 & w28558 ;
  assign w28560 = ~w28160 & w28244 ;
  assign w28561 = w28245 ^ w28560 ;
  assign w28562 = ~w28349 & w28561 ;
  assign w28563 = ( w28153 & w28347 ) | ( w28153 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28564 = ~w28348 & w28563 ;
  assign w28565 = w28562 | w28564 ;
  assign w28566 = ~\pi076 & w28565 ;
  assign w28567 = ~w28166 & w28241 ;
  assign w28568 = w28242 ^ w28567 ;
  assign w28569 = ~w28349 & w28568 ;
  assign w28570 = ( w28159 & w28347 ) | ( w28159 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28571 = ~w28348 & w28570 ;
  assign w28572 = w28569 | w28571 ;
  assign w28573 = ~\pi075 & w28572 ;
  assign w28574 = ~w28172 & w28238 ;
  assign w28575 = w28239 ^ w28574 ;
  assign w28576 = ~w28349 & w28575 ;
  assign w28577 = ( w28165 & w28347 ) | ( w28165 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28578 = ~w28348 & w28577 ;
  assign w28579 = w28576 | w28578 ;
  assign w28580 = ~\pi074 & w28579 ;
  assign w28581 = ~w28178 & w28235 ;
  assign w28582 = w28236 ^ w28581 ;
  assign w28583 = ~w28349 & w28582 ;
  assign w28584 = ( w28171 & w28347 ) | ( w28171 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28585 = ~w28348 & w28584 ;
  assign w28586 = w28583 | w28585 ;
  assign w28587 = ~\pi073 & w28586 ;
  assign w28588 = ~w28184 & w28232 ;
  assign w28589 = w28233 ^ w28588 ;
  assign w28590 = ~w28349 & w28589 ;
  assign w28591 = ( w28177 & w28347 ) | ( w28177 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28592 = ~w28348 & w28591 ;
  assign w28593 = w28590 | w28592 ;
  assign w28594 = ~\pi072 & w28593 ;
  assign w28595 = ~w28190 & w28229 ;
  assign w28596 = w28230 ^ w28595 ;
  assign w28597 = ~w28349 & w28596 ;
  assign w28598 = ( w28183 & w28347 ) | ( w28183 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28599 = ~w28348 & w28598 ;
  assign w28600 = w28597 | w28599 ;
  assign w28601 = ~\pi071 & w28600 ;
  assign w28602 = ~w28196 & w28226 ;
  assign w28603 = w28227 ^ w28602 ;
  assign w28604 = ~w28349 & w28603 ;
  assign w28605 = ( w28189 & w28347 ) | ( w28189 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28606 = ~w28348 & w28605 ;
  assign w28607 = w28604 | w28606 ;
  assign w28608 = ~\pi070 & w28607 ;
  assign w28609 = ~w28202 & w28223 ;
  assign w28610 = w28224 ^ w28609 ;
  assign w28611 = ~w28349 & w28610 ;
  assign w28612 = ( w28195 & w28347 ) | ( w28195 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28613 = ~w28348 & w28612 ;
  assign w28614 = w28611 | w28613 ;
  assign w28615 = ~\pi069 & w28614 ;
  assign w28616 = ~w28210 & w28220 ;
  assign w28617 = w28221 ^ w28616 ;
  assign w28618 = ~w28349 & w28617 ;
  assign w28619 = ( w28201 & w28347 ) | ( w28201 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28620 = ~w28348 & w28619 ;
  assign w28621 = w28618 | w28620 ;
  assign w28622 = ~\pi068 & w28621 ;
  assign w28623 = ( \pi065 & w28214 ) | ( \pi065 & ~w28349 ) | ( w28214 & ~w28349 ) ;
  assign w28624 = ( \pi065 & w28216 ) | ( \pi065 & ~w28623 ) | ( w28216 & ~w28623 ) ;
  assign w28625 = w28217 ^ w28624 ;
  assign w28626 = ~w28349 & w28625 ;
  assign w28627 = ( w28209 & w28347 ) | ( w28209 & w28348 ) | ( w28347 & w28348 ) ;
  assign w28628 = ~w28348 & w28627 ;
  assign w28629 = w28626 | w28628 ;
  assign w28630 = ~\pi067 & w28629 ;
  assign w28631 = w8792 ^ w28214 ;
  assign w28632 = \pi065 ^ w28631 ;
  assign w28633 = w28349 ^ w28632 ;
  assign w28634 = ( w28214 & w28632 ) | ( w28214 & w28633 ) | ( w28632 & w28633 ) ;
  assign w28635 = ~\pi066 & w28634 ;
  assign w28636 = w28214 ^ w28349 ;
  assign w28637 = ( w28214 & w28632 ) | ( w28214 & ~w28636 ) | ( w28632 & ~w28636 ) ;
  assign w28638 = \pi066 ^ w28637 ;
  assign w28639 = ( \pi064 & ~w28349 ) | ( \pi064 & w28638 ) | ( ~w28349 & w28638 ) ;
  assign w28640 = \pi022 ^ w28639 ;
  assign w28641 = ( \pi065 & w9218 ) | ( \pi065 & ~w28640 ) | ( w9218 & ~w28640 ) ;
  assign w28642 = w28638 | w28641 ;
  assign w28643 = \pi067 ^ w28629 ;
  assign w28644 = ( ~w28635 & w28642 ) | ( ~w28635 & w28643 ) | ( w28642 & w28643 ) ;
  assign w28645 = w28643 | w28644 ;
  assign w28646 = \pi068 ^ w28621 ;
  assign w28647 = ( ~w28630 & w28645 ) | ( ~w28630 & w28646 ) | ( w28645 & w28646 ) ;
  assign w28648 = w28646 | w28647 ;
  assign w28649 = \pi069 ^ w28614 ;
  assign w28650 = ( ~w28622 & w28648 ) | ( ~w28622 & w28649 ) | ( w28648 & w28649 ) ;
  assign w28651 = w28649 | w28650 ;
  assign w28652 = \pi070 ^ w28607 ;
  assign w28653 = ( ~w28615 & w28651 ) | ( ~w28615 & w28652 ) | ( w28651 & w28652 ) ;
  assign w28654 = w28652 | w28653 ;
  assign w28655 = \pi071 ^ w28600 ;
  assign w28656 = ( ~w28608 & w28654 ) | ( ~w28608 & w28655 ) | ( w28654 & w28655 ) ;
  assign w28657 = w28655 | w28656 ;
  assign w28658 = \pi072 ^ w28593 ;
  assign w28659 = ( ~w28601 & w28657 ) | ( ~w28601 & w28658 ) | ( w28657 & w28658 ) ;
  assign w28660 = w28658 | w28659 ;
  assign w28661 = \pi073 ^ w28586 ;
  assign w28662 = ( ~w28594 & w28660 ) | ( ~w28594 & w28661 ) | ( w28660 & w28661 ) ;
  assign w28663 = w28661 | w28662 ;
  assign w28664 = \pi074 ^ w28579 ;
  assign w28665 = ( ~w28587 & w28663 ) | ( ~w28587 & w28664 ) | ( w28663 & w28664 ) ;
  assign w28666 = w28664 | w28665 ;
  assign w28667 = \pi075 ^ w28572 ;
  assign w28668 = ( ~w28580 & w28666 ) | ( ~w28580 & w28667 ) | ( w28666 & w28667 ) ;
  assign w28669 = w28667 | w28668 ;
  assign w28670 = \pi076 ^ w28565 ;
  assign w28671 = ( ~w28573 & w28669 ) | ( ~w28573 & w28670 ) | ( w28669 & w28670 ) ;
  assign w28672 = w28670 | w28671 ;
  assign w28673 = \pi077 ^ w28558 ;
  assign w28674 = ( ~w28566 & w28672 ) | ( ~w28566 & w28673 ) | ( w28672 & w28673 ) ;
  assign w28675 = w28673 | w28674 ;
  assign w28676 = \pi078 ^ w28551 ;
  assign w28677 = ( ~w28559 & w28675 ) | ( ~w28559 & w28676 ) | ( w28675 & w28676 ) ;
  assign w28678 = w28676 | w28677 ;
  assign w28679 = \pi079 ^ w28544 ;
  assign w28680 = ( ~w28552 & w28678 ) | ( ~w28552 & w28679 ) | ( w28678 & w28679 ) ;
  assign w28681 = w28679 | w28680 ;
  assign w28682 = \pi080 ^ w28537 ;
  assign w28683 = ( ~w28545 & w28681 ) | ( ~w28545 & w28682 ) | ( w28681 & w28682 ) ;
  assign w28684 = w28682 | w28683 ;
  assign w28685 = \pi081 ^ w28530 ;
  assign w28686 = ( ~w28538 & w28684 ) | ( ~w28538 & w28685 ) | ( w28684 & w28685 ) ;
  assign w28687 = w28685 | w28686 ;
  assign w28688 = \pi082 ^ w28523 ;
  assign w28689 = ( ~w28531 & w28687 ) | ( ~w28531 & w28688 ) | ( w28687 & w28688 ) ;
  assign w28690 = w28688 | w28689 ;
  assign w28691 = \pi083 ^ w28516 ;
  assign w28692 = ( ~w28524 & w28690 ) | ( ~w28524 & w28691 ) | ( w28690 & w28691 ) ;
  assign w28693 = w28691 | w28692 ;
  assign w28694 = \pi084 ^ w28509 ;
  assign w28695 = ( ~w28517 & w28693 ) | ( ~w28517 & w28694 ) | ( w28693 & w28694 ) ;
  assign w28696 = w28694 | w28695 ;
  assign w28697 = \pi085 ^ w28502 ;
  assign w28698 = ( ~w28510 & w28696 ) | ( ~w28510 & w28697 ) | ( w28696 & w28697 ) ;
  assign w28699 = w28697 | w28698 ;
  assign w28700 = \pi086 ^ w28495 ;
  assign w28701 = ( ~w28503 & w28699 ) | ( ~w28503 & w28700 ) | ( w28699 & w28700 ) ;
  assign w28702 = w28700 | w28701 ;
  assign w28703 = \pi087 ^ w28488 ;
  assign w28704 = ( ~w28496 & w28702 ) | ( ~w28496 & w28703 ) | ( w28702 & w28703 ) ;
  assign w28705 = w28703 | w28704 ;
  assign w28706 = \pi088 ^ w28481 ;
  assign w28707 = ( ~w28489 & w28705 ) | ( ~w28489 & w28706 ) | ( w28705 & w28706 ) ;
  assign w28708 = w28706 | w28707 ;
  assign w28709 = \pi089 ^ w28474 ;
  assign w28710 = ( ~w28482 & w28708 ) | ( ~w28482 & w28709 ) | ( w28708 & w28709 ) ;
  assign w28711 = w28709 | w28710 ;
  assign w28712 = \pi090 ^ w28467 ;
  assign w28713 = ( ~w28475 & w28711 ) | ( ~w28475 & w28712 ) | ( w28711 & w28712 ) ;
  assign w28714 = w28712 | w28713 ;
  assign w28715 = \pi091 ^ w28460 ;
  assign w28716 = ( ~w28468 & w28714 ) | ( ~w28468 & w28715 ) | ( w28714 & w28715 ) ;
  assign w28717 = w28715 | w28716 ;
  assign w28718 = \pi092 ^ w28453 ;
  assign w28719 = ( ~w28461 & w28717 ) | ( ~w28461 & w28718 ) | ( w28717 & w28718 ) ;
  assign w28720 = w28718 | w28719 ;
  assign w28721 = \pi093 ^ w28446 ;
  assign w28722 = ( ~w28454 & w28720 ) | ( ~w28454 & w28721 ) | ( w28720 & w28721 ) ;
  assign w28723 = w28721 | w28722 ;
  assign w28724 = \pi094 ^ w28439 ;
  assign w28725 = ( ~w28447 & w28723 ) | ( ~w28447 & w28724 ) | ( w28723 & w28724 ) ;
  assign w28726 = w28724 | w28725 ;
  assign w28727 = \pi095 ^ w28432 ;
  assign w28728 = ( ~w28440 & w28726 ) | ( ~w28440 & w28727 ) | ( w28726 & w28727 ) ;
  assign w28729 = w28727 | w28728 ;
  assign w28730 = \pi096 ^ w28425 ;
  assign w28731 = ( ~w28433 & w28729 ) | ( ~w28433 & w28730 ) | ( w28729 & w28730 ) ;
  assign w28732 = w28730 | w28731 ;
  assign w28733 = \pi097 ^ w28418 ;
  assign w28734 = ( ~w28426 & w28732 ) | ( ~w28426 & w28733 ) | ( w28732 & w28733 ) ;
  assign w28735 = w28733 | w28734 ;
  assign w28736 = \pi098 ^ w28411 ;
  assign w28737 = ( ~w28419 & w28735 ) | ( ~w28419 & w28736 ) | ( w28735 & w28736 ) ;
  assign w28738 = w28736 | w28737 ;
  assign w28739 = \pi099 ^ w28404 ;
  assign w28740 = ( ~w28412 & w28738 ) | ( ~w28412 & w28739 ) | ( w28738 & w28739 ) ;
  assign w28741 = w28739 | w28740 ;
  assign w28742 = \pi100 ^ w28397 ;
  assign w28743 = ( ~w28405 & w28741 ) | ( ~w28405 & w28742 ) | ( w28741 & w28742 ) ;
  assign w28744 = w28742 | w28743 ;
  assign w28745 = \pi101 ^ w28390 ;
  assign w28746 = ( ~w28398 & w28744 ) | ( ~w28398 & w28745 ) | ( w28744 & w28745 ) ;
  assign w28747 = w28745 | w28746 ;
  assign w28748 = \pi102 ^ w28383 ;
  assign w28749 = ( ~w28391 & w28747 ) | ( ~w28391 & w28748 ) | ( w28747 & w28748 ) ;
  assign w28750 = w28748 | w28749 ;
  assign w28751 = \pi103 ^ w28376 ;
  assign w28752 = ( ~w28384 & w28750 ) | ( ~w28384 & w28751 ) | ( w28750 & w28751 ) ;
  assign w28753 = w28751 | w28752 ;
  assign w28754 = \pi104 ^ w28369 ;
  assign w28755 = ( ~w28377 & w28753 ) | ( ~w28377 & w28754 ) | ( w28753 & w28754 ) ;
  assign w28756 = w28754 | w28755 ;
  assign w28757 = \pi105 ^ w28355 ;
  assign w28758 = ( ~w28370 & w28756 ) | ( ~w28370 & w28757 ) | ( w28756 & w28757 ) ;
  assign w28759 = w28757 | w28758 ;
  assign w28760 = \pi106 ^ w28362 ;
  assign w28761 = w28363 & ~w28760 ;
  assign w28762 = ( w28759 & w28760 ) | ( w28759 & ~w28761 ) | ( w28760 & ~w28761 ) ;
  assign w28763 = ~\pi106 & w28362 ;
  assign w28764 = w28762 & ~w28763 ;
  assign w28765 = w9351 | w28764 ;
  assign w28766 = w28355 & w28765 ;
  assign w28767 = ~w28370 & w28756 ;
  assign w28768 = w28757 ^ w28767 ;
  assign w28769 = ~w28765 & w28768 ;
  assign w28770 = w28766 | w28769 ;
  assign w28771 = ~\pi106 & w28770 ;
  assign w28772 = w28369 & w28765 ;
  assign w28773 = ~w28377 & w28753 ;
  assign w28774 = w28754 ^ w28773 ;
  assign w28775 = ~w28765 & w28774 ;
  assign w28776 = w28772 | w28775 ;
  assign w28777 = ~\pi105 & w28776 ;
  assign w28778 = w28376 & w28765 ;
  assign w28779 = ~w28384 & w28750 ;
  assign w28780 = w28751 ^ w28779 ;
  assign w28781 = ~w28765 & w28780 ;
  assign w28782 = w28778 | w28781 ;
  assign w28783 = ~\pi104 & w28782 ;
  assign w28784 = w28383 & w28765 ;
  assign w28785 = ~w28391 & w28747 ;
  assign w28786 = w28748 ^ w28785 ;
  assign w28787 = ~w28765 & w28786 ;
  assign w28788 = w28784 | w28787 ;
  assign w28789 = ~\pi103 & w28788 ;
  assign w28790 = w28390 & w28765 ;
  assign w28791 = ~w28398 & w28744 ;
  assign w28792 = w28745 ^ w28791 ;
  assign w28793 = ~w28765 & w28792 ;
  assign w28794 = w28790 | w28793 ;
  assign w28795 = ~\pi102 & w28794 ;
  assign w28796 = w28397 & w28765 ;
  assign w28797 = ~w28405 & w28741 ;
  assign w28798 = w28742 ^ w28797 ;
  assign w28799 = ~w28765 & w28798 ;
  assign w28800 = w28796 | w28799 ;
  assign w28801 = ~\pi101 & w28800 ;
  assign w28802 = w28404 & w28765 ;
  assign w28803 = ~w28412 & w28738 ;
  assign w28804 = w28739 ^ w28803 ;
  assign w28805 = ~w28765 & w28804 ;
  assign w28806 = w28802 | w28805 ;
  assign w28807 = ~\pi100 & w28806 ;
  assign w28808 = w28411 & w28765 ;
  assign w28809 = ~w28419 & w28735 ;
  assign w28810 = w28736 ^ w28809 ;
  assign w28811 = ~w28765 & w28810 ;
  assign w28812 = w28808 | w28811 ;
  assign w28813 = ~\pi099 & w28812 ;
  assign w28814 = w28418 & w28765 ;
  assign w28815 = ~w28426 & w28732 ;
  assign w28816 = w28733 ^ w28815 ;
  assign w28817 = ~w28765 & w28816 ;
  assign w28818 = w28814 | w28817 ;
  assign w28819 = ~\pi098 & w28818 ;
  assign w28820 = w28425 & w28765 ;
  assign w28821 = ~w28433 & w28729 ;
  assign w28822 = w28730 ^ w28821 ;
  assign w28823 = ~w28765 & w28822 ;
  assign w28824 = w28820 | w28823 ;
  assign w28825 = ~\pi097 & w28824 ;
  assign w28826 = w28432 & w28765 ;
  assign w28827 = ~w28440 & w28726 ;
  assign w28828 = w28727 ^ w28827 ;
  assign w28829 = ~w28765 & w28828 ;
  assign w28830 = w28826 | w28829 ;
  assign w28831 = ~\pi096 & w28830 ;
  assign w28832 = w28439 & w28765 ;
  assign w28833 = ~w28447 & w28723 ;
  assign w28834 = w28724 ^ w28833 ;
  assign w28835 = ~w28765 & w28834 ;
  assign w28836 = w28832 | w28835 ;
  assign w28837 = ~\pi095 & w28836 ;
  assign w28838 = w28446 & w28765 ;
  assign w28839 = ~w28454 & w28720 ;
  assign w28840 = w28721 ^ w28839 ;
  assign w28841 = ~w28765 & w28840 ;
  assign w28842 = w28838 | w28841 ;
  assign w28843 = ~\pi094 & w28842 ;
  assign w28844 = w28453 & w28765 ;
  assign w28845 = ~w28461 & w28717 ;
  assign w28846 = w28718 ^ w28845 ;
  assign w28847 = ~w28765 & w28846 ;
  assign w28848 = w28844 | w28847 ;
  assign w28849 = ~\pi093 & w28848 ;
  assign w28850 = w28460 & w28765 ;
  assign w28851 = ~w28468 & w28714 ;
  assign w28852 = w28715 ^ w28851 ;
  assign w28853 = ~w28765 & w28852 ;
  assign w28854 = w28850 | w28853 ;
  assign w28855 = ~\pi092 & w28854 ;
  assign w28856 = w28467 & w28765 ;
  assign w28857 = ~w28475 & w28711 ;
  assign w28858 = w28712 ^ w28857 ;
  assign w28859 = ~w28765 & w28858 ;
  assign w28860 = w28856 | w28859 ;
  assign w28861 = ~\pi091 & w28860 ;
  assign w28862 = w28474 & w28765 ;
  assign w28863 = ~w28482 & w28708 ;
  assign w28864 = w28709 ^ w28863 ;
  assign w28865 = ~w28765 & w28864 ;
  assign w28866 = w28862 | w28865 ;
  assign w28867 = ~\pi090 & w28866 ;
  assign w28868 = w28481 & w28765 ;
  assign w28869 = ~w28489 & w28705 ;
  assign w28870 = w28706 ^ w28869 ;
  assign w28871 = ~w28765 & w28870 ;
  assign w28872 = w28868 | w28871 ;
  assign w28873 = ~\pi089 & w28872 ;
  assign w28874 = w28488 & w28765 ;
  assign w28875 = ~w28496 & w28702 ;
  assign w28876 = w28703 ^ w28875 ;
  assign w28877 = ~w28765 & w28876 ;
  assign w28878 = w28874 | w28877 ;
  assign w28879 = ~\pi088 & w28878 ;
  assign w28880 = w28495 & w28765 ;
  assign w28881 = ~w28503 & w28699 ;
  assign w28882 = w28700 ^ w28881 ;
  assign w28883 = ~w28765 & w28882 ;
  assign w28884 = w28880 | w28883 ;
  assign w28885 = ~\pi087 & w28884 ;
  assign w28886 = w28502 & w28765 ;
  assign w28887 = ~w28510 & w28696 ;
  assign w28888 = w28697 ^ w28887 ;
  assign w28889 = ~w28765 & w28888 ;
  assign w28890 = w28886 | w28889 ;
  assign w28891 = ~\pi086 & w28890 ;
  assign w28892 = w28509 & w28765 ;
  assign w28893 = ~w28517 & w28693 ;
  assign w28894 = w28694 ^ w28893 ;
  assign w28895 = ~w28765 & w28894 ;
  assign w28896 = w28892 | w28895 ;
  assign w28897 = ~\pi085 & w28896 ;
  assign w28898 = w28516 & w28765 ;
  assign w28899 = ~w28524 & w28690 ;
  assign w28900 = w28691 ^ w28899 ;
  assign w28901 = ~w28765 & w28900 ;
  assign w28902 = w28898 | w28901 ;
  assign w28903 = ~\pi084 & w28902 ;
  assign w28904 = w28523 & w28765 ;
  assign w28905 = ~w28531 & w28687 ;
  assign w28906 = w28688 ^ w28905 ;
  assign w28907 = ~w28765 & w28906 ;
  assign w28908 = w28904 | w28907 ;
  assign w28909 = ~\pi083 & w28908 ;
  assign w28910 = w28530 & w28765 ;
  assign w28911 = ~w28538 & w28684 ;
  assign w28912 = w28685 ^ w28911 ;
  assign w28913 = ~w28765 & w28912 ;
  assign w28914 = w28910 | w28913 ;
  assign w28915 = ~\pi082 & w28914 ;
  assign w28916 = w28537 & w28765 ;
  assign w28917 = ~w28545 & w28681 ;
  assign w28918 = w28682 ^ w28917 ;
  assign w28919 = ~w28765 & w28918 ;
  assign w28920 = w28916 | w28919 ;
  assign w28921 = ~\pi081 & w28920 ;
  assign w28922 = w28544 & w28765 ;
  assign w28923 = ~w28552 & w28678 ;
  assign w28924 = w28679 ^ w28923 ;
  assign w28925 = ~w28765 & w28924 ;
  assign w28926 = w28922 | w28925 ;
  assign w28927 = ~\pi080 & w28926 ;
  assign w28928 = w28551 & w28765 ;
  assign w28929 = ~w28559 & w28675 ;
  assign w28930 = w28676 ^ w28929 ;
  assign w28931 = ~w28765 & w28930 ;
  assign w28932 = w28928 | w28931 ;
  assign w28933 = ~\pi079 & w28932 ;
  assign w28934 = w28558 & w28765 ;
  assign w28935 = ~w28566 & w28672 ;
  assign w28936 = w28673 ^ w28935 ;
  assign w28937 = ~w28765 & w28936 ;
  assign w28938 = w28934 | w28937 ;
  assign w28939 = ~\pi078 & w28938 ;
  assign w28940 = w28565 & w28765 ;
  assign w28941 = ~w28573 & w28669 ;
  assign w28942 = w28670 ^ w28941 ;
  assign w28943 = ~w28765 & w28942 ;
  assign w28944 = w28940 | w28943 ;
  assign w28945 = ~\pi077 & w28944 ;
  assign w28946 = w28572 & w28765 ;
  assign w28947 = ~w28580 & w28666 ;
  assign w28948 = w28667 ^ w28947 ;
  assign w28949 = ~w28765 & w28948 ;
  assign w28950 = w28946 | w28949 ;
  assign w28951 = ~\pi076 & w28950 ;
  assign w28952 = w28579 & w28765 ;
  assign w28953 = ~w28587 & w28663 ;
  assign w28954 = w28664 ^ w28953 ;
  assign w28955 = ~w28765 & w28954 ;
  assign w28956 = w28952 | w28955 ;
  assign w28957 = ~\pi075 & w28956 ;
  assign w28958 = w28586 & w28765 ;
  assign w28959 = ~w28594 & w28660 ;
  assign w28960 = w28661 ^ w28959 ;
  assign w28961 = ~w28765 & w28960 ;
  assign w28962 = w28958 | w28961 ;
  assign w28963 = ~\pi074 & w28962 ;
  assign w28964 = w28593 & w28765 ;
  assign w28965 = ~w28601 & w28657 ;
  assign w28966 = w28658 ^ w28965 ;
  assign w28967 = ~w28765 & w28966 ;
  assign w28968 = w28964 | w28967 ;
  assign w28969 = ~\pi073 & w28968 ;
  assign w28970 = w28600 & w28765 ;
  assign w28971 = ~w28608 & w28654 ;
  assign w28972 = w28655 ^ w28971 ;
  assign w28973 = ~w28765 & w28972 ;
  assign w28974 = w28970 | w28973 ;
  assign w28975 = ~\pi072 & w28974 ;
  assign w28976 = w28607 & w28765 ;
  assign w28977 = ~w28615 & w28651 ;
  assign w28978 = w28652 ^ w28977 ;
  assign w28979 = ~w28765 & w28978 ;
  assign w28980 = w28976 | w28979 ;
  assign w28981 = ~\pi071 & w28980 ;
  assign w28982 = w28614 & w28765 ;
  assign w28983 = ~w28622 & w28648 ;
  assign w28984 = w28649 ^ w28983 ;
  assign w28985 = ~w28765 & w28984 ;
  assign w28986 = w28982 | w28985 ;
  assign w28987 = ~\pi070 & w28986 ;
  assign w28988 = w28621 & w28765 ;
  assign w28989 = ~w28630 & w28645 ;
  assign w28990 = w28646 ^ w28989 ;
  assign w28991 = ~w28765 & w28990 ;
  assign w28992 = w28988 | w28991 ;
  assign w28993 = ~\pi069 & w28992 ;
  assign w28994 = w28629 & w28765 ;
  assign w28995 = ~w28635 & w28642 ;
  assign w28996 = w28643 ^ w28995 ;
  assign w28997 = ~w28765 & w28996 ;
  assign w28998 = w28994 | w28997 ;
  assign w28999 = ~\pi068 & w28998 ;
  assign w29000 = w28634 & w28765 ;
  assign w29001 = \pi064 & ~w28349 ;
  assign w29002 = \pi022 ^ w29001 ;
  assign w29003 = ( \pi065 & w9218 ) | ( \pi065 & ~w29002 ) | ( w9218 & ~w29002 ) ;
  assign w29004 = w28638 ^ w29003 ;
  assign w29005 = ( w9351 & w28764 ) | ( w9351 & w29004 ) | ( w28764 & w29004 ) ;
  assign w29006 = w29004 & ~w29005 ;
  assign w29007 = w29000 | w29006 ;
  assign w29008 = ~\pi067 & w29007 ;
  assign w29009 = \pi021 ^ w28349 ;
  assign w29010 = ( \pi064 & w9351 ) | ( \pi064 & w29009 ) | ( w9351 & w29009 ) ;
  assign w29011 = w9594 ^ w29010 ;
  assign w29012 = ~w9351 & w29011 ;
  assign w29013 = ~w28764 & w29012 ;
  assign w29014 = ( ~\pi064 & w28349 ) | ( ~\pi064 & w28765 ) | ( w28349 & w28765 ) ;
  assign w29015 = \pi022 ^ w29014 ;
  assign w29016 = w28765 & ~w29015 ;
  assign w29017 = w29013 | w29016 ;
  assign w29018 = ~\pi066 & w29017 ;
  assign w29019 = ( \pi064 & w9607 ) | ( \pi064 & w28764 ) | ( w9607 & w28764 ) ;
  assign w29020 = ( \pi021 & ~\pi064 ) | ( \pi021 & w29019 ) | ( ~\pi064 & w29019 ) ;
  assign w29021 = w275 | w28764 ;
  assign w29022 = w9612 | w29021 ;
  assign w29023 = w9610 & ~w29022 ;
  assign w29024 = w28765 | w29013 ;
  assign w29025 = ( w29002 & w29013 ) | ( w29002 & w29024 ) | ( w29013 & w29024 ) ;
  assign w29026 = \pi066 ^ w29025 ;
  assign w29027 = w29020 | w29023 ;
  assign w29028 = ( \pi065 & w9615 ) | ( \pi065 & ~w29027 ) | ( w9615 & ~w29027 ) ;
  assign w29029 = w29026 | w29028 ;
  assign w29030 = \pi067 ^ w29007 ;
  assign w29031 = ( ~w29018 & w29029 ) | ( ~w29018 & w29030 ) | ( w29029 & w29030 ) ;
  assign w29032 = w29030 | w29031 ;
  assign w29033 = \pi068 ^ w28998 ;
  assign w29034 = ( ~w29008 & w29032 ) | ( ~w29008 & w29033 ) | ( w29032 & w29033 ) ;
  assign w29035 = w29033 | w29034 ;
  assign w29036 = \pi069 ^ w28992 ;
  assign w29037 = ( ~w28999 & w29035 ) | ( ~w28999 & w29036 ) | ( w29035 & w29036 ) ;
  assign w29038 = w29036 | w29037 ;
  assign w29039 = \pi070 ^ w28986 ;
  assign w29040 = ( ~w28993 & w29038 ) | ( ~w28993 & w29039 ) | ( w29038 & w29039 ) ;
  assign w29041 = w29039 | w29040 ;
  assign w29042 = \pi071 ^ w28980 ;
  assign w29043 = ( ~w28987 & w29041 ) | ( ~w28987 & w29042 ) | ( w29041 & w29042 ) ;
  assign w29044 = w29042 | w29043 ;
  assign w29045 = \pi072 ^ w28974 ;
  assign w29046 = ( ~w28981 & w29044 ) | ( ~w28981 & w29045 ) | ( w29044 & w29045 ) ;
  assign w29047 = w29045 | w29046 ;
  assign w29048 = \pi073 ^ w28968 ;
  assign w29049 = ( ~w28975 & w29047 ) | ( ~w28975 & w29048 ) | ( w29047 & w29048 ) ;
  assign w29050 = w29048 | w29049 ;
  assign w29051 = \pi074 ^ w28962 ;
  assign w29052 = ( ~w28969 & w29050 ) | ( ~w28969 & w29051 ) | ( w29050 & w29051 ) ;
  assign w29053 = w29051 | w29052 ;
  assign w29054 = \pi075 ^ w28956 ;
  assign w29055 = ( ~w28963 & w29053 ) | ( ~w28963 & w29054 ) | ( w29053 & w29054 ) ;
  assign w29056 = w29054 | w29055 ;
  assign w29057 = \pi076 ^ w28950 ;
  assign w29058 = ( ~w28957 & w29056 ) | ( ~w28957 & w29057 ) | ( w29056 & w29057 ) ;
  assign w29059 = w29057 | w29058 ;
  assign w29060 = \pi077 ^ w28944 ;
  assign w29061 = ( ~w28951 & w29059 ) | ( ~w28951 & w29060 ) | ( w29059 & w29060 ) ;
  assign w29062 = w29060 | w29061 ;
  assign w29063 = \pi078 ^ w28938 ;
  assign w29064 = ( ~w28945 & w29062 ) | ( ~w28945 & w29063 ) | ( w29062 & w29063 ) ;
  assign w29065 = w29063 | w29064 ;
  assign w29066 = \pi079 ^ w28932 ;
  assign w29067 = ( ~w28939 & w29065 ) | ( ~w28939 & w29066 ) | ( w29065 & w29066 ) ;
  assign w29068 = w29066 | w29067 ;
  assign w29069 = \pi080 ^ w28926 ;
  assign w29070 = ( ~w28933 & w29068 ) | ( ~w28933 & w29069 ) | ( w29068 & w29069 ) ;
  assign w29071 = w29069 | w29070 ;
  assign w29072 = \pi081 ^ w28920 ;
  assign w29073 = ( ~w28927 & w29071 ) | ( ~w28927 & w29072 ) | ( w29071 & w29072 ) ;
  assign w29074 = w29072 | w29073 ;
  assign w29075 = \pi082 ^ w28914 ;
  assign w29076 = ( ~w28921 & w29074 ) | ( ~w28921 & w29075 ) | ( w29074 & w29075 ) ;
  assign w29077 = w29075 | w29076 ;
  assign w29078 = \pi083 ^ w28908 ;
  assign w29079 = ( ~w28915 & w29077 ) | ( ~w28915 & w29078 ) | ( w29077 & w29078 ) ;
  assign w29080 = w29078 | w29079 ;
  assign w29081 = \pi084 ^ w28902 ;
  assign w29082 = ( ~w28909 & w29080 ) | ( ~w28909 & w29081 ) | ( w29080 & w29081 ) ;
  assign w29083 = w29081 | w29082 ;
  assign w29084 = \pi085 ^ w28896 ;
  assign w29085 = ( ~w28903 & w29083 ) | ( ~w28903 & w29084 ) | ( w29083 & w29084 ) ;
  assign w29086 = w29084 | w29085 ;
  assign w29087 = \pi086 ^ w28890 ;
  assign w29088 = ( ~w28897 & w29086 ) | ( ~w28897 & w29087 ) | ( w29086 & w29087 ) ;
  assign w29089 = w29087 | w29088 ;
  assign w29090 = \pi087 ^ w28884 ;
  assign w29091 = ( ~w28891 & w29089 ) | ( ~w28891 & w29090 ) | ( w29089 & w29090 ) ;
  assign w29092 = w29090 | w29091 ;
  assign w29093 = \pi088 ^ w28878 ;
  assign w29094 = ( ~w28885 & w29092 ) | ( ~w28885 & w29093 ) | ( w29092 & w29093 ) ;
  assign w29095 = w29093 | w29094 ;
  assign w29096 = \pi089 ^ w28872 ;
  assign w29097 = ( ~w28879 & w29095 ) | ( ~w28879 & w29096 ) | ( w29095 & w29096 ) ;
  assign w29098 = w29096 | w29097 ;
  assign w29099 = \pi090 ^ w28866 ;
  assign w29100 = ( ~w28873 & w29098 ) | ( ~w28873 & w29099 ) | ( w29098 & w29099 ) ;
  assign w29101 = w29099 | w29100 ;
  assign w29102 = \pi091 ^ w28860 ;
  assign w29103 = ( ~w28867 & w29101 ) | ( ~w28867 & w29102 ) | ( w29101 & w29102 ) ;
  assign w29104 = w29102 | w29103 ;
  assign w29105 = \pi092 ^ w28854 ;
  assign w29106 = ( ~w28861 & w29104 ) | ( ~w28861 & w29105 ) | ( w29104 & w29105 ) ;
  assign w29107 = w29105 | w29106 ;
  assign w29108 = \pi093 ^ w28848 ;
  assign w29109 = ( ~w28855 & w29107 ) | ( ~w28855 & w29108 ) | ( w29107 & w29108 ) ;
  assign w29110 = w29108 | w29109 ;
  assign w29111 = \pi094 ^ w28842 ;
  assign w29112 = ( ~w28849 & w29110 ) | ( ~w28849 & w29111 ) | ( w29110 & w29111 ) ;
  assign w29113 = w29111 | w29112 ;
  assign w29114 = \pi095 ^ w28836 ;
  assign w29115 = ( ~w28843 & w29113 ) | ( ~w28843 & w29114 ) | ( w29113 & w29114 ) ;
  assign w29116 = w29114 | w29115 ;
  assign w29117 = \pi096 ^ w28830 ;
  assign w29118 = ( ~w28837 & w29116 ) | ( ~w28837 & w29117 ) | ( w29116 & w29117 ) ;
  assign w29119 = w29117 | w29118 ;
  assign w29120 = \pi097 ^ w28824 ;
  assign w29121 = ( ~w28831 & w29119 ) | ( ~w28831 & w29120 ) | ( w29119 & w29120 ) ;
  assign w29122 = w29120 | w29121 ;
  assign w29123 = \pi098 ^ w28818 ;
  assign w29124 = ( ~w28825 & w29122 ) | ( ~w28825 & w29123 ) | ( w29122 & w29123 ) ;
  assign w29125 = w29123 | w29124 ;
  assign w29126 = \pi099 ^ w28812 ;
  assign w29127 = ( ~w28819 & w29125 ) | ( ~w28819 & w29126 ) | ( w29125 & w29126 ) ;
  assign w29128 = w29126 | w29127 ;
  assign w29129 = \pi100 ^ w28806 ;
  assign w29130 = ( ~w28813 & w29128 ) | ( ~w28813 & w29129 ) | ( w29128 & w29129 ) ;
  assign w29131 = w29129 | w29130 ;
  assign w29132 = \pi101 ^ w28800 ;
  assign w29133 = ( ~w28807 & w29131 ) | ( ~w28807 & w29132 ) | ( w29131 & w29132 ) ;
  assign w29134 = w29132 | w29133 ;
  assign w29135 = \pi102 ^ w28794 ;
  assign w29136 = ( ~w28801 & w29134 ) | ( ~w28801 & w29135 ) | ( w29134 & w29135 ) ;
  assign w29137 = w29135 | w29136 ;
  assign w29138 = \pi103 ^ w28788 ;
  assign w29139 = ( ~w28795 & w29137 ) | ( ~w28795 & w29138 ) | ( w29137 & w29138 ) ;
  assign w29140 = w29138 | w29139 ;
  assign w29141 = \pi104 ^ w28782 ;
  assign w29142 = ( ~w28789 & w29140 ) | ( ~w28789 & w29141 ) | ( w29140 & w29141 ) ;
  assign w29143 = w29141 | w29142 ;
  assign w29144 = \pi105 ^ w28776 ;
  assign w29145 = ( ~w28783 & w29143 ) | ( ~w28783 & w29144 ) | ( w29143 & w29144 ) ;
  assign w29146 = w29144 | w29145 ;
  assign w29147 = \pi106 ^ w28770 ;
  assign w29148 = ( ~w28777 & w29146 ) | ( ~w28777 & w29147 ) | ( w29146 & w29147 ) ;
  assign w29149 = w29147 | w29148 ;
  assign w29150 = w28362 & w28765 ;
  assign w29151 = ~w28363 & w28759 ;
  assign w29152 = w28760 ^ w29151 ;
  assign w29153 = ~w28765 & w29152 ;
  assign w29154 = w29150 | w29153 ;
  assign w29155 = ~\pi107 & w29154 ;
  assign w29156 = ( \pi107 & ~w29150 ) | ( \pi107 & w29153 ) | ( ~w29150 & w29153 ) ;
  assign w29157 = ~w29153 & w29156 ;
  assign w29158 = ( ~w28771 & w29149 ) | ( ~w28771 & w29155 ) | ( w29149 & w29155 ) ;
  assign w29159 = ( w168 & w29155 ) | ( w168 & ~w29158 ) | ( w29155 & ~w29158 ) ;
  assign w29160 = ( w155 & w29157 ) | ( w155 & ~w29158 ) | ( w29157 & ~w29158 ) ;
  assign w29161 = ( w29158 & ~w29159 ) | ( w29158 & w29160 ) | ( ~w29159 & w29160 ) ;
  assign w29162 = w29159 | w29161 ;
  assign w29163 = ~w9351 & w29154 ;
  assign w29164 = w29162 & ~w29163 ;
  assign w29165 = ~w28777 & w29146 ;
  assign w29166 = w29147 ^ w29165 ;
  assign w29167 = ~w29164 & w29166 ;
  assign w29168 = ( w28770 & w29162 ) | ( w28770 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29169 = ~w29163 & w29168 ;
  assign w29170 = w29167 | w29169 ;
  assign w29171 = ~\pi107 & w29170 ;
  assign w29172 = ~w28783 & w29143 ;
  assign w29173 = w29144 ^ w29172 ;
  assign w29174 = ~w29164 & w29173 ;
  assign w29175 = ( w28776 & w29162 ) | ( w28776 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29176 = ~w29163 & w29175 ;
  assign w29177 = w29174 | w29176 ;
  assign w29178 = ~\pi106 & w29177 ;
  assign w29179 = ~w28789 & w29140 ;
  assign w29180 = w29141 ^ w29179 ;
  assign w29181 = ~w29164 & w29180 ;
  assign w29182 = ( w28782 & w29162 ) | ( w28782 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29183 = ~w29163 & w29182 ;
  assign w29184 = w29181 | w29183 ;
  assign w29185 = ~\pi105 & w29184 ;
  assign w29186 = ~w28795 & w29137 ;
  assign w29187 = w29138 ^ w29186 ;
  assign w29188 = ~w29164 & w29187 ;
  assign w29189 = ( w28788 & w29162 ) | ( w28788 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29190 = ~w29163 & w29189 ;
  assign w29191 = w29188 | w29190 ;
  assign w29192 = ~\pi104 & w29191 ;
  assign w29193 = ~w28801 & w29134 ;
  assign w29194 = w29135 ^ w29193 ;
  assign w29195 = ~w29164 & w29194 ;
  assign w29196 = ( w28794 & w29162 ) | ( w28794 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29197 = ~w29163 & w29196 ;
  assign w29198 = w29195 | w29197 ;
  assign w29199 = ~\pi103 & w29198 ;
  assign w29200 = ~w28807 & w29131 ;
  assign w29201 = w29132 ^ w29200 ;
  assign w29202 = ~w29164 & w29201 ;
  assign w29203 = ( w28800 & w29162 ) | ( w28800 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29204 = ~w29163 & w29203 ;
  assign w29205 = w29202 | w29204 ;
  assign w29206 = ~\pi102 & w29205 ;
  assign w29207 = ~w28813 & w29128 ;
  assign w29208 = w29129 ^ w29207 ;
  assign w29209 = ~w29164 & w29208 ;
  assign w29210 = ( w28806 & w29162 ) | ( w28806 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29211 = ~w29163 & w29210 ;
  assign w29212 = w29209 | w29211 ;
  assign w29213 = ~\pi101 & w29212 ;
  assign w29214 = ~w28819 & w29125 ;
  assign w29215 = w29126 ^ w29214 ;
  assign w29216 = ~w29164 & w29215 ;
  assign w29217 = ( w28812 & w29162 ) | ( w28812 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29218 = ~w29163 & w29217 ;
  assign w29219 = w29216 | w29218 ;
  assign w29220 = ~\pi100 & w29219 ;
  assign w29221 = ~w28825 & w29122 ;
  assign w29222 = w29123 ^ w29221 ;
  assign w29223 = ~w29164 & w29222 ;
  assign w29224 = ( w28818 & w29162 ) | ( w28818 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29225 = ~w29163 & w29224 ;
  assign w29226 = w29223 | w29225 ;
  assign w29227 = ~\pi099 & w29226 ;
  assign w29228 = ~w28831 & w29119 ;
  assign w29229 = w29120 ^ w29228 ;
  assign w29230 = ~w29164 & w29229 ;
  assign w29231 = ( w28824 & w29162 ) | ( w28824 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29232 = ~w29163 & w29231 ;
  assign w29233 = w29230 | w29232 ;
  assign w29234 = ~\pi098 & w29233 ;
  assign w29235 = ~w28837 & w29116 ;
  assign w29236 = w29117 ^ w29235 ;
  assign w29237 = ~w29164 & w29236 ;
  assign w29238 = ( w28830 & w29162 ) | ( w28830 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29239 = ~w29163 & w29238 ;
  assign w29240 = w29237 | w29239 ;
  assign w29241 = ~\pi097 & w29240 ;
  assign w29242 = ~w28843 & w29113 ;
  assign w29243 = w29114 ^ w29242 ;
  assign w29244 = ~w29164 & w29243 ;
  assign w29245 = ( w28836 & w29162 ) | ( w28836 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29246 = ~w29163 & w29245 ;
  assign w29247 = w29244 | w29246 ;
  assign w29248 = ~\pi096 & w29247 ;
  assign w29249 = ~w28849 & w29110 ;
  assign w29250 = w29111 ^ w29249 ;
  assign w29251 = ~w29164 & w29250 ;
  assign w29252 = ( w28842 & w29162 ) | ( w28842 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29253 = ~w29163 & w29252 ;
  assign w29254 = w29251 | w29253 ;
  assign w29255 = ~\pi095 & w29254 ;
  assign w29256 = ~w28855 & w29107 ;
  assign w29257 = w29108 ^ w29256 ;
  assign w29258 = ~w29164 & w29257 ;
  assign w29259 = ( w28848 & w29162 ) | ( w28848 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29260 = ~w29163 & w29259 ;
  assign w29261 = w29258 | w29260 ;
  assign w29262 = ~\pi094 & w29261 ;
  assign w29263 = ~w28861 & w29104 ;
  assign w29264 = w29105 ^ w29263 ;
  assign w29265 = ~w29164 & w29264 ;
  assign w29266 = ( w28854 & w29162 ) | ( w28854 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29267 = ~w29163 & w29266 ;
  assign w29268 = w29265 | w29267 ;
  assign w29269 = ~\pi093 & w29268 ;
  assign w29270 = ~w28867 & w29101 ;
  assign w29271 = w29102 ^ w29270 ;
  assign w29272 = ~w29164 & w29271 ;
  assign w29273 = ( w28860 & w29162 ) | ( w28860 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29274 = ~w29163 & w29273 ;
  assign w29275 = w29272 | w29274 ;
  assign w29276 = ~\pi092 & w29275 ;
  assign w29277 = ~w28873 & w29098 ;
  assign w29278 = w29099 ^ w29277 ;
  assign w29279 = ~w29164 & w29278 ;
  assign w29280 = ( w28866 & w29162 ) | ( w28866 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29281 = ~w29163 & w29280 ;
  assign w29282 = w29279 | w29281 ;
  assign w29283 = ~\pi091 & w29282 ;
  assign w29284 = ~w28879 & w29095 ;
  assign w29285 = w29096 ^ w29284 ;
  assign w29286 = ~w29164 & w29285 ;
  assign w29287 = ( w28872 & w29162 ) | ( w28872 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29288 = ~w29163 & w29287 ;
  assign w29289 = w29286 | w29288 ;
  assign w29290 = ~\pi090 & w29289 ;
  assign w29291 = ~w28885 & w29092 ;
  assign w29292 = w29093 ^ w29291 ;
  assign w29293 = ~w29164 & w29292 ;
  assign w29294 = ( w28878 & w29162 ) | ( w28878 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29295 = ~w29163 & w29294 ;
  assign w29296 = w29293 | w29295 ;
  assign w29297 = ~\pi089 & w29296 ;
  assign w29298 = ~w28891 & w29089 ;
  assign w29299 = w29090 ^ w29298 ;
  assign w29300 = ~w29164 & w29299 ;
  assign w29301 = ( w28884 & w29162 ) | ( w28884 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29302 = ~w29163 & w29301 ;
  assign w29303 = w29300 | w29302 ;
  assign w29304 = ~\pi088 & w29303 ;
  assign w29305 = ~w28897 & w29086 ;
  assign w29306 = w29087 ^ w29305 ;
  assign w29307 = ~w29164 & w29306 ;
  assign w29308 = ( w28890 & w29162 ) | ( w28890 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29309 = ~w29163 & w29308 ;
  assign w29310 = w29307 | w29309 ;
  assign w29311 = ~\pi087 & w29310 ;
  assign w29312 = ~w28903 & w29083 ;
  assign w29313 = w29084 ^ w29312 ;
  assign w29314 = ~w29164 & w29313 ;
  assign w29315 = ( w28896 & w29162 ) | ( w28896 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29316 = ~w29163 & w29315 ;
  assign w29317 = w29314 | w29316 ;
  assign w29318 = ~\pi086 & w29317 ;
  assign w29319 = ~w28909 & w29080 ;
  assign w29320 = w29081 ^ w29319 ;
  assign w29321 = ~w29164 & w29320 ;
  assign w29322 = ( w28902 & w29162 ) | ( w28902 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29323 = ~w29163 & w29322 ;
  assign w29324 = w29321 | w29323 ;
  assign w29325 = ~\pi085 & w29324 ;
  assign w29326 = ~w28915 & w29077 ;
  assign w29327 = w29078 ^ w29326 ;
  assign w29328 = ~w29164 & w29327 ;
  assign w29329 = ( w28908 & w29162 ) | ( w28908 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29330 = ~w29163 & w29329 ;
  assign w29331 = w29328 | w29330 ;
  assign w29332 = ~\pi084 & w29331 ;
  assign w29333 = ~w28921 & w29074 ;
  assign w29334 = w29075 ^ w29333 ;
  assign w29335 = ~w29164 & w29334 ;
  assign w29336 = ( w28914 & w29162 ) | ( w28914 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29337 = ~w29163 & w29336 ;
  assign w29338 = w29335 | w29337 ;
  assign w29339 = ~\pi083 & w29338 ;
  assign w29340 = ~w28927 & w29071 ;
  assign w29341 = w29072 ^ w29340 ;
  assign w29342 = ~w29164 & w29341 ;
  assign w29343 = ( w28920 & w29162 ) | ( w28920 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29344 = ~w29163 & w29343 ;
  assign w29345 = w29342 | w29344 ;
  assign w29346 = ~\pi082 & w29345 ;
  assign w29347 = ~w28933 & w29068 ;
  assign w29348 = w29069 ^ w29347 ;
  assign w29349 = ~w29164 & w29348 ;
  assign w29350 = ( w28926 & w29162 ) | ( w28926 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29351 = ~w29163 & w29350 ;
  assign w29352 = w29349 | w29351 ;
  assign w29353 = ~\pi081 & w29352 ;
  assign w29354 = ~w28939 & w29065 ;
  assign w29355 = w29066 ^ w29354 ;
  assign w29356 = ~w29164 & w29355 ;
  assign w29357 = ( w28932 & w29162 ) | ( w28932 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29358 = ~w29163 & w29357 ;
  assign w29359 = w29356 | w29358 ;
  assign w29360 = ~\pi080 & w29359 ;
  assign w29361 = ~w28945 & w29062 ;
  assign w29362 = w29063 ^ w29361 ;
  assign w29363 = ~w29164 & w29362 ;
  assign w29364 = ( w28938 & w29162 ) | ( w28938 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29365 = ~w29163 & w29364 ;
  assign w29366 = w29363 | w29365 ;
  assign w29367 = ~\pi079 & w29366 ;
  assign w29368 = ~w28951 & w29059 ;
  assign w29369 = w29060 ^ w29368 ;
  assign w29370 = ~w29164 & w29369 ;
  assign w29371 = ( w28944 & w29162 ) | ( w28944 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29372 = ~w29163 & w29371 ;
  assign w29373 = w29370 | w29372 ;
  assign w29374 = ~\pi078 & w29373 ;
  assign w29375 = ~w28957 & w29056 ;
  assign w29376 = w29057 ^ w29375 ;
  assign w29377 = ~w29164 & w29376 ;
  assign w29378 = ( w28950 & w29162 ) | ( w28950 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29379 = ~w29163 & w29378 ;
  assign w29380 = w29377 | w29379 ;
  assign w29381 = ~\pi077 & w29380 ;
  assign w29382 = ~w28963 & w29053 ;
  assign w29383 = w29054 ^ w29382 ;
  assign w29384 = ~w29164 & w29383 ;
  assign w29385 = ( w28956 & w29162 ) | ( w28956 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29386 = ~w29163 & w29385 ;
  assign w29387 = w29384 | w29386 ;
  assign w29388 = ~\pi076 & w29387 ;
  assign w29389 = ~w28969 & w29050 ;
  assign w29390 = w29051 ^ w29389 ;
  assign w29391 = ~w29164 & w29390 ;
  assign w29392 = ( w28962 & w29162 ) | ( w28962 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29393 = ~w29163 & w29392 ;
  assign w29394 = w29391 | w29393 ;
  assign w29395 = ~\pi075 & w29394 ;
  assign w29396 = ~w28975 & w29047 ;
  assign w29397 = w29048 ^ w29396 ;
  assign w29398 = ~w29164 & w29397 ;
  assign w29399 = ( w28968 & w29162 ) | ( w28968 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29400 = ~w29163 & w29399 ;
  assign w29401 = w29398 | w29400 ;
  assign w29402 = ~\pi074 & w29401 ;
  assign w29403 = ~w28981 & w29044 ;
  assign w29404 = w29045 ^ w29403 ;
  assign w29405 = ~w29164 & w29404 ;
  assign w29406 = ( w28974 & w29162 ) | ( w28974 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29407 = ~w29163 & w29406 ;
  assign w29408 = w29405 | w29407 ;
  assign w29409 = ~\pi073 & w29408 ;
  assign w29410 = ~w28987 & w29041 ;
  assign w29411 = w29042 ^ w29410 ;
  assign w29412 = ~w29164 & w29411 ;
  assign w29413 = ( w28980 & w29162 ) | ( w28980 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29414 = ~w29163 & w29413 ;
  assign w29415 = w29412 | w29414 ;
  assign w29416 = ~\pi072 & w29415 ;
  assign w29417 = ~w28993 & w29038 ;
  assign w29418 = w29039 ^ w29417 ;
  assign w29419 = ~w29164 & w29418 ;
  assign w29420 = ( w28986 & w29162 ) | ( w28986 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29421 = ~w29163 & w29420 ;
  assign w29422 = w29419 | w29421 ;
  assign w29423 = ~\pi071 & w29422 ;
  assign w29424 = ~w28999 & w29035 ;
  assign w29425 = w29036 ^ w29424 ;
  assign w29426 = ~w29164 & w29425 ;
  assign w29427 = ( w28992 & w29162 ) | ( w28992 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29428 = ~w29163 & w29427 ;
  assign w29429 = w29426 | w29428 ;
  assign w29430 = ~\pi070 & w29429 ;
  assign w29431 = ~w29008 & w29032 ;
  assign w29432 = w29033 ^ w29431 ;
  assign w29433 = ~w29164 & w29432 ;
  assign w29434 = ( w28998 & w29162 ) | ( w28998 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29435 = ~w29163 & w29434 ;
  assign w29436 = w29433 | w29435 ;
  assign w29437 = ~\pi069 & w29436 ;
  assign w29438 = ~w29018 & w29029 ;
  assign w29439 = w29030 ^ w29438 ;
  assign w29440 = ~w29164 & w29439 ;
  assign w29441 = ( w29007 & w29162 ) | ( w29007 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29442 = ~w29163 & w29441 ;
  assign w29443 = w29440 | w29442 ;
  assign w29444 = ~\pi068 & w29443 ;
  assign w29445 = w29026 ^ w29028 ;
  assign w29446 = ~w29164 & w29445 ;
  assign w29447 = ( w29017 & w29162 ) | ( w29017 & w29163 ) | ( w29162 & w29163 ) ;
  assign w29448 = ~w29163 & w29447 ;
  assign w29449 = w29446 | w29448 ;
  assign w29450 = ~\pi067 & w29449 ;
  assign w29451 = w9615 ^ w29027 ;
  assign w29452 = \pi065 ^ w29451 ;
  assign w29453 = w29164 ^ w29452 ;
  assign w29454 = ( w29027 & w29452 ) | ( w29027 & w29453 ) | ( w29452 & w29453 ) ;
  assign w29455 = ~\pi066 & w29454 ;
  assign w29456 = w29027 ^ w29164 ;
  assign w29457 = ( w29027 & w29452 ) | ( w29027 & ~w29456 ) | ( w29452 & ~w29456 ) ;
  assign w29458 = \pi066 ^ w29457 ;
  assign w29459 = ( \pi064 & ~w29164 ) | ( \pi064 & w29458 ) | ( ~w29164 & w29458 ) ;
  assign w29460 = \pi020 ^ w29459 ;
  assign w29461 = ( \pi065 & w10495 ) | ( \pi065 & ~w29460 ) | ( w10495 & ~w29460 ) ;
  assign w29462 = w29458 | w29461 ;
  assign w29463 = \pi067 ^ w29449 ;
  assign w29464 = ( ~w29455 & w29462 ) | ( ~w29455 & w29463 ) | ( w29462 & w29463 ) ;
  assign w29465 = w29463 | w29464 ;
  assign w29466 = \pi068 ^ w29443 ;
  assign w29467 = ( ~w29450 & w29465 ) | ( ~w29450 & w29466 ) | ( w29465 & w29466 ) ;
  assign w29468 = w29466 | w29467 ;
  assign w29469 = \pi069 ^ w29436 ;
  assign w29470 = ( ~w29444 & w29468 ) | ( ~w29444 & w29469 ) | ( w29468 & w29469 ) ;
  assign w29471 = w29469 | w29470 ;
  assign w29472 = \pi070 ^ w29429 ;
  assign w29473 = ( ~w29437 & w29471 ) | ( ~w29437 & w29472 ) | ( w29471 & w29472 ) ;
  assign w29474 = w29472 | w29473 ;
  assign w29475 = \pi071 ^ w29422 ;
  assign w29476 = ( ~w29430 & w29474 ) | ( ~w29430 & w29475 ) | ( w29474 & w29475 ) ;
  assign w29477 = w29475 | w29476 ;
  assign w29478 = \pi072 ^ w29415 ;
  assign w29479 = ( ~w29423 & w29477 ) | ( ~w29423 & w29478 ) | ( w29477 & w29478 ) ;
  assign w29480 = w29478 | w29479 ;
  assign w29481 = \pi073 ^ w29408 ;
  assign w29482 = ( ~w29416 & w29480 ) | ( ~w29416 & w29481 ) | ( w29480 & w29481 ) ;
  assign w29483 = w29481 | w29482 ;
  assign w29484 = \pi074 ^ w29401 ;
  assign w29485 = ( ~w29409 & w29483 ) | ( ~w29409 & w29484 ) | ( w29483 & w29484 ) ;
  assign w29486 = w29484 | w29485 ;
  assign w29487 = \pi075 ^ w29394 ;
  assign w29488 = ( ~w29402 & w29486 ) | ( ~w29402 & w29487 ) | ( w29486 & w29487 ) ;
  assign w29489 = w29487 | w29488 ;
  assign w29490 = \pi076 ^ w29387 ;
  assign w29491 = ( ~w29395 & w29489 ) | ( ~w29395 & w29490 ) | ( w29489 & w29490 ) ;
  assign w29492 = w29490 | w29491 ;
  assign w29493 = \pi077 ^ w29380 ;
  assign w29494 = ( ~w29388 & w29492 ) | ( ~w29388 & w29493 ) | ( w29492 & w29493 ) ;
  assign w29495 = w29493 | w29494 ;
  assign w29496 = \pi078 ^ w29373 ;
  assign w29497 = ( ~w29381 & w29495 ) | ( ~w29381 & w29496 ) | ( w29495 & w29496 ) ;
  assign w29498 = w29496 | w29497 ;
  assign w29499 = \pi079 ^ w29366 ;
  assign w29500 = ( ~w29374 & w29498 ) | ( ~w29374 & w29499 ) | ( w29498 & w29499 ) ;
  assign w29501 = w29499 | w29500 ;
  assign w29502 = \pi080 ^ w29359 ;
  assign w29503 = ( ~w29367 & w29501 ) | ( ~w29367 & w29502 ) | ( w29501 & w29502 ) ;
  assign w29504 = w29502 | w29503 ;
  assign w29505 = \pi081 ^ w29352 ;
  assign w29506 = ( ~w29360 & w29504 ) | ( ~w29360 & w29505 ) | ( w29504 & w29505 ) ;
  assign w29507 = w29505 | w29506 ;
  assign w29508 = \pi082 ^ w29345 ;
  assign w29509 = ( ~w29353 & w29507 ) | ( ~w29353 & w29508 ) | ( w29507 & w29508 ) ;
  assign w29510 = w29508 | w29509 ;
  assign w29511 = \pi083 ^ w29338 ;
  assign w29512 = ( ~w29346 & w29510 ) | ( ~w29346 & w29511 ) | ( w29510 & w29511 ) ;
  assign w29513 = w29511 | w29512 ;
  assign w29514 = \pi084 ^ w29331 ;
  assign w29515 = ( ~w29339 & w29513 ) | ( ~w29339 & w29514 ) | ( w29513 & w29514 ) ;
  assign w29516 = w29514 | w29515 ;
  assign w29517 = \pi085 ^ w29324 ;
  assign w29518 = ( ~w29332 & w29516 ) | ( ~w29332 & w29517 ) | ( w29516 & w29517 ) ;
  assign w29519 = w29517 | w29518 ;
  assign w29520 = \pi086 ^ w29317 ;
  assign w29521 = ( ~w29325 & w29519 ) | ( ~w29325 & w29520 ) | ( w29519 & w29520 ) ;
  assign w29522 = w29520 | w29521 ;
  assign w29523 = \pi087 ^ w29310 ;
  assign w29524 = ( ~w29318 & w29522 ) | ( ~w29318 & w29523 ) | ( w29522 & w29523 ) ;
  assign w29525 = w29523 | w29524 ;
  assign w29526 = \pi088 ^ w29303 ;
  assign w29527 = ( ~w29311 & w29525 ) | ( ~w29311 & w29526 ) | ( w29525 & w29526 ) ;
  assign w29528 = w29526 | w29527 ;
  assign w29529 = \pi089 ^ w29296 ;
  assign w29530 = ( ~w29304 & w29528 ) | ( ~w29304 & w29529 ) | ( w29528 & w29529 ) ;
  assign w29531 = w29529 | w29530 ;
  assign w29532 = \pi090 ^ w29289 ;
  assign w29533 = ( ~w29297 & w29531 ) | ( ~w29297 & w29532 ) | ( w29531 & w29532 ) ;
  assign w29534 = w29532 | w29533 ;
  assign w29535 = \pi091 ^ w29282 ;
  assign w29536 = ( ~w29290 & w29534 ) | ( ~w29290 & w29535 ) | ( w29534 & w29535 ) ;
  assign w29537 = w29535 | w29536 ;
  assign w29538 = \pi092 ^ w29275 ;
  assign w29539 = ( ~w29283 & w29537 ) | ( ~w29283 & w29538 ) | ( w29537 & w29538 ) ;
  assign w29540 = w29538 | w29539 ;
  assign w29541 = \pi093 ^ w29268 ;
  assign w29542 = ( ~w29276 & w29540 ) | ( ~w29276 & w29541 ) | ( w29540 & w29541 ) ;
  assign w29543 = w29541 | w29542 ;
  assign w29544 = \pi094 ^ w29261 ;
  assign w29545 = ( ~w29269 & w29543 ) | ( ~w29269 & w29544 ) | ( w29543 & w29544 ) ;
  assign w29546 = w29544 | w29545 ;
  assign w29547 = \pi095 ^ w29254 ;
  assign w29548 = ( ~w29262 & w29546 ) | ( ~w29262 & w29547 ) | ( w29546 & w29547 ) ;
  assign w29549 = w29547 | w29548 ;
  assign w29550 = \pi096 ^ w29247 ;
  assign w29551 = ( ~w29255 & w29549 ) | ( ~w29255 & w29550 ) | ( w29549 & w29550 ) ;
  assign w29552 = w29550 | w29551 ;
  assign w29553 = \pi097 ^ w29240 ;
  assign w29554 = ( ~w29248 & w29552 ) | ( ~w29248 & w29553 ) | ( w29552 & w29553 ) ;
  assign w29555 = w29553 | w29554 ;
  assign w29556 = \pi098 ^ w29233 ;
  assign w29557 = ( ~w29241 & w29555 ) | ( ~w29241 & w29556 ) | ( w29555 & w29556 ) ;
  assign w29558 = w29556 | w29557 ;
  assign w29559 = \pi099 ^ w29226 ;
  assign w29560 = ( ~w29234 & w29558 ) | ( ~w29234 & w29559 ) | ( w29558 & w29559 ) ;
  assign w29561 = w29559 | w29560 ;
  assign w29562 = \pi100 ^ w29219 ;
  assign w29563 = ( ~w29227 & w29561 ) | ( ~w29227 & w29562 ) | ( w29561 & w29562 ) ;
  assign w29564 = w29562 | w29563 ;
  assign w29565 = \pi101 ^ w29212 ;
  assign w29566 = ( ~w29220 & w29564 ) | ( ~w29220 & w29565 ) | ( w29564 & w29565 ) ;
  assign w29567 = w29565 | w29566 ;
  assign w29568 = \pi102 ^ w29205 ;
  assign w29569 = ( ~w29213 & w29567 ) | ( ~w29213 & w29568 ) | ( w29567 & w29568 ) ;
  assign w29570 = w29568 | w29569 ;
  assign w29571 = \pi103 ^ w29198 ;
  assign w29572 = ( ~w29206 & w29570 ) | ( ~w29206 & w29571 ) | ( w29570 & w29571 ) ;
  assign w29573 = w29571 | w29572 ;
  assign w29574 = \pi104 ^ w29191 ;
  assign w29575 = ( ~w29199 & w29573 ) | ( ~w29199 & w29574 ) | ( w29573 & w29574 ) ;
  assign w29576 = w29574 | w29575 ;
  assign w29577 = \pi105 ^ w29184 ;
  assign w29578 = ( ~w29192 & w29576 ) | ( ~w29192 & w29577 ) | ( w29576 & w29577 ) ;
  assign w29579 = w29577 | w29578 ;
  assign w29580 = \pi106 ^ w29177 ;
  assign w29581 = ( ~w29185 & w29579 ) | ( ~w29185 & w29580 ) | ( w29579 & w29580 ) ;
  assign w29582 = w29580 | w29581 ;
  assign w29583 = \pi107 ^ w29170 ;
  assign w29584 = ( ~w29178 & w29582 ) | ( ~w29178 & w29583 ) | ( w29582 & w29583 ) ;
  assign w29585 = w29583 | w29584 ;
  assign w29586 = w29155 | w29157 ;
  assign w29587 = ( ~w28771 & w29149 ) | ( ~w28771 & w29164 ) | ( w29149 & w29164 ) ;
  assign w29588 = w29586 ^ w29587 ;
  assign w29589 = ~w29164 & w29588 ;
  assign w29590 = ( w9351 & ~w29154 ) | ( w9351 & w29162 ) | ( ~w29154 & w29162 ) ;
  assign w29591 = w29154 & w29590 ;
  assign w29592 = w29589 | w29591 ;
  assign w29593 = ~\pi108 & w29592 ;
  assign w29594 = ( \pi108 & ~w29589 ) | ( \pi108 & w29591 ) | ( ~w29589 & w29591 ) ;
  assign w29595 = ~w29591 & w29594 ;
  assign w29596 = ( ~w29171 & w29585 ) | ( ~w29171 & w29593 ) | ( w29585 & w29593 ) ;
  assign w29597 = ( w449 & w29593 ) | ( w449 & ~w29596 ) | ( w29593 & ~w29596 ) ;
  assign w29598 = ( w448 & w29595 ) | ( w448 & ~w29596 ) | ( w29595 & ~w29596 ) ;
  assign w29599 = ( w29596 & ~w29597 ) | ( w29596 & w29598 ) | ( ~w29597 & w29598 ) ;
  assign w29600 = w29597 | w29599 ;
  assign w29601 = ( w155 & ~w168 ) | ( w155 & w29592 ) | ( ~w168 & w29592 ) ;
  assign w29602 = ~w155 & w29601 ;
  assign w29603 = w29600 & ~w29602 ;
  assign w29604 = ~w29178 & w29582 ;
  assign w29605 = w29583 ^ w29604 ;
  assign w29606 = ~w29603 & w29605 ;
  assign w29607 = ( w29170 & w29600 ) | ( w29170 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29608 = ~w29602 & w29607 ;
  assign w29609 = w29606 | w29608 ;
  assign w29610 = w29593 | w29595 ;
  assign w29611 = ( ~w29171 & w29585 ) | ( ~w29171 & w29603 ) | ( w29585 & w29603 ) ;
  assign w29612 = w29610 ^ w29611 ;
  assign w29613 = ~w29603 & w29612 ;
  assign w29614 = ( w29592 & w29600 ) | ( w29592 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29615 = ~w29602 & w29614 ;
  assign w29616 = w29613 | w29615 ;
  assign w29617 = ~\pi108 & w29609 ;
  assign w29618 = ~w29185 & w29579 ;
  assign w29619 = w29580 ^ w29618 ;
  assign w29620 = ~w29603 & w29619 ;
  assign w29621 = ( w29177 & w29600 ) | ( w29177 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29622 = ~w29602 & w29621 ;
  assign w29623 = w29620 | w29622 ;
  assign w29624 = ~\pi107 & w29623 ;
  assign w29625 = ~w29192 & w29576 ;
  assign w29626 = w29577 ^ w29625 ;
  assign w29627 = ~w29603 & w29626 ;
  assign w29628 = ( w29184 & w29600 ) | ( w29184 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29629 = ~w29602 & w29628 ;
  assign w29630 = w29627 | w29629 ;
  assign w29631 = ~\pi106 & w29630 ;
  assign w29632 = ~w29199 & w29573 ;
  assign w29633 = w29574 ^ w29632 ;
  assign w29634 = ~w29603 & w29633 ;
  assign w29635 = ( w29191 & w29600 ) | ( w29191 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29636 = ~w29602 & w29635 ;
  assign w29637 = w29634 | w29636 ;
  assign w29638 = ~\pi105 & w29637 ;
  assign w29639 = ~w29206 & w29570 ;
  assign w29640 = w29571 ^ w29639 ;
  assign w29641 = ~w29603 & w29640 ;
  assign w29642 = ( w29198 & w29600 ) | ( w29198 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29643 = ~w29602 & w29642 ;
  assign w29644 = w29641 | w29643 ;
  assign w29645 = ~\pi104 & w29644 ;
  assign w29646 = ~w29213 & w29567 ;
  assign w29647 = w29568 ^ w29646 ;
  assign w29648 = ~w29603 & w29647 ;
  assign w29649 = ( w29205 & w29600 ) | ( w29205 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29650 = ~w29602 & w29649 ;
  assign w29651 = w29648 | w29650 ;
  assign w29652 = ~\pi103 & w29651 ;
  assign w29653 = ~w29220 & w29564 ;
  assign w29654 = w29565 ^ w29653 ;
  assign w29655 = ~w29603 & w29654 ;
  assign w29656 = ( w29212 & w29600 ) | ( w29212 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29657 = ~w29602 & w29656 ;
  assign w29658 = w29655 | w29657 ;
  assign w29659 = ~\pi102 & w29658 ;
  assign w29660 = ~w29227 & w29561 ;
  assign w29661 = w29562 ^ w29660 ;
  assign w29662 = ~w29603 & w29661 ;
  assign w29663 = ( w29219 & w29600 ) | ( w29219 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29664 = ~w29602 & w29663 ;
  assign w29665 = w29662 | w29664 ;
  assign w29666 = ~\pi101 & w29665 ;
  assign w29667 = ~w29234 & w29558 ;
  assign w29668 = w29559 ^ w29667 ;
  assign w29669 = ~w29603 & w29668 ;
  assign w29670 = ( w29226 & w29600 ) | ( w29226 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29671 = ~w29602 & w29670 ;
  assign w29672 = w29669 | w29671 ;
  assign w29673 = ~\pi100 & w29672 ;
  assign w29674 = ~w29241 & w29555 ;
  assign w29675 = w29556 ^ w29674 ;
  assign w29676 = ~w29603 & w29675 ;
  assign w29677 = ( w29233 & w29600 ) | ( w29233 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29678 = ~w29602 & w29677 ;
  assign w29679 = w29676 | w29678 ;
  assign w29680 = ~\pi099 & w29679 ;
  assign w29681 = ~w29248 & w29552 ;
  assign w29682 = w29553 ^ w29681 ;
  assign w29683 = ~w29603 & w29682 ;
  assign w29684 = ( w29240 & w29600 ) | ( w29240 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29685 = ~w29602 & w29684 ;
  assign w29686 = w29683 | w29685 ;
  assign w29687 = ~\pi098 & w29686 ;
  assign w29688 = ~w29255 & w29549 ;
  assign w29689 = w29550 ^ w29688 ;
  assign w29690 = ~w29603 & w29689 ;
  assign w29691 = ( w29247 & w29600 ) | ( w29247 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29692 = ~w29602 & w29691 ;
  assign w29693 = w29690 | w29692 ;
  assign w29694 = ~\pi097 & w29693 ;
  assign w29695 = ~w29262 & w29546 ;
  assign w29696 = w29547 ^ w29695 ;
  assign w29697 = ~w29603 & w29696 ;
  assign w29698 = ( w29254 & w29600 ) | ( w29254 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29699 = ~w29602 & w29698 ;
  assign w29700 = w29697 | w29699 ;
  assign w29701 = ~\pi096 & w29700 ;
  assign w29702 = ~w29269 & w29543 ;
  assign w29703 = w29544 ^ w29702 ;
  assign w29704 = ~w29603 & w29703 ;
  assign w29705 = ( w29261 & w29600 ) | ( w29261 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29706 = ~w29602 & w29705 ;
  assign w29707 = w29704 | w29706 ;
  assign w29708 = ~\pi095 & w29707 ;
  assign w29709 = ~w29276 & w29540 ;
  assign w29710 = w29541 ^ w29709 ;
  assign w29711 = ~w29603 & w29710 ;
  assign w29712 = ( w29268 & w29600 ) | ( w29268 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29713 = ~w29602 & w29712 ;
  assign w29714 = w29711 | w29713 ;
  assign w29715 = ~\pi094 & w29714 ;
  assign w29716 = ~w29283 & w29537 ;
  assign w29717 = w29538 ^ w29716 ;
  assign w29718 = ~w29603 & w29717 ;
  assign w29719 = ( w29275 & w29600 ) | ( w29275 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29720 = ~w29602 & w29719 ;
  assign w29721 = w29718 | w29720 ;
  assign w29722 = ~\pi093 & w29721 ;
  assign w29723 = ~w29290 & w29534 ;
  assign w29724 = w29535 ^ w29723 ;
  assign w29725 = ~w29603 & w29724 ;
  assign w29726 = ( w29282 & w29600 ) | ( w29282 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29727 = ~w29602 & w29726 ;
  assign w29728 = w29725 | w29727 ;
  assign w29729 = ~\pi092 & w29728 ;
  assign w29730 = ~w29297 & w29531 ;
  assign w29731 = w29532 ^ w29730 ;
  assign w29732 = ~w29603 & w29731 ;
  assign w29733 = ( w29289 & w29600 ) | ( w29289 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29734 = ~w29602 & w29733 ;
  assign w29735 = w29732 | w29734 ;
  assign w29736 = ~\pi091 & w29735 ;
  assign w29737 = ~w29304 & w29528 ;
  assign w29738 = w29529 ^ w29737 ;
  assign w29739 = ~w29603 & w29738 ;
  assign w29740 = ( w29296 & w29600 ) | ( w29296 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29741 = ~w29602 & w29740 ;
  assign w29742 = w29739 | w29741 ;
  assign w29743 = ~\pi090 & w29742 ;
  assign w29744 = ~w29311 & w29525 ;
  assign w29745 = w29526 ^ w29744 ;
  assign w29746 = ~w29603 & w29745 ;
  assign w29747 = ( w29303 & w29600 ) | ( w29303 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29748 = ~w29602 & w29747 ;
  assign w29749 = w29746 | w29748 ;
  assign w29750 = ~\pi089 & w29749 ;
  assign w29751 = ~w29318 & w29522 ;
  assign w29752 = w29523 ^ w29751 ;
  assign w29753 = ~w29603 & w29752 ;
  assign w29754 = ( w29310 & w29600 ) | ( w29310 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29755 = ~w29602 & w29754 ;
  assign w29756 = w29753 | w29755 ;
  assign w29757 = ~\pi088 & w29756 ;
  assign w29758 = ~w29325 & w29519 ;
  assign w29759 = w29520 ^ w29758 ;
  assign w29760 = ~w29603 & w29759 ;
  assign w29761 = ( w29317 & w29600 ) | ( w29317 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29762 = ~w29602 & w29761 ;
  assign w29763 = w29760 | w29762 ;
  assign w29764 = ~\pi087 & w29763 ;
  assign w29765 = ~w29332 & w29516 ;
  assign w29766 = w29517 ^ w29765 ;
  assign w29767 = ~w29603 & w29766 ;
  assign w29768 = ( w29324 & w29600 ) | ( w29324 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29769 = ~w29602 & w29768 ;
  assign w29770 = w29767 | w29769 ;
  assign w29771 = ~\pi086 & w29770 ;
  assign w29772 = ~w29339 & w29513 ;
  assign w29773 = w29514 ^ w29772 ;
  assign w29774 = ~w29603 & w29773 ;
  assign w29775 = ( w29331 & w29600 ) | ( w29331 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29776 = ~w29602 & w29775 ;
  assign w29777 = w29774 | w29776 ;
  assign w29778 = ~\pi085 & w29777 ;
  assign w29779 = ~w29346 & w29510 ;
  assign w29780 = w29511 ^ w29779 ;
  assign w29781 = ~w29603 & w29780 ;
  assign w29782 = ( w29338 & w29600 ) | ( w29338 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29783 = ~w29602 & w29782 ;
  assign w29784 = w29781 | w29783 ;
  assign w29785 = ~\pi084 & w29784 ;
  assign w29786 = ~w29353 & w29507 ;
  assign w29787 = w29508 ^ w29786 ;
  assign w29788 = ~w29603 & w29787 ;
  assign w29789 = ( w29345 & w29600 ) | ( w29345 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29790 = ~w29602 & w29789 ;
  assign w29791 = w29788 | w29790 ;
  assign w29792 = ~\pi083 & w29791 ;
  assign w29793 = ~w29360 & w29504 ;
  assign w29794 = w29505 ^ w29793 ;
  assign w29795 = ~w29603 & w29794 ;
  assign w29796 = ( w29352 & w29600 ) | ( w29352 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29797 = ~w29602 & w29796 ;
  assign w29798 = w29795 | w29797 ;
  assign w29799 = ~\pi082 & w29798 ;
  assign w29800 = ~w29367 & w29501 ;
  assign w29801 = w29502 ^ w29800 ;
  assign w29802 = ~w29603 & w29801 ;
  assign w29803 = ( w29359 & w29600 ) | ( w29359 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29804 = ~w29602 & w29803 ;
  assign w29805 = w29802 | w29804 ;
  assign w29806 = ~\pi081 & w29805 ;
  assign w29807 = ~w29374 & w29498 ;
  assign w29808 = w29499 ^ w29807 ;
  assign w29809 = ~w29603 & w29808 ;
  assign w29810 = ( w29366 & w29600 ) | ( w29366 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29811 = ~w29602 & w29810 ;
  assign w29812 = w29809 | w29811 ;
  assign w29813 = ~\pi080 & w29812 ;
  assign w29814 = ~w29381 & w29495 ;
  assign w29815 = w29496 ^ w29814 ;
  assign w29816 = ~w29603 & w29815 ;
  assign w29817 = ( w29373 & w29600 ) | ( w29373 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29818 = ~w29602 & w29817 ;
  assign w29819 = w29816 | w29818 ;
  assign w29820 = ~\pi079 & w29819 ;
  assign w29821 = ~w29388 & w29492 ;
  assign w29822 = w29493 ^ w29821 ;
  assign w29823 = ~w29603 & w29822 ;
  assign w29824 = ( w29380 & w29600 ) | ( w29380 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29825 = ~w29602 & w29824 ;
  assign w29826 = w29823 | w29825 ;
  assign w29827 = ~\pi078 & w29826 ;
  assign w29828 = ~w29395 & w29489 ;
  assign w29829 = w29490 ^ w29828 ;
  assign w29830 = ~w29603 & w29829 ;
  assign w29831 = ( w29387 & w29600 ) | ( w29387 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29832 = ~w29602 & w29831 ;
  assign w29833 = w29830 | w29832 ;
  assign w29834 = ~\pi077 & w29833 ;
  assign w29835 = ~w29402 & w29486 ;
  assign w29836 = w29487 ^ w29835 ;
  assign w29837 = ~w29603 & w29836 ;
  assign w29838 = ( w29394 & w29600 ) | ( w29394 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29839 = ~w29602 & w29838 ;
  assign w29840 = w29837 | w29839 ;
  assign w29841 = ~\pi076 & w29840 ;
  assign w29842 = ~w29409 & w29483 ;
  assign w29843 = w29484 ^ w29842 ;
  assign w29844 = ~w29603 & w29843 ;
  assign w29845 = ( w29401 & w29600 ) | ( w29401 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29846 = ~w29602 & w29845 ;
  assign w29847 = w29844 | w29846 ;
  assign w29848 = ~\pi075 & w29847 ;
  assign w29849 = ~w29416 & w29480 ;
  assign w29850 = w29481 ^ w29849 ;
  assign w29851 = ~w29603 & w29850 ;
  assign w29852 = ( w29408 & w29600 ) | ( w29408 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29853 = ~w29602 & w29852 ;
  assign w29854 = w29851 | w29853 ;
  assign w29855 = ~\pi074 & w29854 ;
  assign w29856 = ~w29423 & w29477 ;
  assign w29857 = w29478 ^ w29856 ;
  assign w29858 = ~w29603 & w29857 ;
  assign w29859 = ( w29415 & w29600 ) | ( w29415 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29860 = ~w29602 & w29859 ;
  assign w29861 = w29858 | w29860 ;
  assign w29862 = ~\pi073 & w29861 ;
  assign w29863 = ~w29430 & w29474 ;
  assign w29864 = w29475 ^ w29863 ;
  assign w29865 = ~w29603 & w29864 ;
  assign w29866 = ( w29422 & w29600 ) | ( w29422 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29867 = ~w29602 & w29866 ;
  assign w29868 = w29865 | w29867 ;
  assign w29869 = ~\pi072 & w29868 ;
  assign w29870 = ~w29437 & w29471 ;
  assign w29871 = w29472 ^ w29870 ;
  assign w29872 = ~w29603 & w29871 ;
  assign w29873 = ( w29429 & w29600 ) | ( w29429 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29874 = ~w29602 & w29873 ;
  assign w29875 = w29872 | w29874 ;
  assign w29876 = ~\pi071 & w29875 ;
  assign w29877 = ~w29444 & w29468 ;
  assign w29878 = w29469 ^ w29877 ;
  assign w29879 = ~w29603 & w29878 ;
  assign w29880 = ( w29436 & w29600 ) | ( w29436 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29881 = ~w29602 & w29880 ;
  assign w29882 = w29879 | w29881 ;
  assign w29883 = ~\pi070 & w29882 ;
  assign w29884 = ~w29450 & w29465 ;
  assign w29885 = w29466 ^ w29884 ;
  assign w29886 = ~w29603 & w29885 ;
  assign w29887 = ( w29443 & w29600 ) | ( w29443 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29888 = ~w29602 & w29887 ;
  assign w29889 = w29886 | w29888 ;
  assign w29890 = ~\pi069 & w29889 ;
  assign w29891 = ~w29455 & w29462 ;
  assign w29892 = w29463 ^ w29891 ;
  assign w29893 = ~w29603 & w29892 ;
  assign w29894 = ( w29449 & w29600 ) | ( w29449 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29895 = ~w29602 & w29894 ;
  assign w29896 = w29893 | w29895 ;
  assign w29897 = ~\pi068 & w29896 ;
  assign w29898 = \pi064 & ~w29164 ;
  assign w29899 = \pi020 ^ w29898 ;
  assign w29900 = ( \pi065 & w10495 ) | ( \pi065 & ~w29899 ) | ( w10495 & ~w29899 ) ;
  assign w29901 = w29458 ^ w29900 ;
  assign w29902 = ~w29603 & w29901 ;
  assign w29903 = ( w29454 & w29600 ) | ( w29454 & w29602 ) | ( w29600 & w29602 ) ;
  assign w29904 = ~w29602 & w29903 ;
  assign w29905 = w29902 | w29904 ;
  assign w29906 = ~\pi067 & w29905 ;
  assign w29907 = \pi019 ^ w29164 ;
  assign w29908 = ( \pi064 & w29603 ) | ( \pi064 & w29907 ) | ( w29603 & w29907 ) ;
  assign w29909 = w10503 ^ w29908 ;
  assign w29910 = ~w29603 & w29909 ;
  assign w29911 = w29603 & w29899 ;
  assign w29912 = w29910 | w29911 ;
  assign w29913 = ~\pi066 & w29912 ;
  assign w29914 = \pi066 ^ w29912 ;
  assign w29915 = ( \pi064 & ~w29603 ) | ( \pi064 & w29914 ) | ( ~w29603 & w29914 ) ;
  assign w29916 = \pi019 ^ w29915 ;
  assign w29917 = ( \pi065 & w10904 ) | ( \pi065 & ~w29916 ) | ( w10904 & ~w29916 ) ;
  assign w29918 = w29914 | w29917 ;
  assign w29919 = \pi067 ^ w29905 ;
  assign w29920 = ( ~w29913 & w29918 ) | ( ~w29913 & w29919 ) | ( w29918 & w29919 ) ;
  assign w29921 = w29919 | w29920 ;
  assign w29922 = \pi068 ^ w29896 ;
  assign w29923 = ( ~w29906 & w29921 ) | ( ~w29906 & w29922 ) | ( w29921 & w29922 ) ;
  assign w29924 = w29922 | w29923 ;
  assign w29925 = \pi069 ^ w29889 ;
  assign w29926 = ( ~w29897 & w29924 ) | ( ~w29897 & w29925 ) | ( w29924 & w29925 ) ;
  assign w29927 = w29925 | w29926 ;
  assign w29928 = \pi070 ^ w29882 ;
  assign w29929 = ( ~w29890 & w29927 ) | ( ~w29890 & w29928 ) | ( w29927 & w29928 ) ;
  assign w29930 = w29928 | w29929 ;
  assign w29931 = \pi071 ^ w29875 ;
  assign w29932 = ( ~w29883 & w29930 ) | ( ~w29883 & w29931 ) | ( w29930 & w29931 ) ;
  assign w29933 = w29931 | w29932 ;
  assign w29934 = \pi072 ^ w29868 ;
  assign w29935 = ( ~w29876 & w29933 ) | ( ~w29876 & w29934 ) | ( w29933 & w29934 ) ;
  assign w29936 = w29934 | w29935 ;
  assign w29937 = \pi073 ^ w29861 ;
  assign w29938 = ( ~w29869 & w29936 ) | ( ~w29869 & w29937 ) | ( w29936 & w29937 ) ;
  assign w29939 = w29937 | w29938 ;
  assign w29940 = \pi074 ^ w29854 ;
  assign w29941 = ( ~w29862 & w29939 ) | ( ~w29862 & w29940 ) | ( w29939 & w29940 ) ;
  assign w29942 = w29940 | w29941 ;
  assign w29943 = \pi075 ^ w29847 ;
  assign w29944 = ( ~w29855 & w29942 ) | ( ~w29855 & w29943 ) | ( w29942 & w29943 ) ;
  assign w29945 = w29943 | w29944 ;
  assign w29946 = \pi076 ^ w29840 ;
  assign w29947 = ( ~w29848 & w29945 ) | ( ~w29848 & w29946 ) | ( w29945 & w29946 ) ;
  assign w29948 = w29946 | w29947 ;
  assign w29949 = \pi077 ^ w29833 ;
  assign w29950 = ( ~w29841 & w29948 ) | ( ~w29841 & w29949 ) | ( w29948 & w29949 ) ;
  assign w29951 = w29949 | w29950 ;
  assign w29952 = \pi078 ^ w29826 ;
  assign w29953 = ( ~w29834 & w29951 ) | ( ~w29834 & w29952 ) | ( w29951 & w29952 ) ;
  assign w29954 = w29952 | w29953 ;
  assign w29955 = \pi079 ^ w29819 ;
  assign w29956 = ( ~w29827 & w29954 ) | ( ~w29827 & w29955 ) | ( w29954 & w29955 ) ;
  assign w29957 = w29955 | w29956 ;
  assign w29958 = \pi080 ^ w29812 ;
  assign w29959 = ( ~w29820 & w29957 ) | ( ~w29820 & w29958 ) | ( w29957 & w29958 ) ;
  assign w29960 = w29958 | w29959 ;
  assign w29961 = \pi081 ^ w29805 ;
  assign w29962 = ( ~w29813 & w29960 ) | ( ~w29813 & w29961 ) | ( w29960 & w29961 ) ;
  assign w29963 = w29961 | w29962 ;
  assign w29964 = \pi082 ^ w29798 ;
  assign w29965 = ( ~w29806 & w29963 ) | ( ~w29806 & w29964 ) | ( w29963 & w29964 ) ;
  assign w29966 = w29964 | w29965 ;
  assign w29967 = \pi083 ^ w29791 ;
  assign w29968 = ( ~w29799 & w29966 ) | ( ~w29799 & w29967 ) | ( w29966 & w29967 ) ;
  assign w29969 = w29967 | w29968 ;
  assign w29970 = \pi084 ^ w29784 ;
  assign w29971 = ( ~w29792 & w29969 ) | ( ~w29792 & w29970 ) | ( w29969 & w29970 ) ;
  assign w29972 = w29970 | w29971 ;
  assign w29973 = \pi085 ^ w29777 ;
  assign w29974 = ( ~w29785 & w29972 ) | ( ~w29785 & w29973 ) | ( w29972 & w29973 ) ;
  assign w29975 = w29973 | w29974 ;
  assign w29976 = \pi086 ^ w29770 ;
  assign w29977 = ( ~w29778 & w29975 ) | ( ~w29778 & w29976 ) | ( w29975 & w29976 ) ;
  assign w29978 = w29976 | w29977 ;
  assign w29979 = \pi087 ^ w29763 ;
  assign w29980 = ( ~w29771 & w29978 ) | ( ~w29771 & w29979 ) | ( w29978 & w29979 ) ;
  assign w29981 = w29979 | w29980 ;
  assign w29982 = \pi088 ^ w29756 ;
  assign w29983 = ( ~w29764 & w29981 ) | ( ~w29764 & w29982 ) | ( w29981 & w29982 ) ;
  assign w29984 = w29982 | w29983 ;
  assign w29985 = \pi089 ^ w29749 ;
  assign w29986 = ( ~w29757 & w29984 ) | ( ~w29757 & w29985 ) | ( w29984 & w29985 ) ;
  assign w29987 = w29985 | w29986 ;
  assign w29988 = \pi090 ^ w29742 ;
  assign w29989 = ( ~w29750 & w29987 ) | ( ~w29750 & w29988 ) | ( w29987 & w29988 ) ;
  assign w29990 = w29988 | w29989 ;
  assign w29991 = \pi091 ^ w29735 ;
  assign w29992 = ( ~w29743 & w29990 ) | ( ~w29743 & w29991 ) | ( w29990 & w29991 ) ;
  assign w29993 = w29991 | w29992 ;
  assign w29994 = \pi092 ^ w29728 ;
  assign w29995 = ( ~w29736 & w29993 ) | ( ~w29736 & w29994 ) | ( w29993 & w29994 ) ;
  assign w29996 = w29994 | w29995 ;
  assign w29997 = \pi093 ^ w29721 ;
  assign w29998 = ( ~w29729 & w29996 ) | ( ~w29729 & w29997 ) | ( w29996 & w29997 ) ;
  assign w29999 = w29997 | w29998 ;
  assign w30000 = \pi094 ^ w29714 ;
  assign w30001 = ( ~w29722 & w29999 ) | ( ~w29722 & w30000 ) | ( w29999 & w30000 ) ;
  assign w30002 = w30000 | w30001 ;
  assign w30003 = \pi095 ^ w29707 ;
  assign w30004 = ( ~w29715 & w30002 ) | ( ~w29715 & w30003 ) | ( w30002 & w30003 ) ;
  assign w30005 = w30003 | w30004 ;
  assign w30006 = \pi096 ^ w29700 ;
  assign w30007 = ( ~w29708 & w30005 ) | ( ~w29708 & w30006 ) | ( w30005 & w30006 ) ;
  assign w30008 = w30006 | w30007 ;
  assign w30009 = \pi097 ^ w29693 ;
  assign w30010 = ( ~w29701 & w30008 ) | ( ~w29701 & w30009 ) | ( w30008 & w30009 ) ;
  assign w30011 = w30009 | w30010 ;
  assign w30012 = \pi098 ^ w29686 ;
  assign w30013 = ( ~w29694 & w30011 ) | ( ~w29694 & w30012 ) | ( w30011 & w30012 ) ;
  assign w30014 = w30012 | w30013 ;
  assign w30015 = \pi099 ^ w29679 ;
  assign w30016 = ( ~w29687 & w30014 ) | ( ~w29687 & w30015 ) | ( w30014 & w30015 ) ;
  assign w30017 = w30015 | w30016 ;
  assign w30018 = \pi100 ^ w29672 ;
  assign w30019 = ( ~w29680 & w30017 ) | ( ~w29680 & w30018 ) | ( w30017 & w30018 ) ;
  assign w30020 = w30018 | w30019 ;
  assign w30021 = \pi101 ^ w29665 ;
  assign w30022 = ( ~w29673 & w30020 ) | ( ~w29673 & w30021 ) | ( w30020 & w30021 ) ;
  assign w30023 = w30021 | w30022 ;
  assign w30024 = \pi102 ^ w29658 ;
  assign w30025 = ( ~w29666 & w30023 ) | ( ~w29666 & w30024 ) | ( w30023 & w30024 ) ;
  assign w30026 = w30024 | w30025 ;
  assign w30027 = \pi103 ^ w29651 ;
  assign w30028 = ( ~w29659 & w30026 ) | ( ~w29659 & w30027 ) | ( w30026 & w30027 ) ;
  assign w30029 = w30027 | w30028 ;
  assign w30030 = \pi104 ^ w29644 ;
  assign w30031 = ( ~w29652 & w30029 ) | ( ~w29652 & w30030 ) | ( w30029 & w30030 ) ;
  assign w30032 = w30030 | w30031 ;
  assign w30033 = \pi105 ^ w29637 ;
  assign w30034 = ( ~w29645 & w30032 ) | ( ~w29645 & w30033 ) | ( w30032 & w30033 ) ;
  assign w30035 = w30033 | w30034 ;
  assign w30036 = \pi106 ^ w29630 ;
  assign w30037 = ( ~w29638 & w30035 ) | ( ~w29638 & w30036 ) | ( w30035 & w30036 ) ;
  assign w30038 = w30036 | w30037 ;
  assign w30039 = \pi107 ^ w29623 ;
  assign w30040 = ( ~w29631 & w30038 ) | ( ~w29631 & w30039 ) | ( w30038 & w30039 ) ;
  assign w30041 = w30039 | w30040 ;
  assign w30042 = \pi108 ^ w29609 ;
  assign w30043 = ( ~w29624 & w30041 ) | ( ~w29624 & w30042 ) | ( w30041 & w30042 ) ;
  assign w30044 = w30042 | w30043 ;
  assign w30045 = \pi109 ^ w29616 ;
  assign w30046 = w29617 & ~w30045 ;
  assign w30047 = ( w30044 & w30045 ) | ( w30044 & ~w30046 ) | ( w30045 & ~w30046 ) ;
  assign w30048 = ~\pi109 & w29616 ;
  assign w30049 = w30047 & ~w30048 ;
  assign w30050 = w10650 | w30049 ;
  assign w30051 = w29609 & w30050 ;
  assign w30052 = ~w29624 & w30041 ;
  assign w30053 = w30042 ^ w30052 ;
  assign w30054 = ~w30050 & w30053 ;
  assign w30055 = w30051 | w30054 ;
  assign w30056 = ~\pi109 & w30055 ;
  assign w30057 = w29623 & w30050 ;
  assign w30058 = ~w29631 & w30038 ;
  assign w30059 = w30039 ^ w30058 ;
  assign w30060 = ~w30050 & w30059 ;
  assign w30061 = w30057 | w30060 ;
  assign w30062 = ~\pi108 & w30061 ;
  assign w30063 = w29630 & w30050 ;
  assign w30064 = ~w29638 & w30035 ;
  assign w30065 = w30036 ^ w30064 ;
  assign w30066 = ~w30050 & w30065 ;
  assign w30067 = w30063 | w30066 ;
  assign w30068 = ~\pi107 & w30067 ;
  assign w30069 = w29637 & w30050 ;
  assign w30070 = ~w29645 & w30032 ;
  assign w30071 = w30033 ^ w30070 ;
  assign w30072 = ~w30050 & w30071 ;
  assign w30073 = w30069 | w30072 ;
  assign w30074 = ~\pi106 & w30073 ;
  assign w30075 = w29644 & w30050 ;
  assign w30076 = ~w29652 & w30029 ;
  assign w30077 = w30030 ^ w30076 ;
  assign w30078 = ~w30050 & w30077 ;
  assign w30079 = w30075 | w30078 ;
  assign w30080 = ~\pi105 & w30079 ;
  assign w30081 = w29651 & w30050 ;
  assign w30082 = ~w29659 & w30026 ;
  assign w30083 = w30027 ^ w30082 ;
  assign w30084 = ~w30050 & w30083 ;
  assign w30085 = w30081 | w30084 ;
  assign w30086 = ~\pi104 & w30085 ;
  assign w30087 = w29658 & w30050 ;
  assign w30088 = ~w29666 & w30023 ;
  assign w30089 = w30024 ^ w30088 ;
  assign w30090 = ~w30050 & w30089 ;
  assign w30091 = w30087 | w30090 ;
  assign w30092 = ~\pi103 & w30091 ;
  assign w30093 = w29665 & w30050 ;
  assign w30094 = ~w29673 & w30020 ;
  assign w30095 = w30021 ^ w30094 ;
  assign w30096 = ~w30050 & w30095 ;
  assign w30097 = w30093 | w30096 ;
  assign w30098 = ~\pi102 & w30097 ;
  assign w30099 = w29672 & w30050 ;
  assign w30100 = ~w29680 & w30017 ;
  assign w30101 = w30018 ^ w30100 ;
  assign w30102 = ~w30050 & w30101 ;
  assign w30103 = w30099 | w30102 ;
  assign w30104 = ~\pi101 & w30103 ;
  assign w30105 = w29679 & w30050 ;
  assign w30106 = ~w29687 & w30014 ;
  assign w30107 = w30015 ^ w30106 ;
  assign w30108 = ~w30050 & w30107 ;
  assign w30109 = w30105 | w30108 ;
  assign w30110 = ~\pi100 & w30109 ;
  assign w30111 = w29686 & w30050 ;
  assign w30112 = ~w29694 & w30011 ;
  assign w30113 = w30012 ^ w30112 ;
  assign w30114 = ~w30050 & w30113 ;
  assign w30115 = w30111 | w30114 ;
  assign w30116 = ~\pi099 & w30115 ;
  assign w30117 = w29693 & w30050 ;
  assign w30118 = ~w29701 & w30008 ;
  assign w30119 = w30009 ^ w30118 ;
  assign w30120 = ~w30050 & w30119 ;
  assign w30121 = w30117 | w30120 ;
  assign w30122 = ~\pi098 & w30121 ;
  assign w30123 = w29700 & w30050 ;
  assign w30124 = ~w29708 & w30005 ;
  assign w30125 = w30006 ^ w30124 ;
  assign w30126 = ~w30050 & w30125 ;
  assign w30127 = w30123 | w30126 ;
  assign w30128 = ~\pi097 & w30127 ;
  assign w30129 = w29707 & w30050 ;
  assign w30130 = ~w29715 & w30002 ;
  assign w30131 = w30003 ^ w30130 ;
  assign w30132 = ~w30050 & w30131 ;
  assign w30133 = w30129 | w30132 ;
  assign w30134 = ~\pi096 & w30133 ;
  assign w30135 = w29714 & w30050 ;
  assign w30136 = ~w29722 & w29999 ;
  assign w30137 = w30000 ^ w30136 ;
  assign w30138 = ~w30050 & w30137 ;
  assign w30139 = w30135 | w30138 ;
  assign w30140 = ~\pi095 & w30139 ;
  assign w30141 = w29721 & w30050 ;
  assign w30142 = ~w29729 & w29996 ;
  assign w30143 = w29997 ^ w30142 ;
  assign w30144 = ~w30050 & w30143 ;
  assign w30145 = w30141 | w30144 ;
  assign w30146 = ~\pi094 & w30145 ;
  assign w30147 = w29728 & w30050 ;
  assign w30148 = ~w29736 & w29993 ;
  assign w30149 = w29994 ^ w30148 ;
  assign w30150 = ~w30050 & w30149 ;
  assign w30151 = w30147 | w30150 ;
  assign w30152 = ~\pi093 & w30151 ;
  assign w30153 = w29735 & w30050 ;
  assign w30154 = ~w29743 & w29990 ;
  assign w30155 = w29991 ^ w30154 ;
  assign w30156 = ~w30050 & w30155 ;
  assign w30157 = w30153 | w30156 ;
  assign w30158 = ~\pi092 & w30157 ;
  assign w30159 = w29742 & w30050 ;
  assign w30160 = ~w29750 & w29987 ;
  assign w30161 = w29988 ^ w30160 ;
  assign w30162 = ~w30050 & w30161 ;
  assign w30163 = w30159 | w30162 ;
  assign w30164 = ~\pi091 & w30163 ;
  assign w30165 = w29749 & w30050 ;
  assign w30166 = ~w29757 & w29984 ;
  assign w30167 = w29985 ^ w30166 ;
  assign w30168 = ~w30050 & w30167 ;
  assign w30169 = w30165 | w30168 ;
  assign w30170 = ~\pi090 & w30169 ;
  assign w30171 = w29756 & w30050 ;
  assign w30172 = ~w29764 & w29981 ;
  assign w30173 = w29982 ^ w30172 ;
  assign w30174 = ~w30050 & w30173 ;
  assign w30175 = w30171 | w30174 ;
  assign w30176 = ~\pi089 & w30175 ;
  assign w30177 = w29763 & w30050 ;
  assign w30178 = ~w29771 & w29978 ;
  assign w30179 = w29979 ^ w30178 ;
  assign w30180 = ~w30050 & w30179 ;
  assign w30181 = w30177 | w30180 ;
  assign w30182 = ~\pi088 & w30181 ;
  assign w30183 = w29770 & w30050 ;
  assign w30184 = ~w29778 & w29975 ;
  assign w30185 = w29976 ^ w30184 ;
  assign w30186 = ~w30050 & w30185 ;
  assign w30187 = w30183 | w30186 ;
  assign w30188 = ~\pi087 & w30187 ;
  assign w30189 = w29777 & w30050 ;
  assign w30190 = ~w29785 & w29972 ;
  assign w30191 = w29973 ^ w30190 ;
  assign w30192 = ~w30050 & w30191 ;
  assign w30193 = w30189 | w30192 ;
  assign w30194 = ~\pi086 & w30193 ;
  assign w30195 = w29784 & w30050 ;
  assign w30196 = ~w29792 & w29969 ;
  assign w30197 = w29970 ^ w30196 ;
  assign w30198 = ~w30050 & w30197 ;
  assign w30199 = w30195 | w30198 ;
  assign w30200 = ~\pi085 & w30199 ;
  assign w30201 = w29791 & w30050 ;
  assign w30202 = ~w29799 & w29966 ;
  assign w30203 = w29967 ^ w30202 ;
  assign w30204 = ~w30050 & w30203 ;
  assign w30205 = w30201 | w30204 ;
  assign w30206 = ~\pi084 & w30205 ;
  assign w30207 = w29798 & w30050 ;
  assign w30208 = ~w29806 & w29963 ;
  assign w30209 = w29964 ^ w30208 ;
  assign w30210 = ~w30050 & w30209 ;
  assign w30211 = w30207 | w30210 ;
  assign w30212 = ~\pi083 & w30211 ;
  assign w30213 = w29805 & w30050 ;
  assign w30214 = ~w29813 & w29960 ;
  assign w30215 = w29961 ^ w30214 ;
  assign w30216 = ~w30050 & w30215 ;
  assign w30217 = w30213 | w30216 ;
  assign w30218 = ~\pi082 & w30217 ;
  assign w30219 = w29812 & w30050 ;
  assign w30220 = ~w29820 & w29957 ;
  assign w30221 = w29958 ^ w30220 ;
  assign w30222 = ~w30050 & w30221 ;
  assign w30223 = w30219 | w30222 ;
  assign w30224 = ~\pi081 & w30223 ;
  assign w30225 = w29819 & w30050 ;
  assign w30226 = ~w29827 & w29954 ;
  assign w30227 = w29955 ^ w30226 ;
  assign w30228 = ~w30050 & w30227 ;
  assign w30229 = w30225 | w30228 ;
  assign w30230 = ~\pi080 & w30229 ;
  assign w30231 = w29826 & w30050 ;
  assign w30232 = ~w29834 & w29951 ;
  assign w30233 = w29952 ^ w30232 ;
  assign w30234 = ~w30050 & w30233 ;
  assign w30235 = w30231 | w30234 ;
  assign w30236 = ~\pi079 & w30235 ;
  assign w30237 = w29833 & w30050 ;
  assign w30238 = ~w29841 & w29948 ;
  assign w30239 = w29949 ^ w30238 ;
  assign w30240 = ~w30050 & w30239 ;
  assign w30241 = w30237 | w30240 ;
  assign w30242 = ~\pi078 & w30241 ;
  assign w30243 = w29840 & w30050 ;
  assign w30244 = ~w29848 & w29945 ;
  assign w30245 = w29946 ^ w30244 ;
  assign w30246 = ~w30050 & w30245 ;
  assign w30247 = w30243 | w30246 ;
  assign w30248 = ~\pi077 & w30247 ;
  assign w30249 = w29847 & w30050 ;
  assign w30250 = ~w29855 & w29942 ;
  assign w30251 = w29943 ^ w30250 ;
  assign w30252 = ~w30050 & w30251 ;
  assign w30253 = w30249 | w30252 ;
  assign w30254 = ~\pi076 & w30253 ;
  assign w30255 = w29854 & w30050 ;
  assign w30256 = ~w29862 & w29939 ;
  assign w30257 = w29940 ^ w30256 ;
  assign w30258 = ~w30050 & w30257 ;
  assign w30259 = w30255 | w30258 ;
  assign w30260 = ~\pi075 & w30259 ;
  assign w30261 = w29861 & w30050 ;
  assign w30262 = ~w29869 & w29936 ;
  assign w30263 = w29937 ^ w30262 ;
  assign w30264 = ~w30050 & w30263 ;
  assign w30265 = w30261 | w30264 ;
  assign w30266 = ~\pi074 & w30265 ;
  assign w30267 = w29868 & w30050 ;
  assign w30268 = ~w29876 & w29933 ;
  assign w30269 = w29934 ^ w30268 ;
  assign w30270 = ~w30050 & w30269 ;
  assign w30271 = w30267 | w30270 ;
  assign w30272 = ~\pi073 & w30271 ;
  assign w30273 = w29875 & w30050 ;
  assign w30274 = ~w29883 & w29930 ;
  assign w30275 = w29931 ^ w30274 ;
  assign w30276 = ~w30050 & w30275 ;
  assign w30277 = w30273 | w30276 ;
  assign w30278 = ~\pi072 & w30277 ;
  assign w30279 = w29882 & w30050 ;
  assign w30280 = ~w29890 & w29927 ;
  assign w30281 = w29928 ^ w30280 ;
  assign w30282 = ~w30050 & w30281 ;
  assign w30283 = w30279 | w30282 ;
  assign w30284 = ~\pi071 & w30283 ;
  assign w30285 = w29889 & w30050 ;
  assign w30286 = ~w29897 & w29924 ;
  assign w30287 = w29925 ^ w30286 ;
  assign w30288 = ~w30050 & w30287 ;
  assign w30289 = w30285 | w30288 ;
  assign w30290 = ~\pi070 & w30289 ;
  assign w30291 = w29896 & w30050 ;
  assign w30292 = ~w29906 & w29921 ;
  assign w30293 = w29922 ^ w30292 ;
  assign w30294 = ~w30050 & w30293 ;
  assign w30295 = w30291 | w30294 ;
  assign w30296 = ~\pi069 & w30295 ;
  assign w30297 = w29905 & w30050 ;
  assign w30298 = ~w29913 & w29918 ;
  assign w30299 = w29919 ^ w30298 ;
  assign w30300 = ~w30050 & w30299 ;
  assign w30301 = w30297 | w30300 ;
  assign w30302 = ~\pi068 & w30301 ;
  assign w30303 = \pi064 & ~w29603 ;
  assign w30304 = \pi019 ^ w30303 ;
  assign w30305 = ( \pi065 & w10904 ) | ( \pi065 & ~w30304 ) | ( w10904 & ~w30304 ) ;
  assign w30306 = w29914 ^ w30305 ;
  assign w30307 = ( w10650 & w30049 ) | ( w10650 & w30306 ) | ( w30049 & w30306 ) ;
  assign w30308 = w30306 & ~w30307 ;
  assign w30309 = ( w29912 & w30050 ) | ( w29912 & w30308 ) | ( w30050 & w30308 ) ;
  assign w30310 = w30308 | w30309 ;
  assign w30311 = ~\pi067 & w30310 ;
  assign w30312 = \pi018 ^ w29603 ;
  assign w30313 = ( \pi064 & w10650 ) | ( \pi064 & w30312 ) | ( w10650 & w30312 ) ;
  assign w30314 = w10912 ^ w30313 ;
  assign w30315 = ~w10650 & w30314 ;
  assign w30316 = ~w30049 & w30315 ;
  assign w30317 = ( ~\pi064 & w29603 ) | ( ~\pi064 & w30050 ) | ( w29603 & w30050 ) ;
  assign w30318 = \pi019 ^ w30317 ;
  assign w30319 = w30050 & ~w30318 ;
  assign w30320 = w30316 | w30319 ;
  assign w30321 = ~\pi066 & w30320 ;
  assign w30322 = ( \pi018 & ~w10927 ) | ( \pi018 & w30049 ) | ( ~w10927 & w30049 ) ;
  assign w30323 = \pi018 & w30322 ;
  assign w30324 = w10934 & ~w30049 ;
  assign w30325 = w30323 | w30324 ;
  assign w30326 = \pi065 ^ w30325 ;
  assign w30327 = w10937 | w30326 ;
  assign w30328 = w30050 | w30316 ;
  assign w30329 = ( w30304 & w30316 ) | ( w30304 & w30328 ) | ( w30316 & w30328 ) ;
  assign w30330 = \pi066 ^ w30329 ;
  assign w30331 = ~\pi065 & w30325 ;
  assign w30332 = w30327 | w30331 ;
  assign w30333 = ( w30330 & ~w30331 ) | ( w30330 & w30332 ) | ( ~w30331 & w30332 ) ;
  assign w30334 = ~w29912 & w30050 ;
  assign w30335 = ( w30050 & w30308 ) | ( w30050 & ~w30334 ) | ( w30308 & ~w30334 ) ;
  assign w30336 = \pi067 ^ w30335 ;
  assign w30337 = ( ~w30321 & w30333 ) | ( ~w30321 & w30336 ) | ( w30333 & w30336 ) ;
  assign w30338 = w30336 | w30337 ;
  assign w30339 = \pi068 ^ w30301 ;
  assign w30340 = ( ~w30311 & w30338 ) | ( ~w30311 & w30339 ) | ( w30338 & w30339 ) ;
  assign w30341 = w30339 | w30340 ;
  assign w30342 = \pi069 ^ w30295 ;
  assign w30343 = ( ~w30302 & w30341 ) | ( ~w30302 & w30342 ) | ( w30341 & w30342 ) ;
  assign w30344 = w30342 | w30343 ;
  assign w30345 = \pi070 ^ w30289 ;
  assign w30346 = ( ~w30296 & w30344 ) | ( ~w30296 & w30345 ) | ( w30344 & w30345 ) ;
  assign w30347 = w30345 | w30346 ;
  assign w30348 = \pi071 ^ w30283 ;
  assign w30349 = ( ~w30290 & w30347 ) | ( ~w30290 & w30348 ) | ( w30347 & w30348 ) ;
  assign w30350 = w30348 | w30349 ;
  assign w30351 = \pi072 ^ w30277 ;
  assign w30352 = ( ~w30284 & w30350 ) | ( ~w30284 & w30351 ) | ( w30350 & w30351 ) ;
  assign w30353 = w30351 | w30352 ;
  assign w30354 = \pi073 ^ w30271 ;
  assign w30355 = ( ~w30278 & w30353 ) | ( ~w30278 & w30354 ) | ( w30353 & w30354 ) ;
  assign w30356 = w30354 | w30355 ;
  assign w30357 = \pi074 ^ w30265 ;
  assign w30358 = ( ~w30272 & w30356 ) | ( ~w30272 & w30357 ) | ( w30356 & w30357 ) ;
  assign w30359 = w30357 | w30358 ;
  assign w30360 = \pi075 ^ w30259 ;
  assign w30361 = ( ~w30266 & w30359 ) | ( ~w30266 & w30360 ) | ( w30359 & w30360 ) ;
  assign w30362 = w30360 | w30361 ;
  assign w30363 = \pi076 ^ w30253 ;
  assign w30364 = ( ~w30260 & w30362 ) | ( ~w30260 & w30363 ) | ( w30362 & w30363 ) ;
  assign w30365 = w30363 | w30364 ;
  assign w30366 = \pi077 ^ w30247 ;
  assign w30367 = ( ~w30254 & w30365 ) | ( ~w30254 & w30366 ) | ( w30365 & w30366 ) ;
  assign w30368 = w30366 | w30367 ;
  assign w30369 = \pi078 ^ w30241 ;
  assign w30370 = ( ~w30248 & w30368 ) | ( ~w30248 & w30369 ) | ( w30368 & w30369 ) ;
  assign w30371 = w30369 | w30370 ;
  assign w30372 = \pi079 ^ w30235 ;
  assign w30373 = ( ~w30242 & w30371 ) | ( ~w30242 & w30372 ) | ( w30371 & w30372 ) ;
  assign w30374 = w30372 | w30373 ;
  assign w30375 = \pi080 ^ w30229 ;
  assign w30376 = ( ~w30236 & w30374 ) | ( ~w30236 & w30375 ) | ( w30374 & w30375 ) ;
  assign w30377 = w30375 | w30376 ;
  assign w30378 = \pi081 ^ w30223 ;
  assign w30379 = ( ~w30230 & w30377 ) | ( ~w30230 & w30378 ) | ( w30377 & w30378 ) ;
  assign w30380 = w30378 | w30379 ;
  assign w30381 = \pi082 ^ w30217 ;
  assign w30382 = ( ~w30224 & w30380 ) | ( ~w30224 & w30381 ) | ( w30380 & w30381 ) ;
  assign w30383 = w30381 | w30382 ;
  assign w30384 = \pi083 ^ w30211 ;
  assign w30385 = ( ~w30218 & w30383 ) | ( ~w30218 & w30384 ) | ( w30383 & w30384 ) ;
  assign w30386 = w30384 | w30385 ;
  assign w30387 = \pi084 ^ w30205 ;
  assign w30388 = ( ~w30212 & w30386 ) | ( ~w30212 & w30387 ) | ( w30386 & w30387 ) ;
  assign w30389 = w30387 | w30388 ;
  assign w30390 = \pi085 ^ w30199 ;
  assign w30391 = ( ~w30206 & w30389 ) | ( ~w30206 & w30390 ) | ( w30389 & w30390 ) ;
  assign w30392 = w30390 | w30391 ;
  assign w30393 = \pi086 ^ w30193 ;
  assign w30394 = ( ~w30200 & w30392 ) | ( ~w30200 & w30393 ) | ( w30392 & w30393 ) ;
  assign w30395 = w30393 | w30394 ;
  assign w30396 = \pi087 ^ w30187 ;
  assign w30397 = ( ~w30194 & w30395 ) | ( ~w30194 & w30396 ) | ( w30395 & w30396 ) ;
  assign w30398 = w30396 | w30397 ;
  assign w30399 = \pi088 ^ w30181 ;
  assign w30400 = ( ~w30188 & w30398 ) | ( ~w30188 & w30399 ) | ( w30398 & w30399 ) ;
  assign w30401 = w30399 | w30400 ;
  assign w30402 = \pi089 ^ w30175 ;
  assign w30403 = ( ~w30182 & w30401 ) | ( ~w30182 & w30402 ) | ( w30401 & w30402 ) ;
  assign w30404 = w30402 | w30403 ;
  assign w30405 = \pi090 ^ w30169 ;
  assign w30406 = ( ~w30176 & w30404 ) | ( ~w30176 & w30405 ) | ( w30404 & w30405 ) ;
  assign w30407 = w30405 | w30406 ;
  assign w30408 = \pi091 ^ w30163 ;
  assign w30409 = ( ~w30170 & w30407 ) | ( ~w30170 & w30408 ) | ( w30407 & w30408 ) ;
  assign w30410 = w30408 | w30409 ;
  assign w30411 = \pi092 ^ w30157 ;
  assign w30412 = ( ~w30164 & w30410 ) | ( ~w30164 & w30411 ) | ( w30410 & w30411 ) ;
  assign w30413 = w30411 | w30412 ;
  assign w30414 = \pi093 ^ w30151 ;
  assign w30415 = ( ~w30158 & w30413 ) | ( ~w30158 & w30414 ) | ( w30413 & w30414 ) ;
  assign w30416 = w30414 | w30415 ;
  assign w30417 = \pi094 ^ w30145 ;
  assign w30418 = ( ~w30152 & w30416 ) | ( ~w30152 & w30417 ) | ( w30416 & w30417 ) ;
  assign w30419 = w30417 | w30418 ;
  assign w30420 = \pi095 ^ w30139 ;
  assign w30421 = ( ~w30146 & w30419 ) | ( ~w30146 & w30420 ) | ( w30419 & w30420 ) ;
  assign w30422 = w30420 | w30421 ;
  assign w30423 = \pi096 ^ w30133 ;
  assign w30424 = ( ~w30140 & w30422 ) | ( ~w30140 & w30423 ) | ( w30422 & w30423 ) ;
  assign w30425 = w30423 | w30424 ;
  assign w30426 = \pi097 ^ w30127 ;
  assign w30427 = ( ~w30134 & w30425 ) | ( ~w30134 & w30426 ) | ( w30425 & w30426 ) ;
  assign w30428 = w30426 | w30427 ;
  assign w30429 = \pi098 ^ w30121 ;
  assign w30430 = ( ~w30128 & w30428 ) | ( ~w30128 & w30429 ) | ( w30428 & w30429 ) ;
  assign w30431 = w30429 | w30430 ;
  assign w30432 = \pi099 ^ w30115 ;
  assign w30433 = ( ~w30122 & w30431 ) | ( ~w30122 & w30432 ) | ( w30431 & w30432 ) ;
  assign w30434 = w30432 | w30433 ;
  assign w30435 = \pi100 ^ w30109 ;
  assign w30436 = ( ~w30116 & w30434 ) | ( ~w30116 & w30435 ) | ( w30434 & w30435 ) ;
  assign w30437 = w30435 | w30436 ;
  assign w30438 = \pi101 ^ w30103 ;
  assign w30439 = ( ~w30110 & w30437 ) | ( ~w30110 & w30438 ) | ( w30437 & w30438 ) ;
  assign w30440 = w30438 | w30439 ;
  assign w30441 = \pi102 ^ w30097 ;
  assign w30442 = ( ~w30104 & w30440 ) | ( ~w30104 & w30441 ) | ( w30440 & w30441 ) ;
  assign w30443 = w30441 | w30442 ;
  assign w30444 = \pi103 ^ w30091 ;
  assign w30445 = ( ~w30098 & w30443 ) | ( ~w30098 & w30444 ) | ( w30443 & w30444 ) ;
  assign w30446 = w30444 | w30445 ;
  assign w30447 = \pi104 ^ w30085 ;
  assign w30448 = ( ~w30092 & w30446 ) | ( ~w30092 & w30447 ) | ( w30446 & w30447 ) ;
  assign w30449 = w30447 | w30448 ;
  assign w30450 = \pi105 ^ w30079 ;
  assign w30451 = ( ~w30086 & w30449 ) | ( ~w30086 & w30450 ) | ( w30449 & w30450 ) ;
  assign w30452 = w30450 | w30451 ;
  assign w30453 = \pi106 ^ w30073 ;
  assign w30454 = ( ~w30080 & w30452 ) | ( ~w30080 & w30453 ) | ( w30452 & w30453 ) ;
  assign w30455 = w30453 | w30454 ;
  assign w30456 = \pi107 ^ w30067 ;
  assign w30457 = ( ~w30074 & w30455 ) | ( ~w30074 & w30456 ) | ( w30455 & w30456 ) ;
  assign w30458 = w30456 | w30457 ;
  assign w30459 = \pi108 ^ w30061 ;
  assign w30460 = ( ~w30068 & w30458 ) | ( ~w30068 & w30459 ) | ( w30458 & w30459 ) ;
  assign w30461 = w30459 | w30460 ;
  assign w30462 = \pi109 ^ w30055 ;
  assign w30463 = ( ~w30062 & w30461 ) | ( ~w30062 & w30462 ) | ( w30461 & w30462 ) ;
  assign w30464 = w30462 | w30463 ;
  assign w30465 = w29616 & w30050 ;
  assign w30466 = ~w29617 & w30044 ;
  assign w30467 = w30045 ^ w30466 ;
  assign w30468 = ~w30050 & w30467 ;
  assign w30469 = w30465 | w30468 ;
  assign w30470 = ~\pi110 & w30469 ;
  assign w30471 = ( \pi110 & ~w30465 ) | ( \pi110 & w30468 ) | ( ~w30465 & w30468 ) ;
  assign w30472 = ~w30468 & w30471 ;
  assign w30473 = w30470 | w30472 ;
  assign w30474 = ( ~w30056 & w30464 ) | ( ~w30056 & w30473 ) | ( w30464 & w30473 ) ;
  assign w30475 = ( w11087 & ~w30473 ) | ( w11087 & w30474 ) | ( ~w30473 & w30474 ) ;
  assign w30476 = w30473 | w30475 ;
  assign w30477 = ~w10650 & w30469 ;
  assign w30478 = w30476 & ~w30477 ;
  assign w30479 = ~w30062 & w30461 ;
  assign w30480 = w30462 ^ w30479 ;
  assign w30481 = ~w30478 & w30480 ;
  assign w30482 = ( w30055 & w30476 ) | ( w30055 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30483 = ~w30477 & w30482 ;
  assign w30484 = w30481 | w30483 ;
  assign w30485 = ~\pi110 & w30484 ;
  assign w30486 = ~w30068 & w30458 ;
  assign w30487 = w30459 ^ w30486 ;
  assign w30488 = ~w30478 & w30487 ;
  assign w30489 = ( w30061 & w30476 ) | ( w30061 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30490 = ~w30477 & w30489 ;
  assign w30491 = w30488 | w30490 ;
  assign w30492 = ~\pi109 & w30491 ;
  assign w30493 = ~w30074 & w30455 ;
  assign w30494 = w30456 ^ w30493 ;
  assign w30495 = ~w30478 & w30494 ;
  assign w30496 = ( w30067 & w30476 ) | ( w30067 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30497 = ~w30477 & w30496 ;
  assign w30498 = w30495 | w30497 ;
  assign w30499 = ~\pi108 & w30498 ;
  assign w30500 = ~w30080 & w30452 ;
  assign w30501 = w30453 ^ w30500 ;
  assign w30502 = ~w30478 & w30501 ;
  assign w30503 = ( w30073 & w30476 ) | ( w30073 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30504 = ~w30477 & w30503 ;
  assign w30505 = w30502 | w30504 ;
  assign w30506 = ~\pi107 & w30505 ;
  assign w30507 = ~w30086 & w30449 ;
  assign w30508 = w30450 ^ w30507 ;
  assign w30509 = ~w30478 & w30508 ;
  assign w30510 = ( w30079 & w30476 ) | ( w30079 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30511 = ~w30477 & w30510 ;
  assign w30512 = w30509 | w30511 ;
  assign w30513 = ~\pi106 & w30512 ;
  assign w30514 = ~w30092 & w30446 ;
  assign w30515 = w30447 ^ w30514 ;
  assign w30516 = ~w30478 & w30515 ;
  assign w30517 = ( w30085 & w30476 ) | ( w30085 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30518 = ~w30477 & w30517 ;
  assign w30519 = w30516 | w30518 ;
  assign w30520 = ~\pi105 & w30519 ;
  assign w30521 = ~w30098 & w30443 ;
  assign w30522 = w30444 ^ w30521 ;
  assign w30523 = ~w30478 & w30522 ;
  assign w30524 = ( w30091 & w30476 ) | ( w30091 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30525 = ~w30477 & w30524 ;
  assign w30526 = w30523 | w30525 ;
  assign w30527 = ~\pi104 & w30526 ;
  assign w30528 = ~w30104 & w30440 ;
  assign w30529 = w30441 ^ w30528 ;
  assign w30530 = ~w30478 & w30529 ;
  assign w30531 = ( w30097 & w30476 ) | ( w30097 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30532 = ~w30477 & w30531 ;
  assign w30533 = w30530 | w30532 ;
  assign w30534 = ~\pi103 & w30533 ;
  assign w30535 = ~w30110 & w30437 ;
  assign w30536 = w30438 ^ w30535 ;
  assign w30537 = ~w30478 & w30536 ;
  assign w30538 = ( w30103 & w30476 ) | ( w30103 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30539 = ~w30477 & w30538 ;
  assign w30540 = w30537 | w30539 ;
  assign w30541 = ~\pi102 & w30540 ;
  assign w30542 = ~w30116 & w30434 ;
  assign w30543 = w30435 ^ w30542 ;
  assign w30544 = ~w30478 & w30543 ;
  assign w30545 = ( w30109 & w30476 ) | ( w30109 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30546 = ~w30477 & w30545 ;
  assign w30547 = w30544 | w30546 ;
  assign w30548 = ~\pi101 & w30547 ;
  assign w30549 = ~w30122 & w30431 ;
  assign w30550 = w30432 ^ w30549 ;
  assign w30551 = ~w30478 & w30550 ;
  assign w30552 = ( w30115 & w30476 ) | ( w30115 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30553 = ~w30477 & w30552 ;
  assign w30554 = w30551 | w30553 ;
  assign w30555 = ~\pi100 & w30554 ;
  assign w30556 = ~w30128 & w30428 ;
  assign w30557 = w30429 ^ w30556 ;
  assign w30558 = ~w30478 & w30557 ;
  assign w30559 = ( w30121 & w30476 ) | ( w30121 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30560 = ~w30477 & w30559 ;
  assign w30561 = w30558 | w30560 ;
  assign w30562 = ~\pi099 & w30561 ;
  assign w30563 = ~w30134 & w30425 ;
  assign w30564 = w30426 ^ w30563 ;
  assign w30565 = ~w30478 & w30564 ;
  assign w30566 = ( w30127 & w30476 ) | ( w30127 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30567 = ~w30477 & w30566 ;
  assign w30568 = w30565 | w30567 ;
  assign w30569 = ~\pi098 & w30568 ;
  assign w30570 = ~w30140 & w30422 ;
  assign w30571 = w30423 ^ w30570 ;
  assign w30572 = ~w30478 & w30571 ;
  assign w30573 = ( w30133 & w30476 ) | ( w30133 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30574 = ~w30477 & w30573 ;
  assign w30575 = w30572 | w30574 ;
  assign w30576 = ~\pi097 & w30575 ;
  assign w30577 = ~w30146 & w30419 ;
  assign w30578 = w30420 ^ w30577 ;
  assign w30579 = ~w30478 & w30578 ;
  assign w30580 = ( w30139 & w30476 ) | ( w30139 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30581 = ~w30477 & w30580 ;
  assign w30582 = w30579 | w30581 ;
  assign w30583 = ~\pi096 & w30582 ;
  assign w30584 = ~w30152 & w30416 ;
  assign w30585 = w30417 ^ w30584 ;
  assign w30586 = ~w30478 & w30585 ;
  assign w30587 = ( w30145 & w30476 ) | ( w30145 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30588 = ~w30477 & w30587 ;
  assign w30589 = w30586 | w30588 ;
  assign w30590 = ~\pi095 & w30589 ;
  assign w30591 = ~w30158 & w30413 ;
  assign w30592 = w30414 ^ w30591 ;
  assign w30593 = ~w30478 & w30592 ;
  assign w30594 = ( w30151 & w30476 ) | ( w30151 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30595 = ~w30477 & w30594 ;
  assign w30596 = w30593 | w30595 ;
  assign w30597 = ~\pi094 & w30596 ;
  assign w30598 = ~w30164 & w30410 ;
  assign w30599 = w30411 ^ w30598 ;
  assign w30600 = ~w30478 & w30599 ;
  assign w30601 = ( w30157 & w30476 ) | ( w30157 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30602 = ~w30477 & w30601 ;
  assign w30603 = w30600 | w30602 ;
  assign w30604 = ~\pi093 & w30603 ;
  assign w30605 = ~w30170 & w30407 ;
  assign w30606 = w30408 ^ w30605 ;
  assign w30607 = ~w30478 & w30606 ;
  assign w30608 = ( w30163 & w30476 ) | ( w30163 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30609 = ~w30477 & w30608 ;
  assign w30610 = w30607 | w30609 ;
  assign w30611 = ~\pi092 & w30610 ;
  assign w30612 = ~w30176 & w30404 ;
  assign w30613 = w30405 ^ w30612 ;
  assign w30614 = ~w30478 & w30613 ;
  assign w30615 = ( w30169 & w30476 ) | ( w30169 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30616 = ~w30477 & w30615 ;
  assign w30617 = w30614 | w30616 ;
  assign w30618 = ~\pi091 & w30617 ;
  assign w30619 = ~w30182 & w30401 ;
  assign w30620 = w30402 ^ w30619 ;
  assign w30621 = ~w30478 & w30620 ;
  assign w30622 = ( w30175 & w30476 ) | ( w30175 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30623 = ~w30477 & w30622 ;
  assign w30624 = w30621 | w30623 ;
  assign w30625 = ~\pi090 & w30624 ;
  assign w30626 = ~w30188 & w30398 ;
  assign w30627 = w30399 ^ w30626 ;
  assign w30628 = ~w30478 & w30627 ;
  assign w30629 = ( w30181 & w30476 ) | ( w30181 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30630 = ~w30477 & w30629 ;
  assign w30631 = w30628 | w30630 ;
  assign w30632 = ~\pi089 & w30631 ;
  assign w30633 = ~w30194 & w30395 ;
  assign w30634 = w30396 ^ w30633 ;
  assign w30635 = ~w30478 & w30634 ;
  assign w30636 = ( w30187 & w30476 ) | ( w30187 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30637 = ~w30477 & w30636 ;
  assign w30638 = w30635 | w30637 ;
  assign w30639 = ~\pi088 & w30638 ;
  assign w30640 = ~w30200 & w30392 ;
  assign w30641 = w30393 ^ w30640 ;
  assign w30642 = ~w30478 & w30641 ;
  assign w30643 = ( w30193 & w30476 ) | ( w30193 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30644 = ~w30477 & w30643 ;
  assign w30645 = w30642 | w30644 ;
  assign w30646 = ~\pi087 & w30645 ;
  assign w30647 = ~w30206 & w30389 ;
  assign w30648 = w30390 ^ w30647 ;
  assign w30649 = ~w30478 & w30648 ;
  assign w30650 = ( w30199 & w30476 ) | ( w30199 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30651 = ~w30477 & w30650 ;
  assign w30652 = w30649 | w30651 ;
  assign w30653 = ~\pi086 & w30652 ;
  assign w30654 = ~w30212 & w30386 ;
  assign w30655 = w30387 ^ w30654 ;
  assign w30656 = ~w30478 & w30655 ;
  assign w30657 = ( w30205 & w30476 ) | ( w30205 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30658 = ~w30477 & w30657 ;
  assign w30659 = w30656 | w30658 ;
  assign w30660 = ~\pi085 & w30659 ;
  assign w30661 = ~w30218 & w30383 ;
  assign w30662 = w30384 ^ w30661 ;
  assign w30663 = ~w30478 & w30662 ;
  assign w30664 = ( w30211 & w30476 ) | ( w30211 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30665 = ~w30477 & w30664 ;
  assign w30666 = w30663 | w30665 ;
  assign w30667 = ~\pi084 & w30666 ;
  assign w30668 = ~w30224 & w30380 ;
  assign w30669 = w30381 ^ w30668 ;
  assign w30670 = ~w30478 & w30669 ;
  assign w30671 = ( w30217 & w30476 ) | ( w30217 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30672 = ~w30477 & w30671 ;
  assign w30673 = w30670 | w30672 ;
  assign w30674 = ~\pi083 & w30673 ;
  assign w30675 = ~w30230 & w30377 ;
  assign w30676 = w30378 ^ w30675 ;
  assign w30677 = ~w30478 & w30676 ;
  assign w30678 = ( w30223 & w30476 ) | ( w30223 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30679 = ~w30477 & w30678 ;
  assign w30680 = w30677 | w30679 ;
  assign w30681 = ~\pi082 & w30680 ;
  assign w30682 = ~w30236 & w30374 ;
  assign w30683 = w30375 ^ w30682 ;
  assign w30684 = ~w30478 & w30683 ;
  assign w30685 = ( w30229 & w30476 ) | ( w30229 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30686 = ~w30477 & w30685 ;
  assign w30687 = w30684 | w30686 ;
  assign w30688 = ~\pi081 & w30687 ;
  assign w30689 = ~w30242 & w30371 ;
  assign w30690 = w30372 ^ w30689 ;
  assign w30691 = ~w30478 & w30690 ;
  assign w30692 = ( w30235 & w30476 ) | ( w30235 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30693 = ~w30477 & w30692 ;
  assign w30694 = w30691 | w30693 ;
  assign w30695 = ~\pi080 & w30694 ;
  assign w30696 = ~w30248 & w30368 ;
  assign w30697 = w30369 ^ w30696 ;
  assign w30698 = ~w30478 & w30697 ;
  assign w30699 = ( w30241 & w30476 ) | ( w30241 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30700 = ~w30477 & w30699 ;
  assign w30701 = w30698 | w30700 ;
  assign w30702 = ~\pi079 & w30701 ;
  assign w30703 = ~w30254 & w30365 ;
  assign w30704 = w30366 ^ w30703 ;
  assign w30705 = ~w30478 & w30704 ;
  assign w30706 = ( w30247 & w30476 ) | ( w30247 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30707 = ~w30477 & w30706 ;
  assign w30708 = w30705 | w30707 ;
  assign w30709 = ~\pi078 & w30708 ;
  assign w30710 = ~w30260 & w30362 ;
  assign w30711 = w30363 ^ w30710 ;
  assign w30712 = ~w30478 & w30711 ;
  assign w30713 = ( w30253 & w30476 ) | ( w30253 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30714 = ~w30477 & w30713 ;
  assign w30715 = w30712 | w30714 ;
  assign w30716 = ~\pi077 & w30715 ;
  assign w30717 = ~w30266 & w30359 ;
  assign w30718 = w30360 ^ w30717 ;
  assign w30719 = ~w30478 & w30718 ;
  assign w30720 = ( w30259 & w30476 ) | ( w30259 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30721 = ~w30477 & w30720 ;
  assign w30722 = w30719 | w30721 ;
  assign w30723 = ~\pi076 & w30722 ;
  assign w30724 = ~w30272 & w30356 ;
  assign w30725 = w30357 ^ w30724 ;
  assign w30726 = ~w30478 & w30725 ;
  assign w30727 = ( w30265 & w30476 ) | ( w30265 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30728 = ~w30477 & w30727 ;
  assign w30729 = w30726 | w30728 ;
  assign w30730 = ~\pi075 & w30729 ;
  assign w30731 = ~w30278 & w30353 ;
  assign w30732 = w30354 ^ w30731 ;
  assign w30733 = ~w30478 & w30732 ;
  assign w30734 = ( w30271 & w30476 ) | ( w30271 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30735 = ~w30477 & w30734 ;
  assign w30736 = w30733 | w30735 ;
  assign w30737 = ~\pi074 & w30736 ;
  assign w30738 = ~w30284 & w30350 ;
  assign w30739 = w30351 ^ w30738 ;
  assign w30740 = ~w30478 & w30739 ;
  assign w30741 = ( w30277 & w30476 ) | ( w30277 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30742 = ~w30477 & w30741 ;
  assign w30743 = w30740 | w30742 ;
  assign w30744 = ~\pi073 & w30743 ;
  assign w30745 = ~w30290 & w30347 ;
  assign w30746 = w30348 ^ w30745 ;
  assign w30747 = ~w30478 & w30746 ;
  assign w30748 = ( w30283 & w30476 ) | ( w30283 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30749 = ~w30477 & w30748 ;
  assign w30750 = w30747 | w30749 ;
  assign w30751 = ~\pi072 & w30750 ;
  assign w30752 = ~w30296 & w30344 ;
  assign w30753 = w30345 ^ w30752 ;
  assign w30754 = ~w30478 & w30753 ;
  assign w30755 = ( w30289 & w30476 ) | ( w30289 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30756 = ~w30477 & w30755 ;
  assign w30757 = w30754 | w30756 ;
  assign w30758 = ~\pi071 & w30757 ;
  assign w30759 = ~w30302 & w30341 ;
  assign w30760 = w30342 ^ w30759 ;
  assign w30761 = ~w30478 & w30760 ;
  assign w30762 = ( w30295 & w30476 ) | ( w30295 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30763 = ~w30477 & w30762 ;
  assign w30764 = w30761 | w30763 ;
  assign w30765 = ~\pi070 & w30764 ;
  assign w30766 = ~w30311 & w30338 ;
  assign w30767 = w30339 ^ w30766 ;
  assign w30768 = ~w30478 & w30767 ;
  assign w30769 = ( w30301 & w30476 ) | ( w30301 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30770 = ~w30477 & w30769 ;
  assign w30771 = w30768 | w30770 ;
  assign w30772 = ~\pi069 & w30771 ;
  assign w30773 = ~w30321 & w30333 ;
  assign w30774 = w30336 ^ w30773 ;
  assign w30775 = ~w30478 & w30774 ;
  assign w30776 = ( w30310 & w30476 ) | ( w30310 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30777 = ~w30477 & w30776 ;
  assign w30778 = w30775 | w30777 ;
  assign w30779 = ~\pi068 & w30778 ;
  assign w30780 = ( \pi065 & w30325 ) | ( \pi065 & ~w30478 ) | ( w30325 & ~w30478 ) ;
  assign w30781 = ( \pi065 & w30327 ) | ( \pi065 & ~w30780 ) | ( w30327 & ~w30780 ) ;
  assign w30782 = w30330 ^ w30781 ;
  assign w30783 = ~w30478 & w30782 ;
  assign w30784 = ( w30320 & w30476 ) | ( w30320 & w30477 ) | ( w30476 & w30477 ) ;
  assign w30785 = ~w30477 & w30784 ;
  assign w30786 = w30783 | w30785 ;
  assign w30787 = ~\pi067 & w30786 ;
  assign w30788 = w10937 ^ w30325 ;
  assign w30789 = \pi065 ^ w30788 ;
  assign w30790 = w30478 ^ w30789 ;
  assign w30791 = ( w30325 & w30789 ) | ( w30325 & w30790 ) | ( w30789 & w30790 ) ;
  assign w30792 = ~\pi066 & w30791 ;
  assign w30793 = w30325 ^ w30478 ;
  assign w30794 = ( w30325 & w30789 ) | ( w30325 & ~w30793 ) | ( w30789 & ~w30793 ) ;
  assign w30795 = \pi066 ^ w30794 ;
  assign w30796 = ( \pi064 & ~w30478 ) | ( \pi064 & w30795 ) | ( ~w30478 & w30795 ) ;
  assign w30797 = \pi017 ^ w30796 ;
  assign w30798 = ( \pi065 & w11877 ) | ( \pi065 & ~w30797 ) | ( w11877 & ~w30797 ) ;
  assign w30799 = w30795 | w30798 ;
  assign w30800 = \pi067 ^ w30786 ;
  assign w30801 = ( ~w30792 & w30799 ) | ( ~w30792 & w30800 ) | ( w30799 & w30800 ) ;
  assign w30802 = w30800 | w30801 ;
  assign w30803 = \pi068 ^ w30778 ;
  assign w30804 = ( ~w30787 & w30802 ) | ( ~w30787 & w30803 ) | ( w30802 & w30803 ) ;
  assign w30805 = w30803 | w30804 ;
  assign w30806 = \pi069 ^ w30771 ;
  assign w30807 = ( ~w30779 & w30805 ) | ( ~w30779 & w30806 ) | ( w30805 & w30806 ) ;
  assign w30808 = w30806 | w30807 ;
  assign w30809 = \pi070 ^ w30764 ;
  assign w30810 = ( ~w30772 & w30808 ) | ( ~w30772 & w30809 ) | ( w30808 & w30809 ) ;
  assign w30811 = w30809 | w30810 ;
  assign w30812 = \pi071 ^ w30757 ;
  assign w30813 = ( ~w30765 & w30811 ) | ( ~w30765 & w30812 ) | ( w30811 & w30812 ) ;
  assign w30814 = w30812 | w30813 ;
  assign w30815 = \pi072 ^ w30750 ;
  assign w30816 = ( ~w30758 & w30814 ) | ( ~w30758 & w30815 ) | ( w30814 & w30815 ) ;
  assign w30817 = w30815 | w30816 ;
  assign w30818 = \pi073 ^ w30743 ;
  assign w30819 = ( ~w30751 & w30817 ) | ( ~w30751 & w30818 ) | ( w30817 & w30818 ) ;
  assign w30820 = w30818 | w30819 ;
  assign w30821 = \pi074 ^ w30736 ;
  assign w30822 = ( ~w30744 & w30820 ) | ( ~w30744 & w30821 ) | ( w30820 & w30821 ) ;
  assign w30823 = w30821 | w30822 ;
  assign w30824 = \pi075 ^ w30729 ;
  assign w30825 = ( ~w30737 & w30823 ) | ( ~w30737 & w30824 ) | ( w30823 & w30824 ) ;
  assign w30826 = w30824 | w30825 ;
  assign w30827 = \pi076 ^ w30722 ;
  assign w30828 = ( ~w30730 & w30826 ) | ( ~w30730 & w30827 ) | ( w30826 & w30827 ) ;
  assign w30829 = w30827 | w30828 ;
  assign w30830 = \pi077 ^ w30715 ;
  assign w30831 = ( ~w30723 & w30829 ) | ( ~w30723 & w30830 ) | ( w30829 & w30830 ) ;
  assign w30832 = w30830 | w30831 ;
  assign w30833 = \pi078 ^ w30708 ;
  assign w30834 = ( ~w30716 & w30832 ) | ( ~w30716 & w30833 ) | ( w30832 & w30833 ) ;
  assign w30835 = w30833 | w30834 ;
  assign w30836 = \pi079 ^ w30701 ;
  assign w30837 = ( ~w30709 & w30835 ) | ( ~w30709 & w30836 ) | ( w30835 & w30836 ) ;
  assign w30838 = w30836 | w30837 ;
  assign w30839 = \pi080 ^ w30694 ;
  assign w30840 = ( ~w30702 & w30838 ) | ( ~w30702 & w30839 ) | ( w30838 & w30839 ) ;
  assign w30841 = w30839 | w30840 ;
  assign w30842 = \pi081 ^ w30687 ;
  assign w30843 = ( ~w30695 & w30841 ) | ( ~w30695 & w30842 ) | ( w30841 & w30842 ) ;
  assign w30844 = w30842 | w30843 ;
  assign w30845 = \pi082 ^ w30680 ;
  assign w30846 = ( ~w30688 & w30844 ) | ( ~w30688 & w30845 ) | ( w30844 & w30845 ) ;
  assign w30847 = w30845 | w30846 ;
  assign w30848 = \pi083 ^ w30673 ;
  assign w30849 = ( ~w30681 & w30847 ) | ( ~w30681 & w30848 ) | ( w30847 & w30848 ) ;
  assign w30850 = w30848 | w30849 ;
  assign w30851 = \pi084 ^ w30666 ;
  assign w30852 = ( ~w30674 & w30850 ) | ( ~w30674 & w30851 ) | ( w30850 & w30851 ) ;
  assign w30853 = w30851 | w30852 ;
  assign w30854 = \pi085 ^ w30659 ;
  assign w30855 = ( ~w30667 & w30853 ) | ( ~w30667 & w30854 ) | ( w30853 & w30854 ) ;
  assign w30856 = w30854 | w30855 ;
  assign w30857 = \pi086 ^ w30652 ;
  assign w30858 = ( ~w30660 & w30856 ) | ( ~w30660 & w30857 ) | ( w30856 & w30857 ) ;
  assign w30859 = w30857 | w30858 ;
  assign w30860 = \pi087 ^ w30645 ;
  assign w30861 = ( ~w30653 & w30859 ) | ( ~w30653 & w30860 ) | ( w30859 & w30860 ) ;
  assign w30862 = w30860 | w30861 ;
  assign w30863 = \pi088 ^ w30638 ;
  assign w30864 = ( ~w30646 & w30862 ) | ( ~w30646 & w30863 ) | ( w30862 & w30863 ) ;
  assign w30865 = w30863 | w30864 ;
  assign w30866 = \pi089 ^ w30631 ;
  assign w30867 = ( ~w30639 & w30865 ) | ( ~w30639 & w30866 ) | ( w30865 & w30866 ) ;
  assign w30868 = w30866 | w30867 ;
  assign w30869 = \pi090 ^ w30624 ;
  assign w30870 = ( ~w30632 & w30868 ) | ( ~w30632 & w30869 ) | ( w30868 & w30869 ) ;
  assign w30871 = w30869 | w30870 ;
  assign w30872 = \pi091 ^ w30617 ;
  assign w30873 = ( ~w30625 & w30871 ) | ( ~w30625 & w30872 ) | ( w30871 & w30872 ) ;
  assign w30874 = w30872 | w30873 ;
  assign w30875 = \pi092 ^ w30610 ;
  assign w30876 = ( ~w30618 & w30874 ) | ( ~w30618 & w30875 ) | ( w30874 & w30875 ) ;
  assign w30877 = w30875 | w30876 ;
  assign w30878 = \pi093 ^ w30603 ;
  assign w30879 = ( ~w30611 & w30877 ) | ( ~w30611 & w30878 ) | ( w30877 & w30878 ) ;
  assign w30880 = w30878 | w30879 ;
  assign w30881 = \pi094 ^ w30596 ;
  assign w30882 = ( ~w30604 & w30880 ) | ( ~w30604 & w30881 ) | ( w30880 & w30881 ) ;
  assign w30883 = w30881 | w30882 ;
  assign w30884 = \pi095 ^ w30589 ;
  assign w30885 = ( ~w30597 & w30883 ) | ( ~w30597 & w30884 ) | ( w30883 & w30884 ) ;
  assign w30886 = w30884 | w30885 ;
  assign w30887 = \pi096 ^ w30582 ;
  assign w30888 = ( ~w30590 & w30886 ) | ( ~w30590 & w30887 ) | ( w30886 & w30887 ) ;
  assign w30889 = w30887 | w30888 ;
  assign w30890 = \pi097 ^ w30575 ;
  assign w30891 = ( ~w30583 & w30889 ) | ( ~w30583 & w30890 ) | ( w30889 & w30890 ) ;
  assign w30892 = w30890 | w30891 ;
  assign w30893 = \pi098 ^ w30568 ;
  assign w30894 = ( ~w30576 & w30892 ) | ( ~w30576 & w30893 ) | ( w30892 & w30893 ) ;
  assign w30895 = w30893 | w30894 ;
  assign w30896 = \pi099 ^ w30561 ;
  assign w30897 = ( ~w30569 & w30895 ) | ( ~w30569 & w30896 ) | ( w30895 & w30896 ) ;
  assign w30898 = w30896 | w30897 ;
  assign w30899 = \pi100 ^ w30554 ;
  assign w30900 = ( ~w30562 & w30898 ) | ( ~w30562 & w30899 ) | ( w30898 & w30899 ) ;
  assign w30901 = w30899 | w30900 ;
  assign w30902 = \pi101 ^ w30547 ;
  assign w30903 = ( ~w30555 & w30901 ) | ( ~w30555 & w30902 ) | ( w30901 & w30902 ) ;
  assign w30904 = w30902 | w30903 ;
  assign w30905 = \pi102 ^ w30540 ;
  assign w30906 = ( ~w30548 & w30904 ) | ( ~w30548 & w30905 ) | ( w30904 & w30905 ) ;
  assign w30907 = w30905 | w30906 ;
  assign w30908 = \pi103 ^ w30533 ;
  assign w30909 = ( ~w30541 & w30907 ) | ( ~w30541 & w30908 ) | ( w30907 & w30908 ) ;
  assign w30910 = w30908 | w30909 ;
  assign w30911 = \pi104 ^ w30526 ;
  assign w30912 = ( ~w30534 & w30910 ) | ( ~w30534 & w30911 ) | ( w30910 & w30911 ) ;
  assign w30913 = w30911 | w30912 ;
  assign w30914 = \pi105 ^ w30519 ;
  assign w30915 = ( ~w30527 & w30913 ) | ( ~w30527 & w30914 ) | ( w30913 & w30914 ) ;
  assign w30916 = w30914 | w30915 ;
  assign w30917 = \pi106 ^ w30512 ;
  assign w30918 = ( ~w30520 & w30916 ) | ( ~w30520 & w30917 ) | ( w30916 & w30917 ) ;
  assign w30919 = w30917 | w30918 ;
  assign w30920 = \pi107 ^ w30505 ;
  assign w30921 = ( ~w30513 & w30919 ) | ( ~w30513 & w30920 ) | ( w30919 & w30920 ) ;
  assign w30922 = w30920 | w30921 ;
  assign w30923 = \pi108 ^ w30498 ;
  assign w30924 = ( ~w30506 & w30922 ) | ( ~w30506 & w30923 ) | ( w30922 & w30923 ) ;
  assign w30925 = w30923 | w30924 ;
  assign w30926 = \pi109 ^ w30491 ;
  assign w30927 = ( ~w30499 & w30925 ) | ( ~w30499 & w30926 ) | ( w30925 & w30926 ) ;
  assign w30928 = w30926 | w30927 ;
  assign w30929 = \pi110 ^ w30484 ;
  assign w30930 = ( ~w30492 & w30928 ) | ( ~w30492 & w30929 ) | ( w30928 & w30929 ) ;
  assign w30931 = w30929 | w30930 ;
  assign w30932 = ( ~w30056 & w30464 ) | ( ~w30056 & w30478 ) | ( w30464 & w30478 ) ;
  assign w30933 = w30473 ^ w30932 ;
  assign w30934 = ~w30478 & w30933 ;
  assign w30935 = ( w10650 & ~w30469 ) | ( w10650 & w30476 ) | ( ~w30469 & w30476 ) ;
  assign w30936 = w30469 & w30935 ;
  assign w30937 = w30934 | w30936 ;
  assign w30938 = ~\pi111 & w30937 ;
  assign w30939 = ( \pi111 & ~w30934 ) | ( \pi111 & w30936 ) | ( ~w30934 & w30936 ) ;
  assign w30940 = ~w30936 & w30939 ;
  assign w30941 = w30938 | w30940 ;
  assign w30942 = ( ~w30485 & w30931 ) | ( ~w30485 & w30941 ) | ( w30931 & w30941 ) ;
  assign w30943 = ( w201 & ~w30941 ) | ( w201 & w30942 ) | ( ~w30941 & w30942 ) ;
  assign w30944 = w30941 | w30943 ;
  assign w30945 = ~w11087 & w30937 ;
  assign w30946 = w30944 & ~w30945 ;
  assign w30947 = ~w30492 & w30928 ;
  assign w30948 = w30929 ^ w30947 ;
  assign w30949 = ~w30946 & w30948 ;
  assign w30950 = ( w30484 & w30944 ) | ( w30484 & w30945 ) | ( w30944 & w30945 ) ;
  assign w30951 = ~w30945 & w30950 ;
  assign w30952 = w30949 | w30951 ;
  assign w30953 = ( ~w30485 & w30931 ) | ( ~w30485 & w30946 ) | ( w30931 & w30946 ) ;
  assign w30954 = w30941 ^ w30953 ;
  assign w30955 = ~w30946 & w30954 ;
  assign w30956 = ( w11087 & ~w30937 ) | ( w11087 & w30944 ) | ( ~w30937 & w30944 ) ;
  assign w30957 = w30937 & w30956 ;
  assign w30958 = w30955 | w30957 ;
  assign w30959 = ~\pi111 & w30952 ;
  assign w30960 = ~w30499 & w30925 ;
  assign w30961 = w30926 ^ w30960 ;
  assign w30962 = ~w30946 & w30961 ;
  assign w30963 = ( w30491 & w30944 ) | ( w30491 & w30945 ) | ( w30944 & w30945 ) ;
  assign w30964 = ~w30945 & w30963 ;
  assign w30965 = w30962 | w30964 ;
  assign w30966 = ~\pi110 & w30965 ;
  assign w30967 = ~w30506 & w30922 ;
  assign w30968 = w30923 ^ w30967 ;
  assign w30969 = ~w30946 & w30968 ;
  assign w30970 = ( w30498 & w30944 ) | ( w30498 & w30945 ) | ( w30944 & w30945 ) ;
  assign w30971 = ~w30945 & w30970 ;
  assign w30972 = w30969 | w30971 ;
  assign w30973 = ~\pi109 & w30972 ;
  assign w30974 = ~w30513 & w30919 ;
  assign w30975 = w30920 ^ w30974 ;
  assign w30976 = ~w30946 & w30975 ;
  assign w30977 = ( w30505 & w30944 ) | ( w30505 & w30945 ) | ( w30944 & w30945 ) ;
  assign w30978 = ~w30945 & w30977 ;
  assign w30979 = w30976 | w30978 ;
  assign w30980 = ~\pi108 & w30979 ;
  assign w30981 = ~w30520 & w30916 ;
  assign w30982 = w30917 ^ w30981 ;
  assign w30983 = ~w30946 & w30982 ;
  assign w30984 = ( w30512 & w30944 ) | ( w30512 & w30945 ) | ( w30944 & w30945 ) ;
  assign w30985 = ~w30945 & w30984 ;
  assign w30986 = w30983 | w30985 ;
  assign w30987 = ~\pi107 & w30986 ;
  assign w30988 = ~w30527 & w30913 ;
  assign w30989 = w30914 ^ w30988 ;
  assign w30990 = ~w30946 & w30989 ;
  assign w30991 = ( w30519 & w30944 ) | ( w30519 & w30945 ) | ( w30944 & w30945 ) ;
  assign w30992 = ~w30945 & w30991 ;
  assign w30993 = w30990 | w30992 ;
  assign w30994 = ~\pi106 & w30993 ;
  assign w30995 = ~w30534 & w30910 ;
  assign w30996 = w30911 ^ w30995 ;
  assign w30997 = ~w30946 & w30996 ;
  assign w30998 = ( w30526 & w30944 ) | ( w30526 & w30945 ) | ( w30944 & w30945 ) ;
  assign w30999 = ~w30945 & w30998 ;
  assign w31000 = w30997 | w30999 ;
  assign w31001 = ~\pi105 & w31000 ;
  assign w31002 = ~w30541 & w30907 ;
  assign w31003 = w30908 ^ w31002 ;
  assign w31004 = ~w30946 & w31003 ;
  assign w31005 = ( w30533 & w30944 ) | ( w30533 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31006 = ~w30945 & w31005 ;
  assign w31007 = w31004 | w31006 ;
  assign w31008 = ~\pi104 & w31007 ;
  assign w31009 = ~w30548 & w30904 ;
  assign w31010 = w30905 ^ w31009 ;
  assign w31011 = ~w30946 & w31010 ;
  assign w31012 = ( w30540 & w30944 ) | ( w30540 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31013 = ~w30945 & w31012 ;
  assign w31014 = w31011 | w31013 ;
  assign w31015 = ~\pi103 & w31014 ;
  assign w31016 = ~w30555 & w30901 ;
  assign w31017 = w30902 ^ w31016 ;
  assign w31018 = ~w30946 & w31017 ;
  assign w31019 = ( w30547 & w30944 ) | ( w30547 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31020 = ~w30945 & w31019 ;
  assign w31021 = w31018 | w31020 ;
  assign w31022 = ~\pi102 & w31021 ;
  assign w31023 = ~w30562 & w30898 ;
  assign w31024 = w30899 ^ w31023 ;
  assign w31025 = ~w30946 & w31024 ;
  assign w31026 = ( w30554 & w30944 ) | ( w30554 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31027 = ~w30945 & w31026 ;
  assign w31028 = w31025 | w31027 ;
  assign w31029 = ~\pi101 & w31028 ;
  assign w31030 = ~w30569 & w30895 ;
  assign w31031 = w30896 ^ w31030 ;
  assign w31032 = ~w30946 & w31031 ;
  assign w31033 = ( w30561 & w30944 ) | ( w30561 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31034 = ~w30945 & w31033 ;
  assign w31035 = w31032 | w31034 ;
  assign w31036 = ~\pi100 & w31035 ;
  assign w31037 = ~w30576 & w30892 ;
  assign w31038 = w30893 ^ w31037 ;
  assign w31039 = ~w30946 & w31038 ;
  assign w31040 = ( w30568 & w30944 ) | ( w30568 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31041 = ~w30945 & w31040 ;
  assign w31042 = w31039 | w31041 ;
  assign w31043 = ~\pi099 & w31042 ;
  assign w31044 = ~w30583 & w30889 ;
  assign w31045 = w30890 ^ w31044 ;
  assign w31046 = ~w30946 & w31045 ;
  assign w31047 = ( w30575 & w30944 ) | ( w30575 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31048 = ~w30945 & w31047 ;
  assign w31049 = w31046 | w31048 ;
  assign w31050 = ~\pi098 & w31049 ;
  assign w31051 = ~w30590 & w30886 ;
  assign w31052 = w30887 ^ w31051 ;
  assign w31053 = ~w30946 & w31052 ;
  assign w31054 = ( w30582 & w30944 ) | ( w30582 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31055 = ~w30945 & w31054 ;
  assign w31056 = w31053 | w31055 ;
  assign w31057 = ~\pi097 & w31056 ;
  assign w31058 = ~w30597 & w30883 ;
  assign w31059 = w30884 ^ w31058 ;
  assign w31060 = ~w30946 & w31059 ;
  assign w31061 = ( w30589 & w30944 ) | ( w30589 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31062 = ~w30945 & w31061 ;
  assign w31063 = w31060 | w31062 ;
  assign w31064 = ~\pi096 & w31063 ;
  assign w31065 = ~w30604 & w30880 ;
  assign w31066 = w30881 ^ w31065 ;
  assign w31067 = ~w30946 & w31066 ;
  assign w31068 = ( w30596 & w30944 ) | ( w30596 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31069 = ~w30945 & w31068 ;
  assign w31070 = w31067 | w31069 ;
  assign w31071 = ~\pi095 & w31070 ;
  assign w31072 = ~w30611 & w30877 ;
  assign w31073 = w30878 ^ w31072 ;
  assign w31074 = ~w30946 & w31073 ;
  assign w31075 = ( w30603 & w30944 ) | ( w30603 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31076 = ~w30945 & w31075 ;
  assign w31077 = w31074 | w31076 ;
  assign w31078 = ~\pi094 & w31077 ;
  assign w31079 = ~w30618 & w30874 ;
  assign w31080 = w30875 ^ w31079 ;
  assign w31081 = ~w30946 & w31080 ;
  assign w31082 = ( w30610 & w30944 ) | ( w30610 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31083 = ~w30945 & w31082 ;
  assign w31084 = w31081 | w31083 ;
  assign w31085 = ~\pi093 & w31084 ;
  assign w31086 = ~w30625 & w30871 ;
  assign w31087 = w30872 ^ w31086 ;
  assign w31088 = ~w30946 & w31087 ;
  assign w31089 = ( w30617 & w30944 ) | ( w30617 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31090 = ~w30945 & w31089 ;
  assign w31091 = w31088 | w31090 ;
  assign w31092 = ~\pi092 & w31091 ;
  assign w31093 = ~w30632 & w30868 ;
  assign w31094 = w30869 ^ w31093 ;
  assign w31095 = ~w30946 & w31094 ;
  assign w31096 = ( w30624 & w30944 ) | ( w30624 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31097 = ~w30945 & w31096 ;
  assign w31098 = w31095 | w31097 ;
  assign w31099 = ~\pi091 & w31098 ;
  assign w31100 = ~w30639 & w30865 ;
  assign w31101 = w30866 ^ w31100 ;
  assign w31102 = ~w30946 & w31101 ;
  assign w31103 = ( w30631 & w30944 ) | ( w30631 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31104 = ~w30945 & w31103 ;
  assign w31105 = w31102 | w31104 ;
  assign w31106 = ~\pi090 & w31105 ;
  assign w31107 = ~w30646 & w30862 ;
  assign w31108 = w30863 ^ w31107 ;
  assign w31109 = ~w30946 & w31108 ;
  assign w31110 = ( w30638 & w30944 ) | ( w30638 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31111 = ~w30945 & w31110 ;
  assign w31112 = w31109 | w31111 ;
  assign w31113 = ~\pi089 & w31112 ;
  assign w31114 = ~w30653 & w30859 ;
  assign w31115 = w30860 ^ w31114 ;
  assign w31116 = ~w30946 & w31115 ;
  assign w31117 = ( w30645 & w30944 ) | ( w30645 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31118 = ~w30945 & w31117 ;
  assign w31119 = w31116 | w31118 ;
  assign w31120 = ~\pi088 & w31119 ;
  assign w31121 = ~w30660 & w30856 ;
  assign w31122 = w30857 ^ w31121 ;
  assign w31123 = ~w30946 & w31122 ;
  assign w31124 = ( w30652 & w30944 ) | ( w30652 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31125 = ~w30945 & w31124 ;
  assign w31126 = w31123 | w31125 ;
  assign w31127 = ~\pi087 & w31126 ;
  assign w31128 = ~w30667 & w30853 ;
  assign w31129 = w30854 ^ w31128 ;
  assign w31130 = ~w30946 & w31129 ;
  assign w31131 = ( w30659 & w30944 ) | ( w30659 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31132 = ~w30945 & w31131 ;
  assign w31133 = w31130 | w31132 ;
  assign w31134 = ~\pi086 & w31133 ;
  assign w31135 = ~w30674 & w30850 ;
  assign w31136 = w30851 ^ w31135 ;
  assign w31137 = ~w30946 & w31136 ;
  assign w31138 = ( w30666 & w30944 ) | ( w30666 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31139 = ~w30945 & w31138 ;
  assign w31140 = w31137 | w31139 ;
  assign w31141 = ~\pi085 & w31140 ;
  assign w31142 = ~w30681 & w30847 ;
  assign w31143 = w30848 ^ w31142 ;
  assign w31144 = ~w30946 & w31143 ;
  assign w31145 = ( w30673 & w30944 ) | ( w30673 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31146 = ~w30945 & w31145 ;
  assign w31147 = w31144 | w31146 ;
  assign w31148 = ~\pi084 & w31147 ;
  assign w31149 = ~w30688 & w30844 ;
  assign w31150 = w30845 ^ w31149 ;
  assign w31151 = ~w30946 & w31150 ;
  assign w31152 = ( w30680 & w30944 ) | ( w30680 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31153 = ~w30945 & w31152 ;
  assign w31154 = w31151 | w31153 ;
  assign w31155 = ~\pi083 & w31154 ;
  assign w31156 = ~w30695 & w30841 ;
  assign w31157 = w30842 ^ w31156 ;
  assign w31158 = ~w30946 & w31157 ;
  assign w31159 = ( w30687 & w30944 ) | ( w30687 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31160 = ~w30945 & w31159 ;
  assign w31161 = w31158 | w31160 ;
  assign w31162 = ~\pi082 & w31161 ;
  assign w31163 = ~w30702 & w30838 ;
  assign w31164 = w30839 ^ w31163 ;
  assign w31165 = ~w30946 & w31164 ;
  assign w31166 = ( w30694 & w30944 ) | ( w30694 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31167 = ~w30945 & w31166 ;
  assign w31168 = w31165 | w31167 ;
  assign w31169 = ~\pi081 & w31168 ;
  assign w31170 = ~w30709 & w30835 ;
  assign w31171 = w30836 ^ w31170 ;
  assign w31172 = ~w30946 & w31171 ;
  assign w31173 = ( w30701 & w30944 ) | ( w30701 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31174 = ~w30945 & w31173 ;
  assign w31175 = w31172 | w31174 ;
  assign w31176 = ~\pi080 & w31175 ;
  assign w31177 = ~w30716 & w30832 ;
  assign w31178 = w30833 ^ w31177 ;
  assign w31179 = ~w30946 & w31178 ;
  assign w31180 = ( w30708 & w30944 ) | ( w30708 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31181 = ~w30945 & w31180 ;
  assign w31182 = w31179 | w31181 ;
  assign w31183 = ~\pi079 & w31182 ;
  assign w31184 = ~w30723 & w30829 ;
  assign w31185 = w30830 ^ w31184 ;
  assign w31186 = ~w30946 & w31185 ;
  assign w31187 = ( w30715 & w30944 ) | ( w30715 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31188 = ~w30945 & w31187 ;
  assign w31189 = w31186 | w31188 ;
  assign w31190 = ~\pi078 & w31189 ;
  assign w31191 = ~w30730 & w30826 ;
  assign w31192 = w30827 ^ w31191 ;
  assign w31193 = ~w30946 & w31192 ;
  assign w31194 = ( w30722 & w30944 ) | ( w30722 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31195 = ~w30945 & w31194 ;
  assign w31196 = w31193 | w31195 ;
  assign w31197 = ~\pi077 & w31196 ;
  assign w31198 = ~w30737 & w30823 ;
  assign w31199 = w30824 ^ w31198 ;
  assign w31200 = ~w30946 & w31199 ;
  assign w31201 = ( w30729 & w30944 ) | ( w30729 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31202 = ~w30945 & w31201 ;
  assign w31203 = w31200 | w31202 ;
  assign w31204 = ~\pi076 & w31203 ;
  assign w31205 = ~w30744 & w30820 ;
  assign w31206 = w30821 ^ w31205 ;
  assign w31207 = ~w30946 & w31206 ;
  assign w31208 = ( w30736 & w30944 ) | ( w30736 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31209 = ~w30945 & w31208 ;
  assign w31210 = w31207 | w31209 ;
  assign w31211 = ~\pi075 & w31210 ;
  assign w31212 = ~w30751 & w30817 ;
  assign w31213 = w30818 ^ w31212 ;
  assign w31214 = ~w30946 & w31213 ;
  assign w31215 = ( w30743 & w30944 ) | ( w30743 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31216 = ~w30945 & w31215 ;
  assign w31217 = w31214 | w31216 ;
  assign w31218 = ~\pi074 & w31217 ;
  assign w31219 = ~w30758 & w30814 ;
  assign w31220 = w30815 ^ w31219 ;
  assign w31221 = ~w30946 & w31220 ;
  assign w31222 = ( w30750 & w30944 ) | ( w30750 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31223 = ~w30945 & w31222 ;
  assign w31224 = w31221 | w31223 ;
  assign w31225 = ~\pi073 & w31224 ;
  assign w31226 = ~w30765 & w30811 ;
  assign w31227 = w30812 ^ w31226 ;
  assign w31228 = ~w30946 & w31227 ;
  assign w31229 = ( w30757 & w30944 ) | ( w30757 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31230 = ~w30945 & w31229 ;
  assign w31231 = w31228 | w31230 ;
  assign w31232 = ~\pi072 & w31231 ;
  assign w31233 = ~w30772 & w30808 ;
  assign w31234 = w30809 ^ w31233 ;
  assign w31235 = ~w30946 & w31234 ;
  assign w31236 = ( w30764 & w30944 ) | ( w30764 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31237 = ~w30945 & w31236 ;
  assign w31238 = w31235 | w31237 ;
  assign w31239 = ~\pi071 & w31238 ;
  assign w31240 = ~w30779 & w30805 ;
  assign w31241 = w30806 ^ w31240 ;
  assign w31242 = ~w30946 & w31241 ;
  assign w31243 = ( w30771 & w30944 ) | ( w30771 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31244 = ~w30945 & w31243 ;
  assign w31245 = w31242 | w31244 ;
  assign w31246 = ~\pi070 & w31245 ;
  assign w31247 = ~w30787 & w30802 ;
  assign w31248 = w30803 ^ w31247 ;
  assign w31249 = ~w30946 & w31248 ;
  assign w31250 = ( w30778 & w30944 ) | ( w30778 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31251 = ~w30945 & w31250 ;
  assign w31252 = w31249 | w31251 ;
  assign w31253 = ~\pi069 & w31252 ;
  assign w31254 = ~w30792 & w30799 ;
  assign w31255 = w30800 ^ w31254 ;
  assign w31256 = ~w30946 & w31255 ;
  assign w31257 = ( w30786 & w30944 ) | ( w30786 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31258 = ~w30945 & w31257 ;
  assign w31259 = w31256 | w31258 ;
  assign w31260 = ~\pi068 & w31259 ;
  assign w31261 = \pi064 & ~w30478 ;
  assign w31262 = \pi017 ^ w31261 ;
  assign w31263 = ( \pi065 & w11877 ) | ( \pi065 & ~w31262 ) | ( w11877 & ~w31262 ) ;
  assign w31264 = w30795 ^ w31263 ;
  assign w31265 = ~w30946 & w31264 ;
  assign w31266 = ( w30791 & w30944 ) | ( w30791 & w30945 ) | ( w30944 & w30945 ) ;
  assign w31267 = ~w30945 & w31266 ;
  assign w31268 = w31265 | w31267 ;
  assign w31269 = ~\pi067 & w31268 ;
  assign w31270 = \pi016 ^ w30478 ;
  assign w31271 = ( \pi064 & w30946 ) | ( \pi064 & w31270 ) | ( w30946 & w31270 ) ;
  assign w31272 = w11885 ^ w31271 ;
  assign w31273 = ~w30946 & w31272 ;
  assign w31274 = w30946 & w31262 ;
  assign w31275 = w31273 | w31274 ;
  assign w31276 = ~\pi066 & w31275 ;
  assign w31277 = \pi066 ^ w31275 ;
  assign w31278 = ( \pi064 & ~w30946 ) | ( \pi064 & w31277 ) | ( ~w30946 & w31277 ) ;
  assign w31279 = \pi016 ^ w31278 ;
  assign w31280 = ( \pi065 & w12310 ) | ( \pi065 & ~w31279 ) | ( w12310 & ~w31279 ) ;
  assign w31281 = w31277 | w31280 ;
  assign w31282 = \pi067 ^ w31268 ;
  assign w31283 = ( ~w31276 & w31281 ) | ( ~w31276 & w31282 ) | ( w31281 & w31282 ) ;
  assign w31284 = w31282 | w31283 ;
  assign w31285 = \pi068 ^ w31259 ;
  assign w31286 = ( ~w31269 & w31284 ) | ( ~w31269 & w31285 ) | ( w31284 & w31285 ) ;
  assign w31287 = w31285 | w31286 ;
  assign w31288 = \pi069 ^ w31252 ;
  assign w31289 = ( ~w31260 & w31287 ) | ( ~w31260 & w31288 ) | ( w31287 & w31288 ) ;
  assign w31290 = w31288 | w31289 ;
  assign w31291 = \pi070 ^ w31245 ;
  assign w31292 = ( ~w31253 & w31290 ) | ( ~w31253 & w31291 ) | ( w31290 & w31291 ) ;
  assign w31293 = w31291 | w31292 ;
  assign w31294 = \pi071 ^ w31238 ;
  assign w31295 = ( ~w31246 & w31293 ) | ( ~w31246 & w31294 ) | ( w31293 & w31294 ) ;
  assign w31296 = w31294 | w31295 ;
  assign w31297 = \pi072 ^ w31231 ;
  assign w31298 = ( ~w31239 & w31296 ) | ( ~w31239 & w31297 ) | ( w31296 & w31297 ) ;
  assign w31299 = w31297 | w31298 ;
  assign w31300 = \pi073 ^ w31224 ;
  assign w31301 = ( ~w31232 & w31299 ) | ( ~w31232 & w31300 ) | ( w31299 & w31300 ) ;
  assign w31302 = w31300 | w31301 ;
  assign w31303 = \pi074 ^ w31217 ;
  assign w31304 = ( ~w31225 & w31302 ) | ( ~w31225 & w31303 ) | ( w31302 & w31303 ) ;
  assign w31305 = w31303 | w31304 ;
  assign w31306 = \pi075 ^ w31210 ;
  assign w31307 = ( ~w31218 & w31305 ) | ( ~w31218 & w31306 ) | ( w31305 & w31306 ) ;
  assign w31308 = w31306 | w31307 ;
  assign w31309 = \pi076 ^ w31203 ;
  assign w31310 = ( ~w31211 & w31308 ) | ( ~w31211 & w31309 ) | ( w31308 & w31309 ) ;
  assign w31311 = w31309 | w31310 ;
  assign w31312 = \pi077 ^ w31196 ;
  assign w31313 = ( ~w31204 & w31311 ) | ( ~w31204 & w31312 ) | ( w31311 & w31312 ) ;
  assign w31314 = w31312 | w31313 ;
  assign w31315 = \pi078 ^ w31189 ;
  assign w31316 = ( ~w31197 & w31314 ) | ( ~w31197 & w31315 ) | ( w31314 & w31315 ) ;
  assign w31317 = w31315 | w31316 ;
  assign w31318 = \pi079 ^ w31182 ;
  assign w31319 = ( ~w31190 & w31317 ) | ( ~w31190 & w31318 ) | ( w31317 & w31318 ) ;
  assign w31320 = w31318 | w31319 ;
  assign w31321 = \pi080 ^ w31175 ;
  assign w31322 = ( ~w31183 & w31320 ) | ( ~w31183 & w31321 ) | ( w31320 & w31321 ) ;
  assign w31323 = w31321 | w31322 ;
  assign w31324 = \pi081 ^ w31168 ;
  assign w31325 = ( ~w31176 & w31323 ) | ( ~w31176 & w31324 ) | ( w31323 & w31324 ) ;
  assign w31326 = w31324 | w31325 ;
  assign w31327 = \pi082 ^ w31161 ;
  assign w31328 = ( ~w31169 & w31326 ) | ( ~w31169 & w31327 ) | ( w31326 & w31327 ) ;
  assign w31329 = w31327 | w31328 ;
  assign w31330 = \pi083 ^ w31154 ;
  assign w31331 = ( ~w31162 & w31329 ) | ( ~w31162 & w31330 ) | ( w31329 & w31330 ) ;
  assign w31332 = w31330 | w31331 ;
  assign w31333 = \pi084 ^ w31147 ;
  assign w31334 = ( ~w31155 & w31332 ) | ( ~w31155 & w31333 ) | ( w31332 & w31333 ) ;
  assign w31335 = w31333 | w31334 ;
  assign w31336 = \pi085 ^ w31140 ;
  assign w31337 = ( ~w31148 & w31335 ) | ( ~w31148 & w31336 ) | ( w31335 & w31336 ) ;
  assign w31338 = w31336 | w31337 ;
  assign w31339 = \pi086 ^ w31133 ;
  assign w31340 = ( ~w31141 & w31338 ) | ( ~w31141 & w31339 ) | ( w31338 & w31339 ) ;
  assign w31341 = w31339 | w31340 ;
  assign w31342 = \pi087 ^ w31126 ;
  assign w31343 = ( ~w31134 & w31341 ) | ( ~w31134 & w31342 ) | ( w31341 & w31342 ) ;
  assign w31344 = w31342 | w31343 ;
  assign w31345 = \pi088 ^ w31119 ;
  assign w31346 = ( ~w31127 & w31344 ) | ( ~w31127 & w31345 ) | ( w31344 & w31345 ) ;
  assign w31347 = w31345 | w31346 ;
  assign w31348 = \pi089 ^ w31112 ;
  assign w31349 = ( ~w31120 & w31347 ) | ( ~w31120 & w31348 ) | ( w31347 & w31348 ) ;
  assign w31350 = w31348 | w31349 ;
  assign w31351 = \pi090 ^ w31105 ;
  assign w31352 = ( ~w31113 & w31350 ) | ( ~w31113 & w31351 ) | ( w31350 & w31351 ) ;
  assign w31353 = w31351 | w31352 ;
  assign w31354 = \pi091 ^ w31098 ;
  assign w31355 = ( ~w31106 & w31353 ) | ( ~w31106 & w31354 ) | ( w31353 & w31354 ) ;
  assign w31356 = w31354 | w31355 ;
  assign w31357 = \pi092 ^ w31091 ;
  assign w31358 = ( ~w31099 & w31356 ) | ( ~w31099 & w31357 ) | ( w31356 & w31357 ) ;
  assign w31359 = w31357 | w31358 ;
  assign w31360 = \pi093 ^ w31084 ;
  assign w31361 = ( ~w31092 & w31359 ) | ( ~w31092 & w31360 ) | ( w31359 & w31360 ) ;
  assign w31362 = w31360 | w31361 ;
  assign w31363 = \pi094 ^ w31077 ;
  assign w31364 = ( ~w31085 & w31362 ) | ( ~w31085 & w31363 ) | ( w31362 & w31363 ) ;
  assign w31365 = w31363 | w31364 ;
  assign w31366 = \pi095 ^ w31070 ;
  assign w31367 = ( ~w31078 & w31365 ) | ( ~w31078 & w31366 ) | ( w31365 & w31366 ) ;
  assign w31368 = w31366 | w31367 ;
  assign w31369 = \pi096 ^ w31063 ;
  assign w31370 = ( ~w31071 & w31368 ) | ( ~w31071 & w31369 ) | ( w31368 & w31369 ) ;
  assign w31371 = w31369 | w31370 ;
  assign w31372 = \pi097 ^ w31056 ;
  assign w31373 = ( ~w31064 & w31371 ) | ( ~w31064 & w31372 ) | ( w31371 & w31372 ) ;
  assign w31374 = w31372 | w31373 ;
  assign w31375 = \pi098 ^ w31049 ;
  assign w31376 = ( ~w31057 & w31374 ) | ( ~w31057 & w31375 ) | ( w31374 & w31375 ) ;
  assign w31377 = w31375 | w31376 ;
  assign w31378 = \pi099 ^ w31042 ;
  assign w31379 = ( ~w31050 & w31377 ) | ( ~w31050 & w31378 ) | ( w31377 & w31378 ) ;
  assign w31380 = w31378 | w31379 ;
  assign w31381 = \pi100 ^ w31035 ;
  assign w31382 = ( ~w31043 & w31380 ) | ( ~w31043 & w31381 ) | ( w31380 & w31381 ) ;
  assign w31383 = w31381 | w31382 ;
  assign w31384 = \pi101 ^ w31028 ;
  assign w31385 = ( ~w31036 & w31383 ) | ( ~w31036 & w31384 ) | ( w31383 & w31384 ) ;
  assign w31386 = w31384 | w31385 ;
  assign w31387 = \pi102 ^ w31021 ;
  assign w31388 = ( ~w31029 & w31386 ) | ( ~w31029 & w31387 ) | ( w31386 & w31387 ) ;
  assign w31389 = w31387 | w31388 ;
  assign w31390 = \pi103 ^ w31014 ;
  assign w31391 = ( ~w31022 & w31389 ) | ( ~w31022 & w31390 ) | ( w31389 & w31390 ) ;
  assign w31392 = w31390 | w31391 ;
  assign w31393 = \pi104 ^ w31007 ;
  assign w31394 = ( ~w31015 & w31392 ) | ( ~w31015 & w31393 ) | ( w31392 & w31393 ) ;
  assign w31395 = w31393 | w31394 ;
  assign w31396 = \pi105 ^ w31000 ;
  assign w31397 = ( ~w31008 & w31395 ) | ( ~w31008 & w31396 ) | ( w31395 & w31396 ) ;
  assign w31398 = w31396 | w31397 ;
  assign w31399 = \pi106 ^ w30993 ;
  assign w31400 = ( ~w31001 & w31398 ) | ( ~w31001 & w31399 ) | ( w31398 & w31399 ) ;
  assign w31401 = w31399 | w31400 ;
  assign w31402 = \pi107 ^ w30986 ;
  assign w31403 = ( ~w30994 & w31401 ) | ( ~w30994 & w31402 ) | ( w31401 & w31402 ) ;
  assign w31404 = w31402 | w31403 ;
  assign w31405 = \pi108 ^ w30979 ;
  assign w31406 = ( ~w30987 & w31404 ) | ( ~w30987 & w31405 ) | ( w31404 & w31405 ) ;
  assign w31407 = w31405 | w31406 ;
  assign w31408 = \pi109 ^ w30972 ;
  assign w31409 = ( ~w30980 & w31407 ) | ( ~w30980 & w31408 ) | ( w31407 & w31408 ) ;
  assign w31410 = w31408 | w31409 ;
  assign w31411 = \pi110 ^ w30965 ;
  assign w31412 = ( ~w30973 & w31410 ) | ( ~w30973 & w31411 ) | ( w31410 & w31411 ) ;
  assign w31413 = w31411 | w31412 ;
  assign w31414 = \pi111 ^ w30952 ;
  assign w31415 = ( ~w30966 & w31413 ) | ( ~w30966 & w31414 ) | ( w31413 & w31414 ) ;
  assign w31416 = w31414 | w31415 ;
  assign w31417 = \pi112 ^ w30958 ;
  assign w31418 = w30959 & ~w31417 ;
  assign w31419 = ( w31416 & w31417 ) | ( w31416 & ~w31418 ) | ( w31417 & ~w31418 ) ;
  assign w31420 = ~\pi112 & w30958 ;
  assign w31421 = w31419 & ~w31420 ;
  assign w31422 = w275 | w31421 ;
  assign w31423 = w30952 & w31422 ;
  assign w31424 = ~w30966 & w31413 ;
  assign w31425 = w31414 ^ w31424 ;
  assign w31426 = ~w31422 & w31425 ;
  assign w31427 = w31423 | w31426 ;
  assign w31428 = ~\pi112 & w31427 ;
  assign w31429 = w30965 & w31422 ;
  assign w31430 = ~w30973 & w31410 ;
  assign w31431 = w31411 ^ w31430 ;
  assign w31432 = ~w31422 & w31431 ;
  assign w31433 = w31429 | w31432 ;
  assign w31434 = ~\pi111 & w31433 ;
  assign w31435 = w30972 & w31422 ;
  assign w31436 = ~w30980 & w31407 ;
  assign w31437 = w31408 ^ w31436 ;
  assign w31438 = ~w31422 & w31437 ;
  assign w31439 = w31435 | w31438 ;
  assign w31440 = ~\pi110 & w31439 ;
  assign w31441 = w30979 & w31422 ;
  assign w31442 = ~w30987 & w31404 ;
  assign w31443 = w31405 ^ w31442 ;
  assign w31444 = ~w31422 & w31443 ;
  assign w31445 = w31441 | w31444 ;
  assign w31446 = ~\pi109 & w31445 ;
  assign w31447 = w30986 & w31422 ;
  assign w31448 = ~w30994 & w31401 ;
  assign w31449 = w31402 ^ w31448 ;
  assign w31450 = ~w31422 & w31449 ;
  assign w31451 = w31447 | w31450 ;
  assign w31452 = ~\pi108 & w31451 ;
  assign w31453 = w30993 & w31422 ;
  assign w31454 = ~w31001 & w31398 ;
  assign w31455 = w31399 ^ w31454 ;
  assign w31456 = ~w31422 & w31455 ;
  assign w31457 = w31453 | w31456 ;
  assign w31458 = ~\pi107 & w31457 ;
  assign w31459 = w31000 & w31422 ;
  assign w31460 = ~w31008 & w31395 ;
  assign w31461 = w31396 ^ w31460 ;
  assign w31462 = ~w31422 & w31461 ;
  assign w31463 = w31459 | w31462 ;
  assign w31464 = ~\pi106 & w31463 ;
  assign w31465 = w31007 & w31422 ;
  assign w31466 = ~w31015 & w31392 ;
  assign w31467 = w31393 ^ w31466 ;
  assign w31468 = ~w31422 & w31467 ;
  assign w31469 = w31465 | w31468 ;
  assign w31470 = ~\pi105 & w31469 ;
  assign w31471 = w31014 & w31422 ;
  assign w31472 = ~w31022 & w31389 ;
  assign w31473 = w31390 ^ w31472 ;
  assign w31474 = ~w31422 & w31473 ;
  assign w31475 = w31471 | w31474 ;
  assign w31476 = ~\pi104 & w31475 ;
  assign w31477 = w31021 & w31422 ;
  assign w31478 = ~w31029 & w31386 ;
  assign w31479 = w31387 ^ w31478 ;
  assign w31480 = ~w31422 & w31479 ;
  assign w31481 = w31477 | w31480 ;
  assign w31482 = ~\pi103 & w31481 ;
  assign w31483 = w31028 & w31422 ;
  assign w31484 = ~w31036 & w31383 ;
  assign w31485 = w31384 ^ w31484 ;
  assign w31486 = ~w31422 & w31485 ;
  assign w31487 = w31483 | w31486 ;
  assign w31488 = ~\pi102 & w31487 ;
  assign w31489 = w31035 & w31422 ;
  assign w31490 = ~w31043 & w31380 ;
  assign w31491 = w31381 ^ w31490 ;
  assign w31492 = ~w31422 & w31491 ;
  assign w31493 = w31489 | w31492 ;
  assign w31494 = ~\pi101 & w31493 ;
  assign w31495 = w31042 & w31422 ;
  assign w31496 = ~w31050 & w31377 ;
  assign w31497 = w31378 ^ w31496 ;
  assign w31498 = ~w31422 & w31497 ;
  assign w31499 = w31495 | w31498 ;
  assign w31500 = ~\pi100 & w31499 ;
  assign w31501 = w31049 & w31422 ;
  assign w31502 = ~w31057 & w31374 ;
  assign w31503 = w31375 ^ w31502 ;
  assign w31504 = ~w31422 & w31503 ;
  assign w31505 = w31501 | w31504 ;
  assign w31506 = ~\pi099 & w31505 ;
  assign w31507 = w31056 & w31422 ;
  assign w31508 = ~w31064 & w31371 ;
  assign w31509 = w31372 ^ w31508 ;
  assign w31510 = ~w31422 & w31509 ;
  assign w31511 = w31507 | w31510 ;
  assign w31512 = ~\pi098 & w31511 ;
  assign w31513 = w31063 & w31422 ;
  assign w31514 = ~w31071 & w31368 ;
  assign w31515 = w31369 ^ w31514 ;
  assign w31516 = ~w31422 & w31515 ;
  assign w31517 = w31513 | w31516 ;
  assign w31518 = ~\pi097 & w31517 ;
  assign w31519 = w31070 & w31422 ;
  assign w31520 = ~w31078 & w31365 ;
  assign w31521 = w31366 ^ w31520 ;
  assign w31522 = ~w31422 & w31521 ;
  assign w31523 = w31519 | w31522 ;
  assign w31524 = ~\pi096 & w31523 ;
  assign w31525 = w31077 & w31422 ;
  assign w31526 = ~w31085 & w31362 ;
  assign w31527 = w31363 ^ w31526 ;
  assign w31528 = ~w31422 & w31527 ;
  assign w31529 = w31525 | w31528 ;
  assign w31530 = ~\pi095 & w31529 ;
  assign w31531 = w31084 & w31422 ;
  assign w31532 = ~w31092 & w31359 ;
  assign w31533 = w31360 ^ w31532 ;
  assign w31534 = ~w31422 & w31533 ;
  assign w31535 = w31531 | w31534 ;
  assign w31536 = ~\pi094 & w31535 ;
  assign w31537 = w31091 & w31422 ;
  assign w31538 = ~w31099 & w31356 ;
  assign w31539 = w31357 ^ w31538 ;
  assign w31540 = ~w31422 & w31539 ;
  assign w31541 = w31537 | w31540 ;
  assign w31542 = ~\pi093 & w31541 ;
  assign w31543 = w31098 & w31422 ;
  assign w31544 = ~w31106 & w31353 ;
  assign w31545 = w31354 ^ w31544 ;
  assign w31546 = ~w31422 & w31545 ;
  assign w31547 = w31543 | w31546 ;
  assign w31548 = ~\pi092 & w31547 ;
  assign w31549 = w31105 & w31422 ;
  assign w31550 = ~w31113 & w31350 ;
  assign w31551 = w31351 ^ w31550 ;
  assign w31552 = ~w31422 & w31551 ;
  assign w31553 = w31549 | w31552 ;
  assign w31554 = ~\pi091 & w31553 ;
  assign w31555 = w31112 & w31422 ;
  assign w31556 = ~w31120 & w31347 ;
  assign w31557 = w31348 ^ w31556 ;
  assign w31558 = ~w31422 & w31557 ;
  assign w31559 = w31555 | w31558 ;
  assign w31560 = ~\pi090 & w31559 ;
  assign w31561 = w31119 & w31422 ;
  assign w31562 = ~w31127 & w31344 ;
  assign w31563 = w31345 ^ w31562 ;
  assign w31564 = ~w31422 & w31563 ;
  assign w31565 = w31561 | w31564 ;
  assign w31566 = ~\pi089 & w31565 ;
  assign w31567 = w31126 & w31422 ;
  assign w31568 = ~w31134 & w31341 ;
  assign w31569 = w31342 ^ w31568 ;
  assign w31570 = ~w31422 & w31569 ;
  assign w31571 = w31567 | w31570 ;
  assign w31572 = ~\pi088 & w31571 ;
  assign w31573 = w31133 & w31422 ;
  assign w31574 = ~w31141 & w31338 ;
  assign w31575 = w31339 ^ w31574 ;
  assign w31576 = ~w31422 & w31575 ;
  assign w31577 = w31573 | w31576 ;
  assign w31578 = ~\pi087 & w31577 ;
  assign w31579 = w31140 & w31422 ;
  assign w31580 = ~w31148 & w31335 ;
  assign w31581 = w31336 ^ w31580 ;
  assign w31582 = ~w31422 & w31581 ;
  assign w31583 = w31579 | w31582 ;
  assign w31584 = ~\pi086 & w31583 ;
  assign w31585 = w31147 & w31422 ;
  assign w31586 = ~w31155 & w31332 ;
  assign w31587 = w31333 ^ w31586 ;
  assign w31588 = ~w31422 & w31587 ;
  assign w31589 = w31585 | w31588 ;
  assign w31590 = ~\pi085 & w31589 ;
  assign w31591 = w31154 & w31422 ;
  assign w31592 = ~w31162 & w31329 ;
  assign w31593 = w31330 ^ w31592 ;
  assign w31594 = ~w31422 & w31593 ;
  assign w31595 = w31591 | w31594 ;
  assign w31596 = ~\pi084 & w31595 ;
  assign w31597 = w31161 & w31422 ;
  assign w31598 = ~w31169 & w31326 ;
  assign w31599 = w31327 ^ w31598 ;
  assign w31600 = ~w31422 & w31599 ;
  assign w31601 = w31597 | w31600 ;
  assign w31602 = ~\pi083 & w31601 ;
  assign w31603 = w31168 & w31422 ;
  assign w31604 = ~w31176 & w31323 ;
  assign w31605 = w31324 ^ w31604 ;
  assign w31606 = ~w31422 & w31605 ;
  assign w31607 = w31603 | w31606 ;
  assign w31608 = ~\pi082 & w31607 ;
  assign w31609 = w31175 & w31422 ;
  assign w31610 = ~w31183 & w31320 ;
  assign w31611 = w31321 ^ w31610 ;
  assign w31612 = ~w31422 & w31611 ;
  assign w31613 = w31609 | w31612 ;
  assign w31614 = ~\pi081 & w31613 ;
  assign w31615 = w31182 & w31422 ;
  assign w31616 = ~w31190 & w31317 ;
  assign w31617 = w31318 ^ w31616 ;
  assign w31618 = ~w31422 & w31617 ;
  assign w31619 = w31615 | w31618 ;
  assign w31620 = ~\pi080 & w31619 ;
  assign w31621 = w31189 & w31422 ;
  assign w31622 = ~w31197 & w31314 ;
  assign w31623 = w31315 ^ w31622 ;
  assign w31624 = ~w31422 & w31623 ;
  assign w31625 = w31621 | w31624 ;
  assign w31626 = ~\pi079 & w31625 ;
  assign w31627 = w31196 & w31422 ;
  assign w31628 = ~w31204 & w31311 ;
  assign w31629 = w31312 ^ w31628 ;
  assign w31630 = ~w31422 & w31629 ;
  assign w31631 = w31627 | w31630 ;
  assign w31632 = ~\pi078 & w31631 ;
  assign w31633 = w31203 & w31422 ;
  assign w31634 = ~w31211 & w31308 ;
  assign w31635 = w31309 ^ w31634 ;
  assign w31636 = ~w31422 & w31635 ;
  assign w31637 = w31633 | w31636 ;
  assign w31638 = ~\pi077 & w31637 ;
  assign w31639 = w31210 & w31422 ;
  assign w31640 = ~w31218 & w31305 ;
  assign w31641 = w31306 ^ w31640 ;
  assign w31642 = ~w31422 & w31641 ;
  assign w31643 = w31639 | w31642 ;
  assign w31644 = ~\pi076 & w31643 ;
  assign w31645 = w31217 & w31422 ;
  assign w31646 = ~w31225 & w31302 ;
  assign w31647 = w31303 ^ w31646 ;
  assign w31648 = ~w31422 & w31647 ;
  assign w31649 = w31645 | w31648 ;
  assign w31650 = ~\pi075 & w31649 ;
  assign w31651 = w31224 & w31422 ;
  assign w31652 = ~w31232 & w31299 ;
  assign w31653 = w31300 ^ w31652 ;
  assign w31654 = ~w31422 & w31653 ;
  assign w31655 = w31651 | w31654 ;
  assign w31656 = ~\pi074 & w31655 ;
  assign w31657 = w31231 & w31422 ;
  assign w31658 = ~w31239 & w31296 ;
  assign w31659 = w31297 ^ w31658 ;
  assign w31660 = ~w31422 & w31659 ;
  assign w31661 = w31657 | w31660 ;
  assign w31662 = ~\pi073 & w31661 ;
  assign w31663 = w31238 & w31422 ;
  assign w31664 = ~w31246 & w31293 ;
  assign w31665 = w31294 ^ w31664 ;
  assign w31666 = ~w31422 & w31665 ;
  assign w31667 = w31663 | w31666 ;
  assign w31668 = ~\pi072 & w31667 ;
  assign w31669 = w31245 & w31422 ;
  assign w31670 = ~w31253 & w31290 ;
  assign w31671 = w31291 ^ w31670 ;
  assign w31672 = ~w31422 & w31671 ;
  assign w31673 = w31669 | w31672 ;
  assign w31674 = ~\pi071 & w31673 ;
  assign w31675 = w31252 & w31422 ;
  assign w31676 = ~w31260 & w31287 ;
  assign w31677 = w31288 ^ w31676 ;
  assign w31678 = ~w31422 & w31677 ;
  assign w31679 = w31675 | w31678 ;
  assign w31680 = ~\pi070 & w31679 ;
  assign w31681 = w31259 & w31422 ;
  assign w31682 = ~w31269 & w31284 ;
  assign w31683 = w31285 ^ w31682 ;
  assign w31684 = ~w31422 & w31683 ;
  assign w31685 = w31681 | w31684 ;
  assign w31686 = ~\pi069 & w31685 ;
  assign w31687 = w31268 & w31422 ;
  assign w31688 = ~w31276 & w31281 ;
  assign w31689 = w31282 ^ w31688 ;
  assign w31690 = ~w31422 & w31689 ;
  assign w31691 = w31687 | w31690 ;
  assign w31692 = ~\pi068 & w31691 ;
  assign w31693 = \pi064 & ~w30946 ;
  assign w31694 = \pi016 ^ w31693 ;
  assign w31695 = ( \pi065 & w12310 ) | ( \pi065 & ~w31694 ) | ( w12310 & ~w31694 ) ;
  assign w31696 = w31277 ^ w31695 ;
  assign w31697 = ( w275 & w31421 ) | ( w275 & w31696 ) | ( w31421 & w31696 ) ;
  assign w31698 = w31696 & ~w31697 ;
  assign w31699 = ( w31275 & w31422 ) | ( w31275 & w31698 ) | ( w31422 & w31698 ) ;
  assign w31700 = w31698 | w31699 ;
  assign w31701 = ~\pi067 & w31700 ;
  assign w31702 = \pi015 ^ w30946 ;
  assign w31703 = ( \pi064 & w275 ) | ( \pi064 & w31702 ) | ( w275 & w31702 ) ;
  assign w31704 = w12318 ^ w31703 ;
  assign w31705 = ~w275 & w31704 ;
  assign w31706 = ~w31421 & w31705 ;
  assign w31707 = ( ~\pi064 & w30946 ) | ( ~\pi064 & w31422 ) | ( w30946 & w31422 ) ;
  assign w31708 = \pi016 ^ w31707 ;
  assign w31709 = w31422 & ~w31708 ;
  assign w31710 = w31706 | w31709 ;
  assign w31711 = ~\pi066 & w31710 ;
  assign w31712 = ( \pi015 & ~w12333 ) | ( \pi015 & w31421 ) | ( ~w12333 & w31421 ) ;
  assign w31713 = \pi015 & w31712 ;
  assign w31714 = ( w267 & ~w448 ) | ( w267 & w31421 ) | ( ~w448 & w31421 ) ;
  assign w31715 = w12336 & ~w31714 ;
  assign w31716 = w31422 | w31706 ;
  assign w31717 = ( w31694 & w31706 ) | ( w31694 & w31716 ) | ( w31706 & w31716 ) ;
  assign w31718 = \pi066 ^ w31717 ;
  assign w31719 = w31713 | w31715 ;
  assign w31720 = ( \pi065 & w12339 ) | ( \pi065 & ~w31719 ) | ( w12339 & ~w31719 ) ;
  assign w31721 = w31718 | w31720 ;
  assign w31722 = ~w31275 & w31422 ;
  assign w31723 = ( w31422 & w31698 ) | ( w31422 & ~w31722 ) | ( w31698 & ~w31722 ) ;
  assign w31724 = \pi067 ^ w31723 ;
  assign w31725 = ( ~w31711 & w31721 ) | ( ~w31711 & w31724 ) | ( w31721 & w31724 ) ;
  assign w31726 = w31724 | w31725 ;
  assign w31727 = \pi068 ^ w31691 ;
  assign w31728 = ( ~w31701 & w31726 ) | ( ~w31701 & w31727 ) | ( w31726 & w31727 ) ;
  assign w31729 = w31727 | w31728 ;
  assign w31730 = \pi069 ^ w31685 ;
  assign w31731 = ( ~w31692 & w31729 ) | ( ~w31692 & w31730 ) | ( w31729 & w31730 ) ;
  assign w31732 = w31730 | w31731 ;
  assign w31733 = \pi070 ^ w31679 ;
  assign w31734 = ( ~w31686 & w31732 ) | ( ~w31686 & w31733 ) | ( w31732 & w31733 ) ;
  assign w31735 = w31733 | w31734 ;
  assign w31736 = \pi071 ^ w31673 ;
  assign w31737 = ( ~w31680 & w31735 ) | ( ~w31680 & w31736 ) | ( w31735 & w31736 ) ;
  assign w31738 = w31736 | w31737 ;
  assign w31739 = \pi072 ^ w31667 ;
  assign w31740 = ( ~w31674 & w31738 ) | ( ~w31674 & w31739 ) | ( w31738 & w31739 ) ;
  assign w31741 = w31739 | w31740 ;
  assign w31742 = \pi073 ^ w31661 ;
  assign w31743 = ( ~w31668 & w31741 ) | ( ~w31668 & w31742 ) | ( w31741 & w31742 ) ;
  assign w31744 = w31742 | w31743 ;
  assign w31745 = \pi074 ^ w31655 ;
  assign w31746 = ( ~w31662 & w31744 ) | ( ~w31662 & w31745 ) | ( w31744 & w31745 ) ;
  assign w31747 = w31745 | w31746 ;
  assign w31748 = \pi075 ^ w31649 ;
  assign w31749 = ( ~w31656 & w31747 ) | ( ~w31656 & w31748 ) | ( w31747 & w31748 ) ;
  assign w31750 = w31748 | w31749 ;
  assign w31751 = \pi076 ^ w31643 ;
  assign w31752 = ( ~w31650 & w31750 ) | ( ~w31650 & w31751 ) | ( w31750 & w31751 ) ;
  assign w31753 = w31751 | w31752 ;
  assign w31754 = \pi077 ^ w31637 ;
  assign w31755 = ( ~w31644 & w31753 ) | ( ~w31644 & w31754 ) | ( w31753 & w31754 ) ;
  assign w31756 = w31754 | w31755 ;
  assign w31757 = \pi078 ^ w31631 ;
  assign w31758 = ( ~w31638 & w31756 ) | ( ~w31638 & w31757 ) | ( w31756 & w31757 ) ;
  assign w31759 = w31757 | w31758 ;
  assign w31760 = \pi079 ^ w31625 ;
  assign w31761 = ( ~w31632 & w31759 ) | ( ~w31632 & w31760 ) | ( w31759 & w31760 ) ;
  assign w31762 = w31760 | w31761 ;
  assign w31763 = \pi080 ^ w31619 ;
  assign w31764 = ( ~w31626 & w31762 ) | ( ~w31626 & w31763 ) | ( w31762 & w31763 ) ;
  assign w31765 = w31763 | w31764 ;
  assign w31766 = \pi081 ^ w31613 ;
  assign w31767 = ( ~w31620 & w31765 ) | ( ~w31620 & w31766 ) | ( w31765 & w31766 ) ;
  assign w31768 = w31766 | w31767 ;
  assign w31769 = \pi082 ^ w31607 ;
  assign w31770 = ( ~w31614 & w31768 ) | ( ~w31614 & w31769 ) | ( w31768 & w31769 ) ;
  assign w31771 = w31769 | w31770 ;
  assign w31772 = \pi083 ^ w31601 ;
  assign w31773 = ( ~w31608 & w31771 ) | ( ~w31608 & w31772 ) | ( w31771 & w31772 ) ;
  assign w31774 = w31772 | w31773 ;
  assign w31775 = \pi084 ^ w31595 ;
  assign w31776 = ( ~w31602 & w31774 ) | ( ~w31602 & w31775 ) | ( w31774 & w31775 ) ;
  assign w31777 = w31775 | w31776 ;
  assign w31778 = \pi085 ^ w31589 ;
  assign w31779 = ( ~w31596 & w31777 ) | ( ~w31596 & w31778 ) | ( w31777 & w31778 ) ;
  assign w31780 = w31778 | w31779 ;
  assign w31781 = \pi086 ^ w31583 ;
  assign w31782 = ( ~w31590 & w31780 ) | ( ~w31590 & w31781 ) | ( w31780 & w31781 ) ;
  assign w31783 = w31781 | w31782 ;
  assign w31784 = \pi087 ^ w31577 ;
  assign w31785 = ( ~w31584 & w31783 ) | ( ~w31584 & w31784 ) | ( w31783 & w31784 ) ;
  assign w31786 = w31784 | w31785 ;
  assign w31787 = \pi088 ^ w31571 ;
  assign w31788 = ( ~w31578 & w31786 ) | ( ~w31578 & w31787 ) | ( w31786 & w31787 ) ;
  assign w31789 = w31787 | w31788 ;
  assign w31790 = \pi089 ^ w31565 ;
  assign w31791 = ( ~w31572 & w31789 ) | ( ~w31572 & w31790 ) | ( w31789 & w31790 ) ;
  assign w31792 = w31790 | w31791 ;
  assign w31793 = \pi090 ^ w31559 ;
  assign w31794 = ( ~w31566 & w31792 ) | ( ~w31566 & w31793 ) | ( w31792 & w31793 ) ;
  assign w31795 = w31793 | w31794 ;
  assign w31796 = \pi091 ^ w31553 ;
  assign w31797 = ( ~w31560 & w31795 ) | ( ~w31560 & w31796 ) | ( w31795 & w31796 ) ;
  assign w31798 = w31796 | w31797 ;
  assign w31799 = \pi092 ^ w31547 ;
  assign w31800 = ( ~w31554 & w31798 ) | ( ~w31554 & w31799 ) | ( w31798 & w31799 ) ;
  assign w31801 = w31799 | w31800 ;
  assign w31802 = \pi093 ^ w31541 ;
  assign w31803 = ( ~w31548 & w31801 ) | ( ~w31548 & w31802 ) | ( w31801 & w31802 ) ;
  assign w31804 = w31802 | w31803 ;
  assign w31805 = \pi094 ^ w31535 ;
  assign w31806 = ( ~w31542 & w31804 ) | ( ~w31542 & w31805 ) | ( w31804 & w31805 ) ;
  assign w31807 = w31805 | w31806 ;
  assign w31808 = \pi095 ^ w31529 ;
  assign w31809 = ( ~w31536 & w31807 ) | ( ~w31536 & w31808 ) | ( w31807 & w31808 ) ;
  assign w31810 = w31808 | w31809 ;
  assign w31811 = \pi096 ^ w31523 ;
  assign w31812 = ( ~w31530 & w31810 ) | ( ~w31530 & w31811 ) | ( w31810 & w31811 ) ;
  assign w31813 = w31811 | w31812 ;
  assign w31814 = \pi097 ^ w31517 ;
  assign w31815 = ( ~w31524 & w31813 ) | ( ~w31524 & w31814 ) | ( w31813 & w31814 ) ;
  assign w31816 = w31814 | w31815 ;
  assign w31817 = \pi098 ^ w31511 ;
  assign w31818 = ( ~w31518 & w31816 ) | ( ~w31518 & w31817 ) | ( w31816 & w31817 ) ;
  assign w31819 = w31817 | w31818 ;
  assign w31820 = \pi099 ^ w31505 ;
  assign w31821 = ( ~w31512 & w31819 ) | ( ~w31512 & w31820 ) | ( w31819 & w31820 ) ;
  assign w31822 = w31820 | w31821 ;
  assign w31823 = \pi100 ^ w31499 ;
  assign w31824 = ( ~w31506 & w31822 ) | ( ~w31506 & w31823 ) | ( w31822 & w31823 ) ;
  assign w31825 = w31823 | w31824 ;
  assign w31826 = \pi101 ^ w31493 ;
  assign w31827 = ( ~w31500 & w31825 ) | ( ~w31500 & w31826 ) | ( w31825 & w31826 ) ;
  assign w31828 = w31826 | w31827 ;
  assign w31829 = \pi102 ^ w31487 ;
  assign w31830 = ( ~w31494 & w31828 ) | ( ~w31494 & w31829 ) | ( w31828 & w31829 ) ;
  assign w31831 = w31829 | w31830 ;
  assign w31832 = \pi103 ^ w31481 ;
  assign w31833 = ( ~w31488 & w31831 ) | ( ~w31488 & w31832 ) | ( w31831 & w31832 ) ;
  assign w31834 = w31832 | w31833 ;
  assign w31835 = \pi104 ^ w31475 ;
  assign w31836 = ( ~w31482 & w31834 ) | ( ~w31482 & w31835 ) | ( w31834 & w31835 ) ;
  assign w31837 = w31835 | w31836 ;
  assign w31838 = \pi105 ^ w31469 ;
  assign w31839 = ( ~w31476 & w31837 ) | ( ~w31476 & w31838 ) | ( w31837 & w31838 ) ;
  assign w31840 = w31838 | w31839 ;
  assign w31841 = \pi106 ^ w31463 ;
  assign w31842 = ( ~w31470 & w31840 ) | ( ~w31470 & w31841 ) | ( w31840 & w31841 ) ;
  assign w31843 = w31841 | w31842 ;
  assign w31844 = \pi107 ^ w31457 ;
  assign w31845 = ( ~w31464 & w31843 ) | ( ~w31464 & w31844 ) | ( w31843 & w31844 ) ;
  assign w31846 = w31844 | w31845 ;
  assign w31847 = \pi108 ^ w31451 ;
  assign w31848 = ( ~w31458 & w31846 ) | ( ~w31458 & w31847 ) | ( w31846 & w31847 ) ;
  assign w31849 = w31847 | w31848 ;
  assign w31850 = \pi109 ^ w31445 ;
  assign w31851 = ( ~w31452 & w31849 ) | ( ~w31452 & w31850 ) | ( w31849 & w31850 ) ;
  assign w31852 = w31850 | w31851 ;
  assign w31853 = \pi110 ^ w31439 ;
  assign w31854 = ( ~w31446 & w31852 ) | ( ~w31446 & w31853 ) | ( w31852 & w31853 ) ;
  assign w31855 = w31853 | w31854 ;
  assign w31856 = \pi111 ^ w31433 ;
  assign w31857 = ( ~w31440 & w31855 ) | ( ~w31440 & w31856 ) | ( w31855 & w31856 ) ;
  assign w31858 = w31856 | w31857 ;
  assign w31859 = \pi112 ^ w31427 ;
  assign w31860 = ( ~w31434 & w31858 ) | ( ~w31434 & w31859 ) | ( w31858 & w31859 ) ;
  assign w31861 = w31859 | w31860 ;
  assign w31862 = w30958 & w31422 ;
  assign w31863 = ~w30959 & w31416 ;
  assign w31864 = w31417 ^ w31863 ;
  assign w31865 = ~w31422 & w31864 ;
  assign w31866 = w31862 | w31865 ;
  assign w31867 = ~\pi113 & w31866 ;
  assign w31868 = ( \pi113 & ~w31862 ) | ( \pi113 & w31865 ) | ( ~w31862 & w31865 ) ;
  assign w31869 = ~w31865 & w31868 ;
  assign w31870 = w31867 | w31869 ;
  assign w31871 = ( ~w31428 & w31861 ) | ( ~w31428 & w31870 ) | ( w31861 & w31870 ) ;
  assign w31872 = ( w12496 & ~w31870 ) | ( w12496 & w31871 ) | ( ~w31870 & w31871 ) ;
  assign w31873 = w31870 | w31872 ;
  assign w31874 = ~w275 & w31866 ;
  assign w31875 = w31873 & ~w31874 ;
  assign w31876 = ~w31434 & w31858 ;
  assign w31877 = w31859 ^ w31876 ;
  assign w31878 = ~w31875 & w31877 ;
  assign w31879 = ( w31427 & w31873 ) | ( w31427 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31880 = ~w31874 & w31879 ;
  assign w31881 = w31878 | w31880 ;
  assign w31882 = ~\pi113 & w31881 ;
  assign w31883 = ~w31440 & w31855 ;
  assign w31884 = w31856 ^ w31883 ;
  assign w31885 = ~w31875 & w31884 ;
  assign w31886 = ( w31433 & w31873 ) | ( w31433 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31887 = ~w31874 & w31886 ;
  assign w31888 = w31885 | w31887 ;
  assign w31889 = ~\pi112 & w31888 ;
  assign w31890 = ~w31446 & w31852 ;
  assign w31891 = w31853 ^ w31890 ;
  assign w31892 = ~w31875 & w31891 ;
  assign w31893 = ( w31439 & w31873 ) | ( w31439 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31894 = ~w31874 & w31893 ;
  assign w31895 = w31892 | w31894 ;
  assign w31896 = ~\pi111 & w31895 ;
  assign w31897 = ~w31452 & w31849 ;
  assign w31898 = w31850 ^ w31897 ;
  assign w31899 = ~w31875 & w31898 ;
  assign w31900 = ( w31445 & w31873 ) | ( w31445 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31901 = ~w31874 & w31900 ;
  assign w31902 = w31899 | w31901 ;
  assign w31903 = ~\pi110 & w31902 ;
  assign w31904 = ~w31458 & w31846 ;
  assign w31905 = w31847 ^ w31904 ;
  assign w31906 = ~w31875 & w31905 ;
  assign w31907 = ( w31451 & w31873 ) | ( w31451 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31908 = ~w31874 & w31907 ;
  assign w31909 = w31906 | w31908 ;
  assign w31910 = ~\pi109 & w31909 ;
  assign w31911 = ~w31464 & w31843 ;
  assign w31912 = w31844 ^ w31911 ;
  assign w31913 = ~w31875 & w31912 ;
  assign w31914 = ( w31457 & w31873 ) | ( w31457 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31915 = ~w31874 & w31914 ;
  assign w31916 = w31913 | w31915 ;
  assign w31917 = ~\pi108 & w31916 ;
  assign w31918 = ~w31470 & w31840 ;
  assign w31919 = w31841 ^ w31918 ;
  assign w31920 = ~w31875 & w31919 ;
  assign w31921 = ( w31463 & w31873 ) | ( w31463 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31922 = ~w31874 & w31921 ;
  assign w31923 = w31920 | w31922 ;
  assign w31924 = ~\pi107 & w31923 ;
  assign w31925 = ~w31476 & w31837 ;
  assign w31926 = w31838 ^ w31925 ;
  assign w31927 = ~w31875 & w31926 ;
  assign w31928 = ( w31469 & w31873 ) | ( w31469 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31929 = ~w31874 & w31928 ;
  assign w31930 = w31927 | w31929 ;
  assign w31931 = ~\pi106 & w31930 ;
  assign w31932 = ~w31482 & w31834 ;
  assign w31933 = w31835 ^ w31932 ;
  assign w31934 = ~w31875 & w31933 ;
  assign w31935 = ( w31475 & w31873 ) | ( w31475 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31936 = ~w31874 & w31935 ;
  assign w31937 = w31934 | w31936 ;
  assign w31938 = ~\pi105 & w31937 ;
  assign w31939 = ~w31488 & w31831 ;
  assign w31940 = w31832 ^ w31939 ;
  assign w31941 = ~w31875 & w31940 ;
  assign w31942 = ( w31481 & w31873 ) | ( w31481 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31943 = ~w31874 & w31942 ;
  assign w31944 = w31941 | w31943 ;
  assign w31945 = ~\pi104 & w31944 ;
  assign w31946 = ~w31494 & w31828 ;
  assign w31947 = w31829 ^ w31946 ;
  assign w31948 = ~w31875 & w31947 ;
  assign w31949 = ( w31487 & w31873 ) | ( w31487 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31950 = ~w31874 & w31949 ;
  assign w31951 = w31948 | w31950 ;
  assign w31952 = ~\pi103 & w31951 ;
  assign w31953 = ~w31500 & w31825 ;
  assign w31954 = w31826 ^ w31953 ;
  assign w31955 = ~w31875 & w31954 ;
  assign w31956 = ( w31493 & w31873 ) | ( w31493 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31957 = ~w31874 & w31956 ;
  assign w31958 = w31955 | w31957 ;
  assign w31959 = ~\pi102 & w31958 ;
  assign w31960 = ~w31506 & w31822 ;
  assign w31961 = w31823 ^ w31960 ;
  assign w31962 = ~w31875 & w31961 ;
  assign w31963 = ( w31499 & w31873 ) | ( w31499 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31964 = ~w31874 & w31963 ;
  assign w31965 = w31962 | w31964 ;
  assign w31966 = ~\pi101 & w31965 ;
  assign w31967 = ~w31512 & w31819 ;
  assign w31968 = w31820 ^ w31967 ;
  assign w31969 = ~w31875 & w31968 ;
  assign w31970 = ( w31505 & w31873 ) | ( w31505 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31971 = ~w31874 & w31970 ;
  assign w31972 = w31969 | w31971 ;
  assign w31973 = ~\pi100 & w31972 ;
  assign w31974 = ~w31518 & w31816 ;
  assign w31975 = w31817 ^ w31974 ;
  assign w31976 = ~w31875 & w31975 ;
  assign w31977 = ( w31511 & w31873 ) | ( w31511 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31978 = ~w31874 & w31977 ;
  assign w31979 = w31976 | w31978 ;
  assign w31980 = ~\pi099 & w31979 ;
  assign w31981 = ~w31524 & w31813 ;
  assign w31982 = w31814 ^ w31981 ;
  assign w31983 = ~w31875 & w31982 ;
  assign w31984 = ( w31517 & w31873 ) | ( w31517 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31985 = ~w31874 & w31984 ;
  assign w31986 = w31983 | w31985 ;
  assign w31987 = ~\pi098 & w31986 ;
  assign w31988 = ~w31530 & w31810 ;
  assign w31989 = w31811 ^ w31988 ;
  assign w31990 = ~w31875 & w31989 ;
  assign w31991 = ( w31523 & w31873 ) | ( w31523 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31992 = ~w31874 & w31991 ;
  assign w31993 = w31990 | w31992 ;
  assign w31994 = ~\pi097 & w31993 ;
  assign w31995 = ~w31536 & w31807 ;
  assign w31996 = w31808 ^ w31995 ;
  assign w31997 = ~w31875 & w31996 ;
  assign w31998 = ( w31529 & w31873 ) | ( w31529 & w31874 ) | ( w31873 & w31874 ) ;
  assign w31999 = ~w31874 & w31998 ;
  assign w32000 = w31997 | w31999 ;
  assign w32001 = ~\pi096 & w32000 ;
  assign w32002 = ~w31542 & w31804 ;
  assign w32003 = w31805 ^ w32002 ;
  assign w32004 = ~w31875 & w32003 ;
  assign w32005 = ( w31535 & w31873 ) | ( w31535 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32006 = ~w31874 & w32005 ;
  assign w32007 = w32004 | w32006 ;
  assign w32008 = ~\pi095 & w32007 ;
  assign w32009 = ~w31548 & w31801 ;
  assign w32010 = w31802 ^ w32009 ;
  assign w32011 = ~w31875 & w32010 ;
  assign w32012 = ( w31541 & w31873 ) | ( w31541 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32013 = ~w31874 & w32012 ;
  assign w32014 = w32011 | w32013 ;
  assign w32015 = ~\pi094 & w32014 ;
  assign w32016 = ~w31554 & w31798 ;
  assign w32017 = w31799 ^ w32016 ;
  assign w32018 = ~w31875 & w32017 ;
  assign w32019 = ( w31547 & w31873 ) | ( w31547 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32020 = ~w31874 & w32019 ;
  assign w32021 = w32018 | w32020 ;
  assign w32022 = ~\pi093 & w32021 ;
  assign w32023 = ~w31560 & w31795 ;
  assign w32024 = w31796 ^ w32023 ;
  assign w32025 = ~w31875 & w32024 ;
  assign w32026 = ( w31553 & w31873 ) | ( w31553 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32027 = ~w31874 & w32026 ;
  assign w32028 = w32025 | w32027 ;
  assign w32029 = ~\pi092 & w32028 ;
  assign w32030 = ~w31566 & w31792 ;
  assign w32031 = w31793 ^ w32030 ;
  assign w32032 = ~w31875 & w32031 ;
  assign w32033 = ( w31559 & w31873 ) | ( w31559 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32034 = ~w31874 & w32033 ;
  assign w32035 = w32032 | w32034 ;
  assign w32036 = ~\pi091 & w32035 ;
  assign w32037 = ~w31572 & w31789 ;
  assign w32038 = w31790 ^ w32037 ;
  assign w32039 = ~w31875 & w32038 ;
  assign w32040 = ( w31565 & w31873 ) | ( w31565 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32041 = ~w31874 & w32040 ;
  assign w32042 = w32039 | w32041 ;
  assign w32043 = ~\pi090 & w32042 ;
  assign w32044 = ~w31578 & w31786 ;
  assign w32045 = w31787 ^ w32044 ;
  assign w32046 = ~w31875 & w32045 ;
  assign w32047 = ( w31571 & w31873 ) | ( w31571 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32048 = ~w31874 & w32047 ;
  assign w32049 = w32046 | w32048 ;
  assign w32050 = ~\pi089 & w32049 ;
  assign w32051 = ~w31584 & w31783 ;
  assign w32052 = w31784 ^ w32051 ;
  assign w32053 = ~w31875 & w32052 ;
  assign w32054 = ( w31577 & w31873 ) | ( w31577 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32055 = ~w31874 & w32054 ;
  assign w32056 = w32053 | w32055 ;
  assign w32057 = ~\pi088 & w32056 ;
  assign w32058 = ~w31590 & w31780 ;
  assign w32059 = w31781 ^ w32058 ;
  assign w32060 = ~w31875 & w32059 ;
  assign w32061 = ( w31583 & w31873 ) | ( w31583 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32062 = ~w31874 & w32061 ;
  assign w32063 = w32060 | w32062 ;
  assign w32064 = ~\pi087 & w32063 ;
  assign w32065 = ~w31596 & w31777 ;
  assign w32066 = w31778 ^ w32065 ;
  assign w32067 = ~w31875 & w32066 ;
  assign w32068 = ( w31589 & w31873 ) | ( w31589 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32069 = ~w31874 & w32068 ;
  assign w32070 = w32067 | w32069 ;
  assign w32071 = ~\pi086 & w32070 ;
  assign w32072 = ~w31602 & w31774 ;
  assign w32073 = w31775 ^ w32072 ;
  assign w32074 = ~w31875 & w32073 ;
  assign w32075 = ( w31595 & w31873 ) | ( w31595 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32076 = ~w31874 & w32075 ;
  assign w32077 = w32074 | w32076 ;
  assign w32078 = ~\pi085 & w32077 ;
  assign w32079 = ~w31608 & w31771 ;
  assign w32080 = w31772 ^ w32079 ;
  assign w32081 = ~w31875 & w32080 ;
  assign w32082 = ( w31601 & w31873 ) | ( w31601 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32083 = ~w31874 & w32082 ;
  assign w32084 = w32081 | w32083 ;
  assign w32085 = ~\pi084 & w32084 ;
  assign w32086 = ~w31614 & w31768 ;
  assign w32087 = w31769 ^ w32086 ;
  assign w32088 = ~w31875 & w32087 ;
  assign w32089 = ( w31607 & w31873 ) | ( w31607 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32090 = ~w31874 & w32089 ;
  assign w32091 = w32088 | w32090 ;
  assign w32092 = ~\pi083 & w32091 ;
  assign w32093 = ~w31620 & w31765 ;
  assign w32094 = w31766 ^ w32093 ;
  assign w32095 = ~w31875 & w32094 ;
  assign w32096 = ( w31613 & w31873 ) | ( w31613 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32097 = ~w31874 & w32096 ;
  assign w32098 = w32095 | w32097 ;
  assign w32099 = ~\pi082 & w32098 ;
  assign w32100 = ~w31626 & w31762 ;
  assign w32101 = w31763 ^ w32100 ;
  assign w32102 = ~w31875 & w32101 ;
  assign w32103 = ( w31619 & w31873 ) | ( w31619 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32104 = ~w31874 & w32103 ;
  assign w32105 = w32102 | w32104 ;
  assign w32106 = ~\pi081 & w32105 ;
  assign w32107 = ~w31632 & w31759 ;
  assign w32108 = w31760 ^ w32107 ;
  assign w32109 = ~w31875 & w32108 ;
  assign w32110 = ( w31625 & w31873 ) | ( w31625 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32111 = ~w31874 & w32110 ;
  assign w32112 = w32109 | w32111 ;
  assign w32113 = ~\pi080 & w32112 ;
  assign w32114 = ~w31638 & w31756 ;
  assign w32115 = w31757 ^ w32114 ;
  assign w32116 = ~w31875 & w32115 ;
  assign w32117 = ( w31631 & w31873 ) | ( w31631 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32118 = ~w31874 & w32117 ;
  assign w32119 = w32116 | w32118 ;
  assign w32120 = ~\pi079 & w32119 ;
  assign w32121 = ~w31644 & w31753 ;
  assign w32122 = w31754 ^ w32121 ;
  assign w32123 = ~w31875 & w32122 ;
  assign w32124 = ( w31637 & w31873 ) | ( w31637 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32125 = ~w31874 & w32124 ;
  assign w32126 = w32123 | w32125 ;
  assign w32127 = ~\pi078 & w32126 ;
  assign w32128 = ~w31650 & w31750 ;
  assign w32129 = w31751 ^ w32128 ;
  assign w32130 = ~w31875 & w32129 ;
  assign w32131 = ( w31643 & w31873 ) | ( w31643 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32132 = ~w31874 & w32131 ;
  assign w32133 = w32130 | w32132 ;
  assign w32134 = ~\pi077 & w32133 ;
  assign w32135 = ~w31656 & w31747 ;
  assign w32136 = w31748 ^ w32135 ;
  assign w32137 = ~w31875 & w32136 ;
  assign w32138 = ( w31649 & w31873 ) | ( w31649 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32139 = ~w31874 & w32138 ;
  assign w32140 = w32137 | w32139 ;
  assign w32141 = ~\pi076 & w32140 ;
  assign w32142 = ~w31662 & w31744 ;
  assign w32143 = w31745 ^ w32142 ;
  assign w32144 = ~w31875 & w32143 ;
  assign w32145 = ( w31655 & w31873 ) | ( w31655 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32146 = ~w31874 & w32145 ;
  assign w32147 = w32144 | w32146 ;
  assign w32148 = ~\pi075 & w32147 ;
  assign w32149 = ~w31668 & w31741 ;
  assign w32150 = w31742 ^ w32149 ;
  assign w32151 = ~w31875 & w32150 ;
  assign w32152 = ( w31661 & w31873 ) | ( w31661 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32153 = ~w31874 & w32152 ;
  assign w32154 = w32151 | w32153 ;
  assign w32155 = ~\pi074 & w32154 ;
  assign w32156 = ~w31674 & w31738 ;
  assign w32157 = w31739 ^ w32156 ;
  assign w32158 = ~w31875 & w32157 ;
  assign w32159 = ( w31667 & w31873 ) | ( w31667 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32160 = ~w31874 & w32159 ;
  assign w32161 = w32158 | w32160 ;
  assign w32162 = ~\pi073 & w32161 ;
  assign w32163 = ~w31680 & w31735 ;
  assign w32164 = w31736 ^ w32163 ;
  assign w32165 = ~w31875 & w32164 ;
  assign w32166 = ( w31673 & w31873 ) | ( w31673 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32167 = ~w31874 & w32166 ;
  assign w32168 = w32165 | w32167 ;
  assign w32169 = ~\pi072 & w32168 ;
  assign w32170 = ~w31686 & w31732 ;
  assign w32171 = w31733 ^ w32170 ;
  assign w32172 = ~w31875 & w32171 ;
  assign w32173 = ( w31679 & w31873 ) | ( w31679 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32174 = ~w31874 & w32173 ;
  assign w32175 = w32172 | w32174 ;
  assign w32176 = ~\pi071 & w32175 ;
  assign w32177 = ~w31692 & w31729 ;
  assign w32178 = w31730 ^ w32177 ;
  assign w32179 = ~w31875 & w32178 ;
  assign w32180 = ( w31685 & w31873 ) | ( w31685 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32181 = ~w31874 & w32180 ;
  assign w32182 = w32179 | w32181 ;
  assign w32183 = ~\pi070 & w32182 ;
  assign w32184 = ~w31701 & w31726 ;
  assign w32185 = w31727 ^ w32184 ;
  assign w32186 = ~w31875 & w32185 ;
  assign w32187 = ( w31691 & w31873 ) | ( w31691 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32188 = ~w31874 & w32187 ;
  assign w32189 = w32186 | w32188 ;
  assign w32190 = ~\pi069 & w32189 ;
  assign w32191 = ~w31711 & w31721 ;
  assign w32192 = w31724 ^ w32191 ;
  assign w32193 = ~w31875 & w32192 ;
  assign w32194 = ( w31700 & w31873 ) | ( w31700 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32195 = ~w31874 & w32194 ;
  assign w32196 = w32193 | w32195 ;
  assign w32197 = ~\pi068 & w32196 ;
  assign w32198 = w31718 ^ w31720 ;
  assign w32199 = ~w31875 & w32198 ;
  assign w32200 = ( w31710 & w31873 ) | ( w31710 & w31874 ) | ( w31873 & w31874 ) ;
  assign w32201 = ~w31874 & w32200 ;
  assign w32202 = w32199 | w32201 ;
  assign w32203 = ~\pi067 & w32202 ;
  assign w32204 = w12339 ^ w31719 ;
  assign w32205 = \pi065 ^ w32204 ;
  assign w32206 = w31875 ^ w32205 ;
  assign w32207 = ( w31719 & w32205 ) | ( w31719 & w32206 ) | ( w32205 & w32206 ) ;
  assign w32208 = ~\pi066 & w32207 ;
  assign w32209 = w31719 ^ w31875 ;
  assign w32210 = ( w31719 & w32205 ) | ( w31719 & ~w32209 ) | ( w32205 & ~w32209 ) ;
  assign w32211 = \pi066 ^ w32210 ;
  assign w32212 = ( \pi064 & ~w31875 ) | ( \pi064 & w32211 ) | ( ~w31875 & w32211 ) ;
  assign w32213 = \pi014 ^ w32212 ;
  assign w32214 = ( \pi065 & w13338 ) | ( \pi065 & ~w32213 ) | ( w13338 & ~w32213 ) ;
  assign w32215 = w32211 | w32214 ;
  assign w32216 = \pi067 ^ w32202 ;
  assign w32217 = ( ~w32208 & w32215 ) | ( ~w32208 & w32216 ) | ( w32215 & w32216 ) ;
  assign w32218 = w32216 | w32217 ;
  assign w32219 = \pi068 ^ w32196 ;
  assign w32220 = ( ~w32203 & w32218 ) | ( ~w32203 & w32219 ) | ( w32218 & w32219 ) ;
  assign w32221 = w32219 | w32220 ;
  assign w32222 = \pi069 ^ w32189 ;
  assign w32223 = ( ~w32197 & w32221 ) | ( ~w32197 & w32222 ) | ( w32221 & w32222 ) ;
  assign w32224 = w32222 | w32223 ;
  assign w32225 = \pi070 ^ w32182 ;
  assign w32226 = ( ~w32190 & w32224 ) | ( ~w32190 & w32225 ) | ( w32224 & w32225 ) ;
  assign w32227 = w32225 | w32226 ;
  assign w32228 = \pi071 ^ w32175 ;
  assign w32229 = ( ~w32183 & w32227 ) | ( ~w32183 & w32228 ) | ( w32227 & w32228 ) ;
  assign w32230 = w32228 | w32229 ;
  assign w32231 = \pi072 ^ w32168 ;
  assign w32232 = ( ~w32176 & w32230 ) | ( ~w32176 & w32231 ) | ( w32230 & w32231 ) ;
  assign w32233 = w32231 | w32232 ;
  assign w32234 = \pi073 ^ w32161 ;
  assign w32235 = ( ~w32169 & w32233 ) | ( ~w32169 & w32234 ) | ( w32233 & w32234 ) ;
  assign w32236 = w32234 | w32235 ;
  assign w32237 = \pi074 ^ w32154 ;
  assign w32238 = ( ~w32162 & w32236 ) | ( ~w32162 & w32237 ) | ( w32236 & w32237 ) ;
  assign w32239 = w32237 | w32238 ;
  assign w32240 = \pi075 ^ w32147 ;
  assign w32241 = ( ~w32155 & w32239 ) | ( ~w32155 & w32240 ) | ( w32239 & w32240 ) ;
  assign w32242 = w32240 | w32241 ;
  assign w32243 = \pi076 ^ w32140 ;
  assign w32244 = ( ~w32148 & w32242 ) | ( ~w32148 & w32243 ) | ( w32242 & w32243 ) ;
  assign w32245 = w32243 | w32244 ;
  assign w32246 = \pi077 ^ w32133 ;
  assign w32247 = ( ~w32141 & w32245 ) | ( ~w32141 & w32246 ) | ( w32245 & w32246 ) ;
  assign w32248 = w32246 | w32247 ;
  assign w32249 = \pi078 ^ w32126 ;
  assign w32250 = ( ~w32134 & w32248 ) | ( ~w32134 & w32249 ) | ( w32248 & w32249 ) ;
  assign w32251 = w32249 | w32250 ;
  assign w32252 = \pi079 ^ w32119 ;
  assign w32253 = ( ~w32127 & w32251 ) | ( ~w32127 & w32252 ) | ( w32251 & w32252 ) ;
  assign w32254 = w32252 | w32253 ;
  assign w32255 = \pi080 ^ w32112 ;
  assign w32256 = ( ~w32120 & w32254 ) | ( ~w32120 & w32255 ) | ( w32254 & w32255 ) ;
  assign w32257 = w32255 | w32256 ;
  assign w32258 = \pi081 ^ w32105 ;
  assign w32259 = ( ~w32113 & w32257 ) | ( ~w32113 & w32258 ) | ( w32257 & w32258 ) ;
  assign w32260 = w32258 | w32259 ;
  assign w32261 = \pi082 ^ w32098 ;
  assign w32262 = ( ~w32106 & w32260 ) | ( ~w32106 & w32261 ) | ( w32260 & w32261 ) ;
  assign w32263 = w32261 | w32262 ;
  assign w32264 = \pi083 ^ w32091 ;
  assign w32265 = ( ~w32099 & w32263 ) | ( ~w32099 & w32264 ) | ( w32263 & w32264 ) ;
  assign w32266 = w32264 | w32265 ;
  assign w32267 = \pi084 ^ w32084 ;
  assign w32268 = ( ~w32092 & w32266 ) | ( ~w32092 & w32267 ) | ( w32266 & w32267 ) ;
  assign w32269 = w32267 | w32268 ;
  assign w32270 = \pi085 ^ w32077 ;
  assign w32271 = ( ~w32085 & w32269 ) | ( ~w32085 & w32270 ) | ( w32269 & w32270 ) ;
  assign w32272 = w32270 | w32271 ;
  assign w32273 = \pi086 ^ w32070 ;
  assign w32274 = ( ~w32078 & w32272 ) | ( ~w32078 & w32273 ) | ( w32272 & w32273 ) ;
  assign w32275 = w32273 | w32274 ;
  assign w32276 = \pi087 ^ w32063 ;
  assign w32277 = ( ~w32071 & w32275 ) | ( ~w32071 & w32276 ) | ( w32275 & w32276 ) ;
  assign w32278 = w32276 | w32277 ;
  assign w32279 = \pi088 ^ w32056 ;
  assign w32280 = ( ~w32064 & w32278 ) | ( ~w32064 & w32279 ) | ( w32278 & w32279 ) ;
  assign w32281 = w32279 | w32280 ;
  assign w32282 = \pi089 ^ w32049 ;
  assign w32283 = ( ~w32057 & w32281 ) | ( ~w32057 & w32282 ) | ( w32281 & w32282 ) ;
  assign w32284 = w32282 | w32283 ;
  assign w32285 = \pi090 ^ w32042 ;
  assign w32286 = ( ~w32050 & w32284 ) | ( ~w32050 & w32285 ) | ( w32284 & w32285 ) ;
  assign w32287 = w32285 | w32286 ;
  assign w32288 = \pi091 ^ w32035 ;
  assign w32289 = ( ~w32043 & w32287 ) | ( ~w32043 & w32288 ) | ( w32287 & w32288 ) ;
  assign w32290 = w32288 | w32289 ;
  assign w32291 = \pi092 ^ w32028 ;
  assign w32292 = ( ~w32036 & w32290 ) | ( ~w32036 & w32291 ) | ( w32290 & w32291 ) ;
  assign w32293 = w32291 | w32292 ;
  assign w32294 = \pi093 ^ w32021 ;
  assign w32295 = ( ~w32029 & w32293 ) | ( ~w32029 & w32294 ) | ( w32293 & w32294 ) ;
  assign w32296 = w32294 | w32295 ;
  assign w32297 = \pi094 ^ w32014 ;
  assign w32298 = ( ~w32022 & w32296 ) | ( ~w32022 & w32297 ) | ( w32296 & w32297 ) ;
  assign w32299 = w32297 | w32298 ;
  assign w32300 = \pi095 ^ w32007 ;
  assign w32301 = ( ~w32015 & w32299 ) | ( ~w32015 & w32300 ) | ( w32299 & w32300 ) ;
  assign w32302 = w32300 | w32301 ;
  assign w32303 = \pi096 ^ w32000 ;
  assign w32304 = ( ~w32008 & w32302 ) | ( ~w32008 & w32303 ) | ( w32302 & w32303 ) ;
  assign w32305 = w32303 | w32304 ;
  assign w32306 = \pi097 ^ w31993 ;
  assign w32307 = ( ~w32001 & w32305 ) | ( ~w32001 & w32306 ) | ( w32305 & w32306 ) ;
  assign w32308 = w32306 | w32307 ;
  assign w32309 = \pi098 ^ w31986 ;
  assign w32310 = ( ~w31994 & w32308 ) | ( ~w31994 & w32309 ) | ( w32308 & w32309 ) ;
  assign w32311 = w32309 | w32310 ;
  assign w32312 = \pi099 ^ w31979 ;
  assign w32313 = ( ~w31987 & w32311 ) | ( ~w31987 & w32312 ) | ( w32311 & w32312 ) ;
  assign w32314 = w32312 | w32313 ;
  assign w32315 = \pi100 ^ w31972 ;
  assign w32316 = ( ~w31980 & w32314 ) | ( ~w31980 & w32315 ) | ( w32314 & w32315 ) ;
  assign w32317 = w32315 | w32316 ;
  assign w32318 = \pi101 ^ w31965 ;
  assign w32319 = ( ~w31973 & w32317 ) | ( ~w31973 & w32318 ) | ( w32317 & w32318 ) ;
  assign w32320 = w32318 | w32319 ;
  assign w32321 = \pi102 ^ w31958 ;
  assign w32322 = ( ~w31966 & w32320 ) | ( ~w31966 & w32321 ) | ( w32320 & w32321 ) ;
  assign w32323 = w32321 | w32322 ;
  assign w32324 = \pi103 ^ w31951 ;
  assign w32325 = ( ~w31959 & w32323 ) | ( ~w31959 & w32324 ) | ( w32323 & w32324 ) ;
  assign w32326 = w32324 | w32325 ;
  assign w32327 = \pi104 ^ w31944 ;
  assign w32328 = ( ~w31952 & w32326 ) | ( ~w31952 & w32327 ) | ( w32326 & w32327 ) ;
  assign w32329 = w32327 | w32328 ;
  assign w32330 = \pi105 ^ w31937 ;
  assign w32331 = ( ~w31945 & w32329 ) | ( ~w31945 & w32330 ) | ( w32329 & w32330 ) ;
  assign w32332 = w32330 | w32331 ;
  assign w32333 = \pi106 ^ w31930 ;
  assign w32334 = ( ~w31938 & w32332 ) | ( ~w31938 & w32333 ) | ( w32332 & w32333 ) ;
  assign w32335 = w32333 | w32334 ;
  assign w32336 = \pi107 ^ w31923 ;
  assign w32337 = ( ~w31931 & w32335 ) | ( ~w31931 & w32336 ) | ( w32335 & w32336 ) ;
  assign w32338 = w32336 | w32337 ;
  assign w32339 = \pi108 ^ w31916 ;
  assign w32340 = ( ~w31924 & w32338 ) | ( ~w31924 & w32339 ) | ( w32338 & w32339 ) ;
  assign w32341 = w32339 | w32340 ;
  assign w32342 = \pi109 ^ w31909 ;
  assign w32343 = ( ~w31917 & w32341 ) | ( ~w31917 & w32342 ) | ( w32341 & w32342 ) ;
  assign w32344 = w32342 | w32343 ;
  assign w32345 = \pi110 ^ w31902 ;
  assign w32346 = ( ~w31910 & w32344 ) | ( ~w31910 & w32345 ) | ( w32344 & w32345 ) ;
  assign w32347 = w32345 | w32346 ;
  assign w32348 = \pi111 ^ w31895 ;
  assign w32349 = ( ~w31903 & w32347 ) | ( ~w31903 & w32348 ) | ( w32347 & w32348 ) ;
  assign w32350 = w32348 | w32349 ;
  assign w32351 = \pi112 ^ w31888 ;
  assign w32352 = ( ~w31896 & w32350 ) | ( ~w31896 & w32351 ) | ( w32350 & w32351 ) ;
  assign w32353 = w32351 | w32352 ;
  assign w32354 = \pi113 ^ w31881 ;
  assign w32355 = ( ~w31889 & w32353 ) | ( ~w31889 & w32354 ) | ( w32353 & w32354 ) ;
  assign w32356 = w32354 | w32355 ;
  assign w32357 = ( ~w31428 & w31861 ) | ( ~w31428 & w31875 ) | ( w31861 & w31875 ) ;
  assign w32358 = w31870 ^ w32357 ;
  assign w32359 = ~w31875 & w32358 ;
  assign w32360 = ( w275 & ~w31866 ) | ( w275 & w31873 ) | ( ~w31866 & w31873 ) ;
  assign w32361 = w31866 & w32360 ;
  assign w32362 = w32359 | w32361 ;
  assign w32363 = ~\pi114 & w32362 ;
  assign w32364 = ( \pi114 & ~w32359 ) | ( \pi114 & w32361 ) | ( ~w32359 & w32361 ) ;
  assign w32365 = ~w32361 & w32364 ;
  assign w32366 = w32363 | w32365 ;
  assign w32367 = ( ~w31882 & w32356 ) | ( ~w31882 & w32366 ) | ( w32356 & w32366 ) ;
  assign w32368 = ( w12996 & ~w32366 ) | ( w12996 & w32367 ) | ( ~w32366 & w32367 ) ;
  assign w32369 = w32366 | w32368 ;
  assign w32370 = ~w12496 & w32362 ;
  assign w32371 = w32369 & ~w32370 ;
  assign w32372 = ~w31889 & w32353 ;
  assign w32373 = w32354 ^ w32372 ;
  assign w32374 = ~w32371 & w32373 ;
  assign w32375 = ( w31881 & w32369 ) | ( w31881 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32376 = ~w32370 & w32375 ;
  assign w32377 = w32374 | w32376 ;
  assign w32378 = ( ~w31882 & w32356 ) | ( ~w31882 & w32371 ) | ( w32356 & w32371 ) ;
  assign w32379 = w32366 ^ w32378 ;
  assign w32380 = ~w32371 & w32379 ;
  assign w32381 = ( w12496 & ~w32362 ) | ( w12496 & w32369 ) | ( ~w32362 & w32369 ) ;
  assign w32382 = w32362 & w32381 ;
  assign w32383 = w32380 | w32382 ;
  assign w32384 = ~\pi114 & w32377 ;
  assign w32385 = ~w31896 & w32350 ;
  assign w32386 = w32351 ^ w32385 ;
  assign w32387 = ~w32371 & w32386 ;
  assign w32388 = ( w31888 & w32369 ) | ( w31888 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32389 = ~w32370 & w32388 ;
  assign w32390 = w32387 | w32389 ;
  assign w32391 = ~\pi113 & w32390 ;
  assign w32392 = ~w31903 & w32347 ;
  assign w32393 = w32348 ^ w32392 ;
  assign w32394 = ~w32371 & w32393 ;
  assign w32395 = ( w31895 & w32369 ) | ( w31895 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32396 = ~w32370 & w32395 ;
  assign w32397 = w32394 | w32396 ;
  assign w32398 = ~\pi112 & w32397 ;
  assign w32399 = ~w31910 & w32344 ;
  assign w32400 = w32345 ^ w32399 ;
  assign w32401 = ~w32371 & w32400 ;
  assign w32402 = ( w31902 & w32369 ) | ( w31902 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32403 = ~w32370 & w32402 ;
  assign w32404 = w32401 | w32403 ;
  assign w32405 = ~\pi111 & w32404 ;
  assign w32406 = ~w31917 & w32341 ;
  assign w32407 = w32342 ^ w32406 ;
  assign w32408 = ~w32371 & w32407 ;
  assign w32409 = ( w31909 & w32369 ) | ( w31909 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32410 = ~w32370 & w32409 ;
  assign w32411 = w32408 | w32410 ;
  assign w32412 = ~\pi110 & w32411 ;
  assign w32413 = ~w31924 & w32338 ;
  assign w32414 = w32339 ^ w32413 ;
  assign w32415 = ~w32371 & w32414 ;
  assign w32416 = ( w31916 & w32369 ) | ( w31916 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32417 = ~w32370 & w32416 ;
  assign w32418 = w32415 | w32417 ;
  assign w32419 = ~\pi109 & w32418 ;
  assign w32420 = ~w31931 & w32335 ;
  assign w32421 = w32336 ^ w32420 ;
  assign w32422 = ~w32371 & w32421 ;
  assign w32423 = ( w31923 & w32369 ) | ( w31923 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32424 = ~w32370 & w32423 ;
  assign w32425 = w32422 | w32424 ;
  assign w32426 = ~\pi108 & w32425 ;
  assign w32427 = ~w31938 & w32332 ;
  assign w32428 = w32333 ^ w32427 ;
  assign w32429 = ~w32371 & w32428 ;
  assign w32430 = ( w31930 & w32369 ) | ( w31930 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32431 = ~w32370 & w32430 ;
  assign w32432 = w32429 | w32431 ;
  assign w32433 = ~\pi107 & w32432 ;
  assign w32434 = ~w31945 & w32329 ;
  assign w32435 = w32330 ^ w32434 ;
  assign w32436 = ~w32371 & w32435 ;
  assign w32437 = ( w31937 & w32369 ) | ( w31937 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32438 = ~w32370 & w32437 ;
  assign w32439 = w32436 | w32438 ;
  assign w32440 = ~\pi106 & w32439 ;
  assign w32441 = ~w31952 & w32326 ;
  assign w32442 = w32327 ^ w32441 ;
  assign w32443 = ~w32371 & w32442 ;
  assign w32444 = ( w31944 & w32369 ) | ( w31944 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32445 = ~w32370 & w32444 ;
  assign w32446 = w32443 | w32445 ;
  assign w32447 = ~\pi105 & w32446 ;
  assign w32448 = ~w31959 & w32323 ;
  assign w32449 = w32324 ^ w32448 ;
  assign w32450 = ~w32371 & w32449 ;
  assign w32451 = ( w31951 & w32369 ) | ( w31951 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32452 = ~w32370 & w32451 ;
  assign w32453 = w32450 | w32452 ;
  assign w32454 = ~\pi104 & w32453 ;
  assign w32455 = ~w31966 & w32320 ;
  assign w32456 = w32321 ^ w32455 ;
  assign w32457 = ~w32371 & w32456 ;
  assign w32458 = ( w31958 & w32369 ) | ( w31958 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32459 = ~w32370 & w32458 ;
  assign w32460 = w32457 | w32459 ;
  assign w32461 = ~\pi103 & w32460 ;
  assign w32462 = ~w31973 & w32317 ;
  assign w32463 = w32318 ^ w32462 ;
  assign w32464 = ~w32371 & w32463 ;
  assign w32465 = ( w31965 & w32369 ) | ( w31965 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32466 = ~w32370 & w32465 ;
  assign w32467 = w32464 | w32466 ;
  assign w32468 = ~\pi102 & w32467 ;
  assign w32469 = ~w31980 & w32314 ;
  assign w32470 = w32315 ^ w32469 ;
  assign w32471 = ~w32371 & w32470 ;
  assign w32472 = ( w31972 & w32369 ) | ( w31972 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32473 = ~w32370 & w32472 ;
  assign w32474 = w32471 | w32473 ;
  assign w32475 = ~\pi101 & w32474 ;
  assign w32476 = ~w31987 & w32311 ;
  assign w32477 = w32312 ^ w32476 ;
  assign w32478 = ~w32371 & w32477 ;
  assign w32479 = ( w31979 & w32369 ) | ( w31979 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32480 = ~w32370 & w32479 ;
  assign w32481 = w32478 | w32480 ;
  assign w32482 = ~\pi100 & w32481 ;
  assign w32483 = ~w31994 & w32308 ;
  assign w32484 = w32309 ^ w32483 ;
  assign w32485 = ~w32371 & w32484 ;
  assign w32486 = ( w31986 & w32369 ) | ( w31986 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32487 = ~w32370 & w32486 ;
  assign w32488 = w32485 | w32487 ;
  assign w32489 = ~\pi099 & w32488 ;
  assign w32490 = ~w32001 & w32305 ;
  assign w32491 = w32306 ^ w32490 ;
  assign w32492 = ~w32371 & w32491 ;
  assign w32493 = ( w31993 & w32369 ) | ( w31993 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32494 = ~w32370 & w32493 ;
  assign w32495 = w32492 | w32494 ;
  assign w32496 = ~\pi098 & w32495 ;
  assign w32497 = ~w32008 & w32302 ;
  assign w32498 = w32303 ^ w32497 ;
  assign w32499 = ~w32371 & w32498 ;
  assign w32500 = ( w32000 & w32369 ) | ( w32000 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32501 = ~w32370 & w32500 ;
  assign w32502 = w32499 | w32501 ;
  assign w32503 = ~\pi097 & w32502 ;
  assign w32504 = ~w32015 & w32299 ;
  assign w32505 = w32300 ^ w32504 ;
  assign w32506 = ~w32371 & w32505 ;
  assign w32507 = ( w32007 & w32369 ) | ( w32007 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32508 = ~w32370 & w32507 ;
  assign w32509 = w32506 | w32508 ;
  assign w32510 = ~\pi096 & w32509 ;
  assign w32511 = ~w32022 & w32296 ;
  assign w32512 = w32297 ^ w32511 ;
  assign w32513 = ~w32371 & w32512 ;
  assign w32514 = ( w32014 & w32369 ) | ( w32014 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32515 = ~w32370 & w32514 ;
  assign w32516 = w32513 | w32515 ;
  assign w32517 = ~\pi095 & w32516 ;
  assign w32518 = ~w32029 & w32293 ;
  assign w32519 = w32294 ^ w32518 ;
  assign w32520 = ~w32371 & w32519 ;
  assign w32521 = ( w32021 & w32369 ) | ( w32021 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32522 = ~w32370 & w32521 ;
  assign w32523 = w32520 | w32522 ;
  assign w32524 = ~\pi094 & w32523 ;
  assign w32525 = ~w32036 & w32290 ;
  assign w32526 = w32291 ^ w32525 ;
  assign w32527 = ~w32371 & w32526 ;
  assign w32528 = ( w32028 & w32369 ) | ( w32028 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32529 = ~w32370 & w32528 ;
  assign w32530 = w32527 | w32529 ;
  assign w32531 = ~\pi093 & w32530 ;
  assign w32532 = ~w32043 & w32287 ;
  assign w32533 = w32288 ^ w32532 ;
  assign w32534 = ~w32371 & w32533 ;
  assign w32535 = ( w32035 & w32369 ) | ( w32035 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32536 = ~w32370 & w32535 ;
  assign w32537 = w32534 | w32536 ;
  assign w32538 = ~\pi092 & w32537 ;
  assign w32539 = ~w32050 & w32284 ;
  assign w32540 = w32285 ^ w32539 ;
  assign w32541 = ~w32371 & w32540 ;
  assign w32542 = ( w32042 & w32369 ) | ( w32042 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32543 = ~w32370 & w32542 ;
  assign w32544 = w32541 | w32543 ;
  assign w32545 = ~\pi091 & w32544 ;
  assign w32546 = ~w32057 & w32281 ;
  assign w32547 = w32282 ^ w32546 ;
  assign w32548 = ~w32371 & w32547 ;
  assign w32549 = ( w32049 & w32369 ) | ( w32049 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32550 = ~w32370 & w32549 ;
  assign w32551 = w32548 | w32550 ;
  assign w32552 = ~\pi090 & w32551 ;
  assign w32553 = ~w32064 & w32278 ;
  assign w32554 = w32279 ^ w32553 ;
  assign w32555 = ~w32371 & w32554 ;
  assign w32556 = ( w32056 & w32369 ) | ( w32056 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32557 = ~w32370 & w32556 ;
  assign w32558 = w32555 | w32557 ;
  assign w32559 = ~\pi089 & w32558 ;
  assign w32560 = ~w32071 & w32275 ;
  assign w32561 = w32276 ^ w32560 ;
  assign w32562 = ~w32371 & w32561 ;
  assign w32563 = ( w32063 & w32369 ) | ( w32063 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32564 = ~w32370 & w32563 ;
  assign w32565 = w32562 | w32564 ;
  assign w32566 = ~\pi088 & w32565 ;
  assign w32567 = ~w32078 & w32272 ;
  assign w32568 = w32273 ^ w32567 ;
  assign w32569 = ~w32371 & w32568 ;
  assign w32570 = ( w32070 & w32369 ) | ( w32070 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32571 = ~w32370 & w32570 ;
  assign w32572 = w32569 | w32571 ;
  assign w32573 = ~\pi087 & w32572 ;
  assign w32574 = ~w32085 & w32269 ;
  assign w32575 = w32270 ^ w32574 ;
  assign w32576 = ~w32371 & w32575 ;
  assign w32577 = ( w32077 & w32369 ) | ( w32077 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32578 = ~w32370 & w32577 ;
  assign w32579 = w32576 | w32578 ;
  assign w32580 = ~\pi086 & w32579 ;
  assign w32581 = ~w32092 & w32266 ;
  assign w32582 = w32267 ^ w32581 ;
  assign w32583 = ~w32371 & w32582 ;
  assign w32584 = ( w32084 & w32369 ) | ( w32084 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32585 = ~w32370 & w32584 ;
  assign w32586 = w32583 | w32585 ;
  assign w32587 = ~\pi085 & w32586 ;
  assign w32588 = ~w32099 & w32263 ;
  assign w32589 = w32264 ^ w32588 ;
  assign w32590 = ~w32371 & w32589 ;
  assign w32591 = ( w32091 & w32369 ) | ( w32091 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32592 = ~w32370 & w32591 ;
  assign w32593 = w32590 | w32592 ;
  assign w32594 = ~\pi084 & w32593 ;
  assign w32595 = ~w32106 & w32260 ;
  assign w32596 = w32261 ^ w32595 ;
  assign w32597 = ~w32371 & w32596 ;
  assign w32598 = ( w32098 & w32369 ) | ( w32098 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32599 = ~w32370 & w32598 ;
  assign w32600 = w32597 | w32599 ;
  assign w32601 = ~\pi083 & w32600 ;
  assign w32602 = ~w32113 & w32257 ;
  assign w32603 = w32258 ^ w32602 ;
  assign w32604 = ~w32371 & w32603 ;
  assign w32605 = ( w32105 & w32369 ) | ( w32105 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32606 = ~w32370 & w32605 ;
  assign w32607 = w32604 | w32606 ;
  assign w32608 = ~\pi082 & w32607 ;
  assign w32609 = ~w32120 & w32254 ;
  assign w32610 = w32255 ^ w32609 ;
  assign w32611 = ~w32371 & w32610 ;
  assign w32612 = ( w32112 & w32369 ) | ( w32112 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32613 = ~w32370 & w32612 ;
  assign w32614 = w32611 | w32613 ;
  assign w32615 = ~\pi081 & w32614 ;
  assign w32616 = ~w32127 & w32251 ;
  assign w32617 = w32252 ^ w32616 ;
  assign w32618 = ~w32371 & w32617 ;
  assign w32619 = ( w32119 & w32369 ) | ( w32119 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32620 = ~w32370 & w32619 ;
  assign w32621 = w32618 | w32620 ;
  assign w32622 = ~\pi080 & w32621 ;
  assign w32623 = ~w32134 & w32248 ;
  assign w32624 = w32249 ^ w32623 ;
  assign w32625 = ~w32371 & w32624 ;
  assign w32626 = ( w32126 & w32369 ) | ( w32126 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32627 = ~w32370 & w32626 ;
  assign w32628 = w32625 | w32627 ;
  assign w32629 = ~\pi079 & w32628 ;
  assign w32630 = ~w32141 & w32245 ;
  assign w32631 = w32246 ^ w32630 ;
  assign w32632 = ~w32371 & w32631 ;
  assign w32633 = ( w32133 & w32369 ) | ( w32133 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32634 = ~w32370 & w32633 ;
  assign w32635 = w32632 | w32634 ;
  assign w32636 = ~\pi078 & w32635 ;
  assign w32637 = ~w32148 & w32242 ;
  assign w32638 = w32243 ^ w32637 ;
  assign w32639 = ~w32371 & w32638 ;
  assign w32640 = ( w32140 & w32369 ) | ( w32140 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32641 = ~w32370 & w32640 ;
  assign w32642 = w32639 | w32641 ;
  assign w32643 = ~\pi077 & w32642 ;
  assign w32644 = ~w32155 & w32239 ;
  assign w32645 = w32240 ^ w32644 ;
  assign w32646 = ~w32371 & w32645 ;
  assign w32647 = ( w32147 & w32369 ) | ( w32147 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32648 = ~w32370 & w32647 ;
  assign w32649 = w32646 | w32648 ;
  assign w32650 = ~\pi076 & w32649 ;
  assign w32651 = ~w32162 & w32236 ;
  assign w32652 = w32237 ^ w32651 ;
  assign w32653 = ~w32371 & w32652 ;
  assign w32654 = ( w32154 & w32369 ) | ( w32154 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32655 = ~w32370 & w32654 ;
  assign w32656 = w32653 | w32655 ;
  assign w32657 = ~\pi075 & w32656 ;
  assign w32658 = ~w32169 & w32233 ;
  assign w32659 = w32234 ^ w32658 ;
  assign w32660 = ~w32371 & w32659 ;
  assign w32661 = ( w32161 & w32369 ) | ( w32161 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32662 = ~w32370 & w32661 ;
  assign w32663 = w32660 | w32662 ;
  assign w32664 = ~\pi074 & w32663 ;
  assign w32665 = ~w32176 & w32230 ;
  assign w32666 = w32231 ^ w32665 ;
  assign w32667 = ~w32371 & w32666 ;
  assign w32668 = ( w32168 & w32369 ) | ( w32168 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32669 = ~w32370 & w32668 ;
  assign w32670 = w32667 | w32669 ;
  assign w32671 = ~\pi073 & w32670 ;
  assign w32672 = ~w32183 & w32227 ;
  assign w32673 = w32228 ^ w32672 ;
  assign w32674 = ~w32371 & w32673 ;
  assign w32675 = ( w32175 & w32369 ) | ( w32175 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32676 = ~w32370 & w32675 ;
  assign w32677 = w32674 | w32676 ;
  assign w32678 = ~\pi072 & w32677 ;
  assign w32679 = ~w32190 & w32224 ;
  assign w32680 = w32225 ^ w32679 ;
  assign w32681 = ~w32371 & w32680 ;
  assign w32682 = ( w32182 & w32369 ) | ( w32182 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32683 = ~w32370 & w32682 ;
  assign w32684 = w32681 | w32683 ;
  assign w32685 = ~\pi071 & w32684 ;
  assign w32686 = ~w32197 & w32221 ;
  assign w32687 = w32222 ^ w32686 ;
  assign w32688 = ~w32371 & w32687 ;
  assign w32689 = ( w32189 & w32369 ) | ( w32189 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32690 = ~w32370 & w32689 ;
  assign w32691 = w32688 | w32690 ;
  assign w32692 = ~\pi070 & w32691 ;
  assign w32693 = ~w32203 & w32218 ;
  assign w32694 = w32219 ^ w32693 ;
  assign w32695 = ~w32371 & w32694 ;
  assign w32696 = ( w32196 & w32369 ) | ( w32196 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32697 = ~w32370 & w32696 ;
  assign w32698 = w32695 | w32697 ;
  assign w32699 = ~\pi069 & w32698 ;
  assign w32700 = ~w32208 & w32215 ;
  assign w32701 = w32216 ^ w32700 ;
  assign w32702 = ~w32371 & w32701 ;
  assign w32703 = ( w32202 & w32369 ) | ( w32202 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32704 = ~w32370 & w32703 ;
  assign w32705 = w32702 | w32704 ;
  assign w32706 = ~\pi068 & w32705 ;
  assign w32707 = \pi064 & ~w31875 ;
  assign w32708 = \pi014 ^ w32707 ;
  assign w32709 = ( \pi065 & w13338 ) | ( \pi065 & ~w32708 ) | ( w13338 & ~w32708 ) ;
  assign w32710 = w32211 ^ w32709 ;
  assign w32711 = ~w32371 & w32710 ;
  assign w32712 = ( w32207 & w32369 ) | ( w32207 & w32370 ) | ( w32369 & w32370 ) ;
  assign w32713 = ~w32370 & w32712 ;
  assign w32714 = w32711 | w32713 ;
  assign w32715 = ~\pi067 & w32714 ;
  assign w32716 = \pi013 ^ w31875 ;
  assign w32717 = ( \pi064 & w32371 ) | ( \pi064 & w32716 ) | ( w32371 & w32716 ) ;
  assign w32718 = w13346 ^ w32717 ;
  assign w32719 = ~w32371 & w32718 ;
  assign w32720 = w32371 & w32708 ;
  assign w32721 = w32719 | w32720 ;
  assign w32722 = ~\pi066 & w32721 ;
  assign w32723 = \pi066 ^ w32721 ;
  assign w32724 = ( \pi064 & ~w32371 ) | ( \pi064 & w32723 ) | ( ~w32371 & w32723 ) ;
  assign w32725 = \pi013 ^ w32724 ;
  assign w32726 = ( \pi065 & w13798 ) | ( \pi065 & ~w32725 ) | ( w13798 & ~w32725 ) ;
  assign w32727 = w32723 | w32726 ;
  assign w32728 = \pi067 ^ w32714 ;
  assign w32729 = ( ~w32722 & w32727 ) | ( ~w32722 & w32728 ) | ( w32727 & w32728 ) ;
  assign w32730 = w32728 | w32729 ;
  assign w32731 = \pi068 ^ w32705 ;
  assign w32732 = ( ~w32715 & w32730 ) | ( ~w32715 & w32731 ) | ( w32730 & w32731 ) ;
  assign w32733 = w32731 | w32732 ;
  assign w32734 = \pi069 ^ w32698 ;
  assign w32735 = ( ~w32706 & w32733 ) | ( ~w32706 & w32734 ) | ( w32733 & w32734 ) ;
  assign w32736 = w32734 | w32735 ;
  assign w32737 = \pi070 ^ w32691 ;
  assign w32738 = ( ~w32699 & w32736 ) | ( ~w32699 & w32737 ) | ( w32736 & w32737 ) ;
  assign w32739 = w32737 | w32738 ;
  assign w32740 = \pi071 ^ w32684 ;
  assign w32741 = ( ~w32692 & w32739 ) | ( ~w32692 & w32740 ) | ( w32739 & w32740 ) ;
  assign w32742 = w32740 | w32741 ;
  assign w32743 = \pi072 ^ w32677 ;
  assign w32744 = ( ~w32685 & w32742 ) | ( ~w32685 & w32743 ) | ( w32742 & w32743 ) ;
  assign w32745 = w32743 | w32744 ;
  assign w32746 = \pi073 ^ w32670 ;
  assign w32747 = ( ~w32678 & w32745 ) | ( ~w32678 & w32746 ) | ( w32745 & w32746 ) ;
  assign w32748 = w32746 | w32747 ;
  assign w32749 = \pi074 ^ w32663 ;
  assign w32750 = ( ~w32671 & w32748 ) | ( ~w32671 & w32749 ) | ( w32748 & w32749 ) ;
  assign w32751 = w32749 | w32750 ;
  assign w32752 = \pi075 ^ w32656 ;
  assign w32753 = ( ~w32664 & w32751 ) | ( ~w32664 & w32752 ) | ( w32751 & w32752 ) ;
  assign w32754 = w32752 | w32753 ;
  assign w32755 = \pi076 ^ w32649 ;
  assign w32756 = ( ~w32657 & w32754 ) | ( ~w32657 & w32755 ) | ( w32754 & w32755 ) ;
  assign w32757 = w32755 | w32756 ;
  assign w32758 = \pi077 ^ w32642 ;
  assign w32759 = ( ~w32650 & w32757 ) | ( ~w32650 & w32758 ) | ( w32757 & w32758 ) ;
  assign w32760 = w32758 | w32759 ;
  assign w32761 = \pi078 ^ w32635 ;
  assign w32762 = ( ~w32643 & w32760 ) | ( ~w32643 & w32761 ) | ( w32760 & w32761 ) ;
  assign w32763 = w32761 | w32762 ;
  assign w32764 = \pi079 ^ w32628 ;
  assign w32765 = ( ~w32636 & w32763 ) | ( ~w32636 & w32764 ) | ( w32763 & w32764 ) ;
  assign w32766 = w32764 | w32765 ;
  assign w32767 = \pi080 ^ w32621 ;
  assign w32768 = ( ~w32629 & w32766 ) | ( ~w32629 & w32767 ) | ( w32766 & w32767 ) ;
  assign w32769 = w32767 | w32768 ;
  assign w32770 = \pi081 ^ w32614 ;
  assign w32771 = ( ~w32622 & w32769 ) | ( ~w32622 & w32770 ) | ( w32769 & w32770 ) ;
  assign w32772 = w32770 | w32771 ;
  assign w32773 = \pi082 ^ w32607 ;
  assign w32774 = ( ~w32615 & w32772 ) | ( ~w32615 & w32773 ) | ( w32772 & w32773 ) ;
  assign w32775 = w32773 | w32774 ;
  assign w32776 = \pi083 ^ w32600 ;
  assign w32777 = ( ~w32608 & w32775 ) | ( ~w32608 & w32776 ) | ( w32775 & w32776 ) ;
  assign w32778 = w32776 | w32777 ;
  assign w32779 = \pi084 ^ w32593 ;
  assign w32780 = ( ~w32601 & w32778 ) | ( ~w32601 & w32779 ) | ( w32778 & w32779 ) ;
  assign w32781 = w32779 | w32780 ;
  assign w32782 = \pi085 ^ w32586 ;
  assign w32783 = ( ~w32594 & w32781 ) | ( ~w32594 & w32782 ) | ( w32781 & w32782 ) ;
  assign w32784 = w32782 | w32783 ;
  assign w32785 = \pi086 ^ w32579 ;
  assign w32786 = ( ~w32587 & w32784 ) | ( ~w32587 & w32785 ) | ( w32784 & w32785 ) ;
  assign w32787 = w32785 | w32786 ;
  assign w32788 = \pi087 ^ w32572 ;
  assign w32789 = ( ~w32580 & w32787 ) | ( ~w32580 & w32788 ) | ( w32787 & w32788 ) ;
  assign w32790 = w32788 | w32789 ;
  assign w32791 = \pi088 ^ w32565 ;
  assign w32792 = ( ~w32573 & w32790 ) | ( ~w32573 & w32791 ) | ( w32790 & w32791 ) ;
  assign w32793 = w32791 | w32792 ;
  assign w32794 = \pi089 ^ w32558 ;
  assign w32795 = ( ~w32566 & w32793 ) | ( ~w32566 & w32794 ) | ( w32793 & w32794 ) ;
  assign w32796 = w32794 | w32795 ;
  assign w32797 = \pi090 ^ w32551 ;
  assign w32798 = ( ~w32559 & w32796 ) | ( ~w32559 & w32797 ) | ( w32796 & w32797 ) ;
  assign w32799 = w32797 | w32798 ;
  assign w32800 = \pi091 ^ w32544 ;
  assign w32801 = ( ~w32552 & w32799 ) | ( ~w32552 & w32800 ) | ( w32799 & w32800 ) ;
  assign w32802 = w32800 | w32801 ;
  assign w32803 = \pi092 ^ w32537 ;
  assign w32804 = ( ~w32545 & w32802 ) | ( ~w32545 & w32803 ) | ( w32802 & w32803 ) ;
  assign w32805 = w32803 | w32804 ;
  assign w32806 = \pi093 ^ w32530 ;
  assign w32807 = ( ~w32538 & w32805 ) | ( ~w32538 & w32806 ) | ( w32805 & w32806 ) ;
  assign w32808 = w32806 | w32807 ;
  assign w32809 = \pi094 ^ w32523 ;
  assign w32810 = ( ~w32531 & w32808 ) | ( ~w32531 & w32809 ) | ( w32808 & w32809 ) ;
  assign w32811 = w32809 | w32810 ;
  assign w32812 = \pi095 ^ w32516 ;
  assign w32813 = ( ~w32524 & w32811 ) | ( ~w32524 & w32812 ) | ( w32811 & w32812 ) ;
  assign w32814 = w32812 | w32813 ;
  assign w32815 = \pi096 ^ w32509 ;
  assign w32816 = ( ~w32517 & w32814 ) | ( ~w32517 & w32815 ) | ( w32814 & w32815 ) ;
  assign w32817 = w32815 | w32816 ;
  assign w32818 = \pi097 ^ w32502 ;
  assign w32819 = ( ~w32510 & w32817 ) | ( ~w32510 & w32818 ) | ( w32817 & w32818 ) ;
  assign w32820 = w32818 | w32819 ;
  assign w32821 = \pi098 ^ w32495 ;
  assign w32822 = ( ~w32503 & w32820 ) | ( ~w32503 & w32821 ) | ( w32820 & w32821 ) ;
  assign w32823 = w32821 | w32822 ;
  assign w32824 = \pi099 ^ w32488 ;
  assign w32825 = ( ~w32496 & w32823 ) | ( ~w32496 & w32824 ) | ( w32823 & w32824 ) ;
  assign w32826 = w32824 | w32825 ;
  assign w32827 = \pi100 ^ w32481 ;
  assign w32828 = ( ~w32489 & w32826 ) | ( ~w32489 & w32827 ) | ( w32826 & w32827 ) ;
  assign w32829 = w32827 | w32828 ;
  assign w32830 = \pi101 ^ w32474 ;
  assign w32831 = ( ~w32482 & w32829 ) | ( ~w32482 & w32830 ) | ( w32829 & w32830 ) ;
  assign w32832 = w32830 | w32831 ;
  assign w32833 = \pi102 ^ w32467 ;
  assign w32834 = ( ~w32475 & w32832 ) | ( ~w32475 & w32833 ) | ( w32832 & w32833 ) ;
  assign w32835 = w32833 | w32834 ;
  assign w32836 = \pi103 ^ w32460 ;
  assign w32837 = ( ~w32468 & w32835 ) | ( ~w32468 & w32836 ) | ( w32835 & w32836 ) ;
  assign w32838 = w32836 | w32837 ;
  assign w32839 = \pi104 ^ w32453 ;
  assign w32840 = ( ~w32461 & w32838 ) | ( ~w32461 & w32839 ) | ( w32838 & w32839 ) ;
  assign w32841 = w32839 | w32840 ;
  assign w32842 = \pi105 ^ w32446 ;
  assign w32843 = ( ~w32454 & w32841 ) | ( ~w32454 & w32842 ) | ( w32841 & w32842 ) ;
  assign w32844 = w32842 | w32843 ;
  assign w32845 = \pi106 ^ w32439 ;
  assign w32846 = ( ~w32447 & w32844 ) | ( ~w32447 & w32845 ) | ( w32844 & w32845 ) ;
  assign w32847 = w32845 | w32846 ;
  assign w32848 = \pi107 ^ w32432 ;
  assign w32849 = ( ~w32440 & w32847 ) | ( ~w32440 & w32848 ) | ( w32847 & w32848 ) ;
  assign w32850 = w32848 | w32849 ;
  assign w32851 = \pi108 ^ w32425 ;
  assign w32852 = ( ~w32433 & w32850 ) | ( ~w32433 & w32851 ) | ( w32850 & w32851 ) ;
  assign w32853 = w32851 | w32852 ;
  assign w32854 = \pi109 ^ w32418 ;
  assign w32855 = ( ~w32426 & w32853 ) | ( ~w32426 & w32854 ) | ( w32853 & w32854 ) ;
  assign w32856 = w32854 | w32855 ;
  assign w32857 = \pi110 ^ w32411 ;
  assign w32858 = ( ~w32419 & w32856 ) | ( ~w32419 & w32857 ) | ( w32856 & w32857 ) ;
  assign w32859 = w32857 | w32858 ;
  assign w32860 = \pi111 ^ w32404 ;
  assign w32861 = ( ~w32412 & w32859 ) | ( ~w32412 & w32860 ) | ( w32859 & w32860 ) ;
  assign w32862 = w32860 | w32861 ;
  assign w32863 = \pi112 ^ w32397 ;
  assign w32864 = ( ~w32405 & w32862 ) | ( ~w32405 & w32863 ) | ( w32862 & w32863 ) ;
  assign w32865 = w32863 | w32864 ;
  assign w32866 = \pi113 ^ w32390 ;
  assign w32867 = ( ~w32398 & w32865 ) | ( ~w32398 & w32866 ) | ( w32865 & w32866 ) ;
  assign w32868 = w32866 | w32867 ;
  assign w32869 = \pi114 ^ w32377 ;
  assign w32870 = ( ~w32391 & w32868 ) | ( ~w32391 & w32869 ) | ( w32868 & w32869 ) ;
  assign w32871 = w32869 | w32870 ;
  assign w32872 = \pi115 ^ w32383 ;
  assign w32873 = w32384 & ~w32872 ;
  assign w32874 = ( w32871 & w32872 ) | ( w32871 & ~w32873 ) | ( w32872 & ~w32873 ) ;
  assign w32875 = ~\pi115 & w32383 ;
  assign w32876 = w32874 & ~w32875 ;
  assign w32877 = w155 | w32876 ;
  assign w32878 = w32377 & w32877 ;
  assign w32879 = ~w32391 & w32868 ;
  assign w32880 = w32869 ^ w32879 ;
  assign w32881 = ~w32877 & w32880 ;
  assign w32882 = w32878 | w32881 ;
  assign w32883 = ~\pi115 & w32882 ;
  assign w32884 = w32390 & w32877 ;
  assign w32885 = ~w32398 & w32865 ;
  assign w32886 = w32866 ^ w32885 ;
  assign w32887 = ~w32877 & w32886 ;
  assign w32888 = w32884 | w32887 ;
  assign w32889 = ~\pi114 & w32888 ;
  assign w32890 = w32397 & w32877 ;
  assign w32891 = ~w32405 & w32862 ;
  assign w32892 = w32863 ^ w32891 ;
  assign w32893 = ~w32877 & w32892 ;
  assign w32894 = w32890 | w32893 ;
  assign w32895 = ~\pi113 & w32894 ;
  assign w32896 = w32404 & w32877 ;
  assign w32897 = ~w32412 & w32859 ;
  assign w32898 = w32860 ^ w32897 ;
  assign w32899 = ~w32877 & w32898 ;
  assign w32900 = w32896 | w32899 ;
  assign w32901 = ~\pi112 & w32900 ;
  assign w32902 = w32411 & w32877 ;
  assign w32903 = ~w32419 & w32856 ;
  assign w32904 = w32857 ^ w32903 ;
  assign w32905 = ~w32877 & w32904 ;
  assign w32906 = w32902 | w32905 ;
  assign w32907 = ~\pi111 & w32906 ;
  assign w32908 = w32418 & w32877 ;
  assign w32909 = ~w32426 & w32853 ;
  assign w32910 = w32854 ^ w32909 ;
  assign w32911 = ~w32877 & w32910 ;
  assign w32912 = w32908 | w32911 ;
  assign w32913 = ~\pi110 & w32912 ;
  assign w32914 = w32425 & w32877 ;
  assign w32915 = ~w32433 & w32850 ;
  assign w32916 = w32851 ^ w32915 ;
  assign w32917 = ~w32877 & w32916 ;
  assign w32918 = w32914 | w32917 ;
  assign w32919 = ~\pi109 & w32918 ;
  assign w32920 = w32432 & w32877 ;
  assign w32921 = ~w32440 & w32847 ;
  assign w32922 = w32848 ^ w32921 ;
  assign w32923 = ~w32877 & w32922 ;
  assign w32924 = w32920 | w32923 ;
  assign w32925 = ~\pi108 & w32924 ;
  assign w32926 = w32439 & w32877 ;
  assign w32927 = ~w32447 & w32844 ;
  assign w32928 = w32845 ^ w32927 ;
  assign w32929 = ~w32877 & w32928 ;
  assign w32930 = w32926 | w32929 ;
  assign w32931 = ~\pi107 & w32930 ;
  assign w32932 = w32446 & w32877 ;
  assign w32933 = ~w32454 & w32841 ;
  assign w32934 = w32842 ^ w32933 ;
  assign w32935 = ~w32877 & w32934 ;
  assign w32936 = w32932 | w32935 ;
  assign w32937 = ~\pi106 & w32936 ;
  assign w32938 = w32453 & w32877 ;
  assign w32939 = ~w32461 & w32838 ;
  assign w32940 = w32839 ^ w32939 ;
  assign w32941 = ~w32877 & w32940 ;
  assign w32942 = w32938 | w32941 ;
  assign w32943 = ~\pi105 & w32942 ;
  assign w32944 = w32460 & w32877 ;
  assign w32945 = ~w32468 & w32835 ;
  assign w32946 = w32836 ^ w32945 ;
  assign w32947 = ~w32877 & w32946 ;
  assign w32948 = w32944 | w32947 ;
  assign w32949 = ~\pi104 & w32948 ;
  assign w32950 = w32467 & w32877 ;
  assign w32951 = ~w32475 & w32832 ;
  assign w32952 = w32833 ^ w32951 ;
  assign w32953 = ~w32877 & w32952 ;
  assign w32954 = w32950 | w32953 ;
  assign w32955 = ~\pi103 & w32954 ;
  assign w32956 = w32474 & w32877 ;
  assign w32957 = ~w32482 & w32829 ;
  assign w32958 = w32830 ^ w32957 ;
  assign w32959 = ~w32877 & w32958 ;
  assign w32960 = w32956 | w32959 ;
  assign w32961 = ~\pi102 & w32960 ;
  assign w32962 = w32481 & w32877 ;
  assign w32963 = ~w32489 & w32826 ;
  assign w32964 = w32827 ^ w32963 ;
  assign w32965 = ~w32877 & w32964 ;
  assign w32966 = w32962 | w32965 ;
  assign w32967 = ~\pi101 & w32966 ;
  assign w32968 = w32488 & w32877 ;
  assign w32969 = ~w32496 & w32823 ;
  assign w32970 = w32824 ^ w32969 ;
  assign w32971 = ~w32877 & w32970 ;
  assign w32972 = w32968 | w32971 ;
  assign w32973 = ~\pi100 & w32972 ;
  assign w32974 = w32495 & w32877 ;
  assign w32975 = ~w32503 & w32820 ;
  assign w32976 = w32821 ^ w32975 ;
  assign w32977 = ~w32877 & w32976 ;
  assign w32978 = w32974 | w32977 ;
  assign w32979 = ~\pi099 & w32978 ;
  assign w32980 = w32502 & w32877 ;
  assign w32981 = ~w32510 & w32817 ;
  assign w32982 = w32818 ^ w32981 ;
  assign w32983 = ~w32877 & w32982 ;
  assign w32984 = w32980 | w32983 ;
  assign w32985 = ~\pi098 & w32984 ;
  assign w32986 = w32509 & w32877 ;
  assign w32987 = ~w32517 & w32814 ;
  assign w32988 = w32815 ^ w32987 ;
  assign w32989 = ~w32877 & w32988 ;
  assign w32990 = w32986 | w32989 ;
  assign w32991 = ~\pi097 & w32990 ;
  assign w32992 = w32516 & w32877 ;
  assign w32993 = ~w32524 & w32811 ;
  assign w32994 = w32812 ^ w32993 ;
  assign w32995 = ~w32877 & w32994 ;
  assign w32996 = w32992 | w32995 ;
  assign w32997 = ~\pi096 & w32996 ;
  assign w32998 = w32523 & w32877 ;
  assign w32999 = ~w32531 & w32808 ;
  assign w33000 = w32809 ^ w32999 ;
  assign w33001 = ~w32877 & w33000 ;
  assign w33002 = w32998 | w33001 ;
  assign w33003 = ~\pi095 & w33002 ;
  assign w33004 = w32530 & w32877 ;
  assign w33005 = ~w32538 & w32805 ;
  assign w33006 = w32806 ^ w33005 ;
  assign w33007 = ~w32877 & w33006 ;
  assign w33008 = w33004 | w33007 ;
  assign w33009 = ~\pi094 & w33008 ;
  assign w33010 = w32537 & w32877 ;
  assign w33011 = ~w32545 & w32802 ;
  assign w33012 = w32803 ^ w33011 ;
  assign w33013 = ~w32877 & w33012 ;
  assign w33014 = w33010 | w33013 ;
  assign w33015 = ~\pi093 & w33014 ;
  assign w33016 = w32544 & w32877 ;
  assign w33017 = ~w32552 & w32799 ;
  assign w33018 = w32800 ^ w33017 ;
  assign w33019 = ~w32877 & w33018 ;
  assign w33020 = w33016 | w33019 ;
  assign w33021 = ~\pi092 & w33020 ;
  assign w33022 = w32551 & w32877 ;
  assign w33023 = ~w32559 & w32796 ;
  assign w33024 = w32797 ^ w33023 ;
  assign w33025 = ~w32877 & w33024 ;
  assign w33026 = w33022 | w33025 ;
  assign w33027 = ~\pi091 & w33026 ;
  assign w33028 = w32558 & w32877 ;
  assign w33029 = ~w32566 & w32793 ;
  assign w33030 = w32794 ^ w33029 ;
  assign w33031 = ~w32877 & w33030 ;
  assign w33032 = w33028 | w33031 ;
  assign w33033 = ~\pi090 & w33032 ;
  assign w33034 = w32565 & w32877 ;
  assign w33035 = ~w32573 & w32790 ;
  assign w33036 = w32791 ^ w33035 ;
  assign w33037 = ~w32877 & w33036 ;
  assign w33038 = w33034 | w33037 ;
  assign w33039 = ~\pi089 & w33038 ;
  assign w33040 = w32572 & w32877 ;
  assign w33041 = ~w32580 & w32787 ;
  assign w33042 = w32788 ^ w33041 ;
  assign w33043 = ~w32877 & w33042 ;
  assign w33044 = w33040 | w33043 ;
  assign w33045 = ~\pi088 & w33044 ;
  assign w33046 = w32579 & w32877 ;
  assign w33047 = ~w32587 & w32784 ;
  assign w33048 = w32785 ^ w33047 ;
  assign w33049 = ~w32877 & w33048 ;
  assign w33050 = w33046 | w33049 ;
  assign w33051 = ~\pi087 & w33050 ;
  assign w33052 = w32586 & w32877 ;
  assign w33053 = ~w32594 & w32781 ;
  assign w33054 = w32782 ^ w33053 ;
  assign w33055 = ~w32877 & w33054 ;
  assign w33056 = w33052 | w33055 ;
  assign w33057 = ~\pi086 & w33056 ;
  assign w33058 = w32593 & w32877 ;
  assign w33059 = ~w32601 & w32778 ;
  assign w33060 = w32779 ^ w33059 ;
  assign w33061 = ~w32877 & w33060 ;
  assign w33062 = w33058 | w33061 ;
  assign w33063 = ~\pi085 & w33062 ;
  assign w33064 = w32600 & w32877 ;
  assign w33065 = ~w32608 & w32775 ;
  assign w33066 = w32776 ^ w33065 ;
  assign w33067 = ~w32877 & w33066 ;
  assign w33068 = w33064 | w33067 ;
  assign w33069 = ~\pi084 & w33068 ;
  assign w33070 = w32607 & w32877 ;
  assign w33071 = ~w32615 & w32772 ;
  assign w33072 = w32773 ^ w33071 ;
  assign w33073 = ~w32877 & w33072 ;
  assign w33074 = w33070 | w33073 ;
  assign w33075 = ~\pi083 & w33074 ;
  assign w33076 = w32614 & w32877 ;
  assign w33077 = ~w32622 & w32769 ;
  assign w33078 = w32770 ^ w33077 ;
  assign w33079 = ~w32877 & w33078 ;
  assign w33080 = w33076 | w33079 ;
  assign w33081 = ~\pi082 & w33080 ;
  assign w33082 = w32621 & w32877 ;
  assign w33083 = ~w32629 & w32766 ;
  assign w33084 = w32767 ^ w33083 ;
  assign w33085 = ~w32877 & w33084 ;
  assign w33086 = w33082 | w33085 ;
  assign w33087 = ~\pi081 & w33086 ;
  assign w33088 = w32628 & w32877 ;
  assign w33089 = ~w32636 & w32763 ;
  assign w33090 = w32764 ^ w33089 ;
  assign w33091 = ~w32877 & w33090 ;
  assign w33092 = w33088 | w33091 ;
  assign w33093 = ~\pi080 & w33092 ;
  assign w33094 = w32635 & w32877 ;
  assign w33095 = ~w32643 & w32760 ;
  assign w33096 = w32761 ^ w33095 ;
  assign w33097 = ~w32877 & w33096 ;
  assign w33098 = w33094 | w33097 ;
  assign w33099 = ~\pi079 & w33098 ;
  assign w33100 = w32642 & w32877 ;
  assign w33101 = ~w32650 & w32757 ;
  assign w33102 = w32758 ^ w33101 ;
  assign w33103 = ~w32877 & w33102 ;
  assign w33104 = w33100 | w33103 ;
  assign w33105 = ~\pi078 & w33104 ;
  assign w33106 = w32649 & w32877 ;
  assign w33107 = ~w32657 & w32754 ;
  assign w33108 = w32755 ^ w33107 ;
  assign w33109 = ~w32877 & w33108 ;
  assign w33110 = w33106 | w33109 ;
  assign w33111 = ~\pi077 & w33110 ;
  assign w33112 = w32656 & w32877 ;
  assign w33113 = ~w32664 & w32751 ;
  assign w33114 = w32752 ^ w33113 ;
  assign w33115 = ~w32877 & w33114 ;
  assign w33116 = w33112 | w33115 ;
  assign w33117 = ~\pi076 & w33116 ;
  assign w33118 = w32663 & w32877 ;
  assign w33119 = ~w32671 & w32748 ;
  assign w33120 = w32749 ^ w33119 ;
  assign w33121 = ~w32877 & w33120 ;
  assign w33122 = w33118 | w33121 ;
  assign w33123 = ~\pi075 & w33122 ;
  assign w33124 = w32670 & w32877 ;
  assign w33125 = ~w32678 & w32745 ;
  assign w33126 = w32746 ^ w33125 ;
  assign w33127 = ~w32877 & w33126 ;
  assign w33128 = w33124 | w33127 ;
  assign w33129 = ~\pi074 & w33128 ;
  assign w33130 = w32677 & w32877 ;
  assign w33131 = ~w32685 & w32742 ;
  assign w33132 = w32743 ^ w33131 ;
  assign w33133 = ~w32877 & w33132 ;
  assign w33134 = w33130 | w33133 ;
  assign w33135 = ~\pi073 & w33134 ;
  assign w33136 = w32684 & w32877 ;
  assign w33137 = ~w32692 & w32739 ;
  assign w33138 = w32740 ^ w33137 ;
  assign w33139 = ~w32877 & w33138 ;
  assign w33140 = w33136 | w33139 ;
  assign w33141 = ~\pi072 & w33140 ;
  assign w33142 = w32691 & w32877 ;
  assign w33143 = ~w32699 & w32736 ;
  assign w33144 = w32737 ^ w33143 ;
  assign w33145 = ~w32877 & w33144 ;
  assign w33146 = w33142 | w33145 ;
  assign w33147 = ~\pi071 & w33146 ;
  assign w33148 = w32698 & w32877 ;
  assign w33149 = ~w32706 & w32733 ;
  assign w33150 = w32734 ^ w33149 ;
  assign w33151 = ~w32877 & w33150 ;
  assign w33152 = w33148 | w33151 ;
  assign w33153 = ~\pi070 & w33152 ;
  assign w33154 = w32705 & w32877 ;
  assign w33155 = ~w32715 & w32730 ;
  assign w33156 = w32731 ^ w33155 ;
  assign w33157 = ~w32877 & w33156 ;
  assign w33158 = w33154 | w33157 ;
  assign w33159 = ~\pi069 & w33158 ;
  assign w33160 = w32714 & w32877 ;
  assign w33161 = ~w32722 & w32727 ;
  assign w33162 = w32728 ^ w33161 ;
  assign w33163 = ~w32877 & w33162 ;
  assign w33164 = w33160 | w33163 ;
  assign w33165 = ~\pi068 & w33164 ;
  assign w33166 = \pi064 & ~w32371 ;
  assign w33167 = \pi013 ^ w33166 ;
  assign w33168 = ( \pi065 & w13798 ) | ( \pi065 & ~w33167 ) | ( w13798 & ~w33167 ) ;
  assign w33169 = w32723 ^ w33168 ;
  assign w33170 = ( w155 & w32876 ) | ( w155 & w33169 ) | ( w32876 & w33169 ) ;
  assign w33171 = w33169 & ~w33170 ;
  assign w33172 = ( w32721 & w32877 ) | ( w32721 & w33171 ) | ( w32877 & w33171 ) ;
  assign w33173 = w33171 | w33172 ;
  assign w33174 = ~\pi067 & w33173 ;
  assign w33175 = \pi012 ^ w32371 ;
  assign w33176 = ( \pi064 & w155 ) | ( \pi064 & w33175 ) | ( w155 & w33175 ) ;
  assign w33177 = w13806 ^ w33176 ;
  assign w33178 = ~w155 & w33177 ;
  assign w33179 = ~w32876 & w33178 ;
  assign w33180 = ( ~\pi064 & w32371 ) | ( ~\pi064 & w32877 ) | ( w32371 & w32877 ) ;
  assign w33181 = \pi013 ^ w33180 ;
  assign w33182 = w32877 & ~w33181 ;
  assign w33183 = w33179 | w33182 ;
  assign w33184 = ~\pi066 & w33183 ;
  assign w33185 = ( \pi064 & w13819 ) | ( \pi064 & w32876 ) | ( w13819 & w32876 ) ;
  assign w33186 = ( \pi012 & ~\pi064 ) | ( \pi012 & w33185 ) | ( ~\pi064 & w33185 ) ;
  assign w33187 = ( w153 & ~w199 ) | ( w153 & w32876 ) | ( ~w199 & w32876 ) ;
  assign w33188 = w13822 & ~w33187 ;
  assign w33189 = w32877 | w33179 ;
  assign w33190 = ( w33167 & w33179 ) | ( w33167 & w33189 ) | ( w33179 & w33189 ) ;
  assign w33191 = \pi066 ^ w33190 ;
  assign w33192 = w33186 | w33188 ;
  assign w33193 = ( \pi065 & w13825 ) | ( \pi065 & ~w33192 ) | ( w13825 & ~w33192 ) ;
  assign w33194 = w33191 | w33193 ;
  assign w33195 = ~w32721 & w32877 ;
  assign w33196 = ( w32877 & w33171 ) | ( w32877 & ~w33195 ) | ( w33171 & ~w33195 ) ;
  assign w33197 = \pi067 ^ w33196 ;
  assign w33198 = ( ~w33184 & w33194 ) | ( ~w33184 & w33197 ) | ( w33194 & w33197 ) ;
  assign w33199 = w33197 | w33198 ;
  assign w33200 = \pi068 ^ w33164 ;
  assign w33201 = ( ~w33174 & w33199 ) | ( ~w33174 & w33200 ) | ( w33199 & w33200 ) ;
  assign w33202 = w33200 | w33201 ;
  assign w33203 = \pi069 ^ w33158 ;
  assign w33204 = ( ~w33165 & w33202 ) | ( ~w33165 & w33203 ) | ( w33202 & w33203 ) ;
  assign w33205 = w33203 | w33204 ;
  assign w33206 = \pi070 ^ w33152 ;
  assign w33207 = ( ~w33159 & w33205 ) | ( ~w33159 & w33206 ) | ( w33205 & w33206 ) ;
  assign w33208 = w33206 | w33207 ;
  assign w33209 = \pi071 ^ w33146 ;
  assign w33210 = ( ~w33153 & w33208 ) | ( ~w33153 & w33209 ) | ( w33208 & w33209 ) ;
  assign w33211 = w33209 | w33210 ;
  assign w33212 = \pi072 ^ w33140 ;
  assign w33213 = ( ~w33147 & w33211 ) | ( ~w33147 & w33212 ) | ( w33211 & w33212 ) ;
  assign w33214 = w33212 | w33213 ;
  assign w33215 = \pi073 ^ w33134 ;
  assign w33216 = ( ~w33141 & w33214 ) | ( ~w33141 & w33215 ) | ( w33214 & w33215 ) ;
  assign w33217 = w33215 | w33216 ;
  assign w33218 = \pi074 ^ w33128 ;
  assign w33219 = ( ~w33135 & w33217 ) | ( ~w33135 & w33218 ) | ( w33217 & w33218 ) ;
  assign w33220 = w33218 | w33219 ;
  assign w33221 = \pi075 ^ w33122 ;
  assign w33222 = ( ~w33129 & w33220 ) | ( ~w33129 & w33221 ) | ( w33220 & w33221 ) ;
  assign w33223 = w33221 | w33222 ;
  assign w33224 = \pi076 ^ w33116 ;
  assign w33225 = ( ~w33123 & w33223 ) | ( ~w33123 & w33224 ) | ( w33223 & w33224 ) ;
  assign w33226 = w33224 | w33225 ;
  assign w33227 = \pi077 ^ w33110 ;
  assign w33228 = ( ~w33117 & w33226 ) | ( ~w33117 & w33227 ) | ( w33226 & w33227 ) ;
  assign w33229 = w33227 | w33228 ;
  assign w33230 = \pi078 ^ w33104 ;
  assign w33231 = ( ~w33111 & w33229 ) | ( ~w33111 & w33230 ) | ( w33229 & w33230 ) ;
  assign w33232 = w33230 | w33231 ;
  assign w33233 = \pi079 ^ w33098 ;
  assign w33234 = ( ~w33105 & w33232 ) | ( ~w33105 & w33233 ) | ( w33232 & w33233 ) ;
  assign w33235 = w33233 | w33234 ;
  assign w33236 = \pi080 ^ w33092 ;
  assign w33237 = ( ~w33099 & w33235 ) | ( ~w33099 & w33236 ) | ( w33235 & w33236 ) ;
  assign w33238 = w33236 | w33237 ;
  assign w33239 = \pi081 ^ w33086 ;
  assign w33240 = ( ~w33093 & w33238 ) | ( ~w33093 & w33239 ) | ( w33238 & w33239 ) ;
  assign w33241 = w33239 | w33240 ;
  assign w33242 = \pi082 ^ w33080 ;
  assign w33243 = ( ~w33087 & w33241 ) | ( ~w33087 & w33242 ) | ( w33241 & w33242 ) ;
  assign w33244 = w33242 | w33243 ;
  assign w33245 = \pi083 ^ w33074 ;
  assign w33246 = ( ~w33081 & w33244 ) | ( ~w33081 & w33245 ) | ( w33244 & w33245 ) ;
  assign w33247 = w33245 | w33246 ;
  assign w33248 = \pi084 ^ w33068 ;
  assign w33249 = ( ~w33075 & w33247 ) | ( ~w33075 & w33248 ) | ( w33247 & w33248 ) ;
  assign w33250 = w33248 | w33249 ;
  assign w33251 = \pi085 ^ w33062 ;
  assign w33252 = ( ~w33069 & w33250 ) | ( ~w33069 & w33251 ) | ( w33250 & w33251 ) ;
  assign w33253 = w33251 | w33252 ;
  assign w33254 = \pi086 ^ w33056 ;
  assign w33255 = ( ~w33063 & w33253 ) | ( ~w33063 & w33254 ) | ( w33253 & w33254 ) ;
  assign w33256 = w33254 | w33255 ;
  assign w33257 = \pi087 ^ w33050 ;
  assign w33258 = ( ~w33057 & w33256 ) | ( ~w33057 & w33257 ) | ( w33256 & w33257 ) ;
  assign w33259 = w33257 | w33258 ;
  assign w33260 = \pi088 ^ w33044 ;
  assign w33261 = ( ~w33051 & w33259 ) | ( ~w33051 & w33260 ) | ( w33259 & w33260 ) ;
  assign w33262 = w33260 | w33261 ;
  assign w33263 = \pi089 ^ w33038 ;
  assign w33264 = ( ~w33045 & w33262 ) | ( ~w33045 & w33263 ) | ( w33262 & w33263 ) ;
  assign w33265 = w33263 | w33264 ;
  assign w33266 = \pi090 ^ w33032 ;
  assign w33267 = ( ~w33039 & w33265 ) | ( ~w33039 & w33266 ) | ( w33265 & w33266 ) ;
  assign w33268 = w33266 | w33267 ;
  assign w33269 = \pi091 ^ w33026 ;
  assign w33270 = ( ~w33033 & w33268 ) | ( ~w33033 & w33269 ) | ( w33268 & w33269 ) ;
  assign w33271 = w33269 | w33270 ;
  assign w33272 = \pi092 ^ w33020 ;
  assign w33273 = ( ~w33027 & w33271 ) | ( ~w33027 & w33272 ) | ( w33271 & w33272 ) ;
  assign w33274 = w33272 | w33273 ;
  assign w33275 = \pi093 ^ w33014 ;
  assign w33276 = ( ~w33021 & w33274 ) | ( ~w33021 & w33275 ) | ( w33274 & w33275 ) ;
  assign w33277 = w33275 | w33276 ;
  assign w33278 = \pi094 ^ w33008 ;
  assign w33279 = ( ~w33015 & w33277 ) | ( ~w33015 & w33278 ) | ( w33277 & w33278 ) ;
  assign w33280 = w33278 | w33279 ;
  assign w33281 = \pi095 ^ w33002 ;
  assign w33282 = ( ~w33009 & w33280 ) | ( ~w33009 & w33281 ) | ( w33280 & w33281 ) ;
  assign w33283 = w33281 | w33282 ;
  assign w33284 = \pi096 ^ w32996 ;
  assign w33285 = ( ~w33003 & w33283 ) | ( ~w33003 & w33284 ) | ( w33283 & w33284 ) ;
  assign w33286 = w33284 | w33285 ;
  assign w33287 = \pi097 ^ w32990 ;
  assign w33288 = ( ~w32997 & w33286 ) | ( ~w32997 & w33287 ) | ( w33286 & w33287 ) ;
  assign w33289 = w33287 | w33288 ;
  assign w33290 = \pi098 ^ w32984 ;
  assign w33291 = ( ~w32991 & w33289 ) | ( ~w32991 & w33290 ) | ( w33289 & w33290 ) ;
  assign w33292 = w33290 | w33291 ;
  assign w33293 = \pi099 ^ w32978 ;
  assign w33294 = ( ~w32985 & w33292 ) | ( ~w32985 & w33293 ) | ( w33292 & w33293 ) ;
  assign w33295 = w33293 | w33294 ;
  assign w33296 = \pi100 ^ w32972 ;
  assign w33297 = ( ~w32979 & w33295 ) | ( ~w32979 & w33296 ) | ( w33295 & w33296 ) ;
  assign w33298 = w33296 | w33297 ;
  assign w33299 = \pi101 ^ w32966 ;
  assign w33300 = ( ~w32973 & w33298 ) | ( ~w32973 & w33299 ) | ( w33298 & w33299 ) ;
  assign w33301 = w33299 | w33300 ;
  assign w33302 = \pi102 ^ w32960 ;
  assign w33303 = ( ~w32967 & w33301 ) | ( ~w32967 & w33302 ) | ( w33301 & w33302 ) ;
  assign w33304 = w33302 | w33303 ;
  assign w33305 = \pi103 ^ w32954 ;
  assign w33306 = ( ~w32961 & w33304 ) | ( ~w32961 & w33305 ) | ( w33304 & w33305 ) ;
  assign w33307 = w33305 | w33306 ;
  assign w33308 = \pi104 ^ w32948 ;
  assign w33309 = ( ~w32955 & w33307 ) | ( ~w32955 & w33308 ) | ( w33307 & w33308 ) ;
  assign w33310 = w33308 | w33309 ;
  assign w33311 = \pi105 ^ w32942 ;
  assign w33312 = ( ~w32949 & w33310 ) | ( ~w32949 & w33311 ) | ( w33310 & w33311 ) ;
  assign w33313 = w33311 | w33312 ;
  assign w33314 = \pi106 ^ w32936 ;
  assign w33315 = ( ~w32943 & w33313 ) | ( ~w32943 & w33314 ) | ( w33313 & w33314 ) ;
  assign w33316 = w33314 | w33315 ;
  assign w33317 = \pi107 ^ w32930 ;
  assign w33318 = ( ~w32937 & w33316 ) | ( ~w32937 & w33317 ) | ( w33316 & w33317 ) ;
  assign w33319 = w33317 | w33318 ;
  assign w33320 = \pi108 ^ w32924 ;
  assign w33321 = ( ~w32931 & w33319 ) | ( ~w32931 & w33320 ) | ( w33319 & w33320 ) ;
  assign w33322 = w33320 | w33321 ;
  assign w33323 = \pi109 ^ w32918 ;
  assign w33324 = ( ~w32925 & w33322 ) | ( ~w32925 & w33323 ) | ( w33322 & w33323 ) ;
  assign w33325 = w33323 | w33324 ;
  assign w33326 = \pi110 ^ w32912 ;
  assign w33327 = ( ~w32919 & w33325 ) | ( ~w32919 & w33326 ) | ( w33325 & w33326 ) ;
  assign w33328 = w33326 | w33327 ;
  assign w33329 = \pi111 ^ w32906 ;
  assign w33330 = ( ~w32913 & w33328 ) | ( ~w32913 & w33329 ) | ( w33328 & w33329 ) ;
  assign w33331 = w33329 | w33330 ;
  assign w33332 = \pi112 ^ w32900 ;
  assign w33333 = ( ~w32907 & w33331 ) | ( ~w32907 & w33332 ) | ( w33331 & w33332 ) ;
  assign w33334 = w33332 | w33333 ;
  assign w33335 = \pi113 ^ w32894 ;
  assign w33336 = ( ~w32901 & w33334 ) | ( ~w32901 & w33335 ) | ( w33334 & w33335 ) ;
  assign w33337 = w33335 | w33336 ;
  assign w33338 = \pi114 ^ w32888 ;
  assign w33339 = ( ~w32895 & w33337 ) | ( ~w32895 & w33338 ) | ( w33337 & w33338 ) ;
  assign w33340 = w33338 | w33339 ;
  assign w33341 = \pi115 ^ w32882 ;
  assign w33342 = ( ~w32889 & w33340 ) | ( ~w32889 & w33341 ) | ( w33340 & w33341 ) ;
  assign w33343 = w33341 | w33342 ;
  assign w33344 = w32383 & w32877 ;
  assign w33345 = ~w32384 & w32871 ;
  assign w33346 = w32872 ^ w33345 ;
  assign w33347 = ~w32877 & w33346 ;
  assign w33348 = w33344 | w33347 ;
  assign w33349 = ~\pi116 & w33348 ;
  assign w33350 = ( \pi116 & ~w33344 ) | ( \pi116 & w33347 ) | ( ~w33344 & w33347 ) ;
  assign w33351 = ~w33347 & w33350 ;
  assign w33352 = w33349 | w33351 ;
  assign w33353 = ( ~w32883 & w33343 ) | ( ~w32883 & w33352 ) | ( w33343 & w33352 ) ;
  assign w33354 = ( w448 & ~w33352 ) | ( w448 & w33353 ) | ( ~w33352 & w33353 ) ;
  assign w33355 = w33352 | w33354 ;
  assign w33356 = ~w155 & w33348 ;
  assign w33357 = w33355 & ~w33356 ;
  assign w33358 = ~w32889 & w33340 ;
  assign w33359 = w33341 ^ w33358 ;
  assign w33360 = ~w33357 & w33359 ;
  assign w33361 = ( w32882 & w33355 ) | ( w32882 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33362 = ~w33356 & w33361 ;
  assign w33363 = w33360 | w33362 ;
  assign w33364 = ~\pi116 & w33363 ;
  assign w33365 = ~w32895 & w33337 ;
  assign w33366 = w33338 ^ w33365 ;
  assign w33367 = ~w33357 & w33366 ;
  assign w33368 = ( w32888 & w33355 ) | ( w32888 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33369 = ~w33356 & w33368 ;
  assign w33370 = w33367 | w33369 ;
  assign w33371 = ~\pi115 & w33370 ;
  assign w33372 = ~w32901 & w33334 ;
  assign w33373 = w33335 ^ w33372 ;
  assign w33374 = ~w33357 & w33373 ;
  assign w33375 = ( w32894 & w33355 ) | ( w32894 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33376 = ~w33356 & w33375 ;
  assign w33377 = w33374 | w33376 ;
  assign w33378 = ~\pi114 & w33377 ;
  assign w33379 = ~w32907 & w33331 ;
  assign w33380 = w33332 ^ w33379 ;
  assign w33381 = ~w33357 & w33380 ;
  assign w33382 = ( w32900 & w33355 ) | ( w32900 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33383 = ~w33356 & w33382 ;
  assign w33384 = w33381 | w33383 ;
  assign w33385 = ~\pi113 & w33384 ;
  assign w33386 = ~w32913 & w33328 ;
  assign w33387 = w33329 ^ w33386 ;
  assign w33388 = ~w33357 & w33387 ;
  assign w33389 = ( w32906 & w33355 ) | ( w32906 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33390 = ~w33356 & w33389 ;
  assign w33391 = w33388 | w33390 ;
  assign w33392 = ~\pi112 & w33391 ;
  assign w33393 = ~w32919 & w33325 ;
  assign w33394 = w33326 ^ w33393 ;
  assign w33395 = ~w33357 & w33394 ;
  assign w33396 = ( w32912 & w33355 ) | ( w32912 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33397 = ~w33356 & w33396 ;
  assign w33398 = w33395 | w33397 ;
  assign w33399 = ~\pi111 & w33398 ;
  assign w33400 = ~w32925 & w33322 ;
  assign w33401 = w33323 ^ w33400 ;
  assign w33402 = ~w33357 & w33401 ;
  assign w33403 = ( w32918 & w33355 ) | ( w32918 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33404 = ~w33356 & w33403 ;
  assign w33405 = w33402 | w33404 ;
  assign w33406 = ~\pi110 & w33405 ;
  assign w33407 = ~w32931 & w33319 ;
  assign w33408 = w33320 ^ w33407 ;
  assign w33409 = ~w33357 & w33408 ;
  assign w33410 = ( w32924 & w33355 ) | ( w32924 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33411 = ~w33356 & w33410 ;
  assign w33412 = w33409 | w33411 ;
  assign w33413 = ~\pi109 & w33412 ;
  assign w33414 = ~w32937 & w33316 ;
  assign w33415 = w33317 ^ w33414 ;
  assign w33416 = ~w33357 & w33415 ;
  assign w33417 = ( w32930 & w33355 ) | ( w32930 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33418 = ~w33356 & w33417 ;
  assign w33419 = w33416 | w33418 ;
  assign w33420 = ~\pi108 & w33419 ;
  assign w33421 = ~w32943 & w33313 ;
  assign w33422 = w33314 ^ w33421 ;
  assign w33423 = ~w33357 & w33422 ;
  assign w33424 = ( w32936 & w33355 ) | ( w32936 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33425 = ~w33356 & w33424 ;
  assign w33426 = w33423 | w33425 ;
  assign w33427 = ~\pi107 & w33426 ;
  assign w33428 = ~w32949 & w33310 ;
  assign w33429 = w33311 ^ w33428 ;
  assign w33430 = ~w33357 & w33429 ;
  assign w33431 = ( w32942 & w33355 ) | ( w32942 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33432 = ~w33356 & w33431 ;
  assign w33433 = w33430 | w33432 ;
  assign w33434 = ~\pi106 & w33433 ;
  assign w33435 = ~w32955 & w33307 ;
  assign w33436 = w33308 ^ w33435 ;
  assign w33437 = ~w33357 & w33436 ;
  assign w33438 = ( w32948 & w33355 ) | ( w32948 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33439 = ~w33356 & w33438 ;
  assign w33440 = w33437 | w33439 ;
  assign w33441 = ~\pi105 & w33440 ;
  assign w33442 = ~w32961 & w33304 ;
  assign w33443 = w33305 ^ w33442 ;
  assign w33444 = ~w33357 & w33443 ;
  assign w33445 = ( w32954 & w33355 ) | ( w32954 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33446 = ~w33356 & w33445 ;
  assign w33447 = w33444 | w33446 ;
  assign w33448 = ~\pi104 & w33447 ;
  assign w33449 = ~w32967 & w33301 ;
  assign w33450 = w33302 ^ w33449 ;
  assign w33451 = ~w33357 & w33450 ;
  assign w33452 = ( w32960 & w33355 ) | ( w32960 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33453 = ~w33356 & w33452 ;
  assign w33454 = w33451 | w33453 ;
  assign w33455 = ~\pi103 & w33454 ;
  assign w33456 = ~w32973 & w33298 ;
  assign w33457 = w33299 ^ w33456 ;
  assign w33458 = ~w33357 & w33457 ;
  assign w33459 = ( w32966 & w33355 ) | ( w32966 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33460 = ~w33356 & w33459 ;
  assign w33461 = w33458 | w33460 ;
  assign w33462 = ~\pi102 & w33461 ;
  assign w33463 = ~w32979 & w33295 ;
  assign w33464 = w33296 ^ w33463 ;
  assign w33465 = ~w33357 & w33464 ;
  assign w33466 = ( w32972 & w33355 ) | ( w32972 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33467 = ~w33356 & w33466 ;
  assign w33468 = w33465 | w33467 ;
  assign w33469 = ~\pi101 & w33468 ;
  assign w33470 = ~w32985 & w33292 ;
  assign w33471 = w33293 ^ w33470 ;
  assign w33472 = ~w33357 & w33471 ;
  assign w33473 = ( w32978 & w33355 ) | ( w32978 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33474 = ~w33356 & w33473 ;
  assign w33475 = w33472 | w33474 ;
  assign w33476 = ~\pi100 & w33475 ;
  assign w33477 = ~w32991 & w33289 ;
  assign w33478 = w33290 ^ w33477 ;
  assign w33479 = ~w33357 & w33478 ;
  assign w33480 = ( w32984 & w33355 ) | ( w32984 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33481 = ~w33356 & w33480 ;
  assign w33482 = w33479 | w33481 ;
  assign w33483 = ~\pi099 & w33482 ;
  assign w33484 = ~w32997 & w33286 ;
  assign w33485 = w33287 ^ w33484 ;
  assign w33486 = ~w33357 & w33485 ;
  assign w33487 = ( w32990 & w33355 ) | ( w32990 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33488 = ~w33356 & w33487 ;
  assign w33489 = w33486 | w33488 ;
  assign w33490 = ~\pi098 & w33489 ;
  assign w33491 = ~w33003 & w33283 ;
  assign w33492 = w33284 ^ w33491 ;
  assign w33493 = ~w33357 & w33492 ;
  assign w33494 = ( w32996 & w33355 ) | ( w32996 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33495 = ~w33356 & w33494 ;
  assign w33496 = w33493 | w33495 ;
  assign w33497 = ~\pi097 & w33496 ;
  assign w33498 = ~w33009 & w33280 ;
  assign w33499 = w33281 ^ w33498 ;
  assign w33500 = ~w33357 & w33499 ;
  assign w33501 = ( w33002 & w33355 ) | ( w33002 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33502 = ~w33356 & w33501 ;
  assign w33503 = w33500 | w33502 ;
  assign w33504 = ~\pi096 & w33503 ;
  assign w33505 = ~w33015 & w33277 ;
  assign w33506 = w33278 ^ w33505 ;
  assign w33507 = ~w33357 & w33506 ;
  assign w33508 = ( w33008 & w33355 ) | ( w33008 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33509 = ~w33356 & w33508 ;
  assign w33510 = w33507 | w33509 ;
  assign w33511 = ~\pi095 & w33510 ;
  assign w33512 = ~w33021 & w33274 ;
  assign w33513 = w33275 ^ w33512 ;
  assign w33514 = ~w33357 & w33513 ;
  assign w33515 = ( w33014 & w33355 ) | ( w33014 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33516 = ~w33356 & w33515 ;
  assign w33517 = w33514 | w33516 ;
  assign w33518 = ~\pi094 & w33517 ;
  assign w33519 = ~w33027 & w33271 ;
  assign w33520 = w33272 ^ w33519 ;
  assign w33521 = ~w33357 & w33520 ;
  assign w33522 = ( w33020 & w33355 ) | ( w33020 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33523 = ~w33356 & w33522 ;
  assign w33524 = w33521 | w33523 ;
  assign w33525 = ~\pi093 & w33524 ;
  assign w33526 = ~w33033 & w33268 ;
  assign w33527 = w33269 ^ w33526 ;
  assign w33528 = ~w33357 & w33527 ;
  assign w33529 = ( w33026 & w33355 ) | ( w33026 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33530 = ~w33356 & w33529 ;
  assign w33531 = w33528 | w33530 ;
  assign w33532 = ~\pi092 & w33531 ;
  assign w33533 = ~w33039 & w33265 ;
  assign w33534 = w33266 ^ w33533 ;
  assign w33535 = ~w33357 & w33534 ;
  assign w33536 = ( w33032 & w33355 ) | ( w33032 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33537 = ~w33356 & w33536 ;
  assign w33538 = w33535 | w33537 ;
  assign w33539 = ~\pi091 & w33538 ;
  assign w33540 = ~w33045 & w33262 ;
  assign w33541 = w33263 ^ w33540 ;
  assign w33542 = ~w33357 & w33541 ;
  assign w33543 = ( w33038 & w33355 ) | ( w33038 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33544 = ~w33356 & w33543 ;
  assign w33545 = w33542 | w33544 ;
  assign w33546 = ~\pi090 & w33545 ;
  assign w33547 = ~w33051 & w33259 ;
  assign w33548 = w33260 ^ w33547 ;
  assign w33549 = ~w33357 & w33548 ;
  assign w33550 = ( w33044 & w33355 ) | ( w33044 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33551 = ~w33356 & w33550 ;
  assign w33552 = w33549 | w33551 ;
  assign w33553 = ~\pi089 & w33552 ;
  assign w33554 = ~w33057 & w33256 ;
  assign w33555 = w33257 ^ w33554 ;
  assign w33556 = ~w33357 & w33555 ;
  assign w33557 = ( w33050 & w33355 ) | ( w33050 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33558 = ~w33356 & w33557 ;
  assign w33559 = w33556 | w33558 ;
  assign w33560 = ~\pi088 & w33559 ;
  assign w33561 = ~w33063 & w33253 ;
  assign w33562 = w33254 ^ w33561 ;
  assign w33563 = ~w33357 & w33562 ;
  assign w33564 = ( w33056 & w33355 ) | ( w33056 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33565 = ~w33356 & w33564 ;
  assign w33566 = w33563 | w33565 ;
  assign w33567 = ~\pi087 & w33566 ;
  assign w33568 = ~w33069 & w33250 ;
  assign w33569 = w33251 ^ w33568 ;
  assign w33570 = ~w33357 & w33569 ;
  assign w33571 = ( w33062 & w33355 ) | ( w33062 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33572 = ~w33356 & w33571 ;
  assign w33573 = w33570 | w33572 ;
  assign w33574 = ~\pi086 & w33573 ;
  assign w33575 = ~w33075 & w33247 ;
  assign w33576 = w33248 ^ w33575 ;
  assign w33577 = ~w33357 & w33576 ;
  assign w33578 = ( w33068 & w33355 ) | ( w33068 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33579 = ~w33356 & w33578 ;
  assign w33580 = w33577 | w33579 ;
  assign w33581 = ~\pi085 & w33580 ;
  assign w33582 = ~w33081 & w33244 ;
  assign w33583 = w33245 ^ w33582 ;
  assign w33584 = ~w33357 & w33583 ;
  assign w33585 = ( w33074 & w33355 ) | ( w33074 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33586 = ~w33356 & w33585 ;
  assign w33587 = w33584 | w33586 ;
  assign w33588 = ~\pi084 & w33587 ;
  assign w33589 = ~w33087 & w33241 ;
  assign w33590 = w33242 ^ w33589 ;
  assign w33591 = ~w33357 & w33590 ;
  assign w33592 = ( w33080 & w33355 ) | ( w33080 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33593 = ~w33356 & w33592 ;
  assign w33594 = w33591 | w33593 ;
  assign w33595 = ~\pi083 & w33594 ;
  assign w33596 = ~w33093 & w33238 ;
  assign w33597 = w33239 ^ w33596 ;
  assign w33598 = ~w33357 & w33597 ;
  assign w33599 = ( w33086 & w33355 ) | ( w33086 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33600 = ~w33356 & w33599 ;
  assign w33601 = w33598 | w33600 ;
  assign w33602 = ~\pi082 & w33601 ;
  assign w33603 = ~w33099 & w33235 ;
  assign w33604 = w33236 ^ w33603 ;
  assign w33605 = ~w33357 & w33604 ;
  assign w33606 = ( w33092 & w33355 ) | ( w33092 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33607 = ~w33356 & w33606 ;
  assign w33608 = w33605 | w33607 ;
  assign w33609 = ~\pi081 & w33608 ;
  assign w33610 = ~w33105 & w33232 ;
  assign w33611 = w33233 ^ w33610 ;
  assign w33612 = ~w33357 & w33611 ;
  assign w33613 = ( w33098 & w33355 ) | ( w33098 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33614 = ~w33356 & w33613 ;
  assign w33615 = w33612 | w33614 ;
  assign w33616 = ~\pi080 & w33615 ;
  assign w33617 = ~w33111 & w33229 ;
  assign w33618 = w33230 ^ w33617 ;
  assign w33619 = ~w33357 & w33618 ;
  assign w33620 = ( w33104 & w33355 ) | ( w33104 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33621 = ~w33356 & w33620 ;
  assign w33622 = w33619 | w33621 ;
  assign w33623 = ~\pi079 & w33622 ;
  assign w33624 = ~w33117 & w33226 ;
  assign w33625 = w33227 ^ w33624 ;
  assign w33626 = ~w33357 & w33625 ;
  assign w33627 = ( w33110 & w33355 ) | ( w33110 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33628 = ~w33356 & w33627 ;
  assign w33629 = w33626 | w33628 ;
  assign w33630 = ~\pi078 & w33629 ;
  assign w33631 = ~w33123 & w33223 ;
  assign w33632 = w33224 ^ w33631 ;
  assign w33633 = ~w33357 & w33632 ;
  assign w33634 = ( w33116 & w33355 ) | ( w33116 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33635 = ~w33356 & w33634 ;
  assign w33636 = w33633 | w33635 ;
  assign w33637 = ~\pi077 & w33636 ;
  assign w33638 = ~w33129 & w33220 ;
  assign w33639 = w33221 ^ w33638 ;
  assign w33640 = ~w33357 & w33639 ;
  assign w33641 = ( w33122 & w33355 ) | ( w33122 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33642 = ~w33356 & w33641 ;
  assign w33643 = w33640 | w33642 ;
  assign w33644 = ~\pi076 & w33643 ;
  assign w33645 = ~w33135 & w33217 ;
  assign w33646 = w33218 ^ w33645 ;
  assign w33647 = ~w33357 & w33646 ;
  assign w33648 = ( w33128 & w33355 ) | ( w33128 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33649 = ~w33356 & w33648 ;
  assign w33650 = w33647 | w33649 ;
  assign w33651 = ~\pi075 & w33650 ;
  assign w33652 = ~w33141 & w33214 ;
  assign w33653 = w33215 ^ w33652 ;
  assign w33654 = ~w33357 & w33653 ;
  assign w33655 = ( w33134 & w33355 ) | ( w33134 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33656 = ~w33356 & w33655 ;
  assign w33657 = w33654 | w33656 ;
  assign w33658 = ~\pi074 & w33657 ;
  assign w33659 = ~w33147 & w33211 ;
  assign w33660 = w33212 ^ w33659 ;
  assign w33661 = ~w33357 & w33660 ;
  assign w33662 = ( w33140 & w33355 ) | ( w33140 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33663 = ~w33356 & w33662 ;
  assign w33664 = w33661 | w33663 ;
  assign w33665 = ~\pi073 & w33664 ;
  assign w33666 = ~w33153 & w33208 ;
  assign w33667 = w33209 ^ w33666 ;
  assign w33668 = ~w33357 & w33667 ;
  assign w33669 = ( w33146 & w33355 ) | ( w33146 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33670 = ~w33356 & w33669 ;
  assign w33671 = w33668 | w33670 ;
  assign w33672 = ~\pi072 & w33671 ;
  assign w33673 = ~w33159 & w33205 ;
  assign w33674 = w33206 ^ w33673 ;
  assign w33675 = ~w33357 & w33674 ;
  assign w33676 = ( w33152 & w33355 ) | ( w33152 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33677 = ~w33356 & w33676 ;
  assign w33678 = w33675 | w33677 ;
  assign w33679 = ~\pi071 & w33678 ;
  assign w33680 = ~w33165 & w33202 ;
  assign w33681 = w33203 ^ w33680 ;
  assign w33682 = ~w33357 & w33681 ;
  assign w33683 = ( w33158 & w33355 ) | ( w33158 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33684 = ~w33356 & w33683 ;
  assign w33685 = w33682 | w33684 ;
  assign w33686 = ~\pi070 & w33685 ;
  assign w33687 = ~w33174 & w33199 ;
  assign w33688 = w33200 ^ w33687 ;
  assign w33689 = ~w33357 & w33688 ;
  assign w33690 = ( w33164 & w33355 ) | ( w33164 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33691 = ~w33356 & w33690 ;
  assign w33692 = w33689 | w33691 ;
  assign w33693 = ~\pi069 & w33692 ;
  assign w33694 = ~w33184 & w33194 ;
  assign w33695 = w33197 ^ w33694 ;
  assign w33696 = ~w33357 & w33695 ;
  assign w33697 = ( w33173 & w33355 ) | ( w33173 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33698 = ~w33356 & w33697 ;
  assign w33699 = w33696 | w33698 ;
  assign w33700 = ~\pi068 & w33699 ;
  assign w33701 = w33191 ^ w33193 ;
  assign w33702 = ~w33357 & w33701 ;
  assign w33703 = ( w33183 & w33355 ) | ( w33183 & w33356 ) | ( w33355 & w33356 ) ;
  assign w33704 = ~w33356 & w33703 ;
  assign w33705 = w33702 | w33704 ;
  assign w33706 = ~\pi067 & w33705 ;
  assign w33707 = w13825 ^ w33192 ;
  assign w33708 = \pi065 ^ w33707 ;
  assign w33709 = w33357 ^ w33708 ;
  assign w33710 = ( w33192 & w33708 ) | ( w33192 & w33709 ) | ( w33708 & w33709 ) ;
  assign w33711 = ~\pi066 & w33710 ;
  assign w33712 = w33192 ^ w33357 ;
  assign w33713 = ( w33192 & w33708 ) | ( w33192 & ~w33712 ) | ( w33708 & ~w33712 ) ;
  assign w33714 = \pi066 ^ w33713 ;
  assign w33715 = ( \pi064 & ~w33357 ) | ( \pi064 & w33714 ) | ( ~w33357 & w33714 ) ;
  assign w33716 = \pi011 ^ w33715 ;
  assign w33717 = ( \pi065 & w14881 ) | ( \pi065 & ~w33716 ) | ( w14881 & ~w33716 ) ;
  assign w33718 = w33714 | w33717 ;
  assign w33719 = \pi067 ^ w33705 ;
  assign w33720 = ( ~w33711 & w33718 ) | ( ~w33711 & w33719 ) | ( w33718 & w33719 ) ;
  assign w33721 = w33719 | w33720 ;
  assign w33722 = \pi068 ^ w33699 ;
  assign w33723 = ( ~w33706 & w33721 ) | ( ~w33706 & w33722 ) | ( w33721 & w33722 ) ;
  assign w33724 = w33722 | w33723 ;
  assign w33725 = \pi069 ^ w33692 ;
  assign w33726 = ( ~w33700 & w33724 ) | ( ~w33700 & w33725 ) | ( w33724 & w33725 ) ;
  assign w33727 = w33725 | w33726 ;
  assign w33728 = \pi070 ^ w33685 ;
  assign w33729 = ( ~w33693 & w33727 ) | ( ~w33693 & w33728 ) | ( w33727 & w33728 ) ;
  assign w33730 = w33728 | w33729 ;
  assign w33731 = \pi071 ^ w33678 ;
  assign w33732 = ( ~w33686 & w33730 ) | ( ~w33686 & w33731 ) | ( w33730 & w33731 ) ;
  assign w33733 = w33731 | w33732 ;
  assign w33734 = \pi072 ^ w33671 ;
  assign w33735 = ( ~w33679 & w33733 ) | ( ~w33679 & w33734 ) | ( w33733 & w33734 ) ;
  assign w33736 = w33734 | w33735 ;
  assign w33737 = \pi073 ^ w33664 ;
  assign w33738 = ( ~w33672 & w33736 ) | ( ~w33672 & w33737 ) | ( w33736 & w33737 ) ;
  assign w33739 = w33737 | w33738 ;
  assign w33740 = \pi074 ^ w33657 ;
  assign w33741 = ( ~w33665 & w33739 ) | ( ~w33665 & w33740 ) | ( w33739 & w33740 ) ;
  assign w33742 = w33740 | w33741 ;
  assign w33743 = \pi075 ^ w33650 ;
  assign w33744 = ( ~w33658 & w33742 ) | ( ~w33658 & w33743 ) | ( w33742 & w33743 ) ;
  assign w33745 = w33743 | w33744 ;
  assign w33746 = \pi076 ^ w33643 ;
  assign w33747 = ( ~w33651 & w33745 ) | ( ~w33651 & w33746 ) | ( w33745 & w33746 ) ;
  assign w33748 = w33746 | w33747 ;
  assign w33749 = \pi077 ^ w33636 ;
  assign w33750 = ( ~w33644 & w33748 ) | ( ~w33644 & w33749 ) | ( w33748 & w33749 ) ;
  assign w33751 = w33749 | w33750 ;
  assign w33752 = \pi078 ^ w33629 ;
  assign w33753 = ( ~w33637 & w33751 ) | ( ~w33637 & w33752 ) | ( w33751 & w33752 ) ;
  assign w33754 = w33752 | w33753 ;
  assign w33755 = \pi079 ^ w33622 ;
  assign w33756 = ( ~w33630 & w33754 ) | ( ~w33630 & w33755 ) | ( w33754 & w33755 ) ;
  assign w33757 = w33755 | w33756 ;
  assign w33758 = \pi080 ^ w33615 ;
  assign w33759 = ( ~w33623 & w33757 ) | ( ~w33623 & w33758 ) | ( w33757 & w33758 ) ;
  assign w33760 = w33758 | w33759 ;
  assign w33761 = \pi081 ^ w33608 ;
  assign w33762 = ( ~w33616 & w33760 ) | ( ~w33616 & w33761 ) | ( w33760 & w33761 ) ;
  assign w33763 = w33761 | w33762 ;
  assign w33764 = \pi082 ^ w33601 ;
  assign w33765 = ( ~w33609 & w33763 ) | ( ~w33609 & w33764 ) | ( w33763 & w33764 ) ;
  assign w33766 = w33764 | w33765 ;
  assign w33767 = \pi083 ^ w33594 ;
  assign w33768 = ( ~w33602 & w33766 ) | ( ~w33602 & w33767 ) | ( w33766 & w33767 ) ;
  assign w33769 = w33767 | w33768 ;
  assign w33770 = \pi084 ^ w33587 ;
  assign w33771 = ( ~w33595 & w33769 ) | ( ~w33595 & w33770 ) | ( w33769 & w33770 ) ;
  assign w33772 = w33770 | w33771 ;
  assign w33773 = \pi085 ^ w33580 ;
  assign w33774 = ( ~w33588 & w33772 ) | ( ~w33588 & w33773 ) | ( w33772 & w33773 ) ;
  assign w33775 = w33773 | w33774 ;
  assign w33776 = \pi086 ^ w33573 ;
  assign w33777 = ( ~w33581 & w33775 ) | ( ~w33581 & w33776 ) | ( w33775 & w33776 ) ;
  assign w33778 = w33776 | w33777 ;
  assign w33779 = \pi087 ^ w33566 ;
  assign w33780 = ( ~w33574 & w33778 ) | ( ~w33574 & w33779 ) | ( w33778 & w33779 ) ;
  assign w33781 = w33779 | w33780 ;
  assign w33782 = \pi088 ^ w33559 ;
  assign w33783 = ( ~w33567 & w33781 ) | ( ~w33567 & w33782 ) | ( w33781 & w33782 ) ;
  assign w33784 = w33782 | w33783 ;
  assign w33785 = \pi089 ^ w33552 ;
  assign w33786 = ( ~w33560 & w33784 ) | ( ~w33560 & w33785 ) | ( w33784 & w33785 ) ;
  assign w33787 = w33785 | w33786 ;
  assign w33788 = \pi090 ^ w33545 ;
  assign w33789 = ( ~w33553 & w33787 ) | ( ~w33553 & w33788 ) | ( w33787 & w33788 ) ;
  assign w33790 = w33788 | w33789 ;
  assign w33791 = \pi091 ^ w33538 ;
  assign w33792 = ( ~w33546 & w33790 ) | ( ~w33546 & w33791 ) | ( w33790 & w33791 ) ;
  assign w33793 = w33791 | w33792 ;
  assign w33794 = \pi092 ^ w33531 ;
  assign w33795 = ( ~w33539 & w33793 ) | ( ~w33539 & w33794 ) | ( w33793 & w33794 ) ;
  assign w33796 = w33794 | w33795 ;
  assign w33797 = \pi093 ^ w33524 ;
  assign w33798 = ( ~w33532 & w33796 ) | ( ~w33532 & w33797 ) | ( w33796 & w33797 ) ;
  assign w33799 = w33797 | w33798 ;
  assign w33800 = \pi094 ^ w33517 ;
  assign w33801 = ( ~w33525 & w33799 ) | ( ~w33525 & w33800 ) | ( w33799 & w33800 ) ;
  assign w33802 = w33800 | w33801 ;
  assign w33803 = \pi095 ^ w33510 ;
  assign w33804 = ( ~w33518 & w33802 ) | ( ~w33518 & w33803 ) | ( w33802 & w33803 ) ;
  assign w33805 = w33803 | w33804 ;
  assign w33806 = \pi096 ^ w33503 ;
  assign w33807 = ( ~w33511 & w33805 ) | ( ~w33511 & w33806 ) | ( w33805 & w33806 ) ;
  assign w33808 = w33806 | w33807 ;
  assign w33809 = \pi097 ^ w33496 ;
  assign w33810 = ( ~w33504 & w33808 ) | ( ~w33504 & w33809 ) | ( w33808 & w33809 ) ;
  assign w33811 = w33809 | w33810 ;
  assign w33812 = \pi098 ^ w33489 ;
  assign w33813 = ( ~w33497 & w33811 ) | ( ~w33497 & w33812 ) | ( w33811 & w33812 ) ;
  assign w33814 = w33812 | w33813 ;
  assign w33815 = \pi099 ^ w33482 ;
  assign w33816 = ( ~w33490 & w33814 ) | ( ~w33490 & w33815 ) | ( w33814 & w33815 ) ;
  assign w33817 = w33815 | w33816 ;
  assign w33818 = \pi100 ^ w33475 ;
  assign w33819 = ( ~w33483 & w33817 ) | ( ~w33483 & w33818 ) | ( w33817 & w33818 ) ;
  assign w33820 = w33818 | w33819 ;
  assign w33821 = \pi101 ^ w33468 ;
  assign w33822 = ( ~w33476 & w33820 ) | ( ~w33476 & w33821 ) | ( w33820 & w33821 ) ;
  assign w33823 = w33821 | w33822 ;
  assign w33824 = \pi102 ^ w33461 ;
  assign w33825 = ( ~w33469 & w33823 ) | ( ~w33469 & w33824 ) | ( w33823 & w33824 ) ;
  assign w33826 = w33824 | w33825 ;
  assign w33827 = \pi103 ^ w33454 ;
  assign w33828 = ( ~w33462 & w33826 ) | ( ~w33462 & w33827 ) | ( w33826 & w33827 ) ;
  assign w33829 = w33827 | w33828 ;
  assign w33830 = \pi104 ^ w33447 ;
  assign w33831 = ( ~w33455 & w33829 ) | ( ~w33455 & w33830 ) | ( w33829 & w33830 ) ;
  assign w33832 = w33830 | w33831 ;
  assign w33833 = \pi105 ^ w33440 ;
  assign w33834 = ( ~w33448 & w33832 ) | ( ~w33448 & w33833 ) | ( w33832 & w33833 ) ;
  assign w33835 = w33833 | w33834 ;
  assign w33836 = \pi106 ^ w33433 ;
  assign w33837 = ( ~w33441 & w33835 ) | ( ~w33441 & w33836 ) | ( w33835 & w33836 ) ;
  assign w33838 = w33836 | w33837 ;
  assign w33839 = \pi107 ^ w33426 ;
  assign w33840 = ( ~w33434 & w33838 ) | ( ~w33434 & w33839 ) | ( w33838 & w33839 ) ;
  assign w33841 = w33839 | w33840 ;
  assign w33842 = \pi108 ^ w33419 ;
  assign w33843 = ( ~w33427 & w33841 ) | ( ~w33427 & w33842 ) | ( w33841 & w33842 ) ;
  assign w33844 = w33842 | w33843 ;
  assign w33845 = \pi109 ^ w33412 ;
  assign w33846 = ( ~w33420 & w33844 ) | ( ~w33420 & w33845 ) | ( w33844 & w33845 ) ;
  assign w33847 = w33845 | w33846 ;
  assign w33848 = \pi110 ^ w33405 ;
  assign w33849 = ( ~w33413 & w33847 ) | ( ~w33413 & w33848 ) | ( w33847 & w33848 ) ;
  assign w33850 = w33848 | w33849 ;
  assign w33851 = \pi111 ^ w33398 ;
  assign w33852 = ( ~w33406 & w33850 ) | ( ~w33406 & w33851 ) | ( w33850 & w33851 ) ;
  assign w33853 = w33851 | w33852 ;
  assign w33854 = \pi112 ^ w33391 ;
  assign w33855 = ( ~w33399 & w33853 ) | ( ~w33399 & w33854 ) | ( w33853 & w33854 ) ;
  assign w33856 = w33854 | w33855 ;
  assign w33857 = \pi113 ^ w33384 ;
  assign w33858 = ( ~w33392 & w33856 ) | ( ~w33392 & w33857 ) | ( w33856 & w33857 ) ;
  assign w33859 = w33857 | w33858 ;
  assign w33860 = \pi114 ^ w33377 ;
  assign w33861 = ( ~w33385 & w33859 ) | ( ~w33385 & w33860 ) | ( w33859 & w33860 ) ;
  assign w33862 = w33860 | w33861 ;
  assign w33863 = \pi115 ^ w33370 ;
  assign w33864 = ( ~w33378 & w33862 ) | ( ~w33378 & w33863 ) | ( w33862 & w33863 ) ;
  assign w33865 = w33863 | w33864 ;
  assign w33866 = \pi116 ^ w33363 ;
  assign w33867 = ( ~w33371 & w33865 ) | ( ~w33371 & w33866 ) | ( w33865 & w33866 ) ;
  assign w33868 = w33866 | w33867 ;
  assign w33869 = ( ~w32883 & w33343 ) | ( ~w32883 & w33357 ) | ( w33343 & w33357 ) ;
  assign w33870 = w33352 ^ w33869 ;
  assign w33871 = ~w33357 & w33870 ;
  assign w33872 = ( w155 & ~w33348 ) | ( w155 & w33355 ) | ( ~w33348 & w33355 ) ;
  assign w33873 = w33348 & w33872 ;
  assign w33874 = w33871 | w33873 ;
  assign w33875 = ~\pi117 & w33874 ;
  assign w33876 = ( \pi117 & ~w33871 ) | ( \pi117 & w33873 ) | ( ~w33871 & w33873 ) ;
  assign w33877 = ~w33873 & w33876 ;
  assign w33878 = w33875 | w33877 ;
  assign w33879 = ( ~w33364 & w33868 ) | ( ~w33364 & w33878 ) | ( w33868 & w33878 ) ;
  assign w33880 = ( w14518 & ~w33878 ) | ( w14518 & w33879 ) | ( ~w33878 & w33879 ) ;
  assign w33881 = w33878 | w33880 ;
  assign w33882 = ~w448 & w33874 ;
  assign w33883 = w33881 & ~w33882 ;
  assign w33884 = ~w33371 & w33865 ;
  assign w33885 = w33866 ^ w33884 ;
  assign w33886 = ~w33883 & w33885 ;
  assign w33887 = ( w33363 & w33881 ) | ( w33363 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33888 = ~w33882 & w33887 ;
  assign w33889 = w33886 | w33888 ;
  assign w33890 = ( ~w33364 & w33868 ) | ( ~w33364 & w33883 ) | ( w33868 & w33883 ) ;
  assign w33891 = w33878 ^ w33890 ;
  assign w33892 = ~w33883 & w33891 ;
  assign w33893 = ( w448 & ~w33874 ) | ( w448 & w33881 ) | ( ~w33874 & w33881 ) ;
  assign w33894 = w33874 & w33893 ;
  assign w33895 = w33892 | w33894 ;
  assign w33896 = ~\pi117 & w33889 ;
  assign w33897 = ~w33378 & w33862 ;
  assign w33898 = w33863 ^ w33897 ;
  assign w33899 = ~w33883 & w33898 ;
  assign w33900 = ( w33370 & w33881 ) | ( w33370 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33901 = ~w33882 & w33900 ;
  assign w33902 = w33899 | w33901 ;
  assign w33903 = ~\pi116 & w33902 ;
  assign w33904 = ~w33385 & w33859 ;
  assign w33905 = w33860 ^ w33904 ;
  assign w33906 = ~w33883 & w33905 ;
  assign w33907 = ( w33377 & w33881 ) | ( w33377 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33908 = ~w33882 & w33907 ;
  assign w33909 = w33906 | w33908 ;
  assign w33910 = ~\pi115 & w33909 ;
  assign w33911 = ~w33392 & w33856 ;
  assign w33912 = w33857 ^ w33911 ;
  assign w33913 = ~w33883 & w33912 ;
  assign w33914 = ( w33384 & w33881 ) | ( w33384 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33915 = ~w33882 & w33914 ;
  assign w33916 = w33913 | w33915 ;
  assign w33917 = ~\pi114 & w33916 ;
  assign w33918 = ~w33399 & w33853 ;
  assign w33919 = w33854 ^ w33918 ;
  assign w33920 = ~w33883 & w33919 ;
  assign w33921 = ( w33391 & w33881 ) | ( w33391 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33922 = ~w33882 & w33921 ;
  assign w33923 = w33920 | w33922 ;
  assign w33924 = ~\pi113 & w33923 ;
  assign w33925 = ~w33406 & w33850 ;
  assign w33926 = w33851 ^ w33925 ;
  assign w33927 = ~w33883 & w33926 ;
  assign w33928 = ( w33398 & w33881 ) | ( w33398 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33929 = ~w33882 & w33928 ;
  assign w33930 = w33927 | w33929 ;
  assign w33931 = ~\pi112 & w33930 ;
  assign w33932 = ~w33413 & w33847 ;
  assign w33933 = w33848 ^ w33932 ;
  assign w33934 = ~w33883 & w33933 ;
  assign w33935 = ( w33405 & w33881 ) | ( w33405 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33936 = ~w33882 & w33935 ;
  assign w33937 = w33934 | w33936 ;
  assign w33938 = ~\pi111 & w33937 ;
  assign w33939 = ~w33420 & w33844 ;
  assign w33940 = w33845 ^ w33939 ;
  assign w33941 = ~w33883 & w33940 ;
  assign w33942 = ( w33412 & w33881 ) | ( w33412 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33943 = ~w33882 & w33942 ;
  assign w33944 = w33941 | w33943 ;
  assign w33945 = ~\pi110 & w33944 ;
  assign w33946 = ~w33427 & w33841 ;
  assign w33947 = w33842 ^ w33946 ;
  assign w33948 = ~w33883 & w33947 ;
  assign w33949 = ( w33419 & w33881 ) | ( w33419 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33950 = ~w33882 & w33949 ;
  assign w33951 = w33948 | w33950 ;
  assign w33952 = ~\pi109 & w33951 ;
  assign w33953 = ~w33434 & w33838 ;
  assign w33954 = w33839 ^ w33953 ;
  assign w33955 = ~w33883 & w33954 ;
  assign w33956 = ( w33426 & w33881 ) | ( w33426 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33957 = ~w33882 & w33956 ;
  assign w33958 = w33955 | w33957 ;
  assign w33959 = ~\pi108 & w33958 ;
  assign w33960 = ~w33441 & w33835 ;
  assign w33961 = w33836 ^ w33960 ;
  assign w33962 = ~w33883 & w33961 ;
  assign w33963 = ( w33433 & w33881 ) | ( w33433 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33964 = ~w33882 & w33963 ;
  assign w33965 = w33962 | w33964 ;
  assign w33966 = ~\pi107 & w33965 ;
  assign w33967 = ~w33448 & w33832 ;
  assign w33968 = w33833 ^ w33967 ;
  assign w33969 = ~w33883 & w33968 ;
  assign w33970 = ( w33440 & w33881 ) | ( w33440 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33971 = ~w33882 & w33970 ;
  assign w33972 = w33969 | w33971 ;
  assign w33973 = ~\pi106 & w33972 ;
  assign w33974 = ~w33455 & w33829 ;
  assign w33975 = w33830 ^ w33974 ;
  assign w33976 = ~w33883 & w33975 ;
  assign w33977 = ( w33447 & w33881 ) | ( w33447 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33978 = ~w33882 & w33977 ;
  assign w33979 = w33976 | w33978 ;
  assign w33980 = ~\pi105 & w33979 ;
  assign w33981 = ~w33462 & w33826 ;
  assign w33982 = w33827 ^ w33981 ;
  assign w33983 = ~w33883 & w33982 ;
  assign w33984 = ( w33454 & w33881 ) | ( w33454 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33985 = ~w33882 & w33984 ;
  assign w33986 = w33983 | w33985 ;
  assign w33987 = ~\pi104 & w33986 ;
  assign w33988 = ~w33469 & w33823 ;
  assign w33989 = w33824 ^ w33988 ;
  assign w33990 = ~w33883 & w33989 ;
  assign w33991 = ( w33461 & w33881 ) | ( w33461 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33992 = ~w33882 & w33991 ;
  assign w33993 = w33990 | w33992 ;
  assign w33994 = ~\pi103 & w33993 ;
  assign w33995 = ~w33476 & w33820 ;
  assign w33996 = w33821 ^ w33995 ;
  assign w33997 = ~w33883 & w33996 ;
  assign w33998 = ( w33468 & w33881 ) | ( w33468 & w33882 ) | ( w33881 & w33882 ) ;
  assign w33999 = ~w33882 & w33998 ;
  assign w34000 = w33997 | w33999 ;
  assign w34001 = ~\pi102 & w34000 ;
  assign w34002 = ~w33483 & w33817 ;
  assign w34003 = w33818 ^ w34002 ;
  assign w34004 = ~w33883 & w34003 ;
  assign w34005 = ( w33475 & w33881 ) | ( w33475 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34006 = ~w33882 & w34005 ;
  assign w34007 = w34004 | w34006 ;
  assign w34008 = ~\pi101 & w34007 ;
  assign w34009 = ~w33490 & w33814 ;
  assign w34010 = w33815 ^ w34009 ;
  assign w34011 = ~w33883 & w34010 ;
  assign w34012 = ( w33482 & w33881 ) | ( w33482 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34013 = ~w33882 & w34012 ;
  assign w34014 = w34011 | w34013 ;
  assign w34015 = ~\pi100 & w34014 ;
  assign w34016 = ~w33497 & w33811 ;
  assign w34017 = w33812 ^ w34016 ;
  assign w34018 = ~w33883 & w34017 ;
  assign w34019 = ( w33489 & w33881 ) | ( w33489 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34020 = ~w33882 & w34019 ;
  assign w34021 = w34018 | w34020 ;
  assign w34022 = ~\pi099 & w34021 ;
  assign w34023 = ~w33504 & w33808 ;
  assign w34024 = w33809 ^ w34023 ;
  assign w34025 = ~w33883 & w34024 ;
  assign w34026 = ( w33496 & w33881 ) | ( w33496 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34027 = ~w33882 & w34026 ;
  assign w34028 = w34025 | w34027 ;
  assign w34029 = ~\pi098 & w34028 ;
  assign w34030 = ~w33511 & w33805 ;
  assign w34031 = w33806 ^ w34030 ;
  assign w34032 = ~w33883 & w34031 ;
  assign w34033 = ( w33503 & w33881 ) | ( w33503 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34034 = ~w33882 & w34033 ;
  assign w34035 = w34032 | w34034 ;
  assign w34036 = ~\pi097 & w34035 ;
  assign w34037 = ~w33518 & w33802 ;
  assign w34038 = w33803 ^ w34037 ;
  assign w34039 = ~w33883 & w34038 ;
  assign w34040 = ( w33510 & w33881 ) | ( w33510 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34041 = ~w33882 & w34040 ;
  assign w34042 = w34039 | w34041 ;
  assign w34043 = ~\pi096 & w34042 ;
  assign w34044 = ~w33525 & w33799 ;
  assign w34045 = w33800 ^ w34044 ;
  assign w34046 = ~w33883 & w34045 ;
  assign w34047 = ( w33517 & w33881 ) | ( w33517 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34048 = ~w33882 & w34047 ;
  assign w34049 = w34046 | w34048 ;
  assign w34050 = ~\pi095 & w34049 ;
  assign w34051 = ~w33532 & w33796 ;
  assign w34052 = w33797 ^ w34051 ;
  assign w34053 = ~w33883 & w34052 ;
  assign w34054 = ( w33524 & w33881 ) | ( w33524 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34055 = ~w33882 & w34054 ;
  assign w34056 = w34053 | w34055 ;
  assign w34057 = ~\pi094 & w34056 ;
  assign w34058 = ~w33539 & w33793 ;
  assign w34059 = w33794 ^ w34058 ;
  assign w34060 = ~w33883 & w34059 ;
  assign w34061 = ( w33531 & w33881 ) | ( w33531 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34062 = ~w33882 & w34061 ;
  assign w34063 = w34060 | w34062 ;
  assign w34064 = ~\pi093 & w34063 ;
  assign w34065 = ~w33546 & w33790 ;
  assign w34066 = w33791 ^ w34065 ;
  assign w34067 = ~w33883 & w34066 ;
  assign w34068 = ( w33538 & w33881 ) | ( w33538 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34069 = ~w33882 & w34068 ;
  assign w34070 = w34067 | w34069 ;
  assign w34071 = ~\pi092 & w34070 ;
  assign w34072 = ~w33553 & w33787 ;
  assign w34073 = w33788 ^ w34072 ;
  assign w34074 = ~w33883 & w34073 ;
  assign w34075 = ( w33545 & w33881 ) | ( w33545 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34076 = ~w33882 & w34075 ;
  assign w34077 = w34074 | w34076 ;
  assign w34078 = ~\pi091 & w34077 ;
  assign w34079 = ~w33560 & w33784 ;
  assign w34080 = w33785 ^ w34079 ;
  assign w34081 = ~w33883 & w34080 ;
  assign w34082 = ( w33552 & w33881 ) | ( w33552 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34083 = ~w33882 & w34082 ;
  assign w34084 = w34081 | w34083 ;
  assign w34085 = ~\pi090 & w34084 ;
  assign w34086 = ~w33567 & w33781 ;
  assign w34087 = w33782 ^ w34086 ;
  assign w34088 = ~w33883 & w34087 ;
  assign w34089 = ( w33559 & w33881 ) | ( w33559 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34090 = ~w33882 & w34089 ;
  assign w34091 = w34088 | w34090 ;
  assign w34092 = ~\pi089 & w34091 ;
  assign w34093 = ~w33574 & w33778 ;
  assign w34094 = w33779 ^ w34093 ;
  assign w34095 = ~w33883 & w34094 ;
  assign w34096 = ( w33566 & w33881 ) | ( w33566 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34097 = ~w33882 & w34096 ;
  assign w34098 = w34095 | w34097 ;
  assign w34099 = ~\pi088 & w34098 ;
  assign w34100 = ~w33581 & w33775 ;
  assign w34101 = w33776 ^ w34100 ;
  assign w34102 = ~w33883 & w34101 ;
  assign w34103 = ( w33573 & w33881 ) | ( w33573 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34104 = ~w33882 & w34103 ;
  assign w34105 = w34102 | w34104 ;
  assign w34106 = ~\pi087 & w34105 ;
  assign w34107 = ~w33588 & w33772 ;
  assign w34108 = w33773 ^ w34107 ;
  assign w34109 = ~w33883 & w34108 ;
  assign w34110 = ( w33580 & w33881 ) | ( w33580 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34111 = ~w33882 & w34110 ;
  assign w34112 = w34109 | w34111 ;
  assign w34113 = ~\pi086 & w34112 ;
  assign w34114 = ~w33595 & w33769 ;
  assign w34115 = w33770 ^ w34114 ;
  assign w34116 = ~w33883 & w34115 ;
  assign w34117 = ( w33587 & w33881 ) | ( w33587 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34118 = ~w33882 & w34117 ;
  assign w34119 = w34116 | w34118 ;
  assign w34120 = ~\pi085 & w34119 ;
  assign w34121 = ~w33602 & w33766 ;
  assign w34122 = w33767 ^ w34121 ;
  assign w34123 = ~w33883 & w34122 ;
  assign w34124 = ( w33594 & w33881 ) | ( w33594 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34125 = ~w33882 & w34124 ;
  assign w34126 = w34123 | w34125 ;
  assign w34127 = ~\pi084 & w34126 ;
  assign w34128 = ~w33609 & w33763 ;
  assign w34129 = w33764 ^ w34128 ;
  assign w34130 = ~w33883 & w34129 ;
  assign w34131 = ( w33601 & w33881 ) | ( w33601 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34132 = ~w33882 & w34131 ;
  assign w34133 = w34130 | w34132 ;
  assign w34134 = ~\pi083 & w34133 ;
  assign w34135 = ~w33616 & w33760 ;
  assign w34136 = w33761 ^ w34135 ;
  assign w34137 = ~w33883 & w34136 ;
  assign w34138 = ( w33608 & w33881 ) | ( w33608 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34139 = ~w33882 & w34138 ;
  assign w34140 = w34137 | w34139 ;
  assign w34141 = ~\pi082 & w34140 ;
  assign w34142 = ~w33623 & w33757 ;
  assign w34143 = w33758 ^ w34142 ;
  assign w34144 = ~w33883 & w34143 ;
  assign w34145 = ( w33615 & w33881 ) | ( w33615 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34146 = ~w33882 & w34145 ;
  assign w34147 = w34144 | w34146 ;
  assign w34148 = ~\pi081 & w34147 ;
  assign w34149 = ~w33630 & w33754 ;
  assign w34150 = w33755 ^ w34149 ;
  assign w34151 = ~w33883 & w34150 ;
  assign w34152 = ( w33622 & w33881 ) | ( w33622 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34153 = ~w33882 & w34152 ;
  assign w34154 = w34151 | w34153 ;
  assign w34155 = ~\pi080 & w34154 ;
  assign w34156 = ~w33637 & w33751 ;
  assign w34157 = w33752 ^ w34156 ;
  assign w34158 = ~w33883 & w34157 ;
  assign w34159 = ( w33629 & w33881 ) | ( w33629 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34160 = ~w33882 & w34159 ;
  assign w34161 = w34158 | w34160 ;
  assign w34162 = ~\pi079 & w34161 ;
  assign w34163 = ~w33644 & w33748 ;
  assign w34164 = w33749 ^ w34163 ;
  assign w34165 = ~w33883 & w34164 ;
  assign w34166 = ( w33636 & w33881 ) | ( w33636 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34167 = ~w33882 & w34166 ;
  assign w34168 = w34165 | w34167 ;
  assign w34169 = ~\pi078 & w34168 ;
  assign w34170 = ~w33651 & w33745 ;
  assign w34171 = w33746 ^ w34170 ;
  assign w34172 = ~w33883 & w34171 ;
  assign w34173 = ( w33643 & w33881 ) | ( w33643 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34174 = ~w33882 & w34173 ;
  assign w34175 = w34172 | w34174 ;
  assign w34176 = ~\pi077 & w34175 ;
  assign w34177 = ~w33658 & w33742 ;
  assign w34178 = w33743 ^ w34177 ;
  assign w34179 = ~w33883 & w34178 ;
  assign w34180 = ( w33650 & w33881 ) | ( w33650 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34181 = ~w33882 & w34180 ;
  assign w34182 = w34179 | w34181 ;
  assign w34183 = ~\pi076 & w34182 ;
  assign w34184 = ~w33665 & w33739 ;
  assign w34185 = w33740 ^ w34184 ;
  assign w34186 = ~w33883 & w34185 ;
  assign w34187 = ( w33657 & w33881 ) | ( w33657 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34188 = ~w33882 & w34187 ;
  assign w34189 = w34186 | w34188 ;
  assign w34190 = ~\pi075 & w34189 ;
  assign w34191 = ~w33672 & w33736 ;
  assign w34192 = w33737 ^ w34191 ;
  assign w34193 = ~w33883 & w34192 ;
  assign w34194 = ( w33664 & w33881 ) | ( w33664 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34195 = ~w33882 & w34194 ;
  assign w34196 = w34193 | w34195 ;
  assign w34197 = ~\pi074 & w34196 ;
  assign w34198 = ~w33679 & w33733 ;
  assign w34199 = w33734 ^ w34198 ;
  assign w34200 = ~w33883 & w34199 ;
  assign w34201 = ( w33671 & w33881 ) | ( w33671 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34202 = ~w33882 & w34201 ;
  assign w34203 = w34200 | w34202 ;
  assign w34204 = ~\pi073 & w34203 ;
  assign w34205 = ~w33686 & w33730 ;
  assign w34206 = w33731 ^ w34205 ;
  assign w34207 = ~w33883 & w34206 ;
  assign w34208 = ( w33678 & w33881 ) | ( w33678 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34209 = ~w33882 & w34208 ;
  assign w34210 = w34207 | w34209 ;
  assign w34211 = ~\pi072 & w34210 ;
  assign w34212 = ~w33693 & w33727 ;
  assign w34213 = w33728 ^ w34212 ;
  assign w34214 = ~w33883 & w34213 ;
  assign w34215 = ( w33685 & w33881 ) | ( w33685 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34216 = ~w33882 & w34215 ;
  assign w34217 = w34214 | w34216 ;
  assign w34218 = ~\pi071 & w34217 ;
  assign w34219 = ~w33700 & w33724 ;
  assign w34220 = w33725 ^ w34219 ;
  assign w34221 = ~w33883 & w34220 ;
  assign w34222 = ( w33692 & w33881 ) | ( w33692 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34223 = ~w33882 & w34222 ;
  assign w34224 = w34221 | w34223 ;
  assign w34225 = ~\pi070 & w34224 ;
  assign w34226 = ~w33706 & w33721 ;
  assign w34227 = w33722 ^ w34226 ;
  assign w34228 = ~w33883 & w34227 ;
  assign w34229 = ( w33699 & w33881 ) | ( w33699 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34230 = ~w33882 & w34229 ;
  assign w34231 = w34228 | w34230 ;
  assign w34232 = ~\pi069 & w34231 ;
  assign w34233 = ~w33711 & w33718 ;
  assign w34234 = w33719 ^ w34233 ;
  assign w34235 = ~w33883 & w34234 ;
  assign w34236 = ( w33705 & w33881 ) | ( w33705 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34237 = ~w33882 & w34236 ;
  assign w34238 = w34235 | w34237 ;
  assign w34239 = ~\pi068 & w34238 ;
  assign w34240 = \pi064 & ~w33357 ;
  assign w34241 = \pi011 ^ w34240 ;
  assign w34242 = ( \pi065 & w14881 ) | ( \pi065 & ~w34241 ) | ( w14881 & ~w34241 ) ;
  assign w34243 = w33714 ^ w34242 ;
  assign w34244 = ~w33883 & w34243 ;
  assign w34245 = ( w33710 & w33881 ) | ( w33710 & w33882 ) | ( w33881 & w33882 ) ;
  assign w34246 = ~w33882 & w34245 ;
  assign w34247 = w34244 | w34246 ;
  assign w34248 = ~\pi067 & w34247 ;
  assign w34249 = \pi010 ^ w33357 ;
  assign w34250 = ( \pi064 & w33883 ) | ( \pi064 & w34249 ) | ( w33883 & w34249 ) ;
  assign w34251 = w14889 ^ w34250 ;
  assign w34252 = ~w33883 & w34251 ;
  assign w34253 = w33883 & w34241 ;
  assign w34254 = w34252 | w34253 ;
  assign w34255 = ~\pi066 & w34254 ;
  assign w34256 = \pi066 ^ w34254 ;
  assign w34257 = ( \pi064 & ~w33883 ) | ( \pi064 & w34256 ) | ( ~w33883 & w34256 ) ;
  assign w34258 = \pi010 ^ w34257 ;
  assign w34259 = ( \pi065 & w15371 ) | ( \pi065 & ~w34258 ) | ( w15371 & ~w34258 ) ;
  assign w34260 = w34256 | w34259 ;
  assign w34261 = \pi067 ^ w34247 ;
  assign w34262 = ( ~w34255 & w34260 ) | ( ~w34255 & w34261 ) | ( w34260 & w34261 ) ;
  assign w34263 = w34261 | w34262 ;
  assign w34264 = \pi068 ^ w34238 ;
  assign w34265 = ( ~w34248 & w34263 ) | ( ~w34248 & w34264 ) | ( w34263 & w34264 ) ;
  assign w34266 = w34264 | w34265 ;
  assign w34267 = \pi069 ^ w34231 ;
  assign w34268 = ( ~w34239 & w34266 ) | ( ~w34239 & w34267 ) | ( w34266 & w34267 ) ;
  assign w34269 = w34267 | w34268 ;
  assign w34270 = \pi070 ^ w34224 ;
  assign w34271 = ( ~w34232 & w34269 ) | ( ~w34232 & w34270 ) | ( w34269 & w34270 ) ;
  assign w34272 = w34270 | w34271 ;
  assign w34273 = \pi071 ^ w34217 ;
  assign w34274 = ( ~w34225 & w34272 ) | ( ~w34225 & w34273 ) | ( w34272 & w34273 ) ;
  assign w34275 = w34273 | w34274 ;
  assign w34276 = \pi072 ^ w34210 ;
  assign w34277 = ( ~w34218 & w34275 ) | ( ~w34218 & w34276 ) | ( w34275 & w34276 ) ;
  assign w34278 = w34276 | w34277 ;
  assign w34279 = \pi073 ^ w34203 ;
  assign w34280 = ( ~w34211 & w34278 ) | ( ~w34211 & w34279 ) | ( w34278 & w34279 ) ;
  assign w34281 = w34279 | w34280 ;
  assign w34282 = \pi074 ^ w34196 ;
  assign w34283 = ( ~w34204 & w34281 ) | ( ~w34204 & w34282 ) | ( w34281 & w34282 ) ;
  assign w34284 = w34282 | w34283 ;
  assign w34285 = \pi075 ^ w34189 ;
  assign w34286 = ( ~w34197 & w34284 ) | ( ~w34197 & w34285 ) | ( w34284 & w34285 ) ;
  assign w34287 = w34285 | w34286 ;
  assign w34288 = \pi076 ^ w34182 ;
  assign w34289 = ( ~w34190 & w34287 ) | ( ~w34190 & w34288 ) | ( w34287 & w34288 ) ;
  assign w34290 = w34288 | w34289 ;
  assign w34291 = \pi077 ^ w34175 ;
  assign w34292 = ( ~w34183 & w34290 ) | ( ~w34183 & w34291 ) | ( w34290 & w34291 ) ;
  assign w34293 = w34291 | w34292 ;
  assign w34294 = \pi078 ^ w34168 ;
  assign w34295 = ( ~w34176 & w34293 ) | ( ~w34176 & w34294 ) | ( w34293 & w34294 ) ;
  assign w34296 = w34294 | w34295 ;
  assign w34297 = \pi079 ^ w34161 ;
  assign w34298 = ( ~w34169 & w34296 ) | ( ~w34169 & w34297 ) | ( w34296 & w34297 ) ;
  assign w34299 = w34297 | w34298 ;
  assign w34300 = \pi080 ^ w34154 ;
  assign w34301 = ( ~w34162 & w34299 ) | ( ~w34162 & w34300 ) | ( w34299 & w34300 ) ;
  assign w34302 = w34300 | w34301 ;
  assign w34303 = \pi081 ^ w34147 ;
  assign w34304 = ( ~w34155 & w34302 ) | ( ~w34155 & w34303 ) | ( w34302 & w34303 ) ;
  assign w34305 = w34303 | w34304 ;
  assign w34306 = \pi082 ^ w34140 ;
  assign w34307 = ( ~w34148 & w34305 ) | ( ~w34148 & w34306 ) | ( w34305 & w34306 ) ;
  assign w34308 = w34306 | w34307 ;
  assign w34309 = \pi083 ^ w34133 ;
  assign w34310 = ( ~w34141 & w34308 ) | ( ~w34141 & w34309 ) | ( w34308 & w34309 ) ;
  assign w34311 = w34309 | w34310 ;
  assign w34312 = \pi084 ^ w34126 ;
  assign w34313 = ( ~w34134 & w34311 ) | ( ~w34134 & w34312 ) | ( w34311 & w34312 ) ;
  assign w34314 = w34312 | w34313 ;
  assign w34315 = \pi085 ^ w34119 ;
  assign w34316 = ( ~w34127 & w34314 ) | ( ~w34127 & w34315 ) | ( w34314 & w34315 ) ;
  assign w34317 = w34315 | w34316 ;
  assign w34318 = \pi086 ^ w34112 ;
  assign w34319 = ( ~w34120 & w34317 ) | ( ~w34120 & w34318 ) | ( w34317 & w34318 ) ;
  assign w34320 = w34318 | w34319 ;
  assign w34321 = \pi087 ^ w34105 ;
  assign w34322 = ( ~w34113 & w34320 ) | ( ~w34113 & w34321 ) | ( w34320 & w34321 ) ;
  assign w34323 = w34321 | w34322 ;
  assign w34324 = \pi088 ^ w34098 ;
  assign w34325 = ( ~w34106 & w34323 ) | ( ~w34106 & w34324 ) | ( w34323 & w34324 ) ;
  assign w34326 = w34324 | w34325 ;
  assign w34327 = \pi089 ^ w34091 ;
  assign w34328 = ( ~w34099 & w34326 ) | ( ~w34099 & w34327 ) | ( w34326 & w34327 ) ;
  assign w34329 = w34327 | w34328 ;
  assign w34330 = \pi090 ^ w34084 ;
  assign w34331 = ( ~w34092 & w34329 ) | ( ~w34092 & w34330 ) | ( w34329 & w34330 ) ;
  assign w34332 = w34330 | w34331 ;
  assign w34333 = \pi091 ^ w34077 ;
  assign w34334 = ( ~w34085 & w34332 ) | ( ~w34085 & w34333 ) | ( w34332 & w34333 ) ;
  assign w34335 = w34333 | w34334 ;
  assign w34336 = \pi092 ^ w34070 ;
  assign w34337 = ( ~w34078 & w34335 ) | ( ~w34078 & w34336 ) | ( w34335 & w34336 ) ;
  assign w34338 = w34336 | w34337 ;
  assign w34339 = \pi093 ^ w34063 ;
  assign w34340 = ( ~w34071 & w34338 ) | ( ~w34071 & w34339 ) | ( w34338 & w34339 ) ;
  assign w34341 = w34339 | w34340 ;
  assign w34342 = \pi094 ^ w34056 ;
  assign w34343 = ( ~w34064 & w34341 ) | ( ~w34064 & w34342 ) | ( w34341 & w34342 ) ;
  assign w34344 = w34342 | w34343 ;
  assign w34345 = \pi095 ^ w34049 ;
  assign w34346 = ( ~w34057 & w34344 ) | ( ~w34057 & w34345 ) | ( w34344 & w34345 ) ;
  assign w34347 = w34345 | w34346 ;
  assign w34348 = \pi096 ^ w34042 ;
  assign w34349 = ( ~w34050 & w34347 ) | ( ~w34050 & w34348 ) | ( w34347 & w34348 ) ;
  assign w34350 = w34348 | w34349 ;
  assign w34351 = \pi097 ^ w34035 ;
  assign w34352 = ( ~w34043 & w34350 ) | ( ~w34043 & w34351 ) | ( w34350 & w34351 ) ;
  assign w34353 = w34351 | w34352 ;
  assign w34354 = \pi098 ^ w34028 ;
  assign w34355 = ( ~w34036 & w34353 ) | ( ~w34036 & w34354 ) | ( w34353 & w34354 ) ;
  assign w34356 = w34354 | w34355 ;
  assign w34357 = \pi099 ^ w34021 ;
  assign w34358 = ( ~w34029 & w34356 ) | ( ~w34029 & w34357 ) | ( w34356 & w34357 ) ;
  assign w34359 = w34357 | w34358 ;
  assign w34360 = \pi100 ^ w34014 ;
  assign w34361 = ( ~w34022 & w34359 ) | ( ~w34022 & w34360 ) | ( w34359 & w34360 ) ;
  assign w34362 = w34360 | w34361 ;
  assign w34363 = \pi101 ^ w34007 ;
  assign w34364 = ( ~w34015 & w34362 ) | ( ~w34015 & w34363 ) | ( w34362 & w34363 ) ;
  assign w34365 = w34363 | w34364 ;
  assign w34366 = \pi102 ^ w34000 ;
  assign w34367 = ( ~w34008 & w34365 ) | ( ~w34008 & w34366 ) | ( w34365 & w34366 ) ;
  assign w34368 = w34366 | w34367 ;
  assign w34369 = \pi103 ^ w33993 ;
  assign w34370 = ( ~w34001 & w34368 ) | ( ~w34001 & w34369 ) | ( w34368 & w34369 ) ;
  assign w34371 = w34369 | w34370 ;
  assign w34372 = \pi104 ^ w33986 ;
  assign w34373 = ( ~w33994 & w34371 ) | ( ~w33994 & w34372 ) | ( w34371 & w34372 ) ;
  assign w34374 = w34372 | w34373 ;
  assign w34375 = \pi105 ^ w33979 ;
  assign w34376 = ( ~w33987 & w34374 ) | ( ~w33987 & w34375 ) | ( w34374 & w34375 ) ;
  assign w34377 = w34375 | w34376 ;
  assign w34378 = \pi106 ^ w33972 ;
  assign w34379 = ( ~w33980 & w34377 ) | ( ~w33980 & w34378 ) | ( w34377 & w34378 ) ;
  assign w34380 = w34378 | w34379 ;
  assign w34381 = \pi107 ^ w33965 ;
  assign w34382 = ( ~w33973 & w34380 ) | ( ~w33973 & w34381 ) | ( w34380 & w34381 ) ;
  assign w34383 = w34381 | w34382 ;
  assign w34384 = \pi108 ^ w33958 ;
  assign w34385 = ( ~w33966 & w34383 ) | ( ~w33966 & w34384 ) | ( w34383 & w34384 ) ;
  assign w34386 = w34384 | w34385 ;
  assign w34387 = \pi109 ^ w33951 ;
  assign w34388 = ( ~w33959 & w34386 ) | ( ~w33959 & w34387 ) | ( w34386 & w34387 ) ;
  assign w34389 = w34387 | w34388 ;
  assign w34390 = \pi110 ^ w33944 ;
  assign w34391 = ( ~w33952 & w34389 ) | ( ~w33952 & w34390 ) | ( w34389 & w34390 ) ;
  assign w34392 = w34390 | w34391 ;
  assign w34393 = \pi111 ^ w33937 ;
  assign w34394 = ( ~w33945 & w34392 ) | ( ~w33945 & w34393 ) | ( w34392 & w34393 ) ;
  assign w34395 = w34393 | w34394 ;
  assign w34396 = \pi112 ^ w33930 ;
  assign w34397 = ( ~w33938 & w34395 ) | ( ~w33938 & w34396 ) | ( w34395 & w34396 ) ;
  assign w34398 = w34396 | w34397 ;
  assign w34399 = \pi113 ^ w33923 ;
  assign w34400 = ( ~w33931 & w34398 ) | ( ~w33931 & w34399 ) | ( w34398 & w34399 ) ;
  assign w34401 = w34399 | w34400 ;
  assign w34402 = \pi114 ^ w33916 ;
  assign w34403 = ( ~w33924 & w34401 ) | ( ~w33924 & w34402 ) | ( w34401 & w34402 ) ;
  assign w34404 = w34402 | w34403 ;
  assign w34405 = \pi115 ^ w33909 ;
  assign w34406 = ( ~w33917 & w34404 ) | ( ~w33917 & w34405 ) | ( w34404 & w34405 ) ;
  assign w34407 = w34405 | w34406 ;
  assign w34408 = \pi116 ^ w33902 ;
  assign w34409 = ( ~w33910 & w34407 ) | ( ~w33910 & w34408 ) | ( w34407 & w34408 ) ;
  assign w34410 = w34408 | w34409 ;
  assign w34411 = \pi117 ^ w33889 ;
  assign w34412 = ( ~w33903 & w34410 ) | ( ~w33903 & w34411 ) | ( w34410 & w34411 ) ;
  assign w34413 = w34411 | w34412 ;
  assign w34414 = \pi118 ^ w33895 ;
  assign w34415 = w33896 & ~w34414 ;
  assign w34416 = ( w34413 & w34414 ) | ( w34413 & ~w34415 ) | ( w34414 & ~w34415 ) ;
  assign w34417 = ~\pi118 & w33895 ;
  assign w34418 = w34416 & ~w34417 ;
  assign w34419 = w15063 | w34418 ;
  assign w34420 = w33889 & w34419 ;
  assign w34421 = ~w33903 & w34410 ;
  assign w34422 = w34411 ^ w34421 ;
  assign w34423 = ~w34419 & w34422 ;
  assign w34424 = w34420 | w34423 ;
  assign w34425 = ~\pi118 & w34424 ;
  assign w34426 = w33902 & w34419 ;
  assign w34427 = ~w33910 & w34407 ;
  assign w34428 = w34408 ^ w34427 ;
  assign w34429 = ~w34419 & w34428 ;
  assign w34430 = w34426 | w34429 ;
  assign w34431 = ~\pi117 & w34430 ;
  assign w34432 = w33909 & w34419 ;
  assign w34433 = ~w33917 & w34404 ;
  assign w34434 = w34405 ^ w34433 ;
  assign w34435 = ~w34419 & w34434 ;
  assign w34436 = w34432 | w34435 ;
  assign w34437 = ~\pi116 & w34436 ;
  assign w34438 = w33916 & w34419 ;
  assign w34439 = ~w33924 & w34401 ;
  assign w34440 = w34402 ^ w34439 ;
  assign w34441 = ~w34419 & w34440 ;
  assign w34442 = w34438 | w34441 ;
  assign w34443 = ~\pi115 & w34442 ;
  assign w34444 = w33923 & w34419 ;
  assign w34445 = ~w33931 & w34398 ;
  assign w34446 = w34399 ^ w34445 ;
  assign w34447 = ~w34419 & w34446 ;
  assign w34448 = w34444 | w34447 ;
  assign w34449 = ~\pi114 & w34448 ;
  assign w34450 = w33930 & w34419 ;
  assign w34451 = ~w33938 & w34395 ;
  assign w34452 = w34396 ^ w34451 ;
  assign w34453 = ~w34419 & w34452 ;
  assign w34454 = w34450 | w34453 ;
  assign w34455 = ~\pi113 & w34454 ;
  assign w34456 = w33937 & w34419 ;
  assign w34457 = ~w33945 & w34392 ;
  assign w34458 = w34393 ^ w34457 ;
  assign w34459 = ~w34419 & w34458 ;
  assign w34460 = w34456 | w34459 ;
  assign w34461 = ~\pi112 & w34460 ;
  assign w34462 = w33944 & w34419 ;
  assign w34463 = ~w33952 & w34389 ;
  assign w34464 = w34390 ^ w34463 ;
  assign w34465 = ~w34419 & w34464 ;
  assign w34466 = w34462 | w34465 ;
  assign w34467 = ~\pi111 & w34466 ;
  assign w34468 = w33951 & w34419 ;
  assign w34469 = ~w33959 & w34386 ;
  assign w34470 = w34387 ^ w34469 ;
  assign w34471 = ~w34419 & w34470 ;
  assign w34472 = w34468 | w34471 ;
  assign w34473 = ~\pi110 & w34472 ;
  assign w34474 = w33958 & w34419 ;
  assign w34475 = ~w33966 & w34383 ;
  assign w34476 = w34384 ^ w34475 ;
  assign w34477 = ~w34419 & w34476 ;
  assign w34478 = w34474 | w34477 ;
  assign w34479 = ~\pi109 & w34478 ;
  assign w34480 = w33965 & w34419 ;
  assign w34481 = ~w33973 & w34380 ;
  assign w34482 = w34381 ^ w34481 ;
  assign w34483 = ~w34419 & w34482 ;
  assign w34484 = w34480 | w34483 ;
  assign w34485 = ~\pi108 & w34484 ;
  assign w34486 = w33972 & w34419 ;
  assign w34487 = ~w33980 & w34377 ;
  assign w34488 = w34378 ^ w34487 ;
  assign w34489 = ~w34419 & w34488 ;
  assign w34490 = w34486 | w34489 ;
  assign w34491 = ~\pi107 & w34490 ;
  assign w34492 = w33979 & w34419 ;
  assign w34493 = ~w33987 & w34374 ;
  assign w34494 = w34375 ^ w34493 ;
  assign w34495 = ~w34419 & w34494 ;
  assign w34496 = w34492 | w34495 ;
  assign w34497 = ~\pi106 & w34496 ;
  assign w34498 = w33986 & w34419 ;
  assign w34499 = ~w33994 & w34371 ;
  assign w34500 = w34372 ^ w34499 ;
  assign w34501 = ~w34419 & w34500 ;
  assign w34502 = w34498 | w34501 ;
  assign w34503 = ~\pi105 & w34502 ;
  assign w34504 = w33993 & w34419 ;
  assign w34505 = ~w34001 & w34368 ;
  assign w34506 = w34369 ^ w34505 ;
  assign w34507 = ~w34419 & w34506 ;
  assign w34508 = w34504 | w34507 ;
  assign w34509 = ~\pi104 & w34508 ;
  assign w34510 = w34000 & w34419 ;
  assign w34511 = ~w34008 & w34365 ;
  assign w34512 = w34366 ^ w34511 ;
  assign w34513 = ~w34419 & w34512 ;
  assign w34514 = w34510 | w34513 ;
  assign w34515 = ~\pi103 & w34514 ;
  assign w34516 = w34007 & w34419 ;
  assign w34517 = ~w34015 & w34362 ;
  assign w34518 = w34363 ^ w34517 ;
  assign w34519 = ~w34419 & w34518 ;
  assign w34520 = w34516 | w34519 ;
  assign w34521 = ~\pi102 & w34520 ;
  assign w34522 = w34014 & w34419 ;
  assign w34523 = ~w34022 & w34359 ;
  assign w34524 = w34360 ^ w34523 ;
  assign w34525 = ~w34419 & w34524 ;
  assign w34526 = w34522 | w34525 ;
  assign w34527 = ~\pi101 & w34526 ;
  assign w34528 = w34021 & w34419 ;
  assign w34529 = ~w34029 & w34356 ;
  assign w34530 = w34357 ^ w34529 ;
  assign w34531 = ~w34419 & w34530 ;
  assign w34532 = w34528 | w34531 ;
  assign w34533 = ~\pi100 & w34532 ;
  assign w34534 = w34028 & w34419 ;
  assign w34535 = ~w34036 & w34353 ;
  assign w34536 = w34354 ^ w34535 ;
  assign w34537 = ~w34419 & w34536 ;
  assign w34538 = w34534 | w34537 ;
  assign w34539 = ~\pi099 & w34538 ;
  assign w34540 = w34035 & w34419 ;
  assign w34541 = ~w34043 & w34350 ;
  assign w34542 = w34351 ^ w34541 ;
  assign w34543 = ~w34419 & w34542 ;
  assign w34544 = w34540 | w34543 ;
  assign w34545 = ~\pi098 & w34544 ;
  assign w34546 = w34042 & w34419 ;
  assign w34547 = ~w34050 & w34347 ;
  assign w34548 = w34348 ^ w34547 ;
  assign w34549 = ~w34419 & w34548 ;
  assign w34550 = w34546 | w34549 ;
  assign w34551 = ~\pi097 & w34550 ;
  assign w34552 = w34049 & w34419 ;
  assign w34553 = ~w34057 & w34344 ;
  assign w34554 = w34345 ^ w34553 ;
  assign w34555 = ~w34419 & w34554 ;
  assign w34556 = w34552 | w34555 ;
  assign w34557 = ~\pi096 & w34556 ;
  assign w34558 = w34056 & w34419 ;
  assign w34559 = ~w34064 & w34341 ;
  assign w34560 = w34342 ^ w34559 ;
  assign w34561 = ~w34419 & w34560 ;
  assign w34562 = w34558 | w34561 ;
  assign w34563 = ~\pi095 & w34562 ;
  assign w34564 = w34063 & w34419 ;
  assign w34565 = ~w34071 & w34338 ;
  assign w34566 = w34339 ^ w34565 ;
  assign w34567 = ~w34419 & w34566 ;
  assign w34568 = w34564 | w34567 ;
  assign w34569 = ~\pi094 & w34568 ;
  assign w34570 = w34070 & w34419 ;
  assign w34571 = ~w34078 & w34335 ;
  assign w34572 = w34336 ^ w34571 ;
  assign w34573 = ~w34419 & w34572 ;
  assign w34574 = w34570 | w34573 ;
  assign w34575 = ~\pi093 & w34574 ;
  assign w34576 = w34077 & w34419 ;
  assign w34577 = ~w34085 & w34332 ;
  assign w34578 = w34333 ^ w34577 ;
  assign w34579 = ~w34419 & w34578 ;
  assign w34580 = w34576 | w34579 ;
  assign w34581 = ~\pi092 & w34580 ;
  assign w34582 = w34084 & w34419 ;
  assign w34583 = ~w34092 & w34329 ;
  assign w34584 = w34330 ^ w34583 ;
  assign w34585 = ~w34419 & w34584 ;
  assign w34586 = w34582 | w34585 ;
  assign w34587 = ~\pi091 & w34586 ;
  assign w34588 = w34091 & w34419 ;
  assign w34589 = ~w34099 & w34326 ;
  assign w34590 = w34327 ^ w34589 ;
  assign w34591 = ~w34419 & w34590 ;
  assign w34592 = w34588 | w34591 ;
  assign w34593 = ~\pi090 & w34592 ;
  assign w34594 = w34098 & w34419 ;
  assign w34595 = ~w34106 & w34323 ;
  assign w34596 = w34324 ^ w34595 ;
  assign w34597 = ~w34419 & w34596 ;
  assign w34598 = w34594 | w34597 ;
  assign w34599 = ~\pi089 & w34598 ;
  assign w34600 = w34105 & w34419 ;
  assign w34601 = ~w34113 & w34320 ;
  assign w34602 = w34321 ^ w34601 ;
  assign w34603 = ~w34419 & w34602 ;
  assign w34604 = w34600 | w34603 ;
  assign w34605 = ~\pi088 & w34604 ;
  assign w34606 = w34112 & w34419 ;
  assign w34607 = ~w34120 & w34317 ;
  assign w34608 = w34318 ^ w34607 ;
  assign w34609 = ~w34419 & w34608 ;
  assign w34610 = w34606 | w34609 ;
  assign w34611 = ~\pi087 & w34610 ;
  assign w34612 = w34119 & w34419 ;
  assign w34613 = ~w34127 & w34314 ;
  assign w34614 = w34315 ^ w34613 ;
  assign w34615 = ~w34419 & w34614 ;
  assign w34616 = w34612 | w34615 ;
  assign w34617 = ~\pi086 & w34616 ;
  assign w34618 = w34126 & w34419 ;
  assign w34619 = ~w34134 & w34311 ;
  assign w34620 = w34312 ^ w34619 ;
  assign w34621 = ~w34419 & w34620 ;
  assign w34622 = w34618 | w34621 ;
  assign w34623 = ~\pi085 & w34622 ;
  assign w34624 = w34133 & w34419 ;
  assign w34625 = ~w34141 & w34308 ;
  assign w34626 = w34309 ^ w34625 ;
  assign w34627 = ~w34419 & w34626 ;
  assign w34628 = w34624 | w34627 ;
  assign w34629 = ~\pi084 & w34628 ;
  assign w34630 = w34140 & w34419 ;
  assign w34631 = ~w34148 & w34305 ;
  assign w34632 = w34306 ^ w34631 ;
  assign w34633 = ~w34419 & w34632 ;
  assign w34634 = w34630 | w34633 ;
  assign w34635 = ~\pi083 & w34634 ;
  assign w34636 = w34147 & w34419 ;
  assign w34637 = ~w34155 & w34302 ;
  assign w34638 = w34303 ^ w34637 ;
  assign w34639 = ~w34419 & w34638 ;
  assign w34640 = w34636 | w34639 ;
  assign w34641 = ~\pi082 & w34640 ;
  assign w34642 = w34154 & w34419 ;
  assign w34643 = ~w34162 & w34299 ;
  assign w34644 = w34300 ^ w34643 ;
  assign w34645 = ~w34419 & w34644 ;
  assign w34646 = w34642 | w34645 ;
  assign w34647 = ~\pi081 & w34646 ;
  assign w34648 = w34161 & w34419 ;
  assign w34649 = ~w34169 & w34296 ;
  assign w34650 = w34297 ^ w34649 ;
  assign w34651 = ~w34419 & w34650 ;
  assign w34652 = w34648 | w34651 ;
  assign w34653 = ~\pi080 & w34652 ;
  assign w34654 = w34168 & w34419 ;
  assign w34655 = ~w34176 & w34293 ;
  assign w34656 = w34294 ^ w34655 ;
  assign w34657 = ~w34419 & w34656 ;
  assign w34658 = w34654 | w34657 ;
  assign w34659 = ~\pi079 & w34658 ;
  assign w34660 = w34175 & w34419 ;
  assign w34661 = ~w34183 & w34290 ;
  assign w34662 = w34291 ^ w34661 ;
  assign w34663 = ~w34419 & w34662 ;
  assign w34664 = w34660 | w34663 ;
  assign w34665 = ~\pi078 & w34664 ;
  assign w34666 = w34182 & w34419 ;
  assign w34667 = ~w34190 & w34287 ;
  assign w34668 = w34288 ^ w34667 ;
  assign w34669 = ~w34419 & w34668 ;
  assign w34670 = w34666 | w34669 ;
  assign w34671 = ~\pi077 & w34670 ;
  assign w34672 = w34189 & w34419 ;
  assign w34673 = ~w34197 & w34284 ;
  assign w34674 = w34285 ^ w34673 ;
  assign w34675 = ~w34419 & w34674 ;
  assign w34676 = w34672 | w34675 ;
  assign w34677 = ~\pi076 & w34676 ;
  assign w34678 = w34196 & w34419 ;
  assign w34679 = ~w34204 & w34281 ;
  assign w34680 = w34282 ^ w34679 ;
  assign w34681 = ~w34419 & w34680 ;
  assign w34682 = w34678 | w34681 ;
  assign w34683 = ~\pi075 & w34682 ;
  assign w34684 = w34203 & w34419 ;
  assign w34685 = ~w34211 & w34278 ;
  assign w34686 = w34279 ^ w34685 ;
  assign w34687 = ~w34419 & w34686 ;
  assign w34688 = w34684 | w34687 ;
  assign w34689 = ~\pi074 & w34688 ;
  assign w34690 = w34210 & w34419 ;
  assign w34691 = ~w34218 & w34275 ;
  assign w34692 = w34276 ^ w34691 ;
  assign w34693 = ~w34419 & w34692 ;
  assign w34694 = w34690 | w34693 ;
  assign w34695 = ~\pi073 & w34694 ;
  assign w34696 = w34217 & w34419 ;
  assign w34697 = ~w34225 & w34272 ;
  assign w34698 = w34273 ^ w34697 ;
  assign w34699 = ~w34419 & w34698 ;
  assign w34700 = w34696 | w34699 ;
  assign w34701 = ~\pi072 & w34700 ;
  assign w34702 = w34224 & w34419 ;
  assign w34703 = ~w34232 & w34269 ;
  assign w34704 = w34270 ^ w34703 ;
  assign w34705 = ~w34419 & w34704 ;
  assign w34706 = w34702 | w34705 ;
  assign w34707 = ~\pi071 & w34706 ;
  assign w34708 = w34231 & w34419 ;
  assign w34709 = ~w34239 & w34266 ;
  assign w34710 = w34267 ^ w34709 ;
  assign w34711 = ~w34419 & w34710 ;
  assign w34712 = w34708 | w34711 ;
  assign w34713 = ~\pi070 & w34712 ;
  assign w34714 = w34238 & w34419 ;
  assign w34715 = ~w34248 & w34263 ;
  assign w34716 = w34264 ^ w34715 ;
  assign w34717 = ~w34419 & w34716 ;
  assign w34718 = w34714 | w34717 ;
  assign w34719 = ~\pi069 & w34718 ;
  assign w34720 = w34247 & w34419 ;
  assign w34721 = ~w34255 & w34260 ;
  assign w34722 = w34261 ^ w34721 ;
  assign w34723 = ~w34419 & w34722 ;
  assign w34724 = w34720 | w34723 ;
  assign w34725 = ~\pi068 & w34724 ;
  assign w34726 = \pi064 & ~w33883 ;
  assign w34727 = \pi010 ^ w34726 ;
  assign w34728 = ( \pi065 & w15371 ) | ( \pi065 & ~w34727 ) | ( w15371 & ~w34727 ) ;
  assign w34729 = w34256 ^ w34728 ;
  assign w34730 = ( w15063 & w34418 ) | ( w15063 & w34729 ) | ( w34418 & w34729 ) ;
  assign w34731 = w34729 & ~w34730 ;
  assign w34732 = ( w34254 & w34419 ) | ( w34254 & w34731 ) | ( w34419 & w34731 ) ;
  assign w34733 = w34731 | w34732 ;
  assign w34734 = ~\pi067 & w34733 ;
  assign w34735 = \pi009 ^ w33883 ;
  assign w34736 = ( \pi064 & w15063 ) | ( \pi064 & w34735 ) | ( w15063 & w34735 ) ;
  assign w34737 = w15379 ^ w34736 ;
  assign w34738 = ~w15063 & w34737 ;
  assign w34739 = ~w34418 & w34738 ;
  assign w34740 = ( ~\pi064 & w33883 ) | ( ~\pi064 & w34419 ) | ( w33883 & w34419 ) ;
  assign w34741 = \pi010 ^ w34740 ;
  assign w34742 = w34419 & ~w34741 ;
  assign w34743 = w34739 | w34742 ;
  assign w34744 = ~\pi066 & w34743 ;
  assign w34745 = ( \pi064 & w15392 ) | ( \pi064 & w34418 ) | ( w15392 & w34418 ) ;
  assign w34746 = ( \pi009 & ~\pi064 ) | ( \pi009 & w34745 ) | ( ~\pi064 & w34745 ) ;
  assign w34747 = w15398 & ~w34418 ;
  assign w34748 = w34419 | w34739 ;
  assign w34749 = ( w34727 & w34739 ) | ( w34727 & w34748 ) | ( w34739 & w34748 ) ;
  assign w34750 = \pi066 ^ w34749 ;
  assign w34751 = w34746 | w34747 ;
  assign w34752 = ( \pi065 & w15400 ) | ( \pi065 & ~w34751 ) | ( w15400 & ~w34751 ) ;
  assign w34753 = w34750 | w34752 ;
  assign w34754 = ~w34254 & w34419 ;
  assign w34755 = ( w34419 & w34731 ) | ( w34419 & ~w34754 ) | ( w34731 & ~w34754 ) ;
  assign w34756 = \pi067 ^ w34755 ;
  assign w34757 = ( ~w34744 & w34753 ) | ( ~w34744 & w34756 ) | ( w34753 & w34756 ) ;
  assign w34758 = w34756 | w34757 ;
  assign w34759 = \pi068 ^ w34724 ;
  assign w34760 = ( ~w34734 & w34758 ) | ( ~w34734 & w34759 ) | ( w34758 & w34759 ) ;
  assign w34761 = w34759 | w34760 ;
  assign w34762 = \pi069 ^ w34718 ;
  assign w34763 = ( ~w34725 & w34761 ) | ( ~w34725 & w34762 ) | ( w34761 & w34762 ) ;
  assign w34764 = w34762 | w34763 ;
  assign w34765 = \pi070 ^ w34712 ;
  assign w34766 = ( ~w34719 & w34764 ) | ( ~w34719 & w34765 ) | ( w34764 & w34765 ) ;
  assign w34767 = w34765 | w34766 ;
  assign w34768 = \pi071 ^ w34706 ;
  assign w34769 = ( ~w34713 & w34767 ) | ( ~w34713 & w34768 ) | ( w34767 & w34768 ) ;
  assign w34770 = w34768 | w34769 ;
  assign w34771 = \pi072 ^ w34700 ;
  assign w34772 = ( ~w34707 & w34770 ) | ( ~w34707 & w34771 ) | ( w34770 & w34771 ) ;
  assign w34773 = w34771 | w34772 ;
  assign w34774 = \pi073 ^ w34694 ;
  assign w34775 = ( ~w34701 & w34773 ) | ( ~w34701 & w34774 ) | ( w34773 & w34774 ) ;
  assign w34776 = w34774 | w34775 ;
  assign w34777 = \pi074 ^ w34688 ;
  assign w34778 = ( ~w34695 & w34776 ) | ( ~w34695 & w34777 ) | ( w34776 & w34777 ) ;
  assign w34779 = w34777 | w34778 ;
  assign w34780 = \pi075 ^ w34682 ;
  assign w34781 = ( ~w34689 & w34779 ) | ( ~w34689 & w34780 ) | ( w34779 & w34780 ) ;
  assign w34782 = w34780 | w34781 ;
  assign w34783 = \pi076 ^ w34676 ;
  assign w34784 = ( ~w34683 & w34782 ) | ( ~w34683 & w34783 ) | ( w34782 & w34783 ) ;
  assign w34785 = w34783 | w34784 ;
  assign w34786 = \pi077 ^ w34670 ;
  assign w34787 = ( ~w34677 & w34785 ) | ( ~w34677 & w34786 ) | ( w34785 & w34786 ) ;
  assign w34788 = w34786 | w34787 ;
  assign w34789 = \pi078 ^ w34664 ;
  assign w34790 = ( ~w34671 & w34788 ) | ( ~w34671 & w34789 ) | ( w34788 & w34789 ) ;
  assign w34791 = w34789 | w34790 ;
  assign w34792 = \pi079 ^ w34658 ;
  assign w34793 = ( ~w34665 & w34791 ) | ( ~w34665 & w34792 ) | ( w34791 & w34792 ) ;
  assign w34794 = w34792 | w34793 ;
  assign w34795 = \pi080 ^ w34652 ;
  assign w34796 = ( ~w34659 & w34794 ) | ( ~w34659 & w34795 ) | ( w34794 & w34795 ) ;
  assign w34797 = w34795 | w34796 ;
  assign w34798 = \pi081 ^ w34646 ;
  assign w34799 = ( ~w34653 & w34797 ) | ( ~w34653 & w34798 ) | ( w34797 & w34798 ) ;
  assign w34800 = w34798 | w34799 ;
  assign w34801 = \pi082 ^ w34640 ;
  assign w34802 = ( ~w34647 & w34800 ) | ( ~w34647 & w34801 ) | ( w34800 & w34801 ) ;
  assign w34803 = w34801 | w34802 ;
  assign w34804 = \pi083 ^ w34634 ;
  assign w34805 = ( ~w34641 & w34803 ) | ( ~w34641 & w34804 ) | ( w34803 & w34804 ) ;
  assign w34806 = w34804 | w34805 ;
  assign w34807 = \pi084 ^ w34628 ;
  assign w34808 = ( ~w34635 & w34806 ) | ( ~w34635 & w34807 ) | ( w34806 & w34807 ) ;
  assign w34809 = w34807 | w34808 ;
  assign w34810 = \pi085 ^ w34622 ;
  assign w34811 = ( ~w34629 & w34809 ) | ( ~w34629 & w34810 ) | ( w34809 & w34810 ) ;
  assign w34812 = w34810 | w34811 ;
  assign w34813 = \pi086 ^ w34616 ;
  assign w34814 = ( ~w34623 & w34812 ) | ( ~w34623 & w34813 ) | ( w34812 & w34813 ) ;
  assign w34815 = w34813 | w34814 ;
  assign w34816 = \pi087 ^ w34610 ;
  assign w34817 = ( ~w34617 & w34815 ) | ( ~w34617 & w34816 ) | ( w34815 & w34816 ) ;
  assign w34818 = w34816 | w34817 ;
  assign w34819 = \pi088 ^ w34604 ;
  assign w34820 = ( ~w34611 & w34818 ) | ( ~w34611 & w34819 ) | ( w34818 & w34819 ) ;
  assign w34821 = w34819 | w34820 ;
  assign w34822 = \pi089 ^ w34598 ;
  assign w34823 = ( ~w34605 & w34821 ) | ( ~w34605 & w34822 ) | ( w34821 & w34822 ) ;
  assign w34824 = w34822 | w34823 ;
  assign w34825 = \pi090 ^ w34592 ;
  assign w34826 = ( ~w34599 & w34824 ) | ( ~w34599 & w34825 ) | ( w34824 & w34825 ) ;
  assign w34827 = w34825 | w34826 ;
  assign w34828 = \pi091 ^ w34586 ;
  assign w34829 = ( ~w34593 & w34827 ) | ( ~w34593 & w34828 ) | ( w34827 & w34828 ) ;
  assign w34830 = w34828 | w34829 ;
  assign w34831 = \pi092 ^ w34580 ;
  assign w34832 = ( ~w34587 & w34830 ) | ( ~w34587 & w34831 ) | ( w34830 & w34831 ) ;
  assign w34833 = w34831 | w34832 ;
  assign w34834 = \pi093 ^ w34574 ;
  assign w34835 = ( ~w34581 & w34833 ) | ( ~w34581 & w34834 ) | ( w34833 & w34834 ) ;
  assign w34836 = w34834 | w34835 ;
  assign w34837 = \pi094 ^ w34568 ;
  assign w34838 = ( ~w34575 & w34836 ) | ( ~w34575 & w34837 ) | ( w34836 & w34837 ) ;
  assign w34839 = w34837 | w34838 ;
  assign w34840 = \pi095 ^ w34562 ;
  assign w34841 = ( ~w34569 & w34839 ) | ( ~w34569 & w34840 ) | ( w34839 & w34840 ) ;
  assign w34842 = w34840 | w34841 ;
  assign w34843 = \pi096 ^ w34556 ;
  assign w34844 = ( ~w34563 & w34842 ) | ( ~w34563 & w34843 ) | ( w34842 & w34843 ) ;
  assign w34845 = w34843 | w34844 ;
  assign w34846 = \pi097 ^ w34550 ;
  assign w34847 = ( ~w34557 & w34845 ) | ( ~w34557 & w34846 ) | ( w34845 & w34846 ) ;
  assign w34848 = w34846 | w34847 ;
  assign w34849 = \pi098 ^ w34544 ;
  assign w34850 = ( ~w34551 & w34848 ) | ( ~w34551 & w34849 ) | ( w34848 & w34849 ) ;
  assign w34851 = w34849 | w34850 ;
  assign w34852 = \pi099 ^ w34538 ;
  assign w34853 = ( ~w34545 & w34851 ) | ( ~w34545 & w34852 ) | ( w34851 & w34852 ) ;
  assign w34854 = w34852 | w34853 ;
  assign w34855 = \pi100 ^ w34532 ;
  assign w34856 = ( ~w34539 & w34854 ) | ( ~w34539 & w34855 ) | ( w34854 & w34855 ) ;
  assign w34857 = w34855 | w34856 ;
  assign w34858 = \pi101 ^ w34526 ;
  assign w34859 = ( ~w34533 & w34857 ) | ( ~w34533 & w34858 ) | ( w34857 & w34858 ) ;
  assign w34860 = w34858 | w34859 ;
  assign w34861 = \pi102 ^ w34520 ;
  assign w34862 = ( ~w34527 & w34860 ) | ( ~w34527 & w34861 ) | ( w34860 & w34861 ) ;
  assign w34863 = w34861 | w34862 ;
  assign w34864 = \pi103 ^ w34514 ;
  assign w34865 = ( ~w34521 & w34863 ) | ( ~w34521 & w34864 ) | ( w34863 & w34864 ) ;
  assign w34866 = w34864 | w34865 ;
  assign w34867 = \pi104 ^ w34508 ;
  assign w34868 = ( ~w34515 & w34866 ) | ( ~w34515 & w34867 ) | ( w34866 & w34867 ) ;
  assign w34869 = w34867 | w34868 ;
  assign w34870 = \pi105 ^ w34502 ;
  assign w34871 = ( ~w34509 & w34869 ) | ( ~w34509 & w34870 ) | ( w34869 & w34870 ) ;
  assign w34872 = w34870 | w34871 ;
  assign w34873 = \pi106 ^ w34496 ;
  assign w34874 = ( ~w34503 & w34872 ) | ( ~w34503 & w34873 ) | ( w34872 & w34873 ) ;
  assign w34875 = w34873 | w34874 ;
  assign w34876 = \pi107 ^ w34490 ;
  assign w34877 = ( ~w34497 & w34875 ) | ( ~w34497 & w34876 ) | ( w34875 & w34876 ) ;
  assign w34878 = w34876 | w34877 ;
  assign w34879 = \pi108 ^ w34484 ;
  assign w34880 = ( ~w34491 & w34878 ) | ( ~w34491 & w34879 ) | ( w34878 & w34879 ) ;
  assign w34881 = w34879 | w34880 ;
  assign w34882 = \pi109 ^ w34478 ;
  assign w34883 = ( ~w34485 & w34881 ) | ( ~w34485 & w34882 ) | ( w34881 & w34882 ) ;
  assign w34884 = w34882 | w34883 ;
  assign w34885 = \pi110 ^ w34472 ;
  assign w34886 = ( ~w34479 & w34884 ) | ( ~w34479 & w34885 ) | ( w34884 & w34885 ) ;
  assign w34887 = w34885 | w34886 ;
  assign w34888 = \pi111 ^ w34466 ;
  assign w34889 = ( ~w34473 & w34887 ) | ( ~w34473 & w34888 ) | ( w34887 & w34888 ) ;
  assign w34890 = w34888 | w34889 ;
  assign w34891 = \pi112 ^ w34460 ;
  assign w34892 = ( ~w34467 & w34890 ) | ( ~w34467 & w34891 ) | ( w34890 & w34891 ) ;
  assign w34893 = w34891 | w34892 ;
  assign w34894 = \pi113 ^ w34454 ;
  assign w34895 = ( ~w34461 & w34893 ) | ( ~w34461 & w34894 ) | ( w34893 & w34894 ) ;
  assign w34896 = w34894 | w34895 ;
  assign w34897 = \pi114 ^ w34448 ;
  assign w34898 = ( ~w34455 & w34896 ) | ( ~w34455 & w34897 ) | ( w34896 & w34897 ) ;
  assign w34899 = w34897 | w34898 ;
  assign w34900 = \pi115 ^ w34442 ;
  assign w34901 = ( ~w34449 & w34899 ) | ( ~w34449 & w34900 ) | ( w34899 & w34900 ) ;
  assign w34902 = w34900 | w34901 ;
  assign w34903 = \pi116 ^ w34436 ;
  assign w34904 = ( ~w34443 & w34902 ) | ( ~w34443 & w34903 ) | ( w34902 & w34903 ) ;
  assign w34905 = w34903 | w34904 ;
  assign w34906 = \pi117 ^ w34430 ;
  assign w34907 = ( ~w34437 & w34905 ) | ( ~w34437 & w34906 ) | ( w34905 & w34906 ) ;
  assign w34908 = w34906 | w34907 ;
  assign w34909 = \pi118 ^ w34424 ;
  assign w34910 = ( ~w34431 & w34908 ) | ( ~w34431 & w34909 ) | ( w34908 & w34909 ) ;
  assign w34911 = w34909 | w34910 ;
  assign w34912 = w33895 & w34419 ;
  assign w34913 = ~w33896 & w34413 ;
  assign w34914 = w34414 ^ w34913 ;
  assign w34915 = ~w34419 & w34914 ;
  assign w34916 = w34912 | w34915 ;
  assign w34917 = ~\pi119 & w34916 ;
  assign w34918 = ( \pi119 & ~w34912 ) | ( \pi119 & w34915 ) | ( ~w34912 & w34915 ) ;
  assign w34919 = ~w34915 & w34918 ;
  assign w34920 = w34917 | w34919 ;
  assign w34921 = ( ~w34425 & w34911 ) | ( ~w34425 & w34920 ) | ( w34911 & w34920 ) ;
  assign w34922 = ( w199 & ~w34920 ) | ( w199 & w34921 ) | ( ~w34920 & w34921 ) ;
  assign w34923 = w34920 | w34922 ;
  assign w34924 = ~w15063 & w34916 ;
  assign w34925 = w34923 & ~w34924 ;
  assign w34926 = ~w34431 & w34908 ;
  assign w34927 = w34909 ^ w34926 ;
  assign w34928 = ~w34925 & w34927 ;
  assign w34929 = ( w34424 & w34923 ) | ( w34424 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34930 = ~w34924 & w34929 ;
  assign w34931 = w34928 | w34930 ;
  assign w34932 = ~\pi119 & w34931 ;
  assign w34933 = ~w34437 & w34905 ;
  assign w34934 = w34906 ^ w34933 ;
  assign w34935 = ~w34925 & w34934 ;
  assign w34936 = ( w34430 & w34923 ) | ( w34430 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34937 = ~w34924 & w34936 ;
  assign w34938 = w34935 | w34937 ;
  assign w34939 = ~\pi118 & w34938 ;
  assign w34940 = ~w34443 & w34902 ;
  assign w34941 = w34903 ^ w34940 ;
  assign w34942 = ~w34925 & w34941 ;
  assign w34943 = ( w34436 & w34923 ) | ( w34436 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34944 = ~w34924 & w34943 ;
  assign w34945 = w34942 | w34944 ;
  assign w34946 = ~\pi117 & w34945 ;
  assign w34947 = ~w34449 & w34899 ;
  assign w34948 = w34900 ^ w34947 ;
  assign w34949 = ~w34925 & w34948 ;
  assign w34950 = ( w34442 & w34923 ) | ( w34442 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34951 = ~w34924 & w34950 ;
  assign w34952 = w34949 | w34951 ;
  assign w34953 = ~\pi116 & w34952 ;
  assign w34954 = ~w34455 & w34896 ;
  assign w34955 = w34897 ^ w34954 ;
  assign w34956 = ~w34925 & w34955 ;
  assign w34957 = ( w34448 & w34923 ) | ( w34448 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34958 = ~w34924 & w34957 ;
  assign w34959 = w34956 | w34958 ;
  assign w34960 = ~\pi115 & w34959 ;
  assign w34961 = ~w34461 & w34893 ;
  assign w34962 = w34894 ^ w34961 ;
  assign w34963 = ~w34925 & w34962 ;
  assign w34964 = ( w34454 & w34923 ) | ( w34454 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34965 = ~w34924 & w34964 ;
  assign w34966 = w34963 | w34965 ;
  assign w34967 = ~\pi114 & w34966 ;
  assign w34968 = ~w34467 & w34890 ;
  assign w34969 = w34891 ^ w34968 ;
  assign w34970 = ~w34925 & w34969 ;
  assign w34971 = ( w34460 & w34923 ) | ( w34460 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34972 = ~w34924 & w34971 ;
  assign w34973 = w34970 | w34972 ;
  assign w34974 = ~\pi113 & w34973 ;
  assign w34975 = ~w34473 & w34887 ;
  assign w34976 = w34888 ^ w34975 ;
  assign w34977 = ~w34925 & w34976 ;
  assign w34978 = ( w34466 & w34923 ) | ( w34466 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34979 = ~w34924 & w34978 ;
  assign w34980 = w34977 | w34979 ;
  assign w34981 = ~\pi112 & w34980 ;
  assign w34982 = ~w34479 & w34884 ;
  assign w34983 = w34885 ^ w34982 ;
  assign w34984 = ~w34925 & w34983 ;
  assign w34985 = ( w34472 & w34923 ) | ( w34472 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34986 = ~w34924 & w34985 ;
  assign w34987 = w34984 | w34986 ;
  assign w34988 = ~\pi111 & w34987 ;
  assign w34989 = ~w34485 & w34881 ;
  assign w34990 = w34882 ^ w34989 ;
  assign w34991 = ~w34925 & w34990 ;
  assign w34992 = ( w34478 & w34923 ) | ( w34478 & w34924 ) | ( w34923 & w34924 ) ;
  assign w34993 = ~w34924 & w34992 ;
  assign w34994 = w34991 | w34993 ;
  assign w34995 = ~\pi110 & w34994 ;
  assign w34996 = ~w34491 & w34878 ;
  assign w34997 = w34879 ^ w34996 ;
  assign w34998 = ~w34925 & w34997 ;
  assign w34999 = ( w34484 & w34923 ) | ( w34484 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35000 = ~w34924 & w34999 ;
  assign w35001 = w34998 | w35000 ;
  assign w35002 = ~\pi109 & w35001 ;
  assign w35003 = ~w34497 & w34875 ;
  assign w35004 = w34876 ^ w35003 ;
  assign w35005 = ~w34925 & w35004 ;
  assign w35006 = ( w34490 & w34923 ) | ( w34490 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35007 = ~w34924 & w35006 ;
  assign w35008 = w35005 | w35007 ;
  assign w35009 = ~\pi108 & w35008 ;
  assign w35010 = ~w34503 & w34872 ;
  assign w35011 = w34873 ^ w35010 ;
  assign w35012 = ~w34925 & w35011 ;
  assign w35013 = ( w34496 & w34923 ) | ( w34496 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35014 = ~w34924 & w35013 ;
  assign w35015 = w35012 | w35014 ;
  assign w35016 = ~\pi107 & w35015 ;
  assign w35017 = ~w34509 & w34869 ;
  assign w35018 = w34870 ^ w35017 ;
  assign w35019 = ~w34925 & w35018 ;
  assign w35020 = ( w34502 & w34923 ) | ( w34502 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35021 = ~w34924 & w35020 ;
  assign w35022 = w35019 | w35021 ;
  assign w35023 = ~\pi106 & w35022 ;
  assign w35024 = ~w34515 & w34866 ;
  assign w35025 = w34867 ^ w35024 ;
  assign w35026 = ~w34925 & w35025 ;
  assign w35027 = ( w34508 & w34923 ) | ( w34508 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35028 = ~w34924 & w35027 ;
  assign w35029 = w35026 | w35028 ;
  assign w35030 = ~\pi105 & w35029 ;
  assign w35031 = ~w34521 & w34863 ;
  assign w35032 = w34864 ^ w35031 ;
  assign w35033 = ~w34925 & w35032 ;
  assign w35034 = ( w34514 & w34923 ) | ( w34514 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35035 = ~w34924 & w35034 ;
  assign w35036 = w35033 | w35035 ;
  assign w35037 = ~\pi104 & w35036 ;
  assign w35038 = ~w34527 & w34860 ;
  assign w35039 = w34861 ^ w35038 ;
  assign w35040 = ~w34925 & w35039 ;
  assign w35041 = ( w34520 & w34923 ) | ( w34520 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35042 = ~w34924 & w35041 ;
  assign w35043 = w35040 | w35042 ;
  assign w35044 = ~\pi103 & w35043 ;
  assign w35045 = ~w34533 & w34857 ;
  assign w35046 = w34858 ^ w35045 ;
  assign w35047 = ~w34925 & w35046 ;
  assign w35048 = ( w34526 & w34923 ) | ( w34526 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35049 = ~w34924 & w35048 ;
  assign w35050 = w35047 | w35049 ;
  assign w35051 = ~\pi102 & w35050 ;
  assign w35052 = ~w34539 & w34854 ;
  assign w35053 = w34855 ^ w35052 ;
  assign w35054 = ~w34925 & w35053 ;
  assign w35055 = ( w34532 & w34923 ) | ( w34532 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35056 = ~w34924 & w35055 ;
  assign w35057 = w35054 | w35056 ;
  assign w35058 = ~\pi101 & w35057 ;
  assign w35059 = ~w34545 & w34851 ;
  assign w35060 = w34852 ^ w35059 ;
  assign w35061 = ~w34925 & w35060 ;
  assign w35062 = ( w34538 & w34923 ) | ( w34538 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35063 = ~w34924 & w35062 ;
  assign w35064 = w35061 | w35063 ;
  assign w35065 = ~\pi100 & w35064 ;
  assign w35066 = ~w34551 & w34848 ;
  assign w35067 = w34849 ^ w35066 ;
  assign w35068 = ~w34925 & w35067 ;
  assign w35069 = ( w34544 & w34923 ) | ( w34544 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35070 = ~w34924 & w35069 ;
  assign w35071 = w35068 | w35070 ;
  assign w35072 = ~\pi099 & w35071 ;
  assign w35073 = ~w34557 & w34845 ;
  assign w35074 = w34846 ^ w35073 ;
  assign w35075 = ~w34925 & w35074 ;
  assign w35076 = ( w34550 & w34923 ) | ( w34550 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35077 = ~w34924 & w35076 ;
  assign w35078 = w35075 | w35077 ;
  assign w35079 = ~\pi098 & w35078 ;
  assign w35080 = ~w34563 & w34842 ;
  assign w35081 = w34843 ^ w35080 ;
  assign w35082 = ~w34925 & w35081 ;
  assign w35083 = ( w34556 & w34923 ) | ( w34556 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35084 = ~w34924 & w35083 ;
  assign w35085 = w35082 | w35084 ;
  assign w35086 = ~\pi097 & w35085 ;
  assign w35087 = ~w34569 & w34839 ;
  assign w35088 = w34840 ^ w35087 ;
  assign w35089 = ~w34925 & w35088 ;
  assign w35090 = ( w34562 & w34923 ) | ( w34562 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35091 = ~w34924 & w35090 ;
  assign w35092 = w35089 | w35091 ;
  assign w35093 = ~\pi096 & w35092 ;
  assign w35094 = ~w34575 & w34836 ;
  assign w35095 = w34837 ^ w35094 ;
  assign w35096 = ~w34925 & w35095 ;
  assign w35097 = ( w34568 & w34923 ) | ( w34568 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35098 = ~w34924 & w35097 ;
  assign w35099 = w35096 | w35098 ;
  assign w35100 = ~\pi095 & w35099 ;
  assign w35101 = ~w34581 & w34833 ;
  assign w35102 = w34834 ^ w35101 ;
  assign w35103 = ~w34925 & w35102 ;
  assign w35104 = ( w34574 & w34923 ) | ( w34574 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35105 = ~w34924 & w35104 ;
  assign w35106 = w35103 | w35105 ;
  assign w35107 = ~\pi094 & w35106 ;
  assign w35108 = ~w34587 & w34830 ;
  assign w35109 = w34831 ^ w35108 ;
  assign w35110 = ~w34925 & w35109 ;
  assign w35111 = ( w34580 & w34923 ) | ( w34580 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35112 = ~w34924 & w35111 ;
  assign w35113 = w35110 | w35112 ;
  assign w35114 = ~\pi093 & w35113 ;
  assign w35115 = ~w34593 & w34827 ;
  assign w35116 = w34828 ^ w35115 ;
  assign w35117 = ~w34925 & w35116 ;
  assign w35118 = ( w34586 & w34923 ) | ( w34586 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35119 = ~w34924 & w35118 ;
  assign w35120 = w35117 | w35119 ;
  assign w35121 = ~\pi092 & w35120 ;
  assign w35122 = ~w34599 & w34824 ;
  assign w35123 = w34825 ^ w35122 ;
  assign w35124 = ~w34925 & w35123 ;
  assign w35125 = ( w34592 & w34923 ) | ( w34592 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35126 = ~w34924 & w35125 ;
  assign w35127 = w35124 | w35126 ;
  assign w35128 = ~\pi091 & w35127 ;
  assign w35129 = ~w34605 & w34821 ;
  assign w35130 = w34822 ^ w35129 ;
  assign w35131 = ~w34925 & w35130 ;
  assign w35132 = ( w34598 & w34923 ) | ( w34598 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35133 = ~w34924 & w35132 ;
  assign w35134 = w35131 | w35133 ;
  assign w35135 = ~\pi090 & w35134 ;
  assign w35136 = ~w34611 & w34818 ;
  assign w35137 = w34819 ^ w35136 ;
  assign w35138 = ~w34925 & w35137 ;
  assign w35139 = ( w34604 & w34923 ) | ( w34604 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35140 = ~w34924 & w35139 ;
  assign w35141 = w35138 | w35140 ;
  assign w35142 = ~\pi089 & w35141 ;
  assign w35143 = ~w34617 & w34815 ;
  assign w35144 = w34816 ^ w35143 ;
  assign w35145 = ~w34925 & w35144 ;
  assign w35146 = ( w34610 & w34923 ) | ( w34610 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35147 = ~w34924 & w35146 ;
  assign w35148 = w35145 | w35147 ;
  assign w35149 = ~\pi088 & w35148 ;
  assign w35150 = ~w34623 & w34812 ;
  assign w35151 = w34813 ^ w35150 ;
  assign w35152 = ~w34925 & w35151 ;
  assign w35153 = ( w34616 & w34923 ) | ( w34616 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35154 = ~w34924 & w35153 ;
  assign w35155 = w35152 | w35154 ;
  assign w35156 = ~\pi087 & w35155 ;
  assign w35157 = ~w34629 & w34809 ;
  assign w35158 = w34810 ^ w35157 ;
  assign w35159 = ~w34925 & w35158 ;
  assign w35160 = ( w34622 & w34923 ) | ( w34622 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35161 = ~w34924 & w35160 ;
  assign w35162 = w35159 | w35161 ;
  assign w35163 = ~\pi086 & w35162 ;
  assign w35164 = ~w34635 & w34806 ;
  assign w35165 = w34807 ^ w35164 ;
  assign w35166 = ~w34925 & w35165 ;
  assign w35167 = ( w34628 & w34923 ) | ( w34628 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35168 = ~w34924 & w35167 ;
  assign w35169 = w35166 | w35168 ;
  assign w35170 = ~\pi085 & w35169 ;
  assign w35171 = ~w34641 & w34803 ;
  assign w35172 = w34804 ^ w35171 ;
  assign w35173 = ~w34925 & w35172 ;
  assign w35174 = ( w34634 & w34923 ) | ( w34634 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35175 = ~w34924 & w35174 ;
  assign w35176 = w35173 | w35175 ;
  assign w35177 = ~\pi084 & w35176 ;
  assign w35178 = ~w34647 & w34800 ;
  assign w35179 = w34801 ^ w35178 ;
  assign w35180 = ~w34925 & w35179 ;
  assign w35181 = ( w34640 & w34923 ) | ( w34640 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35182 = ~w34924 & w35181 ;
  assign w35183 = w35180 | w35182 ;
  assign w35184 = ~\pi083 & w35183 ;
  assign w35185 = ~w34653 & w34797 ;
  assign w35186 = w34798 ^ w35185 ;
  assign w35187 = ~w34925 & w35186 ;
  assign w35188 = ( w34646 & w34923 ) | ( w34646 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35189 = ~w34924 & w35188 ;
  assign w35190 = w35187 | w35189 ;
  assign w35191 = ~\pi082 & w35190 ;
  assign w35192 = ~w34659 & w34794 ;
  assign w35193 = w34795 ^ w35192 ;
  assign w35194 = ~w34925 & w35193 ;
  assign w35195 = ( w34652 & w34923 ) | ( w34652 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35196 = ~w34924 & w35195 ;
  assign w35197 = w35194 | w35196 ;
  assign w35198 = ~\pi081 & w35197 ;
  assign w35199 = ~w34665 & w34791 ;
  assign w35200 = w34792 ^ w35199 ;
  assign w35201 = ~w34925 & w35200 ;
  assign w35202 = ( w34658 & w34923 ) | ( w34658 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35203 = ~w34924 & w35202 ;
  assign w35204 = w35201 | w35203 ;
  assign w35205 = ~\pi080 & w35204 ;
  assign w35206 = ~w34671 & w34788 ;
  assign w35207 = w34789 ^ w35206 ;
  assign w35208 = ~w34925 & w35207 ;
  assign w35209 = ( w34664 & w34923 ) | ( w34664 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35210 = ~w34924 & w35209 ;
  assign w35211 = w35208 | w35210 ;
  assign w35212 = ~\pi079 & w35211 ;
  assign w35213 = ~w34677 & w34785 ;
  assign w35214 = w34786 ^ w35213 ;
  assign w35215 = ~w34925 & w35214 ;
  assign w35216 = ( w34670 & w34923 ) | ( w34670 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35217 = ~w34924 & w35216 ;
  assign w35218 = w35215 | w35217 ;
  assign w35219 = ~\pi078 & w35218 ;
  assign w35220 = ~w34683 & w34782 ;
  assign w35221 = w34783 ^ w35220 ;
  assign w35222 = ~w34925 & w35221 ;
  assign w35223 = ( w34676 & w34923 ) | ( w34676 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35224 = ~w34924 & w35223 ;
  assign w35225 = w35222 | w35224 ;
  assign w35226 = ~\pi077 & w35225 ;
  assign w35227 = ~w34689 & w34779 ;
  assign w35228 = w34780 ^ w35227 ;
  assign w35229 = ~w34925 & w35228 ;
  assign w35230 = ( w34682 & w34923 ) | ( w34682 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35231 = ~w34924 & w35230 ;
  assign w35232 = w35229 | w35231 ;
  assign w35233 = ~\pi076 & w35232 ;
  assign w35234 = ~w34695 & w34776 ;
  assign w35235 = w34777 ^ w35234 ;
  assign w35236 = ~w34925 & w35235 ;
  assign w35237 = ( w34688 & w34923 ) | ( w34688 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35238 = ~w34924 & w35237 ;
  assign w35239 = w35236 | w35238 ;
  assign w35240 = ~\pi075 & w35239 ;
  assign w35241 = ~w34701 & w34773 ;
  assign w35242 = w34774 ^ w35241 ;
  assign w35243 = ~w34925 & w35242 ;
  assign w35244 = ( w34694 & w34923 ) | ( w34694 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35245 = ~w34924 & w35244 ;
  assign w35246 = w35243 | w35245 ;
  assign w35247 = ~\pi074 & w35246 ;
  assign w35248 = ~w34707 & w34770 ;
  assign w35249 = w34771 ^ w35248 ;
  assign w35250 = ~w34925 & w35249 ;
  assign w35251 = ( w34700 & w34923 ) | ( w34700 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35252 = ~w34924 & w35251 ;
  assign w35253 = w35250 | w35252 ;
  assign w35254 = ~\pi073 & w35253 ;
  assign w35255 = ~w34713 & w34767 ;
  assign w35256 = w34768 ^ w35255 ;
  assign w35257 = ~w34925 & w35256 ;
  assign w35258 = ( w34706 & w34923 ) | ( w34706 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35259 = ~w34924 & w35258 ;
  assign w35260 = w35257 | w35259 ;
  assign w35261 = ~\pi072 & w35260 ;
  assign w35262 = ~w34719 & w34764 ;
  assign w35263 = w34765 ^ w35262 ;
  assign w35264 = ~w34925 & w35263 ;
  assign w35265 = ( w34712 & w34923 ) | ( w34712 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35266 = ~w34924 & w35265 ;
  assign w35267 = w35264 | w35266 ;
  assign w35268 = ~\pi071 & w35267 ;
  assign w35269 = ~w34725 & w34761 ;
  assign w35270 = w34762 ^ w35269 ;
  assign w35271 = ~w34925 & w35270 ;
  assign w35272 = ( w34718 & w34923 ) | ( w34718 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35273 = ~w34924 & w35272 ;
  assign w35274 = w35271 | w35273 ;
  assign w35275 = ~\pi070 & w35274 ;
  assign w35276 = ~w34734 & w34758 ;
  assign w35277 = w34759 ^ w35276 ;
  assign w35278 = ~w34925 & w35277 ;
  assign w35279 = ( w34724 & w34923 ) | ( w34724 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35280 = ~w34924 & w35279 ;
  assign w35281 = w35278 | w35280 ;
  assign w35282 = ~\pi069 & w35281 ;
  assign w35283 = ~w34744 & w34753 ;
  assign w35284 = w34756 ^ w35283 ;
  assign w35285 = ~w34925 & w35284 ;
  assign w35286 = ( w34733 & w34923 ) | ( w34733 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35287 = ~w34924 & w35286 ;
  assign w35288 = w35285 | w35287 ;
  assign w35289 = ~\pi068 & w35288 ;
  assign w35290 = w34750 ^ w34752 ;
  assign w35291 = ~w34925 & w35290 ;
  assign w35292 = ( w34743 & w34923 ) | ( w34743 & w34924 ) | ( w34923 & w34924 ) ;
  assign w35293 = ~w34924 & w35292 ;
  assign w35294 = w35291 | w35293 ;
  assign w35295 = ~\pi067 & w35294 ;
  assign w35296 = w15400 ^ w34751 ;
  assign w35297 = \pi065 ^ w35296 ;
  assign w35298 = ~w34925 & w35297 ;
  assign w35299 = ( w34746 & w34747 ) | ( w34746 & ~w34924 ) | ( w34747 & ~w34924 ) ;
  assign w35300 = w34924 & w35299 ;
  assign w35301 = ( ~w34923 & w35299 ) | ( ~w34923 & w35300 ) | ( w35299 & w35300 ) ;
  assign w35302 = ( w35298 & w35299 ) | ( w35298 & ~w35301 ) | ( w35299 & ~w35301 ) ;
  assign w35303 = ~\pi066 & w35302 ;
  assign w35304 = w34923 | w34924 ;
  assign w35305 = ( w35298 & w35299 ) | ( w35298 & w35304 ) | ( w35299 & w35304 ) ;
  assign w35306 = ( ~w34924 & w35298 ) | ( ~w34924 & w35305 ) | ( w35298 & w35305 ) ;
  assign w35307 = \pi066 ^ w35306 ;
  assign w35308 = ( \pi064 & ~w34925 ) | ( \pi064 & w35307 ) | ( ~w34925 & w35307 ) ;
  assign w35309 = \pi008 ^ w35308 ;
  assign w35310 = ( \pi065 & w16517 ) | ( \pi065 & ~w35309 ) | ( w16517 & ~w35309 ) ;
  assign w35311 = w35307 | w35310 ;
  assign w35312 = \pi067 ^ w35294 ;
  assign w35313 = ( ~w35303 & w35311 ) | ( ~w35303 & w35312 ) | ( w35311 & w35312 ) ;
  assign w35314 = w35312 | w35313 ;
  assign w35315 = \pi068 ^ w35288 ;
  assign w35316 = ( ~w35295 & w35314 ) | ( ~w35295 & w35315 ) | ( w35314 & w35315 ) ;
  assign w35317 = w35315 | w35316 ;
  assign w35318 = \pi069 ^ w35281 ;
  assign w35319 = ( ~w35289 & w35317 ) | ( ~w35289 & w35318 ) | ( w35317 & w35318 ) ;
  assign w35320 = w35318 | w35319 ;
  assign w35321 = \pi070 ^ w35274 ;
  assign w35322 = ( ~w35282 & w35320 ) | ( ~w35282 & w35321 ) | ( w35320 & w35321 ) ;
  assign w35323 = w35321 | w35322 ;
  assign w35324 = \pi071 ^ w35267 ;
  assign w35325 = ( ~w35275 & w35323 ) | ( ~w35275 & w35324 ) | ( w35323 & w35324 ) ;
  assign w35326 = w35324 | w35325 ;
  assign w35327 = \pi072 ^ w35260 ;
  assign w35328 = ( ~w35268 & w35326 ) | ( ~w35268 & w35327 ) | ( w35326 & w35327 ) ;
  assign w35329 = w35327 | w35328 ;
  assign w35330 = \pi073 ^ w35253 ;
  assign w35331 = ( ~w35261 & w35329 ) | ( ~w35261 & w35330 ) | ( w35329 & w35330 ) ;
  assign w35332 = w35330 | w35331 ;
  assign w35333 = \pi074 ^ w35246 ;
  assign w35334 = ( ~w35254 & w35332 ) | ( ~w35254 & w35333 ) | ( w35332 & w35333 ) ;
  assign w35335 = w35333 | w35334 ;
  assign w35336 = \pi075 ^ w35239 ;
  assign w35337 = ( ~w35247 & w35335 ) | ( ~w35247 & w35336 ) | ( w35335 & w35336 ) ;
  assign w35338 = w35336 | w35337 ;
  assign w35339 = \pi076 ^ w35232 ;
  assign w35340 = ( ~w35240 & w35338 ) | ( ~w35240 & w35339 ) | ( w35338 & w35339 ) ;
  assign w35341 = w35339 | w35340 ;
  assign w35342 = \pi077 ^ w35225 ;
  assign w35343 = ( ~w35233 & w35341 ) | ( ~w35233 & w35342 ) | ( w35341 & w35342 ) ;
  assign w35344 = w35342 | w35343 ;
  assign w35345 = \pi078 ^ w35218 ;
  assign w35346 = ( ~w35226 & w35344 ) | ( ~w35226 & w35345 ) | ( w35344 & w35345 ) ;
  assign w35347 = w35345 | w35346 ;
  assign w35348 = \pi079 ^ w35211 ;
  assign w35349 = ( ~w35219 & w35347 ) | ( ~w35219 & w35348 ) | ( w35347 & w35348 ) ;
  assign w35350 = w35348 | w35349 ;
  assign w35351 = \pi080 ^ w35204 ;
  assign w35352 = ( ~w35212 & w35350 ) | ( ~w35212 & w35351 ) | ( w35350 & w35351 ) ;
  assign w35353 = w35351 | w35352 ;
  assign w35354 = \pi081 ^ w35197 ;
  assign w35355 = ( ~w35205 & w35353 ) | ( ~w35205 & w35354 ) | ( w35353 & w35354 ) ;
  assign w35356 = w35354 | w35355 ;
  assign w35357 = \pi082 ^ w35190 ;
  assign w35358 = ( ~w35198 & w35356 ) | ( ~w35198 & w35357 ) | ( w35356 & w35357 ) ;
  assign w35359 = w35357 | w35358 ;
  assign w35360 = \pi083 ^ w35183 ;
  assign w35361 = ( ~w35191 & w35359 ) | ( ~w35191 & w35360 ) | ( w35359 & w35360 ) ;
  assign w35362 = w35360 | w35361 ;
  assign w35363 = \pi084 ^ w35176 ;
  assign w35364 = ( ~w35184 & w35362 ) | ( ~w35184 & w35363 ) | ( w35362 & w35363 ) ;
  assign w35365 = w35363 | w35364 ;
  assign w35366 = \pi085 ^ w35169 ;
  assign w35367 = ( ~w35177 & w35365 ) | ( ~w35177 & w35366 ) | ( w35365 & w35366 ) ;
  assign w35368 = w35366 | w35367 ;
  assign w35369 = \pi086 ^ w35162 ;
  assign w35370 = ( ~w35170 & w35368 ) | ( ~w35170 & w35369 ) | ( w35368 & w35369 ) ;
  assign w35371 = w35369 | w35370 ;
  assign w35372 = \pi087 ^ w35155 ;
  assign w35373 = ( ~w35163 & w35371 ) | ( ~w35163 & w35372 ) | ( w35371 & w35372 ) ;
  assign w35374 = w35372 | w35373 ;
  assign w35375 = \pi088 ^ w35148 ;
  assign w35376 = ( ~w35156 & w35374 ) | ( ~w35156 & w35375 ) | ( w35374 & w35375 ) ;
  assign w35377 = w35375 | w35376 ;
  assign w35378 = \pi089 ^ w35141 ;
  assign w35379 = ( ~w35149 & w35377 ) | ( ~w35149 & w35378 ) | ( w35377 & w35378 ) ;
  assign w35380 = w35378 | w35379 ;
  assign w35381 = \pi090 ^ w35134 ;
  assign w35382 = ( ~w35142 & w35380 ) | ( ~w35142 & w35381 ) | ( w35380 & w35381 ) ;
  assign w35383 = w35381 | w35382 ;
  assign w35384 = \pi091 ^ w35127 ;
  assign w35385 = ( ~w35135 & w35383 ) | ( ~w35135 & w35384 ) | ( w35383 & w35384 ) ;
  assign w35386 = w35384 | w35385 ;
  assign w35387 = \pi092 ^ w35120 ;
  assign w35388 = ( ~w35128 & w35386 ) | ( ~w35128 & w35387 ) | ( w35386 & w35387 ) ;
  assign w35389 = w35387 | w35388 ;
  assign w35390 = \pi093 ^ w35113 ;
  assign w35391 = ( ~w35121 & w35389 ) | ( ~w35121 & w35390 ) | ( w35389 & w35390 ) ;
  assign w35392 = w35390 | w35391 ;
  assign w35393 = \pi094 ^ w35106 ;
  assign w35394 = ( ~w35114 & w35392 ) | ( ~w35114 & w35393 ) | ( w35392 & w35393 ) ;
  assign w35395 = w35393 | w35394 ;
  assign w35396 = \pi095 ^ w35099 ;
  assign w35397 = ( ~w35107 & w35395 ) | ( ~w35107 & w35396 ) | ( w35395 & w35396 ) ;
  assign w35398 = w35396 | w35397 ;
  assign w35399 = \pi096 ^ w35092 ;
  assign w35400 = ( ~w35100 & w35398 ) | ( ~w35100 & w35399 ) | ( w35398 & w35399 ) ;
  assign w35401 = w35399 | w35400 ;
  assign w35402 = \pi097 ^ w35085 ;
  assign w35403 = ( ~w35093 & w35401 ) | ( ~w35093 & w35402 ) | ( w35401 & w35402 ) ;
  assign w35404 = w35402 | w35403 ;
  assign w35405 = \pi098 ^ w35078 ;
  assign w35406 = ( ~w35086 & w35404 ) | ( ~w35086 & w35405 ) | ( w35404 & w35405 ) ;
  assign w35407 = w35405 | w35406 ;
  assign w35408 = \pi099 ^ w35071 ;
  assign w35409 = ( ~w35079 & w35407 ) | ( ~w35079 & w35408 ) | ( w35407 & w35408 ) ;
  assign w35410 = w35408 | w35409 ;
  assign w35411 = \pi100 ^ w35064 ;
  assign w35412 = ( ~w35072 & w35410 ) | ( ~w35072 & w35411 ) | ( w35410 & w35411 ) ;
  assign w35413 = w35411 | w35412 ;
  assign w35414 = \pi101 ^ w35057 ;
  assign w35415 = ( ~w35065 & w35413 ) | ( ~w35065 & w35414 ) | ( w35413 & w35414 ) ;
  assign w35416 = w35414 | w35415 ;
  assign w35417 = \pi102 ^ w35050 ;
  assign w35418 = ( ~w35058 & w35416 ) | ( ~w35058 & w35417 ) | ( w35416 & w35417 ) ;
  assign w35419 = w35417 | w35418 ;
  assign w35420 = \pi103 ^ w35043 ;
  assign w35421 = ( ~w35051 & w35419 ) | ( ~w35051 & w35420 ) | ( w35419 & w35420 ) ;
  assign w35422 = w35420 | w35421 ;
  assign w35423 = \pi104 ^ w35036 ;
  assign w35424 = ( ~w35044 & w35422 ) | ( ~w35044 & w35423 ) | ( w35422 & w35423 ) ;
  assign w35425 = w35423 | w35424 ;
  assign w35426 = \pi105 ^ w35029 ;
  assign w35427 = ( ~w35037 & w35425 ) | ( ~w35037 & w35426 ) | ( w35425 & w35426 ) ;
  assign w35428 = w35426 | w35427 ;
  assign w35429 = \pi106 ^ w35022 ;
  assign w35430 = ( ~w35030 & w35428 ) | ( ~w35030 & w35429 ) | ( w35428 & w35429 ) ;
  assign w35431 = w35429 | w35430 ;
  assign w35432 = \pi107 ^ w35015 ;
  assign w35433 = ( ~w35023 & w35431 ) | ( ~w35023 & w35432 ) | ( w35431 & w35432 ) ;
  assign w35434 = w35432 | w35433 ;
  assign w35435 = \pi108 ^ w35008 ;
  assign w35436 = ( ~w35016 & w35434 ) | ( ~w35016 & w35435 ) | ( w35434 & w35435 ) ;
  assign w35437 = w35435 | w35436 ;
  assign w35438 = \pi109 ^ w35001 ;
  assign w35439 = ( ~w35009 & w35437 ) | ( ~w35009 & w35438 ) | ( w35437 & w35438 ) ;
  assign w35440 = w35438 | w35439 ;
  assign w35441 = \pi110 ^ w34994 ;
  assign w35442 = ( ~w35002 & w35440 ) | ( ~w35002 & w35441 ) | ( w35440 & w35441 ) ;
  assign w35443 = w35441 | w35442 ;
  assign w35444 = \pi111 ^ w34987 ;
  assign w35445 = ( ~w34995 & w35443 ) | ( ~w34995 & w35444 ) | ( w35443 & w35444 ) ;
  assign w35446 = w35444 | w35445 ;
  assign w35447 = \pi112 ^ w34980 ;
  assign w35448 = ( ~w34988 & w35446 ) | ( ~w34988 & w35447 ) | ( w35446 & w35447 ) ;
  assign w35449 = w35447 | w35448 ;
  assign w35450 = \pi113 ^ w34973 ;
  assign w35451 = ( ~w34981 & w35449 ) | ( ~w34981 & w35450 ) | ( w35449 & w35450 ) ;
  assign w35452 = w35450 | w35451 ;
  assign w35453 = \pi114 ^ w34966 ;
  assign w35454 = ( ~w34974 & w35452 ) | ( ~w34974 & w35453 ) | ( w35452 & w35453 ) ;
  assign w35455 = w35453 | w35454 ;
  assign w35456 = \pi115 ^ w34959 ;
  assign w35457 = ( ~w34967 & w35455 ) | ( ~w34967 & w35456 ) | ( w35455 & w35456 ) ;
  assign w35458 = w35456 | w35457 ;
  assign w35459 = \pi116 ^ w34952 ;
  assign w35460 = ( ~w34960 & w35458 ) | ( ~w34960 & w35459 ) | ( w35458 & w35459 ) ;
  assign w35461 = w35459 | w35460 ;
  assign w35462 = \pi117 ^ w34945 ;
  assign w35463 = ( ~w34953 & w35461 ) | ( ~w34953 & w35462 ) | ( w35461 & w35462 ) ;
  assign w35464 = w35462 | w35463 ;
  assign w35465 = \pi118 ^ w34938 ;
  assign w35466 = ( ~w34946 & w35464 ) | ( ~w34946 & w35465 ) | ( w35464 & w35465 ) ;
  assign w35467 = w35465 | w35466 ;
  assign w35468 = \pi119 ^ w34931 ;
  assign w35469 = ( ~w34939 & w35467 ) | ( ~w34939 & w35468 ) | ( w35467 & w35468 ) ;
  assign w35470 = w35468 | w35469 ;
  assign w35471 = ( ~w34425 & w34911 ) | ( ~w34425 & w34925 ) | ( w34911 & w34925 ) ;
  assign w35472 = w34920 ^ w35471 ;
  assign w35473 = ~w34925 & w35472 ;
  assign w35474 = ( w15063 & ~w34916 ) | ( w15063 & w34923 ) | ( ~w34916 & w34923 ) ;
  assign w35475 = w34916 & w35474 ;
  assign w35476 = w35473 | w35475 ;
  assign w35477 = ~\pi120 & w35476 ;
  assign w35478 = ( \pi120 & ~w35473 ) | ( \pi120 & w35475 ) | ( ~w35473 & w35475 ) ;
  assign w35479 = ~w35475 & w35478 ;
  assign w35480 = w35477 | w35479 ;
  assign w35481 = ( ~w34932 & w35470 ) | ( ~w34932 & w35480 ) | ( w35470 & w35480 ) ;
  assign w35482 = ( w273 & ~w35480 ) | ( w273 & w35481 ) | ( ~w35480 & w35481 ) ;
  assign w35483 = w35480 | w35482 ;
  assign w35484 = ~w199 & w35476 ;
  assign w35485 = w35483 & ~w35484 ;
  assign w35486 = ~w34939 & w35467 ;
  assign w35487 = w35468 ^ w35486 ;
  assign w35488 = ~w35485 & w35487 ;
  assign w35489 = ( w34931 & w35483 ) | ( w34931 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35490 = ~w35484 & w35489 ;
  assign w35491 = w35488 | w35490 ;
  assign w35492 = ( ~w34932 & w35470 ) | ( ~w34932 & w35485 ) | ( w35470 & w35485 ) ;
  assign w35493 = w35480 ^ w35492 ;
  assign w35494 = ~w35485 & w35493 ;
  assign w35495 = ( w199 & ~w35476 ) | ( w199 & w35483 ) | ( ~w35476 & w35483 ) ;
  assign w35496 = w35476 & w35495 ;
  assign w35497 = w35494 | w35496 ;
  assign w35498 = ~\pi120 & w35491 ;
  assign w35499 = ~w34946 & w35464 ;
  assign w35500 = w35465 ^ w35499 ;
  assign w35501 = ~w35485 & w35500 ;
  assign w35502 = ( w34938 & w35483 ) | ( w34938 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35503 = ~w35484 & w35502 ;
  assign w35504 = w35501 | w35503 ;
  assign w35505 = ~\pi119 & w35504 ;
  assign w35506 = ~w34953 & w35461 ;
  assign w35507 = w35462 ^ w35506 ;
  assign w35508 = ~w35485 & w35507 ;
  assign w35509 = ( w34945 & w35483 ) | ( w34945 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35510 = ~w35484 & w35509 ;
  assign w35511 = w35508 | w35510 ;
  assign w35512 = ~\pi118 & w35511 ;
  assign w35513 = ~w34960 & w35458 ;
  assign w35514 = w35459 ^ w35513 ;
  assign w35515 = ~w35485 & w35514 ;
  assign w35516 = ( w34952 & w35483 ) | ( w34952 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35517 = ~w35484 & w35516 ;
  assign w35518 = w35515 | w35517 ;
  assign w35519 = ~\pi117 & w35518 ;
  assign w35520 = ~w34967 & w35455 ;
  assign w35521 = w35456 ^ w35520 ;
  assign w35522 = ~w35485 & w35521 ;
  assign w35523 = ( w34959 & w35483 ) | ( w34959 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35524 = ~w35484 & w35523 ;
  assign w35525 = w35522 | w35524 ;
  assign w35526 = ~\pi116 & w35525 ;
  assign w35527 = ~w34974 & w35452 ;
  assign w35528 = w35453 ^ w35527 ;
  assign w35529 = ~w35485 & w35528 ;
  assign w35530 = ( w34966 & w35483 ) | ( w34966 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35531 = ~w35484 & w35530 ;
  assign w35532 = w35529 | w35531 ;
  assign w35533 = ~\pi115 & w35532 ;
  assign w35534 = ~w34981 & w35449 ;
  assign w35535 = w35450 ^ w35534 ;
  assign w35536 = ~w35485 & w35535 ;
  assign w35537 = ( w34973 & w35483 ) | ( w34973 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35538 = ~w35484 & w35537 ;
  assign w35539 = w35536 | w35538 ;
  assign w35540 = ~\pi114 & w35539 ;
  assign w35541 = ~w34988 & w35446 ;
  assign w35542 = w35447 ^ w35541 ;
  assign w35543 = ~w35485 & w35542 ;
  assign w35544 = ( w34980 & w35483 ) | ( w34980 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35545 = ~w35484 & w35544 ;
  assign w35546 = w35543 | w35545 ;
  assign w35547 = ~\pi113 & w35546 ;
  assign w35548 = ~w34995 & w35443 ;
  assign w35549 = w35444 ^ w35548 ;
  assign w35550 = ~w35485 & w35549 ;
  assign w35551 = ( w34987 & w35483 ) | ( w34987 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35552 = ~w35484 & w35551 ;
  assign w35553 = w35550 | w35552 ;
  assign w35554 = ~\pi112 & w35553 ;
  assign w35555 = ~w35002 & w35440 ;
  assign w35556 = w35441 ^ w35555 ;
  assign w35557 = ~w35485 & w35556 ;
  assign w35558 = ( w34994 & w35483 ) | ( w34994 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35559 = ~w35484 & w35558 ;
  assign w35560 = w35557 | w35559 ;
  assign w35561 = ~\pi111 & w35560 ;
  assign w35562 = ~w35009 & w35437 ;
  assign w35563 = w35438 ^ w35562 ;
  assign w35564 = ~w35485 & w35563 ;
  assign w35565 = ( w35001 & w35483 ) | ( w35001 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35566 = ~w35484 & w35565 ;
  assign w35567 = w35564 | w35566 ;
  assign w35568 = ~\pi110 & w35567 ;
  assign w35569 = ~w35016 & w35434 ;
  assign w35570 = w35435 ^ w35569 ;
  assign w35571 = ~w35485 & w35570 ;
  assign w35572 = ( w35008 & w35483 ) | ( w35008 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35573 = ~w35484 & w35572 ;
  assign w35574 = w35571 | w35573 ;
  assign w35575 = ~\pi109 & w35574 ;
  assign w35576 = ~w35023 & w35431 ;
  assign w35577 = w35432 ^ w35576 ;
  assign w35578 = ~w35485 & w35577 ;
  assign w35579 = ( w35015 & w35483 ) | ( w35015 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35580 = ~w35484 & w35579 ;
  assign w35581 = w35578 | w35580 ;
  assign w35582 = ~\pi108 & w35581 ;
  assign w35583 = ~w35030 & w35428 ;
  assign w35584 = w35429 ^ w35583 ;
  assign w35585 = ~w35485 & w35584 ;
  assign w35586 = ( w35022 & w35483 ) | ( w35022 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35587 = ~w35484 & w35586 ;
  assign w35588 = w35585 | w35587 ;
  assign w35589 = ~\pi107 & w35588 ;
  assign w35590 = ~w35037 & w35425 ;
  assign w35591 = w35426 ^ w35590 ;
  assign w35592 = ~w35485 & w35591 ;
  assign w35593 = ( w35029 & w35483 ) | ( w35029 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35594 = ~w35484 & w35593 ;
  assign w35595 = w35592 | w35594 ;
  assign w35596 = ~\pi106 & w35595 ;
  assign w35597 = ~w35044 & w35422 ;
  assign w35598 = w35423 ^ w35597 ;
  assign w35599 = ~w35485 & w35598 ;
  assign w35600 = ( w35036 & w35483 ) | ( w35036 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35601 = ~w35484 & w35600 ;
  assign w35602 = w35599 | w35601 ;
  assign w35603 = ~\pi105 & w35602 ;
  assign w35604 = ~w35051 & w35419 ;
  assign w35605 = w35420 ^ w35604 ;
  assign w35606 = ~w35485 & w35605 ;
  assign w35607 = ( w35043 & w35483 ) | ( w35043 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35608 = ~w35484 & w35607 ;
  assign w35609 = w35606 | w35608 ;
  assign w35610 = ~\pi104 & w35609 ;
  assign w35611 = ~w35058 & w35416 ;
  assign w35612 = w35417 ^ w35611 ;
  assign w35613 = ~w35485 & w35612 ;
  assign w35614 = ( w35050 & w35483 ) | ( w35050 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35615 = ~w35484 & w35614 ;
  assign w35616 = w35613 | w35615 ;
  assign w35617 = ~\pi103 & w35616 ;
  assign w35618 = ~w35065 & w35413 ;
  assign w35619 = w35414 ^ w35618 ;
  assign w35620 = ~w35485 & w35619 ;
  assign w35621 = ( w35057 & w35483 ) | ( w35057 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35622 = ~w35484 & w35621 ;
  assign w35623 = w35620 | w35622 ;
  assign w35624 = ~\pi102 & w35623 ;
  assign w35625 = ~w35072 & w35410 ;
  assign w35626 = w35411 ^ w35625 ;
  assign w35627 = ~w35485 & w35626 ;
  assign w35628 = ( w35064 & w35483 ) | ( w35064 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35629 = ~w35484 & w35628 ;
  assign w35630 = w35627 | w35629 ;
  assign w35631 = ~\pi101 & w35630 ;
  assign w35632 = ~w35079 & w35407 ;
  assign w35633 = w35408 ^ w35632 ;
  assign w35634 = ~w35485 & w35633 ;
  assign w35635 = ( w35071 & w35483 ) | ( w35071 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35636 = ~w35484 & w35635 ;
  assign w35637 = w35634 | w35636 ;
  assign w35638 = ~\pi100 & w35637 ;
  assign w35639 = ~w35086 & w35404 ;
  assign w35640 = w35405 ^ w35639 ;
  assign w35641 = ~w35485 & w35640 ;
  assign w35642 = ( w35078 & w35483 ) | ( w35078 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35643 = ~w35484 & w35642 ;
  assign w35644 = w35641 | w35643 ;
  assign w35645 = ~\pi099 & w35644 ;
  assign w35646 = ~w35093 & w35401 ;
  assign w35647 = w35402 ^ w35646 ;
  assign w35648 = ~w35485 & w35647 ;
  assign w35649 = ( w35085 & w35483 ) | ( w35085 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35650 = ~w35484 & w35649 ;
  assign w35651 = w35648 | w35650 ;
  assign w35652 = ~\pi098 & w35651 ;
  assign w35653 = ~w35100 & w35398 ;
  assign w35654 = w35399 ^ w35653 ;
  assign w35655 = ~w35485 & w35654 ;
  assign w35656 = ( w35092 & w35483 ) | ( w35092 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35657 = ~w35484 & w35656 ;
  assign w35658 = w35655 | w35657 ;
  assign w35659 = ~\pi097 & w35658 ;
  assign w35660 = ~w35107 & w35395 ;
  assign w35661 = w35396 ^ w35660 ;
  assign w35662 = ~w35485 & w35661 ;
  assign w35663 = ( w35099 & w35483 ) | ( w35099 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35664 = ~w35484 & w35663 ;
  assign w35665 = w35662 | w35664 ;
  assign w35666 = ~\pi096 & w35665 ;
  assign w35667 = ~w35114 & w35392 ;
  assign w35668 = w35393 ^ w35667 ;
  assign w35669 = ~w35485 & w35668 ;
  assign w35670 = ( w35106 & w35483 ) | ( w35106 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35671 = ~w35484 & w35670 ;
  assign w35672 = w35669 | w35671 ;
  assign w35673 = ~\pi095 & w35672 ;
  assign w35674 = ~w35121 & w35389 ;
  assign w35675 = w35390 ^ w35674 ;
  assign w35676 = ~w35485 & w35675 ;
  assign w35677 = ( w35113 & w35483 ) | ( w35113 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35678 = ~w35484 & w35677 ;
  assign w35679 = w35676 | w35678 ;
  assign w35680 = ~\pi094 & w35679 ;
  assign w35681 = ~w35128 & w35386 ;
  assign w35682 = w35387 ^ w35681 ;
  assign w35683 = ~w35485 & w35682 ;
  assign w35684 = ( w35120 & w35483 ) | ( w35120 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35685 = ~w35484 & w35684 ;
  assign w35686 = w35683 | w35685 ;
  assign w35687 = ~\pi093 & w35686 ;
  assign w35688 = ~w35135 & w35383 ;
  assign w35689 = w35384 ^ w35688 ;
  assign w35690 = ~w35485 & w35689 ;
  assign w35691 = ( w35127 & w35483 ) | ( w35127 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35692 = ~w35484 & w35691 ;
  assign w35693 = w35690 | w35692 ;
  assign w35694 = ~\pi092 & w35693 ;
  assign w35695 = ~w35142 & w35380 ;
  assign w35696 = w35381 ^ w35695 ;
  assign w35697 = ~w35485 & w35696 ;
  assign w35698 = ( w35134 & w35483 ) | ( w35134 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35699 = ~w35484 & w35698 ;
  assign w35700 = w35697 | w35699 ;
  assign w35701 = ~\pi091 & w35700 ;
  assign w35702 = ~w35149 & w35377 ;
  assign w35703 = w35378 ^ w35702 ;
  assign w35704 = ~w35485 & w35703 ;
  assign w35705 = ( w35141 & w35483 ) | ( w35141 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35706 = ~w35484 & w35705 ;
  assign w35707 = w35704 | w35706 ;
  assign w35708 = ~\pi090 & w35707 ;
  assign w35709 = ~w35156 & w35374 ;
  assign w35710 = w35375 ^ w35709 ;
  assign w35711 = ~w35485 & w35710 ;
  assign w35712 = ( w35148 & w35483 ) | ( w35148 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35713 = ~w35484 & w35712 ;
  assign w35714 = w35711 | w35713 ;
  assign w35715 = ~\pi089 & w35714 ;
  assign w35716 = ~w35163 & w35371 ;
  assign w35717 = w35372 ^ w35716 ;
  assign w35718 = ~w35485 & w35717 ;
  assign w35719 = ( w35155 & w35483 ) | ( w35155 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35720 = ~w35484 & w35719 ;
  assign w35721 = w35718 | w35720 ;
  assign w35722 = ~\pi088 & w35721 ;
  assign w35723 = ~w35170 & w35368 ;
  assign w35724 = w35369 ^ w35723 ;
  assign w35725 = ~w35485 & w35724 ;
  assign w35726 = ( w35162 & w35483 ) | ( w35162 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35727 = ~w35484 & w35726 ;
  assign w35728 = w35725 | w35727 ;
  assign w35729 = ~\pi087 & w35728 ;
  assign w35730 = ~w35177 & w35365 ;
  assign w35731 = w35366 ^ w35730 ;
  assign w35732 = ~w35485 & w35731 ;
  assign w35733 = ( w35169 & w35483 ) | ( w35169 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35734 = ~w35484 & w35733 ;
  assign w35735 = w35732 | w35734 ;
  assign w35736 = ~\pi086 & w35735 ;
  assign w35737 = ~w35184 & w35362 ;
  assign w35738 = w35363 ^ w35737 ;
  assign w35739 = ~w35485 & w35738 ;
  assign w35740 = ( w35176 & w35483 ) | ( w35176 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35741 = ~w35484 & w35740 ;
  assign w35742 = w35739 | w35741 ;
  assign w35743 = ~\pi085 & w35742 ;
  assign w35744 = ~w35191 & w35359 ;
  assign w35745 = w35360 ^ w35744 ;
  assign w35746 = ~w35485 & w35745 ;
  assign w35747 = ( w35183 & w35483 ) | ( w35183 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35748 = ~w35484 & w35747 ;
  assign w35749 = w35746 | w35748 ;
  assign w35750 = ~\pi084 & w35749 ;
  assign w35751 = ~w35198 & w35356 ;
  assign w35752 = w35357 ^ w35751 ;
  assign w35753 = ~w35485 & w35752 ;
  assign w35754 = ( w35190 & w35483 ) | ( w35190 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35755 = ~w35484 & w35754 ;
  assign w35756 = w35753 | w35755 ;
  assign w35757 = ~\pi083 & w35756 ;
  assign w35758 = ~w35205 & w35353 ;
  assign w35759 = w35354 ^ w35758 ;
  assign w35760 = ~w35485 & w35759 ;
  assign w35761 = ( w35197 & w35483 ) | ( w35197 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35762 = ~w35484 & w35761 ;
  assign w35763 = w35760 | w35762 ;
  assign w35764 = ~\pi082 & w35763 ;
  assign w35765 = ~w35212 & w35350 ;
  assign w35766 = w35351 ^ w35765 ;
  assign w35767 = ~w35485 & w35766 ;
  assign w35768 = ( w35204 & w35483 ) | ( w35204 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35769 = ~w35484 & w35768 ;
  assign w35770 = w35767 | w35769 ;
  assign w35771 = ~\pi081 & w35770 ;
  assign w35772 = ~w35219 & w35347 ;
  assign w35773 = w35348 ^ w35772 ;
  assign w35774 = ~w35485 & w35773 ;
  assign w35775 = ( w35211 & w35483 ) | ( w35211 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35776 = ~w35484 & w35775 ;
  assign w35777 = w35774 | w35776 ;
  assign w35778 = ~\pi080 & w35777 ;
  assign w35779 = ~w35226 & w35344 ;
  assign w35780 = w35345 ^ w35779 ;
  assign w35781 = ~w35485 & w35780 ;
  assign w35782 = ( w35218 & w35483 ) | ( w35218 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35783 = ~w35484 & w35782 ;
  assign w35784 = w35781 | w35783 ;
  assign w35785 = ~\pi079 & w35784 ;
  assign w35786 = ~w35233 & w35341 ;
  assign w35787 = w35342 ^ w35786 ;
  assign w35788 = ~w35485 & w35787 ;
  assign w35789 = ( w35225 & w35483 ) | ( w35225 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35790 = ~w35484 & w35789 ;
  assign w35791 = w35788 | w35790 ;
  assign w35792 = ~\pi078 & w35791 ;
  assign w35793 = ~w35240 & w35338 ;
  assign w35794 = w35339 ^ w35793 ;
  assign w35795 = ~w35485 & w35794 ;
  assign w35796 = ( w35232 & w35483 ) | ( w35232 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35797 = ~w35484 & w35796 ;
  assign w35798 = w35795 | w35797 ;
  assign w35799 = ~\pi077 & w35798 ;
  assign w35800 = ~w35247 & w35335 ;
  assign w35801 = w35336 ^ w35800 ;
  assign w35802 = ~w35485 & w35801 ;
  assign w35803 = ( w35239 & w35483 ) | ( w35239 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35804 = ~w35484 & w35803 ;
  assign w35805 = w35802 | w35804 ;
  assign w35806 = ~\pi076 & w35805 ;
  assign w35807 = ~w35254 & w35332 ;
  assign w35808 = w35333 ^ w35807 ;
  assign w35809 = ~w35485 & w35808 ;
  assign w35810 = ( w35246 & w35483 ) | ( w35246 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35811 = ~w35484 & w35810 ;
  assign w35812 = w35809 | w35811 ;
  assign w35813 = ~\pi075 & w35812 ;
  assign w35814 = ~w35261 & w35329 ;
  assign w35815 = w35330 ^ w35814 ;
  assign w35816 = ~w35485 & w35815 ;
  assign w35817 = ( w35253 & w35483 ) | ( w35253 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35818 = ~w35484 & w35817 ;
  assign w35819 = w35816 | w35818 ;
  assign w35820 = ~\pi074 & w35819 ;
  assign w35821 = ~w35268 & w35326 ;
  assign w35822 = w35327 ^ w35821 ;
  assign w35823 = ~w35485 & w35822 ;
  assign w35824 = ( w35260 & w35483 ) | ( w35260 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35825 = ~w35484 & w35824 ;
  assign w35826 = w35823 | w35825 ;
  assign w35827 = ~\pi073 & w35826 ;
  assign w35828 = ~w35275 & w35323 ;
  assign w35829 = w35324 ^ w35828 ;
  assign w35830 = ~w35485 & w35829 ;
  assign w35831 = ( w35267 & w35483 ) | ( w35267 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35832 = ~w35484 & w35831 ;
  assign w35833 = w35830 | w35832 ;
  assign w35834 = ~\pi072 & w35833 ;
  assign w35835 = ~w35282 & w35320 ;
  assign w35836 = w35321 ^ w35835 ;
  assign w35837 = ~w35485 & w35836 ;
  assign w35838 = ( w35274 & w35483 ) | ( w35274 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35839 = ~w35484 & w35838 ;
  assign w35840 = w35837 | w35839 ;
  assign w35841 = ~\pi071 & w35840 ;
  assign w35842 = ~w35289 & w35317 ;
  assign w35843 = w35318 ^ w35842 ;
  assign w35844 = ~w35485 & w35843 ;
  assign w35845 = ( w35281 & w35483 ) | ( w35281 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35846 = ~w35484 & w35845 ;
  assign w35847 = w35844 | w35846 ;
  assign w35848 = ~\pi070 & w35847 ;
  assign w35849 = ~w35295 & w35314 ;
  assign w35850 = w35315 ^ w35849 ;
  assign w35851 = ~w35485 & w35850 ;
  assign w35852 = ( w35288 & w35483 ) | ( w35288 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35853 = ~w35484 & w35852 ;
  assign w35854 = w35851 | w35853 ;
  assign w35855 = ~\pi069 & w35854 ;
  assign w35856 = ~w35303 & w35311 ;
  assign w35857 = w35312 ^ w35856 ;
  assign w35858 = ~w35485 & w35857 ;
  assign w35859 = ( w35294 & w35483 ) | ( w35294 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35860 = ~w35484 & w35859 ;
  assign w35861 = w35858 | w35860 ;
  assign w35862 = ~\pi068 & w35861 ;
  assign w35863 = \pi064 & ~w34925 ;
  assign w35864 = \pi008 ^ w35863 ;
  assign w35865 = ( \pi065 & w16517 ) | ( \pi065 & ~w35864 ) | ( w16517 & ~w35864 ) ;
  assign w35866 = w35307 ^ w35865 ;
  assign w35867 = ~w35485 & w35866 ;
  assign w35868 = ( w35302 & w35483 ) | ( w35302 & w35484 ) | ( w35483 & w35484 ) ;
  assign w35869 = ~w35484 & w35868 ;
  assign w35870 = w35867 | w35869 ;
  assign w35871 = ~\pi067 & w35870 ;
  assign w35872 = \pi007 ^ w34925 ;
  assign w35873 = ( \pi064 & w35485 ) | ( \pi064 & w35872 ) | ( w35485 & w35872 ) ;
  assign w35874 = w16525 ^ w35873 ;
  assign w35875 = ~w35485 & w35874 ;
  assign w35876 = w35485 & w35864 ;
  assign w35877 = w35875 | w35876 ;
  assign w35878 = ~\pi066 & w35877 ;
  assign w35879 = \pi066 ^ w35877 ;
  assign w35880 = ( \pi064 & ~w35485 ) | ( \pi064 & w35879 ) | ( ~w35485 & w35879 ) ;
  assign w35881 = \pi007 ^ w35880 ;
  assign w35882 = ( \pi065 & w17033 ) | ( \pi065 & ~w35881 ) | ( w17033 & ~w35881 ) ;
  assign w35883 = w35879 | w35882 ;
  assign w35884 = \pi067 ^ w35870 ;
  assign w35885 = ( ~w35878 & w35883 ) | ( ~w35878 & w35884 ) | ( w35883 & w35884 ) ;
  assign w35886 = w35884 | w35885 ;
  assign w35887 = \pi068 ^ w35861 ;
  assign w35888 = ( ~w35871 & w35886 ) | ( ~w35871 & w35887 ) | ( w35886 & w35887 ) ;
  assign w35889 = w35887 | w35888 ;
  assign w35890 = \pi069 ^ w35854 ;
  assign w35891 = ( ~w35862 & w35889 ) | ( ~w35862 & w35890 ) | ( w35889 & w35890 ) ;
  assign w35892 = w35890 | w35891 ;
  assign w35893 = \pi070 ^ w35847 ;
  assign w35894 = ( ~w35855 & w35892 ) | ( ~w35855 & w35893 ) | ( w35892 & w35893 ) ;
  assign w35895 = w35893 | w35894 ;
  assign w35896 = \pi071 ^ w35840 ;
  assign w35897 = ( ~w35848 & w35895 ) | ( ~w35848 & w35896 ) | ( w35895 & w35896 ) ;
  assign w35898 = w35896 | w35897 ;
  assign w35899 = \pi072 ^ w35833 ;
  assign w35900 = ( ~w35841 & w35898 ) | ( ~w35841 & w35899 ) | ( w35898 & w35899 ) ;
  assign w35901 = w35899 | w35900 ;
  assign w35902 = \pi073 ^ w35826 ;
  assign w35903 = ( ~w35834 & w35901 ) | ( ~w35834 & w35902 ) | ( w35901 & w35902 ) ;
  assign w35904 = w35902 | w35903 ;
  assign w35905 = \pi074 ^ w35819 ;
  assign w35906 = ( ~w35827 & w35904 ) | ( ~w35827 & w35905 ) | ( w35904 & w35905 ) ;
  assign w35907 = w35905 | w35906 ;
  assign w35908 = \pi075 ^ w35812 ;
  assign w35909 = ( ~w35820 & w35907 ) | ( ~w35820 & w35908 ) | ( w35907 & w35908 ) ;
  assign w35910 = w35908 | w35909 ;
  assign w35911 = \pi076 ^ w35805 ;
  assign w35912 = ( ~w35813 & w35910 ) | ( ~w35813 & w35911 ) | ( w35910 & w35911 ) ;
  assign w35913 = w35911 | w35912 ;
  assign w35914 = \pi077 ^ w35798 ;
  assign w35915 = ( ~w35806 & w35913 ) | ( ~w35806 & w35914 ) | ( w35913 & w35914 ) ;
  assign w35916 = w35914 | w35915 ;
  assign w35917 = \pi078 ^ w35791 ;
  assign w35918 = ( ~w35799 & w35916 ) | ( ~w35799 & w35917 ) | ( w35916 & w35917 ) ;
  assign w35919 = w35917 | w35918 ;
  assign w35920 = \pi079 ^ w35784 ;
  assign w35921 = ( ~w35792 & w35919 ) | ( ~w35792 & w35920 ) | ( w35919 & w35920 ) ;
  assign w35922 = w35920 | w35921 ;
  assign w35923 = \pi080 ^ w35777 ;
  assign w35924 = ( ~w35785 & w35922 ) | ( ~w35785 & w35923 ) | ( w35922 & w35923 ) ;
  assign w35925 = w35923 | w35924 ;
  assign w35926 = \pi081 ^ w35770 ;
  assign w35927 = ( ~w35778 & w35925 ) | ( ~w35778 & w35926 ) | ( w35925 & w35926 ) ;
  assign w35928 = w35926 | w35927 ;
  assign w35929 = \pi082 ^ w35763 ;
  assign w35930 = ( ~w35771 & w35928 ) | ( ~w35771 & w35929 ) | ( w35928 & w35929 ) ;
  assign w35931 = w35929 | w35930 ;
  assign w35932 = \pi083 ^ w35756 ;
  assign w35933 = ( ~w35764 & w35931 ) | ( ~w35764 & w35932 ) | ( w35931 & w35932 ) ;
  assign w35934 = w35932 | w35933 ;
  assign w35935 = \pi084 ^ w35749 ;
  assign w35936 = ( ~w35757 & w35934 ) | ( ~w35757 & w35935 ) | ( w35934 & w35935 ) ;
  assign w35937 = w35935 | w35936 ;
  assign w35938 = \pi085 ^ w35742 ;
  assign w35939 = ( ~w35750 & w35937 ) | ( ~w35750 & w35938 ) | ( w35937 & w35938 ) ;
  assign w35940 = w35938 | w35939 ;
  assign w35941 = \pi086 ^ w35735 ;
  assign w35942 = ( ~w35743 & w35940 ) | ( ~w35743 & w35941 ) | ( w35940 & w35941 ) ;
  assign w35943 = w35941 | w35942 ;
  assign w35944 = \pi087 ^ w35728 ;
  assign w35945 = ( ~w35736 & w35943 ) | ( ~w35736 & w35944 ) | ( w35943 & w35944 ) ;
  assign w35946 = w35944 | w35945 ;
  assign w35947 = \pi088 ^ w35721 ;
  assign w35948 = ( ~w35729 & w35946 ) | ( ~w35729 & w35947 ) | ( w35946 & w35947 ) ;
  assign w35949 = w35947 | w35948 ;
  assign w35950 = \pi089 ^ w35714 ;
  assign w35951 = ( ~w35722 & w35949 ) | ( ~w35722 & w35950 ) | ( w35949 & w35950 ) ;
  assign w35952 = w35950 | w35951 ;
  assign w35953 = \pi090 ^ w35707 ;
  assign w35954 = ( ~w35715 & w35952 ) | ( ~w35715 & w35953 ) | ( w35952 & w35953 ) ;
  assign w35955 = w35953 | w35954 ;
  assign w35956 = \pi091 ^ w35700 ;
  assign w35957 = ( ~w35708 & w35955 ) | ( ~w35708 & w35956 ) | ( w35955 & w35956 ) ;
  assign w35958 = w35956 | w35957 ;
  assign w35959 = \pi092 ^ w35693 ;
  assign w35960 = ( ~w35701 & w35958 ) | ( ~w35701 & w35959 ) | ( w35958 & w35959 ) ;
  assign w35961 = w35959 | w35960 ;
  assign w35962 = \pi093 ^ w35686 ;
  assign w35963 = ( ~w35694 & w35961 ) | ( ~w35694 & w35962 ) | ( w35961 & w35962 ) ;
  assign w35964 = w35962 | w35963 ;
  assign w35965 = \pi094 ^ w35679 ;
  assign w35966 = ( ~w35687 & w35964 ) | ( ~w35687 & w35965 ) | ( w35964 & w35965 ) ;
  assign w35967 = w35965 | w35966 ;
  assign w35968 = \pi095 ^ w35672 ;
  assign w35969 = ( ~w35680 & w35967 ) | ( ~w35680 & w35968 ) | ( w35967 & w35968 ) ;
  assign w35970 = w35968 | w35969 ;
  assign w35971 = \pi096 ^ w35665 ;
  assign w35972 = ( ~w35673 & w35970 ) | ( ~w35673 & w35971 ) | ( w35970 & w35971 ) ;
  assign w35973 = w35971 | w35972 ;
  assign w35974 = \pi097 ^ w35658 ;
  assign w35975 = ( ~w35666 & w35973 ) | ( ~w35666 & w35974 ) | ( w35973 & w35974 ) ;
  assign w35976 = w35974 | w35975 ;
  assign w35977 = \pi098 ^ w35651 ;
  assign w35978 = ( ~w35659 & w35976 ) | ( ~w35659 & w35977 ) | ( w35976 & w35977 ) ;
  assign w35979 = w35977 | w35978 ;
  assign w35980 = \pi099 ^ w35644 ;
  assign w35981 = ( ~w35652 & w35979 ) | ( ~w35652 & w35980 ) | ( w35979 & w35980 ) ;
  assign w35982 = w35980 | w35981 ;
  assign w35983 = \pi100 ^ w35637 ;
  assign w35984 = ( ~w35645 & w35982 ) | ( ~w35645 & w35983 ) | ( w35982 & w35983 ) ;
  assign w35985 = w35983 | w35984 ;
  assign w35986 = \pi101 ^ w35630 ;
  assign w35987 = ( ~w35638 & w35985 ) | ( ~w35638 & w35986 ) | ( w35985 & w35986 ) ;
  assign w35988 = w35986 | w35987 ;
  assign w35989 = \pi102 ^ w35623 ;
  assign w35990 = ( ~w35631 & w35988 ) | ( ~w35631 & w35989 ) | ( w35988 & w35989 ) ;
  assign w35991 = w35989 | w35990 ;
  assign w35992 = \pi103 ^ w35616 ;
  assign w35993 = ( ~w35624 & w35991 ) | ( ~w35624 & w35992 ) | ( w35991 & w35992 ) ;
  assign w35994 = w35992 | w35993 ;
  assign w35995 = \pi104 ^ w35609 ;
  assign w35996 = ( ~w35617 & w35994 ) | ( ~w35617 & w35995 ) | ( w35994 & w35995 ) ;
  assign w35997 = w35995 | w35996 ;
  assign w35998 = \pi105 ^ w35602 ;
  assign w35999 = ( ~w35610 & w35997 ) | ( ~w35610 & w35998 ) | ( w35997 & w35998 ) ;
  assign w36000 = w35998 | w35999 ;
  assign w36001 = \pi106 ^ w35595 ;
  assign w36002 = ( ~w35603 & w36000 ) | ( ~w35603 & w36001 ) | ( w36000 & w36001 ) ;
  assign w36003 = w36001 | w36002 ;
  assign w36004 = \pi107 ^ w35588 ;
  assign w36005 = ( ~w35596 & w36003 ) | ( ~w35596 & w36004 ) | ( w36003 & w36004 ) ;
  assign w36006 = w36004 | w36005 ;
  assign w36007 = \pi108 ^ w35581 ;
  assign w36008 = ( ~w35589 & w36006 ) | ( ~w35589 & w36007 ) | ( w36006 & w36007 ) ;
  assign w36009 = w36007 | w36008 ;
  assign w36010 = \pi109 ^ w35574 ;
  assign w36011 = ( ~w35582 & w36009 ) | ( ~w35582 & w36010 ) | ( w36009 & w36010 ) ;
  assign w36012 = w36010 | w36011 ;
  assign w36013 = \pi110 ^ w35567 ;
  assign w36014 = ( ~w35575 & w36012 ) | ( ~w35575 & w36013 ) | ( w36012 & w36013 ) ;
  assign w36015 = w36013 | w36014 ;
  assign w36016 = \pi111 ^ w35560 ;
  assign w36017 = ( ~w35568 & w36015 ) | ( ~w35568 & w36016 ) | ( w36015 & w36016 ) ;
  assign w36018 = w36016 | w36017 ;
  assign w36019 = \pi112 ^ w35553 ;
  assign w36020 = ( ~w35561 & w36018 ) | ( ~w35561 & w36019 ) | ( w36018 & w36019 ) ;
  assign w36021 = w36019 | w36020 ;
  assign w36022 = \pi113 ^ w35546 ;
  assign w36023 = ( ~w35554 & w36021 ) | ( ~w35554 & w36022 ) | ( w36021 & w36022 ) ;
  assign w36024 = w36022 | w36023 ;
  assign w36025 = \pi114 ^ w35539 ;
  assign w36026 = ( ~w35547 & w36024 ) | ( ~w35547 & w36025 ) | ( w36024 & w36025 ) ;
  assign w36027 = w36025 | w36026 ;
  assign w36028 = \pi115 ^ w35532 ;
  assign w36029 = ( ~w35540 & w36027 ) | ( ~w35540 & w36028 ) | ( w36027 & w36028 ) ;
  assign w36030 = w36028 | w36029 ;
  assign w36031 = \pi116 ^ w35525 ;
  assign w36032 = ( ~w35533 & w36030 ) | ( ~w35533 & w36031 ) | ( w36030 & w36031 ) ;
  assign w36033 = w36031 | w36032 ;
  assign w36034 = \pi117 ^ w35518 ;
  assign w36035 = ( ~w35526 & w36033 ) | ( ~w35526 & w36034 ) | ( w36033 & w36034 ) ;
  assign w36036 = w36034 | w36035 ;
  assign w36037 = \pi118 ^ w35511 ;
  assign w36038 = ( ~w35519 & w36036 ) | ( ~w35519 & w36037 ) | ( w36036 & w36037 ) ;
  assign w36039 = w36037 | w36038 ;
  assign w36040 = \pi119 ^ w35504 ;
  assign w36041 = ( ~w35512 & w36039 ) | ( ~w35512 & w36040 ) | ( w36039 & w36040 ) ;
  assign w36042 = w36040 | w36041 ;
  assign w36043 = \pi120 ^ w35491 ;
  assign w36044 = ( ~w35505 & w36042 ) | ( ~w35505 & w36043 ) | ( w36042 & w36043 ) ;
  assign w36045 = w36043 | w36044 ;
  assign w36046 = \pi121 ^ w35497 ;
  assign w36047 = w35498 & ~w36046 ;
  assign w36048 = ( w36045 & w36046 ) | ( w36045 & ~w36047 ) | ( w36046 & ~w36047 ) ;
  assign w36049 = ~\pi121 & w35497 ;
  assign w36050 = w36048 & ~w36049 ;
  assign w36051 = w16707 | w36050 ;
  assign w36052 = w35491 & w36051 ;
  assign w36053 = ~w35505 & w36042 ;
  assign w36054 = w36043 ^ w36053 ;
  assign w36055 = ~w36051 & w36054 ;
  assign w36056 = w36052 | w36055 ;
  assign w36057 = ~\pi121 & w36056 ;
  assign w36058 = w35504 & w36051 ;
  assign w36059 = ~w35512 & w36039 ;
  assign w36060 = w36040 ^ w36059 ;
  assign w36061 = ~w36051 & w36060 ;
  assign w36062 = w36058 | w36061 ;
  assign w36063 = ~\pi120 & w36062 ;
  assign w36064 = w35511 & w36051 ;
  assign w36065 = ~w35519 & w36036 ;
  assign w36066 = w36037 ^ w36065 ;
  assign w36067 = ~w36051 & w36066 ;
  assign w36068 = w36064 | w36067 ;
  assign w36069 = ~\pi119 & w36068 ;
  assign w36070 = w35518 & w36051 ;
  assign w36071 = ~w35526 & w36033 ;
  assign w36072 = w36034 ^ w36071 ;
  assign w36073 = ~w36051 & w36072 ;
  assign w36074 = w36070 | w36073 ;
  assign w36075 = ~\pi118 & w36074 ;
  assign w36076 = w35525 & w36051 ;
  assign w36077 = ~w35533 & w36030 ;
  assign w36078 = w36031 ^ w36077 ;
  assign w36079 = ~w36051 & w36078 ;
  assign w36080 = w36076 | w36079 ;
  assign w36081 = ~\pi117 & w36080 ;
  assign w36082 = w35532 & w36051 ;
  assign w36083 = ~w35540 & w36027 ;
  assign w36084 = w36028 ^ w36083 ;
  assign w36085 = ~w36051 & w36084 ;
  assign w36086 = w36082 | w36085 ;
  assign w36087 = ~\pi116 & w36086 ;
  assign w36088 = w35539 & w36051 ;
  assign w36089 = ~w35547 & w36024 ;
  assign w36090 = w36025 ^ w36089 ;
  assign w36091 = ~w36051 & w36090 ;
  assign w36092 = w36088 | w36091 ;
  assign w36093 = ~\pi115 & w36092 ;
  assign w36094 = w35546 & w36051 ;
  assign w36095 = ~w35554 & w36021 ;
  assign w36096 = w36022 ^ w36095 ;
  assign w36097 = ~w36051 & w36096 ;
  assign w36098 = w36094 | w36097 ;
  assign w36099 = ~\pi114 & w36098 ;
  assign w36100 = w35553 & w36051 ;
  assign w36101 = ~w35561 & w36018 ;
  assign w36102 = w36019 ^ w36101 ;
  assign w36103 = ~w36051 & w36102 ;
  assign w36104 = w36100 | w36103 ;
  assign w36105 = ~\pi113 & w36104 ;
  assign w36106 = w35560 & w36051 ;
  assign w36107 = ~w35568 & w36015 ;
  assign w36108 = w36016 ^ w36107 ;
  assign w36109 = ~w36051 & w36108 ;
  assign w36110 = w36106 | w36109 ;
  assign w36111 = ~\pi112 & w36110 ;
  assign w36112 = w35567 & w36051 ;
  assign w36113 = ~w35575 & w36012 ;
  assign w36114 = w36013 ^ w36113 ;
  assign w36115 = ~w36051 & w36114 ;
  assign w36116 = w36112 | w36115 ;
  assign w36117 = ~\pi111 & w36116 ;
  assign w36118 = w35574 & w36051 ;
  assign w36119 = ~w35582 & w36009 ;
  assign w36120 = w36010 ^ w36119 ;
  assign w36121 = ~w36051 & w36120 ;
  assign w36122 = w36118 | w36121 ;
  assign w36123 = ~\pi110 & w36122 ;
  assign w36124 = w35581 & w36051 ;
  assign w36125 = ~w35589 & w36006 ;
  assign w36126 = w36007 ^ w36125 ;
  assign w36127 = ~w36051 & w36126 ;
  assign w36128 = w36124 | w36127 ;
  assign w36129 = ~\pi109 & w36128 ;
  assign w36130 = w35588 & w36051 ;
  assign w36131 = ~w35596 & w36003 ;
  assign w36132 = w36004 ^ w36131 ;
  assign w36133 = ~w36051 & w36132 ;
  assign w36134 = w36130 | w36133 ;
  assign w36135 = ~\pi108 & w36134 ;
  assign w36136 = w35595 & w36051 ;
  assign w36137 = ~w35603 & w36000 ;
  assign w36138 = w36001 ^ w36137 ;
  assign w36139 = ~w36051 & w36138 ;
  assign w36140 = w36136 | w36139 ;
  assign w36141 = ~\pi107 & w36140 ;
  assign w36142 = w35602 & w36051 ;
  assign w36143 = ~w35610 & w35997 ;
  assign w36144 = w35998 ^ w36143 ;
  assign w36145 = ~w36051 & w36144 ;
  assign w36146 = w36142 | w36145 ;
  assign w36147 = ~\pi106 & w36146 ;
  assign w36148 = w35609 & w36051 ;
  assign w36149 = ~w35617 & w35994 ;
  assign w36150 = w35995 ^ w36149 ;
  assign w36151 = ~w36051 & w36150 ;
  assign w36152 = w36148 | w36151 ;
  assign w36153 = ~\pi105 & w36152 ;
  assign w36154 = w35616 & w36051 ;
  assign w36155 = ~w35624 & w35991 ;
  assign w36156 = w35992 ^ w36155 ;
  assign w36157 = ~w36051 & w36156 ;
  assign w36158 = w36154 | w36157 ;
  assign w36159 = ~\pi104 & w36158 ;
  assign w36160 = w35623 & w36051 ;
  assign w36161 = ~w35631 & w35988 ;
  assign w36162 = w35989 ^ w36161 ;
  assign w36163 = ~w36051 & w36162 ;
  assign w36164 = w36160 | w36163 ;
  assign w36165 = ~\pi103 & w36164 ;
  assign w36166 = w35630 & w36051 ;
  assign w36167 = ~w35638 & w35985 ;
  assign w36168 = w35986 ^ w36167 ;
  assign w36169 = ~w36051 & w36168 ;
  assign w36170 = w36166 | w36169 ;
  assign w36171 = ~\pi102 & w36170 ;
  assign w36172 = w35637 & w36051 ;
  assign w36173 = ~w35645 & w35982 ;
  assign w36174 = w35983 ^ w36173 ;
  assign w36175 = ~w36051 & w36174 ;
  assign w36176 = w36172 | w36175 ;
  assign w36177 = ~\pi101 & w36176 ;
  assign w36178 = w35644 & w36051 ;
  assign w36179 = ~w35652 & w35979 ;
  assign w36180 = w35980 ^ w36179 ;
  assign w36181 = ~w36051 & w36180 ;
  assign w36182 = w36178 | w36181 ;
  assign w36183 = ~\pi100 & w36182 ;
  assign w36184 = w35651 & w36051 ;
  assign w36185 = ~w35659 & w35976 ;
  assign w36186 = w35977 ^ w36185 ;
  assign w36187 = ~w36051 & w36186 ;
  assign w36188 = w36184 | w36187 ;
  assign w36189 = ~\pi099 & w36188 ;
  assign w36190 = w35658 & w36051 ;
  assign w36191 = ~w35666 & w35973 ;
  assign w36192 = w35974 ^ w36191 ;
  assign w36193 = ~w36051 & w36192 ;
  assign w36194 = w36190 | w36193 ;
  assign w36195 = ~\pi098 & w36194 ;
  assign w36196 = w35665 & w36051 ;
  assign w36197 = ~w35673 & w35970 ;
  assign w36198 = w35971 ^ w36197 ;
  assign w36199 = ~w36051 & w36198 ;
  assign w36200 = w36196 | w36199 ;
  assign w36201 = ~\pi097 & w36200 ;
  assign w36202 = w35672 & w36051 ;
  assign w36203 = ~w35680 & w35967 ;
  assign w36204 = w35968 ^ w36203 ;
  assign w36205 = ~w36051 & w36204 ;
  assign w36206 = w36202 | w36205 ;
  assign w36207 = ~\pi096 & w36206 ;
  assign w36208 = w35679 & w36051 ;
  assign w36209 = ~w35687 & w35964 ;
  assign w36210 = w35965 ^ w36209 ;
  assign w36211 = ~w36051 & w36210 ;
  assign w36212 = w36208 | w36211 ;
  assign w36213 = ~\pi095 & w36212 ;
  assign w36214 = w35686 & w36051 ;
  assign w36215 = ~w35694 & w35961 ;
  assign w36216 = w35962 ^ w36215 ;
  assign w36217 = ~w36051 & w36216 ;
  assign w36218 = w36214 | w36217 ;
  assign w36219 = ~\pi094 & w36218 ;
  assign w36220 = w35693 & w36051 ;
  assign w36221 = ~w35701 & w35958 ;
  assign w36222 = w35959 ^ w36221 ;
  assign w36223 = ~w36051 & w36222 ;
  assign w36224 = w36220 | w36223 ;
  assign w36225 = ~\pi093 & w36224 ;
  assign w36226 = w35700 & w36051 ;
  assign w36227 = ~w35708 & w35955 ;
  assign w36228 = w35956 ^ w36227 ;
  assign w36229 = ~w36051 & w36228 ;
  assign w36230 = w36226 | w36229 ;
  assign w36231 = ~\pi092 & w36230 ;
  assign w36232 = w35707 & w36051 ;
  assign w36233 = ~w35715 & w35952 ;
  assign w36234 = w35953 ^ w36233 ;
  assign w36235 = ~w36051 & w36234 ;
  assign w36236 = w36232 | w36235 ;
  assign w36237 = ~\pi091 & w36236 ;
  assign w36238 = w35714 & w36051 ;
  assign w36239 = ~w35722 & w35949 ;
  assign w36240 = w35950 ^ w36239 ;
  assign w36241 = ~w36051 & w36240 ;
  assign w36242 = w36238 | w36241 ;
  assign w36243 = ~\pi090 & w36242 ;
  assign w36244 = w35721 & w36051 ;
  assign w36245 = ~w35729 & w35946 ;
  assign w36246 = w35947 ^ w36245 ;
  assign w36247 = ~w36051 & w36246 ;
  assign w36248 = w36244 | w36247 ;
  assign w36249 = ~\pi089 & w36248 ;
  assign w36250 = w35728 & w36051 ;
  assign w36251 = ~w35736 & w35943 ;
  assign w36252 = w35944 ^ w36251 ;
  assign w36253 = ~w36051 & w36252 ;
  assign w36254 = w36250 | w36253 ;
  assign w36255 = ~\pi088 & w36254 ;
  assign w36256 = w35735 & w36051 ;
  assign w36257 = ~w35743 & w35940 ;
  assign w36258 = w35941 ^ w36257 ;
  assign w36259 = ~w36051 & w36258 ;
  assign w36260 = w36256 | w36259 ;
  assign w36261 = ~\pi087 & w36260 ;
  assign w36262 = w35742 & w36051 ;
  assign w36263 = ~w35750 & w35937 ;
  assign w36264 = w35938 ^ w36263 ;
  assign w36265 = ~w36051 & w36264 ;
  assign w36266 = w36262 | w36265 ;
  assign w36267 = ~\pi086 & w36266 ;
  assign w36268 = w35749 & w36051 ;
  assign w36269 = ~w35757 & w35934 ;
  assign w36270 = w35935 ^ w36269 ;
  assign w36271 = ~w36051 & w36270 ;
  assign w36272 = w36268 | w36271 ;
  assign w36273 = ~\pi085 & w36272 ;
  assign w36274 = w35756 & w36051 ;
  assign w36275 = ~w35764 & w35931 ;
  assign w36276 = w35932 ^ w36275 ;
  assign w36277 = ~w36051 & w36276 ;
  assign w36278 = w36274 | w36277 ;
  assign w36279 = ~\pi084 & w36278 ;
  assign w36280 = w35763 & w36051 ;
  assign w36281 = ~w35771 & w35928 ;
  assign w36282 = w35929 ^ w36281 ;
  assign w36283 = ~w36051 & w36282 ;
  assign w36284 = w36280 | w36283 ;
  assign w36285 = ~\pi083 & w36284 ;
  assign w36286 = w35770 & w36051 ;
  assign w36287 = ~w35778 & w35925 ;
  assign w36288 = w35926 ^ w36287 ;
  assign w36289 = ~w36051 & w36288 ;
  assign w36290 = w36286 | w36289 ;
  assign w36291 = ~\pi082 & w36290 ;
  assign w36292 = w35777 & w36051 ;
  assign w36293 = ~w35785 & w35922 ;
  assign w36294 = w35923 ^ w36293 ;
  assign w36295 = ~w36051 & w36294 ;
  assign w36296 = w36292 | w36295 ;
  assign w36297 = ~\pi081 & w36296 ;
  assign w36298 = w35784 & w36051 ;
  assign w36299 = ~w35792 & w35919 ;
  assign w36300 = w35920 ^ w36299 ;
  assign w36301 = ~w36051 & w36300 ;
  assign w36302 = w36298 | w36301 ;
  assign w36303 = ~\pi080 & w36302 ;
  assign w36304 = w35791 & w36051 ;
  assign w36305 = ~w35799 & w35916 ;
  assign w36306 = w35917 ^ w36305 ;
  assign w36307 = ~w36051 & w36306 ;
  assign w36308 = w36304 | w36307 ;
  assign w36309 = ~\pi079 & w36308 ;
  assign w36310 = w35798 & w36051 ;
  assign w36311 = ~w35806 & w35913 ;
  assign w36312 = w35914 ^ w36311 ;
  assign w36313 = ~w36051 & w36312 ;
  assign w36314 = w36310 | w36313 ;
  assign w36315 = ~\pi078 & w36314 ;
  assign w36316 = w35805 & w36051 ;
  assign w36317 = ~w35813 & w35910 ;
  assign w36318 = w35911 ^ w36317 ;
  assign w36319 = ~w36051 & w36318 ;
  assign w36320 = w36316 | w36319 ;
  assign w36321 = ~\pi077 & w36320 ;
  assign w36322 = w35812 & w36051 ;
  assign w36323 = ~w35820 & w35907 ;
  assign w36324 = w35908 ^ w36323 ;
  assign w36325 = ~w36051 & w36324 ;
  assign w36326 = w36322 | w36325 ;
  assign w36327 = ~\pi076 & w36326 ;
  assign w36328 = w35819 & w36051 ;
  assign w36329 = ~w35827 & w35904 ;
  assign w36330 = w35905 ^ w36329 ;
  assign w36331 = ~w36051 & w36330 ;
  assign w36332 = w36328 | w36331 ;
  assign w36333 = ~\pi075 & w36332 ;
  assign w36334 = w35826 & w36051 ;
  assign w36335 = ~w35834 & w35901 ;
  assign w36336 = w35902 ^ w36335 ;
  assign w36337 = ~w36051 & w36336 ;
  assign w36338 = w36334 | w36337 ;
  assign w36339 = ~\pi074 & w36338 ;
  assign w36340 = w35833 & w36051 ;
  assign w36341 = ~w35841 & w35898 ;
  assign w36342 = w35899 ^ w36341 ;
  assign w36343 = ~w36051 & w36342 ;
  assign w36344 = w36340 | w36343 ;
  assign w36345 = ~\pi073 & w36344 ;
  assign w36346 = w35840 & w36051 ;
  assign w36347 = ~w35848 & w35895 ;
  assign w36348 = w35896 ^ w36347 ;
  assign w36349 = ~w36051 & w36348 ;
  assign w36350 = w36346 | w36349 ;
  assign w36351 = ~\pi072 & w36350 ;
  assign w36352 = w35847 & w36051 ;
  assign w36353 = ~w35855 & w35892 ;
  assign w36354 = w35893 ^ w36353 ;
  assign w36355 = ~w36051 & w36354 ;
  assign w36356 = w36352 | w36355 ;
  assign w36357 = ~\pi071 & w36356 ;
  assign w36358 = w35854 & w36051 ;
  assign w36359 = ~w35862 & w35889 ;
  assign w36360 = w35890 ^ w36359 ;
  assign w36361 = ~w36051 & w36360 ;
  assign w36362 = w36358 | w36361 ;
  assign w36363 = ~\pi070 & w36362 ;
  assign w36364 = w35861 & w36051 ;
  assign w36365 = ~w35871 & w35886 ;
  assign w36366 = w35887 ^ w36365 ;
  assign w36367 = ~w36051 & w36366 ;
  assign w36368 = w36364 | w36367 ;
  assign w36369 = ~\pi069 & w36368 ;
  assign w36370 = w35870 & w36051 ;
  assign w36371 = ~w35878 & w35883 ;
  assign w36372 = w35884 ^ w36371 ;
  assign w36373 = ~w36051 & w36372 ;
  assign w36374 = w36370 | w36373 ;
  assign w36375 = ~\pi068 & w36374 ;
  assign w36376 = \pi064 & ~w35485 ;
  assign w36377 = \pi007 ^ w36376 ;
  assign w36378 = ( \pi065 & w17033 ) | ( \pi065 & ~w36377 ) | ( w17033 & ~w36377 ) ;
  assign w36379 = w35879 ^ w36378 ;
  assign w36380 = ( w16707 & w36050 ) | ( w16707 & w36379 ) | ( w36050 & w36379 ) ;
  assign w36381 = w36379 & ~w36380 ;
  assign w36382 = ( w35877 & w36051 ) | ( w35877 & w36381 ) | ( w36051 & w36381 ) ;
  assign w36383 = w36381 | w36382 ;
  assign w36384 = ~\pi067 & w36383 ;
  assign w36385 = \pi006 ^ w35485 ;
  assign w36386 = ( \pi064 & w16707 ) | ( \pi064 & w36385 ) | ( w16707 & w36385 ) ;
  assign w36387 = w17041 ^ w36386 ;
  assign w36388 = ~w16707 & w36387 ;
  assign w36389 = ~w36050 & w36388 ;
  assign w36390 = ( ~\pi064 & w35485 ) | ( ~\pi064 & w36051 ) | ( w35485 & w36051 ) ;
  assign w36391 = \pi007 ^ w36390 ;
  assign w36392 = w36051 & ~w36391 ;
  assign w36393 = w36389 | w36392 ;
  assign w36394 = ~\pi066 & w36393 ;
  assign w36395 = ( \pi064 & w17054 ) | ( \pi064 & w36050 ) | ( w17054 & w36050 ) ;
  assign w36396 = ( \pi006 & ~\pi064 ) | ( \pi006 & w36395 ) | ( ~\pi064 & w36395 ) ;
  assign w36397 = w147 | w36050 ;
  assign w36398 = w17059 | w36397 ;
  assign w36399 = w17057 & ~w36398 ;
  assign w36400 = w36051 | w36389 ;
  assign w36401 = ( w36377 & w36389 ) | ( w36377 & w36400 ) | ( w36389 & w36400 ) ;
  assign w36402 = \pi066 ^ w36401 ;
  assign w36403 = w36396 | w36399 ;
  assign w36404 = ( \pi065 & w17062 ) | ( \pi065 & ~w36403 ) | ( w17062 & ~w36403 ) ;
  assign w36405 = w36402 | w36404 ;
  assign w36406 = ~w35877 & w36051 ;
  assign w36407 = ( w36051 & w36381 ) | ( w36051 & ~w36406 ) | ( w36381 & ~w36406 ) ;
  assign w36408 = \pi067 ^ w36407 ;
  assign w36409 = ( ~w36394 & w36405 ) | ( ~w36394 & w36408 ) | ( w36405 & w36408 ) ;
  assign w36410 = w36408 | w36409 ;
  assign w36411 = \pi068 ^ w36374 ;
  assign w36412 = ( ~w36384 & w36410 ) | ( ~w36384 & w36411 ) | ( w36410 & w36411 ) ;
  assign w36413 = w36411 | w36412 ;
  assign w36414 = \pi069 ^ w36368 ;
  assign w36415 = ( ~w36375 & w36413 ) | ( ~w36375 & w36414 ) | ( w36413 & w36414 ) ;
  assign w36416 = w36414 | w36415 ;
  assign w36417 = \pi070 ^ w36362 ;
  assign w36418 = ( ~w36369 & w36416 ) | ( ~w36369 & w36417 ) | ( w36416 & w36417 ) ;
  assign w36419 = w36417 | w36418 ;
  assign w36420 = \pi071 ^ w36356 ;
  assign w36421 = ( ~w36363 & w36419 ) | ( ~w36363 & w36420 ) | ( w36419 & w36420 ) ;
  assign w36422 = w36420 | w36421 ;
  assign w36423 = \pi072 ^ w36350 ;
  assign w36424 = ( ~w36357 & w36422 ) | ( ~w36357 & w36423 ) | ( w36422 & w36423 ) ;
  assign w36425 = w36423 | w36424 ;
  assign w36426 = \pi073 ^ w36344 ;
  assign w36427 = ( ~w36351 & w36425 ) | ( ~w36351 & w36426 ) | ( w36425 & w36426 ) ;
  assign w36428 = w36426 | w36427 ;
  assign w36429 = \pi074 ^ w36338 ;
  assign w36430 = ( ~w36345 & w36428 ) | ( ~w36345 & w36429 ) | ( w36428 & w36429 ) ;
  assign w36431 = w36429 | w36430 ;
  assign w36432 = \pi075 ^ w36332 ;
  assign w36433 = ( ~w36339 & w36431 ) | ( ~w36339 & w36432 ) | ( w36431 & w36432 ) ;
  assign w36434 = w36432 | w36433 ;
  assign w36435 = \pi076 ^ w36326 ;
  assign w36436 = ( ~w36333 & w36434 ) | ( ~w36333 & w36435 ) | ( w36434 & w36435 ) ;
  assign w36437 = w36435 | w36436 ;
  assign w36438 = \pi077 ^ w36320 ;
  assign w36439 = ( ~w36327 & w36437 ) | ( ~w36327 & w36438 ) | ( w36437 & w36438 ) ;
  assign w36440 = w36438 | w36439 ;
  assign w36441 = \pi078 ^ w36314 ;
  assign w36442 = ( ~w36321 & w36440 ) | ( ~w36321 & w36441 ) | ( w36440 & w36441 ) ;
  assign w36443 = w36441 | w36442 ;
  assign w36444 = \pi079 ^ w36308 ;
  assign w36445 = ( ~w36315 & w36443 ) | ( ~w36315 & w36444 ) | ( w36443 & w36444 ) ;
  assign w36446 = w36444 | w36445 ;
  assign w36447 = \pi080 ^ w36302 ;
  assign w36448 = ( ~w36309 & w36446 ) | ( ~w36309 & w36447 ) | ( w36446 & w36447 ) ;
  assign w36449 = w36447 | w36448 ;
  assign w36450 = \pi081 ^ w36296 ;
  assign w36451 = ( ~w36303 & w36449 ) | ( ~w36303 & w36450 ) | ( w36449 & w36450 ) ;
  assign w36452 = w36450 | w36451 ;
  assign w36453 = \pi082 ^ w36290 ;
  assign w36454 = ( ~w36297 & w36452 ) | ( ~w36297 & w36453 ) | ( w36452 & w36453 ) ;
  assign w36455 = w36453 | w36454 ;
  assign w36456 = \pi083 ^ w36284 ;
  assign w36457 = ( ~w36291 & w36455 ) | ( ~w36291 & w36456 ) | ( w36455 & w36456 ) ;
  assign w36458 = w36456 | w36457 ;
  assign w36459 = \pi084 ^ w36278 ;
  assign w36460 = ( ~w36285 & w36458 ) | ( ~w36285 & w36459 ) | ( w36458 & w36459 ) ;
  assign w36461 = w36459 | w36460 ;
  assign w36462 = \pi085 ^ w36272 ;
  assign w36463 = ( ~w36279 & w36461 ) | ( ~w36279 & w36462 ) | ( w36461 & w36462 ) ;
  assign w36464 = w36462 | w36463 ;
  assign w36465 = \pi086 ^ w36266 ;
  assign w36466 = ( ~w36273 & w36464 ) | ( ~w36273 & w36465 ) | ( w36464 & w36465 ) ;
  assign w36467 = w36465 | w36466 ;
  assign w36468 = \pi087 ^ w36260 ;
  assign w36469 = ( ~w36267 & w36467 ) | ( ~w36267 & w36468 ) | ( w36467 & w36468 ) ;
  assign w36470 = w36468 | w36469 ;
  assign w36471 = \pi088 ^ w36254 ;
  assign w36472 = ( ~w36261 & w36470 ) | ( ~w36261 & w36471 ) | ( w36470 & w36471 ) ;
  assign w36473 = w36471 | w36472 ;
  assign w36474 = \pi089 ^ w36248 ;
  assign w36475 = ( ~w36255 & w36473 ) | ( ~w36255 & w36474 ) | ( w36473 & w36474 ) ;
  assign w36476 = w36474 | w36475 ;
  assign w36477 = \pi090 ^ w36242 ;
  assign w36478 = ( ~w36249 & w36476 ) | ( ~w36249 & w36477 ) | ( w36476 & w36477 ) ;
  assign w36479 = w36477 | w36478 ;
  assign w36480 = \pi091 ^ w36236 ;
  assign w36481 = ( ~w36243 & w36479 ) | ( ~w36243 & w36480 ) | ( w36479 & w36480 ) ;
  assign w36482 = w36480 | w36481 ;
  assign w36483 = \pi092 ^ w36230 ;
  assign w36484 = ( ~w36237 & w36482 ) | ( ~w36237 & w36483 ) | ( w36482 & w36483 ) ;
  assign w36485 = w36483 | w36484 ;
  assign w36486 = \pi093 ^ w36224 ;
  assign w36487 = ( ~w36231 & w36485 ) | ( ~w36231 & w36486 ) | ( w36485 & w36486 ) ;
  assign w36488 = w36486 | w36487 ;
  assign w36489 = \pi094 ^ w36218 ;
  assign w36490 = ( ~w36225 & w36488 ) | ( ~w36225 & w36489 ) | ( w36488 & w36489 ) ;
  assign w36491 = w36489 | w36490 ;
  assign w36492 = \pi095 ^ w36212 ;
  assign w36493 = ( ~w36219 & w36491 ) | ( ~w36219 & w36492 ) | ( w36491 & w36492 ) ;
  assign w36494 = w36492 | w36493 ;
  assign w36495 = \pi096 ^ w36206 ;
  assign w36496 = ( ~w36213 & w36494 ) | ( ~w36213 & w36495 ) | ( w36494 & w36495 ) ;
  assign w36497 = w36495 | w36496 ;
  assign w36498 = \pi097 ^ w36200 ;
  assign w36499 = ( ~w36207 & w36497 ) | ( ~w36207 & w36498 ) | ( w36497 & w36498 ) ;
  assign w36500 = w36498 | w36499 ;
  assign w36501 = \pi098 ^ w36194 ;
  assign w36502 = ( ~w36201 & w36500 ) | ( ~w36201 & w36501 ) | ( w36500 & w36501 ) ;
  assign w36503 = w36501 | w36502 ;
  assign w36504 = \pi099 ^ w36188 ;
  assign w36505 = ( ~w36195 & w36503 ) | ( ~w36195 & w36504 ) | ( w36503 & w36504 ) ;
  assign w36506 = w36504 | w36505 ;
  assign w36507 = \pi100 ^ w36182 ;
  assign w36508 = ( ~w36189 & w36506 ) | ( ~w36189 & w36507 ) | ( w36506 & w36507 ) ;
  assign w36509 = w36507 | w36508 ;
  assign w36510 = \pi101 ^ w36176 ;
  assign w36511 = ( ~w36183 & w36509 ) | ( ~w36183 & w36510 ) | ( w36509 & w36510 ) ;
  assign w36512 = w36510 | w36511 ;
  assign w36513 = \pi102 ^ w36170 ;
  assign w36514 = ( ~w36177 & w36512 ) | ( ~w36177 & w36513 ) | ( w36512 & w36513 ) ;
  assign w36515 = w36513 | w36514 ;
  assign w36516 = \pi103 ^ w36164 ;
  assign w36517 = ( ~w36171 & w36515 ) | ( ~w36171 & w36516 ) | ( w36515 & w36516 ) ;
  assign w36518 = w36516 | w36517 ;
  assign w36519 = \pi104 ^ w36158 ;
  assign w36520 = ( ~w36165 & w36518 ) | ( ~w36165 & w36519 ) | ( w36518 & w36519 ) ;
  assign w36521 = w36519 | w36520 ;
  assign w36522 = \pi105 ^ w36152 ;
  assign w36523 = ( ~w36159 & w36521 ) | ( ~w36159 & w36522 ) | ( w36521 & w36522 ) ;
  assign w36524 = w36522 | w36523 ;
  assign w36525 = \pi106 ^ w36146 ;
  assign w36526 = ( ~w36153 & w36524 ) | ( ~w36153 & w36525 ) | ( w36524 & w36525 ) ;
  assign w36527 = w36525 | w36526 ;
  assign w36528 = \pi107 ^ w36140 ;
  assign w36529 = ( ~w36147 & w36527 ) | ( ~w36147 & w36528 ) | ( w36527 & w36528 ) ;
  assign w36530 = w36528 | w36529 ;
  assign w36531 = \pi108 ^ w36134 ;
  assign w36532 = ( ~w36141 & w36530 ) | ( ~w36141 & w36531 ) | ( w36530 & w36531 ) ;
  assign w36533 = w36531 | w36532 ;
  assign w36534 = \pi109 ^ w36128 ;
  assign w36535 = ( ~w36135 & w36533 ) | ( ~w36135 & w36534 ) | ( w36533 & w36534 ) ;
  assign w36536 = w36534 | w36535 ;
  assign w36537 = \pi110 ^ w36122 ;
  assign w36538 = ( ~w36129 & w36536 ) | ( ~w36129 & w36537 ) | ( w36536 & w36537 ) ;
  assign w36539 = w36537 | w36538 ;
  assign w36540 = \pi111 ^ w36116 ;
  assign w36541 = ( ~w36123 & w36539 ) | ( ~w36123 & w36540 ) | ( w36539 & w36540 ) ;
  assign w36542 = w36540 | w36541 ;
  assign w36543 = \pi112 ^ w36110 ;
  assign w36544 = ( ~w36117 & w36542 ) | ( ~w36117 & w36543 ) | ( w36542 & w36543 ) ;
  assign w36545 = w36543 | w36544 ;
  assign w36546 = \pi113 ^ w36104 ;
  assign w36547 = ( ~w36111 & w36545 ) | ( ~w36111 & w36546 ) | ( w36545 & w36546 ) ;
  assign w36548 = w36546 | w36547 ;
  assign w36549 = \pi114 ^ w36098 ;
  assign w36550 = ( ~w36105 & w36548 ) | ( ~w36105 & w36549 ) | ( w36548 & w36549 ) ;
  assign w36551 = w36549 | w36550 ;
  assign w36552 = \pi115 ^ w36092 ;
  assign w36553 = ( ~w36099 & w36551 ) | ( ~w36099 & w36552 ) | ( w36551 & w36552 ) ;
  assign w36554 = w36552 | w36553 ;
  assign w36555 = \pi116 ^ w36086 ;
  assign w36556 = ( ~w36093 & w36554 ) | ( ~w36093 & w36555 ) | ( w36554 & w36555 ) ;
  assign w36557 = w36555 | w36556 ;
  assign w36558 = \pi117 ^ w36080 ;
  assign w36559 = ( ~w36087 & w36557 ) | ( ~w36087 & w36558 ) | ( w36557 & w36558 ) ;
  assign w36560 = w36558 | w36559 ;
  assign w36561 = \pi118 ^ w36074 ;
  assign w36562 = ( ~w36081 & w36560 ) | ( ~w36081 & w36561 ) | ( w36560 & w36561 ) ;
  assign w36563 = w36561 | w36562 ;
  assign w36564 = \pi119 ^ w36068 ;
  assign w36565 = ( ~w36075 & w36563 ) | ( ~w36075 & w36564 ) | ( w36563 & w36564 ) ;
  assign w36566 = w36564 | w36565 ;
  assign w36567 = \pi120 ^ w36062 ;
  assign w36568 = ( ~w36069 & w36566 ) | ( ~w36069 & w36567 ) | ( w36566 & w36567 ) ;
  assign w36569 = w36567 | w36568 ;
  assign w36570 = \pi121 ^ w36056 ;
  assign w36571 = ( ~w36063 & w36569 ) | ( ~w36063 & w36570 ) | ( w36569 & w36570 ) ;
  assign w36572 = w36570 | w36571 ;
  assign w36573 = w35497 & w36051 ;
  assign w36574 = ~w35498 & w36045 ;
  assign w36575 = w36046 ^ w36574 ;
  assign w36576 = ~w36051 & w36575 ;
  assign w36577 = w36573 | w36576 ;
  assign w36578 = ~\pi122 & w36577 ;
  assign w36579 = ( \pi122 & ~w36573 ) | ( \pi122 & w36576 ) | ( ~w36573 & w36576 ) ;
  assign w36580 = ~w36576 & w36579 ;
  assign w36581 = ( ~w36057 & w36572 ) | ( ~w36057 & w36578 ) | ( w36572 & w36578 ) ;
  assign w36582 = ( w270 & w36578 ) | ( w270 & ~w36581 ) | ( w36578 & ~w36581 ) ;
  assign w36583 = ( w269 & w36580 ) | ( w269 & ~w36581 ) | ( w36580 & ~w36581 ) ;
  assign w36584 = ( w36581 & ~w36582 ) | ( w36581 & w36583 ) | ( ~w36582 & w36583 ) ;
  assign w36585 = w36582 | w36584 ;
  assign w36586 = ~w16707 & w36577 ;
  assign w36587 = w36585 & ~w36586 ;
  assign w36588 = ~w36063 & w36569 ;
  assign w36589 = w36570 ^ w36588 ;
  assign w36590 = ~w36587 & w36589 ;
  assign w36591 = ( w36056 & w36585 ) | ( w36056 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36592 = ~w36586 & w36591 ;
  assign w36593 = w36590 | w36592 ;
  assign w36594 = ~\pi122 & w36593 ;
  assign w36595 = ~w36069 & w36566 ;
  assign w36596 = w36567 ^ w36595 ;
  assign w36597 = ~w36587 & w36596 ;
  assign w36598 = ( w36062 & w36585 ) | ( w36062 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36599 = ~w36586 & w36598 ;
  assign w36600 = w36597 | w36599 ;
  assign w36601 = ~\pi121 & w36600 ;
  assign w36602 = ~w36075 & w36563 ;
  assign w36603 = w36564 ^ w36602 ;
  assign w36604 = ~w36587 & w36603 ;
  assign w36605 = ( w36068 & w36585 ) | ( w36068 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36606 = ~w36586 & w36605 ;
  assign w36607 = w36604 | w36606 ;
  assign w36608 = ~\pi120 & w36607 ;
  assign w36609 = ~w36081 & w36560 ;
  assign w36610 = w36561 ^ w36609 ;
  assign w36611 = ~w36587 & w36610 ;
  assign w36612 = ( w36074 & w36585 ) | ( w36074 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36613 = ~w36586 & w36612 ;
  assign w36614 = w36611 | w36613 ;
  assign w36615 = ~\pi119 & w36614 ;
  assign w36616 = ~w36087 & w36557 ;
  assign w36617 = w36558 ^ w36616 ;
  assign w36618 = ~w36587 & w36617 ;
  assign w36619 = ( w36080 & w36585 ) | ( w36080 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36620 = ~w36586 & w36619 ;
  assign w36621 = w36618 | w36620 ;
  assign w36622 = ~\pi118 & w36621 ;
  assign w36623 = ~w36093 & w36554 ;
  assign w36624 = w36555 ^ w36623 ;
  assign w36625 = ~w36587 & w36624 ;
  assign w36626 = ( w36086 & w36585 ) | ( w36086 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36627 = ~w36586 & w36626 ;
  assign w36628 = w36625 | w36627 ;
  assign w36629 = ~\pi117 & w36628 ;
  assign w36630 = ~w36099 & w36551 ;
  assign w36631 = w36552 ^ w36630 ;
  assign w36632 = ~w36587 & w36631 ;
  assign w36633 = ( w36092 & w36585 ) | ( w36092 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36634 = ~w36586 & w36633 ;
  assign w36635 = w36632 | w36634 ;
  assign w36636 = ~\pi116 & w36635 ;
  assign w36637 = ~w36105 & w36548 ;
  assign w36638 = w36549 ^ w36637 ;
  assign w36639 = ~w36587 & w36638 ;
  assign w36640 = ( w36098 & w36585 ) | ( w36098 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36641 = ~w36586 & w36640 ;
  assign w36642 = w36639 | w36641 ;
  assign w36643 = ~\pi115 & w36642 ;
  assign w36644 = ~w36111 & w36545 ;
  assign w36645 = w36546 ^ w36644 ;
  assign w36646 = ~w36587 & w36645 ;
  assign w36647 = ( w36104 & w36585 ) | ( w36104 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36648 = ~w36586 & w36647 ;
  assign w36649 = w36646 | w36648 ;
  assign w36650 = ~\pi114 & w36649 ;
  assign w36651 = ~w36117 & w36542 ;
  assign w36652 = w36543 ^ w36651 ;
  assign w36653 = ~w36587 & w36652 ;
  assign w36654 = ( w36110 & w36585 ) | ( w36110 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36655 = ~w36586 & w36654 ;
  assign w36656 = w36653 | w36655 ;
  assign w36657 = ~\pi113 & w36656 ;
  assign w36658 = ~w36123 & w36539 ;
  assign w36659 = w36540 ^ w36658 ;
  assign w36660 = ~w36587 & w36659 ;
  assign w36661 = ( w36116 & w36585 ) | ( w36116 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36662 = ~w36586 & w36661 ;
  assign w36663 = w36660 | w36662 ;
  assign w36664 = ~\pi112 & w36663 ;
  assign w36665 = ~w36129 & w36536 ;
  assign w36666 = w36537 ^ w36665 ;
  assign w36667 = ~w36587 & w36666 ;
  assign w36668 = ( w36122 & w36585 ) | ( w36122 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36669 = ~w36586 & w36668 ;
  assign w36670 = w36667 | w36669 ;
  assign w36671 = ~\pi111 & w36670 ;
  assign w36672 = ~w36135 & w36533 ;
  assign w36673 = w36534 ^ w36672 ;
  assign w36674 = ~w36587 & w36673 ;
  assign w36675 = ( w36128 & w36585 ) | ( w36128 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36676 = ~w36586 & w36675 ;
  assign w36677 = w36674 | w36676 ;
  assign w36678 = ~\pi110 & w36677 ;
  assign w36679 = ~w36141 & w36530 ;
  assign w36680 = w36531 ^ w36679 ;
  assign w36681 = ~w36587 & w36680 ;
  assign w36682 = ( w36134 & w36585 ) | ( w36134 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36683 = ~w36586 & w36682 ;
  assign w36684 = w36681 | w36683 ;
  assign w36685 = ~\pi109 & w36684 ;
  assign w36686 = ~w36147 & w36527 ;
  assign w36687 = w36528 ^ w36686 ;
  assign w36688 = ~w36587 & w36687 ;
  assign w36689 = ( w36140 & w36585 ) | ( w36140 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36690 = ~w36586 & w36689 ;
  assign w36691 = w36688 | w36690 ;
  assign w36692 = ~\pi108 & w36691 ;
  assign w36693 = ~w36153 & w36524 ;
  assign w36694 = w36525 ^ w36693 ;
  assign w36695 = ~w36587 & w36694 ;
  assign w36696 = ( w36146 & w36585 ) | ( w36146 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36697 = ~w36586 & w36696 ;
  assign w36698 = w36695 | w36697 ;
  assign w36699 = ~\pi107 & w36698 ;
  assign w36700 = ~w36159 & w36521 ;
  assign w36701 = w36522 ^ w36700 ;
  assign w36702 = ~w36587 & w36701 ;
  assign w36703 = ( w36152 & w36585 ) | ( w36152 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36704 = ~w36586 & w36703 ;
  assign w36705 = w36702 | w36704 ;
  assign w36706 = ~\pi106 & w36705 ;
  assign w36707 = ~w36165 & w36518 ;
  assign w36708 = w36519 ^ w36707 ;
  assign w36709 = ~w36587 & w36708 ;
  assign w36710 = ( w36158 & w36585 ) | ( w36158 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36711 = ~w36586 & w36710 ;
  assign w36712 = w36709 | w36711 ;
  assign w36713 = ~\pi105 & w36712 ;
  assign w36714 = ~w36171 & w36515 ;
  assign w36715 = w36516 ^ w36714 ;
  assign w36716 = ~w36587 & w36715 ;
  assign w36717 = ( w36164 & w36585 ) | ( w36164 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36718 = ~w36586 & w36717 ;
  assign w36719 = w36716 | w36718 ;
  assign w36720 = ~\pi104 & w36719 ;
  assign w36721 = ~w36177 & w36512 ;
  assign w36722 = w36513 ^ w36721 ;
  assign w36723 = ~w36587 & w36722 ;
  assign w36724 = ( w36170 & w36585 ) | ( w36170 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36725 = ~w36586 & w36724 ;
  assign w36726 = w36723 | w36725 ;
  assign w36727 = ~\pi103 & w36726 ;
  assign w36728 = ~w36183 & w36509 ;
  assign w36729 = w36510 ^ w36728 ;
  assign w36730 = ~w36587 & w36729 ;
  assign w36731 = ( w36176 & w36585 ) | ( w36176 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36732 = ~w36586 & w36731 ;
  assign w36733 = w36730 | w36732 ;
  assign w36734 = ~\pi102 & w36733 ;
  assign w36735 = ~w36189 & w36506 ;
  assign w36736 = w36507 ^ w36735 ;
  assign w36737 = ~w36587 & w36736 ;
  assign w36738 = ( w36182 & w36585 ) | ( w36182 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36739 = ~w36586 & w36738 ;
  assign w36740 = w36737 | w36739 ;
  assign w36741 = ~\pi101 & w36740 ;
  assign w36742 = ~w36195 & w36503 ;
  assign w36743 = w36504 ^ w36742 ;
  assign w36744 = ~w36587 & w36743 ;
  assign w36745 = ( w36188 & w36585 ) | ( w36188 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36746 = ~w36586 & w36745 ;
  assign w36747 = w36744 | w36746 ;
  assign w36748 = ~\pi100 & w36747 ;
  assign w36749 = ~w36201 & w36500 ;
  assign w36750 = w36501 ^ w36749 ;
  assign w36751 = ~w36587 & w36750 ;
  assign w36752 = ( w36194 & w36585 ) | ( w36194 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36753 = ~w36586 & w36752 ;
  assign w36754 = w36751 | w36753 ;
  assign w36755 = ~\pi099 & w36754 ;
  assign w36756 = ~w36207 & w36497 ;
  assign w36757 = w36498 ^ w36756 ;
  assign w36758 = ~w36587 & w36757 ;
  assign w36759 = ( w36200 & w36585 ) | ( w36200 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36760 = ~w36586 & w36759 ;
  assign w36761 = w36758 | w36760 ;
  assign w36762 = ~\pi098 & w36761 ;
  assign w36763 = ~w36213 & w36494 ;
  assign w36764 = w36495 ^ w36763 ;
  assign w36765 = ~w36587 & w36764 ;
  assign w36766 = ( w36206 & w36585 ) | ( w36206 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36767 = ~w36586 & w36766 ;
  assign w36768 = w36765 | w36767 ;
  assign w36769 = ~\pi097 & w36768 ;
  assign w36770 = ~w36219 & w36491 ;
  assign w36771 = w36492 ^ w36770 ;
  assign w36772 = ~w36587 & w36771 ;
  assign w36773 = ( w36212 & w36585 ) | ( w36212 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36774 = ~w36586 & w36773 ;
  assign w36775 = w36772 | w36774 ;
  assign w36776 = ~\pi096 & w36775 ;
  assign w36777 = ~w36225 & w36488 ;
  assign w36778 = w36489 ^ w36777 ;
  assign w36779 = ~w36587 & w36778 ;
  assign w36780 = ( w36218 & w36585 ) | ( w36218 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36781 = ~w36586 & w36780 ;
  assign w36782 = w36779 | w36781 ;
  assign w36783 = ~\pi095 & w36782 ;
  assign w36784 = ~w36231 & w36485 ;
  assign w36785 = w36486 ^ w36784 ;
  assign w36786 = ~w36587 & w36785 ;
  assign w36787 = ( w36224 & w36585 ) | ( w36224 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36788 = ~w36586 & w36787 ;
  assign w36789 = w36786 | w36788 ;
  assign w36790 = ~\pi094 & w36789 ;
  assign w36791 = ~w36237 & w36482 ;
  assign w36792 = w36483 ^ w36791 ;
  assign w36793 = ~w36587 & w36792 ;
  assign w36794 = ( w36230 & w36585 ) | ( w36230 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36795 = ~w36586 & w36794 ;
  assign w36796 = w36793 | w36795 ;
  assign w36797 = ~\pi093 & w36796 ;
  assign w36798 = ~w36243 & w36479 ;
  assign w36799 = w36480 ^ w36798 ;
  assign w36800 = ~w36587 & w36799 ;
  assign w36801 = ( w36236 & w36585 ) | ( w36236 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36802 = ~w36586 & w36801 ;
  assign w36803 = w36800 | w36802 ;
  assign w36804 = ~\pi092 & w36803 ;
  assign w36805 = ~w36249 & w36476 ;
  assign w36806 = w36477 ^ w36805 ;
  assign w36807 = ~w36587 & w36806 ;
  assign w36808 = ( w36242 & w36585 ) | ( w36242 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36809 = ~w36586 & w36808 ;
  assign w36810 = w36807 | w36809 ;
  assign w36811 = ~\pi091 & w36810 ;
  assign w36812 = ~w36255 & w36473 ;
  assign w36813 = w36474 ^ w36812 ;
  assign w36814 = ~w36587 & w36813 ;
  assign w36815 = ( w36248 & w36585 ) | ( w36248 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36816 = ~w36586 & w36815 ;
  assign w36817 = w36814 | w36816 ;
  assign w36818 = ~\pi090 & w36817 ;
  assign w36819 = ~w36261 & w36470 ;
  assign w36820 = w36471 ^ w36819 ;
  assign w36821 = ~w36587 & w36820 ;
  assign w36822 = ( w36254 & w36585 ) | ( w36254 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36823 = ~w36586 & w36822 ;
  assign w36824 = w36821 | w36823 ;
  assign w36825 = ~\pi089 & w36824 ;
  assign w36826 = ~w36267 & w36467 ;
  assign w36827 = w36468 ^ w36826 ;
  assign w36828 = ~w36587 & w36827 ;
  assign w36829 = ( w36260 & w36585 ) | ( w36260 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36830 = ~w36586 & w36829 ;
  assign w36831 = w36828 | w36830 ;
  assign w36832 = ~\pi088 & w36831 ;
  assign w36833 = ~w36273 & w36464 ;
  assign w36834 = w36465 ^ w36833 ;
  assign w36835 = ~w36587 & w36834 ;
  assign w36836 = ( w36266 & w36585 ) | ( w36266 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36837 = ~w36586 & w36836 ;
  assign w36838 = w36835 | w36837 ;
  assign w36839 = ~\pi087 & w36838 ;
  assign w36840 = ~w36279 & w36461 ;
  assign w36841 = w36462 ^ w36840 ;
  assign w36842 = ~w36587 & w36841 ;
  assign w36843 = ( w36272 & w36585 ) | ( w36272 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36844 = ~w36586 & w36843 ;
  assign w36845 = w36842 | w36844 ;
  assign w36846 = ~\pi086 & w36845 ;
  assign w36847 = ~w36285 & w36458 ;
  assign w36848 = w36459 ^ w36847 ;
  assign w36849 = ~w36587 & w36848 ;
  assign w36850 = ( w36278 & w36585 ) | ( w36278 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36851 = ~w36586 & w36850 ;
  assign w36852 = w36849 | w36851 ;
  assign w36853 = ~\pi085 & w36852 ;
  assign w36854 = ~w36291 & w36455 ;
  assign w36855 = w36456 ^ w36854 ;
  assign w36856 = ~w36587 & w36855 ;
  assign w36857 = ( w36284 & w36585 ) | ( w36284 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36858 = ~w36586 & w36857 ;
  assign w36859 = w36856 | w36858 ;
  assign w36860 = ~\pi084 & w36859 ;
  assign w36861 = ~w36297 & w36452 ;
  assign w36862 = w36453 ^ w36861 ;
  assign w36863 = ~w36587 & w36862 ;
  assign w36864 = ( w36290 & w36585 ) | ( w36290 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36865 = ~w36586 & w36864 ;
  assign w36866 = w36863 | w36865 ;
  assign w36867 = ~\pi083 & w36866 ;
  assign w36868 = ~w36303 & w36449 ;
  assign w36869 = w36450 ^ w36868 ;
  assign w36870 = ~w36587 & w36869 ;
  assign w36871 = ( w36296 & w36585 ) | ( w36296 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36872 = ~w36586 & w36871 ;
  assign w36873 = w36870 | w36872 ;
  assign w36874 = ~\pi082 & w36873 ;
  assign w36875 = ~w36309 & w36446 ;
  assign w36876 = w36447 ^ w36875 ;
  assign w36877 = ~w36587 & w36876 ;
  assign w36878 = ( w36302 & w36585 ) | ( w36302 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36879 = ~w36586 & w36878 ;
  assign w36880 = w36877 | w36879 ;
  assign w36881 = ~\pi081 & w36880 ;
  assign w36882 = ~w36315 & w36443 ;
  assign w36883 = w36444 ^ w36882 ;
  assign w36884 = ~w36587 & w36883 ;
  assign w36885 = ( w36308 & w36585 ) | ( w36308 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36886 = ~w36586 & w36885 ;
  assign w36887 = w36884 | w36886 ;
  assign w36888 = ~\pi080 & w36887 ;
  assign w36889 = ~w36321 & w36440 ;
  assign w36890 = w36441 ^ w36889 ;
  assign w36891 = ~w36587 & w36890 ;
  assign w36892 = ( w36314 & w36585 ) | ( w36314 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36893 = ~w36586 & w36892 ;
  assign w36894 = w36891 | w36893 ;
  assign w36895 = ~\pi079 & w36894 ;
  assign w36896 = ~w36327 & w36437 ;
  assign w36897 = w36438 ^ w36896 ;
  assign w36898 = ~w36587 & w36897 ;
  assign w36899 = ( w36320 & w36585 ) | ( w36320 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36900 = ~w36586 & w36899 ;
  assign w36901 = w36898 | w36900 ;
  assign w36902 = ~\pi078 & w36901 ;
  assign w36903 = ~w36333 & w36434 ;
  assign w36904 = w36435 ^ w36903 ;
  assign w36905 = ~w36587 & w36904 ;
  assign w36906 = ( w36326 & w36585 ) | ( w36326 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36907 = ~w36586 & w36906 ;
  assign w36908 = w36905 | w36907 ;
  assign w36909 = ~\pi077 & w36908 ;
  assign w36910 = ~w36339 & w36431 ;
  assign w36911 = w36432 ^ w36910 ;
  assign w36912 = ~w36587 & w36911 ;
  assign w36913 = ( w36332 & w36585 ) | ( w36332 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36914 = ~w36586 & w36913 ;
  assign w36915 = w36912 | w36914 ;
  assign w36916 = ~\pi076 & w36915 ;
  assign w36917 = ~w36345 & w36428 ;
  assign w36918 = w36429 ^ w36917 ;
  assign w36919 = ~w36587 & w36918 ;
  assign w36920 = ( w36338 & w36585 ) | ( w36338 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36921 = ~w36586 & w36920 ;
  assign w36922 = w36919 | w36921 ;
  assign w36923 = ~\pi075 & w36922 ;
  assign w36924 = ~w36351 & w36425 ;
  assign w36925 = w36426 ^ w36924 ;
  assign w36926 = ~w36587 & w36925 ;
  assign w36927 = ( w36344 & w36585 ) | ( w36344 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36928 = ~w36586 & w36927 ;
  assign w36929 = w36926 | w36928 ;
  assign w36930 = ~\pi074 & w36929 ;
  assign w36931 = ~w36357 & w36422 ;
  assign w36932 = w36423 ^ w36931 ;
  assign w36933 = ~w36587 & w36932 ;
  assign w36934 = ( w36350 & w36585 ) | ( w36350 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36935 = ~w36586 & w36934 ;
  assign w36936 = w36933 | w36935 ;
  assign w36937 = ~\pi073 & w36936 ;
  assign w36938 = ~w36363 & w36419 ;
  assign w36939 = w36420 ^ w36938 ;
  assign w36940 = ~w36587 & w36939 ;
  assign w36941 = ( w36356 & w36585 ) | ( w36356 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36942 = ~w36586 & w36941 ;
  assign w36943 = w36940 | w36942 ;
  assign w36944 = ~\pi072 & w36943 ;
  assign w36945 = ~w36369 & w36416 ;
  assign w36946 = w36417 ^ w36945 ;
  assign w36947 = ~w36587 & w36946 ;
  assign w36948 = ( w36362 & w36585 ) | ( w36362 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36949 = ~w36586 & w36948 ;
  assign w36950 = w36947 | w36949 ;
  assign w36951 = ~\pi071 & w36950 ;
  assign w36952 = ~w36375 & w36413 ;
  assign w36953 = w36414 ^ w36952 ;
  assign w36954 = ~w36587 & w36953 ;
  assign w36955 = ( w36368 & w36585 ) | ( w36368 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36956 = ~w36586 & w36955 ;
  assign w36957 = w36954 | w36956 ;
  assign w36958 = ~\pi070 & w36957 ;
  assign w36959 = ~w36384 & w36410 ;
  assign w36960 = w36411 ^ w36959 ;
  assign w36961 = ~w36587 & w36960 ;
  assign w36962 = ( w36374 & w36585 ) | ( w36374 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36963 = ~w36586 & w36962 ;
  assign w36964 = w36961 | w36963 ;
  assign w36965 = ~\pi069 & w36964 ;
  assign w36966 = ~w36394 & w36405 ;
  assign w36967 = w36408 ^ w36966 ;
  assign w36968 = ~w36587 & w36967 ;
  assign w36969 = ( w36383 & w36585 ) | ( w36383 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36970 = ~w36586 & w36969 ;
  assign w36971 = w36968 | w36970 ;
  assign w36972 = ~\pi068 & w36971 ;
  assign w36973 = w36402 ^ w36404 ;
  assign w36974 = ~w36587 & w36973 ;
  assign w36975 = ( w36393 & w36585 ) | ( w36393 & w36586 ) | ( w36585 & w36586 ) ;
  assign w36976 = ~w36586 & w36975 ;
  assign w36977 = w36974 | w36976 ;
  assign w36978 = ~\pi067 & w36977 ;
  assign w36979 = w17062 ^ w36403 ;
  assign w36980 = \pi065 ^ w36979 ;
  assign w36981 = ~w36587 & w36980 ;
  assign w36982 = ( w36396 & w36399 ) | ( w36396 & ~w36586 ) | ( w36399 & ~w36586 ) ;
  assign w36983 = w36586 & w36982 ;
  assign w36984 = ( ~w36585 & w36982 ) | ( ~w36585 & w36983 ) | ( w36982 & w36983 ) ;
  assign w36985 = ( w36981 & w36982 ) | ( w36981 & ~w36984 ) | ( w36982 & ~w36984 ) ;
  assign w36986 = ~\pi066 & w36985 ;
  assign w36987 = w36585 | w36586 ;
  assign w36988 = ( w36981 & w36982 ) | ( w36981 & w36987 ) | ( w36982 & w36987 ) ;
  assign w36989 = ( ~w36586 & w36981 ) | ( ~w36586 & w36988 ) | ( w36981 & w36988 ) ;
  assign w36990 = \pi066 ^ w36989 ;
  assign w36991 = ( \pi064 & ~w36587 ) | ( \pi064 & w36990 ) | ( ~w36587 & w36990 ) ;
  assign w36992 = \pi005 ^ w36991 ;
  assign w36993 = ( \pi065 & w18236 ) | ( \pi065 & ~w36992 ) | ( w18236 & ~w36992 ) ;
  assign w36994 = w36990 | w36993 ;
  assign w36995 = \pi067 ^ w36977 ;
  assign w36996 = ( ~w36986 & w36994 ) | ( ~w36986 & w36995 ) | ( w36994 & w36995 ) ;
  assign w36997 = w36995 | w36996 ;
  assign w36998 = \pi068 ^ w36971 ;
  assign w36999 = ( ~w36978 & w36997 ) | ( ~w36978 & w36998 ) | ( w36997 & w36998 ) ;
  assign w37000 = w36998 | w36999 ;
  assign w37001 = \pi069 ^ w36964 ;
  assign w37002 = ( ~w36972 & w37000 ) | ( ~w36972 & w37001 ) | ( w37000 & w37001 ) ;
  assign w37003 = w37001 | w37002 ;
  assign w37004 = \pi070 ^ w36957 ;
  assign w37005 = ( ~w36965 & w37003 ) | ( ~w36965 & w37004 ) | ( w37003 & w37004 ) ;
  assign w37006 = w37004 | w37005 ;
  assign w37007 = \pi071 ^ w36950 ;
  assign w37008 = ( ~w36958 & w37006 ) | ( ~w36958 & w37007 ) | ( w37006 & w37007 ) ;
  assign w37009 = w37007 | w37008 ;
  assign w37010 = \pi072 ^ w36943 ;
  assign w37011 = ( ~w36951 & w37009 ) | ( ~w36951 & w37010 ) | ( w37009 & w37010 ) ;
  assign w37012 = w37010 | w37011 ;
  assign w37013 = \pi073 ^ w36936 ;
  assign w37014 = ( ~w36944 & w37012 ) | ( ~w36944 & w37013 ) | ( w37012 & w37013 ) ;
  assign w37015 = w37013 | w37014 ;
  assign w37016 = \pi074 ^ w36929 ;
  assign w37017 = ( ~w36937 & w37015 ) | ( ~w36937 & w37016 ) | ( w37015 & w37016 ) ;
  assign w37018 = w37016 | w37017 ;
  assign w37019 = \pi075 ^ w36922 ;
  assign w37020 = ( ~w36930 & w37018 ) | ( ~w36930 & w37019 ) | ( w37018 & w37019 ) ;
  assign w37021 = w37019 | w37020 ;
  assign w37022 = \pi076 ^ w36915 ;
  assign w37023 = ( ~w36923 & w37021 ) | ( ~w36923 & w37022 ) | ( w37021 & w37022 ) ;
  assign w37024 = w37022 | w37023 ;
  assign w37025 = \pi077 ^ w36908 ;
  assign w37026 = ( ~w36916 & w37024 ) | ( ~w36916 & w37025 ) | ( w37024 & w37025 ) ;
  assign w37027 = w37025 | w37026 ;
  assign w37028 = \pi078 ^ w36901 ;
  assign w37029 = ( ~w36909 & w37027 ) | ( ~w36909 & w37028 ) | ( w37027 & w37028 ) ;
  assign w37030 = w37028 | w37029 ;
  assign w37031 = \pi079 ^ w36894 ;
  assign w37032 = ( ~w36902 & w37030 ) | ( ~w36902 & w37031 ) | ( w37030 & w37031 ) ;
  assign w37033 = w37031 | w37032 ;
  assign w37034 = \pi080 ^ w36887 ;
  assign w37035 = ( ~w36895 & w37033 ) | ( ~w36895 & w37034 ) | ( w37033 & w37034 ) ;
  assign w37036 = w37034 | w37035 ;
  assign w37037 = \pi081 ^ w36880 ;
  assign w37038 = ( ~w36888 & w37036 ) | ( ~w36888 & w37037 ) | ( w37036 & w37037 ) ;
  assign w37039 = w37037 | w37038 ;
  assign w37040 = \pi082 ^ w36873 ;
  assign w37041 = ( ~w36881 & w37039 ) | ( ~w36881 & w37040 ) | ( w37039 & w37040 ) ;
  assign w37042 = w37040 | w37041 ;
  assign w37043 = \pi083 ^ w36866 ;
  assign w37044 = ( ~w36874 & w37042 ) | ( ~w36874 & w37043 ) | ( w37042 & w37043 ) ;
  assign w37045 = w37043 | w37044 ;
  assign w37046 = \pi084 ^ w36859 ;
  assign w37047 = ( ~w36867 & w37045 ) | ( ~w36867 & w37046 ) | ( w37045 & w37046 ) ;
  assign w37048 = w37046 | w37047 ;
  assign w37049 = \pi085 ^ w36852 ;
  assign w37050 = ( ~w36860 & w37048 ) | ( ~w36860 & w37049 ) | ( w37048 & w37049 ) ;
  assign w37051 = w37049 | w37050 ;
  assign w37052 = \pi086 ^ w36845 ;
  assign w37053 = ( ~w36853 & w37051 ) | ( ~w36853 & w37052 ) | ( w37051 & w37052 ) ;
  assign w37054 = w37052 | w37053 ;
  assign w37055 = \pi087 ^ w36838 ;
  assign w37056 = ( ~w36846 & w37054 ) | ( ~w36846 & w37055 ) | ( w37054 & w37055 ) ;
  assign w37057 = w37055 | w37056 ;
  assign w37058 = \pi088 ^ w36831 ;
  assign w37059 = ( ~w36839 & w37057 ) | ( ~w36839 & w37058 ) | ( w37057 & w37058 ) ;
  assign w37060 = w37058 | w37059 ;
  assign w37061 = \pi089 ^ w36824 ;
  assign w37062 = ( ~w36832 & w37060 ) | ( ~w36832 & w37061 ) | ( w37060 & w37061 ) ;
  assign w37063 = w37061 | w37062 ;
  assign w37064 = \pi090 ^ w36817 ;
  assign w37065 = ( ~w36825 & w37063 ) | ( ~w36825 & w37064 ) | ( w37063 & w37064 ) ;
  assign w37066 = w37064 | w37065 ;
  assign w37067 = \pi091 ^ w36810 ;
  assign w37068 = ( ~w36818 & w37066 ) | ( ~w36818 & w37067 ) | ( w37066 & w37067 ) ;
  assign w37069 = w37067 | w37068 ;
  assign w37070 = \pi092 ^ w36803 ;
  assign w37071 = ( ~w36811 & w37069 ) | ( ~w36811 & w37070 ) | ( w37069 & w37070 ) ;
  assign w37072 = w37070 | w37071 ;
  assign w37073 = \pi093 ^ w36796 ;
  assign w37074 = ( ~w36804 & w37072 ) | ( ~w36804 & w37073 ) | ( w37072 & w37073 ) ;
  assign w37075 = w37073 | w37074 ;
  assign w37076 = \pi094 ^ w36789 ;
  assign w37077 = ( ~w36797 & w37075 ) | ( ~w36797 & w37076 ) | ( w37075 & w37076 ) ;
  assign w37078 = w37076 | w37077 ;
  assign w37079 = \pi095 ^ w36782 ;
  assign w37080 = ( ~w36790 & w37078 ) | ( ~w36790 & w37079 ) | ( w37078 & w37079 ) ;
  assign w37081 = w37079 | w37080 ;
  assign w37082 = \pi096 ^ w36775 ;
  assign w37083 = ( ~w36783 & w37081 ) | ( ~w36783 & w37082 ) | ( w37081 & w37082 ) ;
  assign w37084 = w37082 | w37083 ;
  assign w37085 = \pi097 ^ w36768 ;
  assign w37086 = ( ~w36776 & w37084 ) | ( ~w36776 & w37085 ) | ( w37084 & w37085 ) ;
  assign w37087 = w37085 | w37086 ;
  assign w37088 = \pi098 ^ w36761 ;
  assign w37089 = ( ~w36769 & w37087 ) | ( ~w36769 & w37088 ) | ( w37087 & w37088 ) ;
  assign w37090 = w37088 | w37089 ;
  assign w37091 = \pi099 ^ w36754 ;
  assign w37092 = ( ~w36762 & w37090 ) | ( ~w36762 & w37091 ) | ( w37090 & w37091 ) ;
  assign w37093 = w37091 | w37092 ;
  assign w37094 = \pi100 ^ w36747 ;
  assign w37095 = ( ~w36755 & w37093 ) | ( ~w36755 & w37094 ) | ( w37093 & w37094 ) ;
  assign w37096 = w37094 | w37095 ;
  assign w37097 = \pi101 ^ w36740 ;
  assign w37098 = ( ~w36748 & w37096 ) | ( ~w36748 & w37097 ) | ( w37096 & w37097 ) ;
  assign w37099 = w37097 | w37098 ;
  assign w37100 = \pi102 ^ w36733 ;
  assign w37101 = ( ~w36741 & w37099 ) | ( ~w36741 & w37100 ) | ( w37099 & w37100 ) ;
  assign w37102 = w37100 | w37101 ;
  assign w37103 = \pi103 ^ w36726 ;
  assign w37104 = ( ~w36734 & w37102 ) | ( ~w36734 & w37103 ) | ( w37102 & w37103 ) ;
  assign w37105 = w37103 | w37104 ;
  assign w37106 = \pi104 ^ w36719 ;
  assign w37107 = ( ~w36727 & w37105 ) | ( ~w36727 & w37106 ) | ( w37105 & w37106 ) ;
  assign w37108 = w37106 | w37107 ;
  assign w37109 = \pi105 ^ w36712 ;
  assign w37110 = ( ~w36720 & w37108 ) | ( ~w36720 & w37109 ) | ( w37108 & w37109 ) ;
  assign w37111 = w37109 | w37110 ;
  assign w37112 = \pi106 ^ w36705 ;
  assign w37113 = ( ~w36713 & w37111 ) | ( ~w36713 & w37112 ) | ( w37111 & w37112 ) ;
  assign w37114 = w37112 | w37113 ;
  assign w37115 = \pi107 ^ w36698 ;
  assign w37116 = ( ~w36706 & w37114 ) | ( ~w36706 & w37115 ) | ( w37114 & w37115 ) ;
  assign w37117 = w37115 | w37116 ;
  assign w37118 = \pi108 ^ w36691 ;
  assign w37119 = ( ~w36699 & w37117 ) | ( ~w36699 & w37118 ) | ( w37117 & w37118 ) ;
  assign w37120 = w37118 | w37119 ;
  assign w37121 = \pi109 ^ w36684 ;
  assign w37122 = ( ~w36692 & w37120 ) | ( ~w36692 & w37121 ) | ( w37120 & w37121 ) ;
  assign w37123 = w37121 | w37122 ;
  assign w37124 = \pi110 ^ w36677 ;
  assign w37125 = ( ~w36685 & w37123 ) | ( ~w36685 & w37124 ) | ( w37123 & w37124 ) ;
  assign w37126 = w37124 | w37125 ;
  assign w37127 = \pi111 ^ w36670 ;
  assign w37128 = ( ~w36678 & w37126 ) | ( ~w36678 & w37127 ) | ( w37126 & w37127 ) ;
  assign w37129 = w37127 | w37128 ;
  assign w37130 = \pi112 ^ w36663 ;
  assign w37131 = ( ~w36671 & w37129 ) | ( ~w36671 & w37130 ) | ( w37129 & w37130 ) ;
  assign w37132 = w37130 | w37131 ;
  assign w37133 = \pi113 ^ w36656 ;
  assign w37134 = ( ~w36664 & w37132 ) | ( ~w36664 & w37133 ) | ( w37132 & w37133 ) ;
  assign w37135 = w37133 | w37134 ;
  assign w37136 = \pi114 ^ w36649 ;
  assign w37137 = ( ~w36657 & w37135 ) | ( ~w36657 & w37136 ) | ( w37135 & w37136 ) ;
  assign w37138 = w37136 | w37137 ;
  assign w37139 = \pi115 ^ w36642 ;
  assign w37140 = ( ~w36650 & w37138 ) | ( ~w36650 & w37139 ) | ( w37138 & w37139 ) ;
  assign w37141 = w37139 | w37140 ;
  assign w37142 = \pi116 ^ w36635 ;
  assign w37143 = ( ~w36643 & w37141 ) | ( ~w36643 & w37142 ) | ( w37141 & w37142 ) ;
  assign w37144 = w37142 | w37143 ;
  assign w37145 = \pi117 ^ w36628 ;
  assign w37146 = ( ~w36636 & w37144 ) | ( ~w36636 & w37145 ) | ( w37144 & w37145 ) ;
  assign w37147 = w37145 | w37146 ;
  assign w37148 = \pi118 ^ w36621 ;
  assign w37149 = ( ~w36629 & w37147 ) | ( ~w36629 & w37148 ) | ( w37147 & w37148 ) ;
  assign w37150 = w37148 | w37149 ;
  assign w37151 = \pi119 ^ w36614 ;
  assign w37152 = ( ~w36622 & w37150 ) | ( ~w36622 & w37151 ) | ( w37150 & w37151 ) ;
  assign w37153 = w37151 | w37152 ;
  assign w37154 = \pi120 ^ w36607 ;
  assign w37155 = ( ~w36615 & w37153 ) | ( ~w36615 & w37154 ) | ( w37153 & w37154 ) ;
  assign w37156 = w37154 | w37155 ;
  assign w37157 = \pi121 ^ w36600 ;
  assign w37158 = ( ~w36608 & w37156 ) | ( ~w36608 & w37157 ) | ( w37156 & w37157 ) ;
  assign w37159 = w37157 | w37158 ;
  assign w37160 = \pi122 ^ w36593 ;
  assign w37161 = ( ~w36601 & w37159 ) | ( ~w36601 & w37160 ) | ( w37159 & w37160 ) ;
  assign w37162 = w37160 | w37161 ;
  assign w37163 = w36578 | w36580 ;
  assign w37164 = ( ~w36057 & w36572 ) | ( ~w36057 & w36587 ) | ( w36572 & w36587 ) ;
  assign w37165 = w37163 ^ w37164 ;
  assign w37166 = ~w36587 & w37165 ;
  assign w37167 = ( w16707 & ~w36577 ) | ( w16707 & w36585 ) | ( ~w36577 & w36585 ) ;
  assign w37168 = w36577 & w37167 ;
  assign w37169 = w37166 | w37168 ;
  assign w37170 = ~\pi123 & w37169 ;
  assign w37171 = ( \pi123 & ~w37166 ) | ( \pi123 & w37168 ) | ( ~w37166 & w37168 ) ;
  assign w37172 = ~w37168 & w37171 ;
  assign w37173 = w37170 | w37172 ;
  assign w37174 = ( ~w36594 & w37162 ) | ( ~w36594 & w37173 ) | ( w37162 & w37173 ) ;
  assign w37175 = ( w147 & ~w37173 ) | ( w147 & w37174 ) | ( ~w37173 & w37174 ) ;
  assign w37176 = w37173 | w37175 ;
  assign w37177 = ( w269 & ~w270 ) | ( w269 & w37169 ) | ( ~w270 & w37169 ) ;
  assign w37178 = ~w269 & w37177 ;
  assign w37179 = w37176 & ~w37178 ;
  assign w37180 = ~w36601 & w37159 ;
  assign w37181 = w37160 ^ w37180 ;
  assign w37182 = ~w37179 & w37181 ;
  assign w37183 = ( w36593 & w37176 ) | ( w36593 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37184 = ~w37178 & w37183 ;
  assign w37185 = w37182 | w37184 ;
  assign w37186 = ~\pi123 & w37185 ;
  assign w37187 = ~w36608 & w37156 ;
  assign w37188 = w37157 ^ w37187 ;
  assign w37189 = ~w37179 & w37188 ;
  assign w37190 = ( w36600 & w37176 ) | ( w36600 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37191 = ~w37178 & w37190 ;
  assign w37192 = w37189 | w37191 ;
  assign w37193 = ~\pi122 & w37192 ;
  assign w37194 = ~w36615 & w37153 ;
  assign w37195 = w37154 ^ w37194 ;
  assign w37196 = ~w37179 & w37195 ;
  assign w37197 = ( w36607 & w37176 ) | ( w36607 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37198 = ~w37178 & w37197 ;
  assign w37199 = w37196 | w37198 ;
  assign w37200 = ~\pi121 & w37199 ;
  assign w37201 = ~w36622 & w37150 ;
  assign w37202 = w37151 ^ w37201 ;
  assign w37203 = ~w37179 & w37202 ;
  assign w37204 = ( w36614 & w37176 ) | ( w36614 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37205 = ~w37178 & w37204 ;
  assign w37206 = w37203 | w37205 ;
  assign w37207 = ~\pi120 & w37206 ;
  assign w37208 = ~w36629 & w37147 ;
  assign w37209 = w37148 ^ w37208 ;
  assign w37210 = ~w37179 & w37209 ;
  assign w37211 = ( w36621 & w37176 ) | ( w36621 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37212 = ~w37178 & w37211 ;
  assign w37213 = w37210 | w37212 ;
  assign w37214 = ~\pi119 & w37213 ;
  assign w37215 = ~w36636 & w37144 ;
  assign w37216 = w37145 ^ w37215 ;
  assign w37217 = ~w37179 & w37216 ;
  assign w37218 = ( w36628 & w37176 ) | ( w36628 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37219 = ~w37178 & w37218 ;
  assign w37220 = w37217 | w37219 ;
  assign w37221 = ~\pi118 & w37220 ;
  assign w37222 = ~w36643 & w37141 ;
  assign w37223 = w37142 ^ w37222 ;
  assign w37224 = ~w37179 & w37223 ;
  assign w37225 = ( w36635 & w37176 ) | ( w36635 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37226 = ~w37178 & w37225 ;
  assign w37227 = w37224 | w37226 ;
  assign w37228 = ~\pi117 & w37227 ;
  assign w37229 = ~w36650 & w37138 ;
  assign w37230 = w37139 ^ w37229 ;
  assign w37231 = ~w37179 & w37230 ;
  assign w37232 = ( w36642 & w37176 ) | ( w36642 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37233 = ~w37178 & w37232 ;
  assign w37234 = w37231 | w37233 ;
  assign w37235 = ~\pi116 & w37234 ;
  assign w37236 = ~w36657 & w37135 ;
  assign w37237 = w37136 ^ w37236 ;
  assign w37238 = ~w37179 & w37237 ;
  assign w37239 = ( w36649 & w37176 ) | ( w36649 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37240 = ~w37178 & w37239 ;
  assign w37241 = w37238 | w37240 ;
  assign w37242 = ~\pi115 & w37241 ;
  assign w37243 = ~w36664 & w37132 ;
  assign w37244 = w37133 ^ w37243 ;
  assign w37245 = ~w37179 & w37244 ;
  assign w37246 = ( w36656 & w37176 ) | ( w36656 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37247 = ~w37178 & w37246 ;
  assign w37248 = w37245 | w37247 ;
  assign w37249 = ~\pi114 & w37248 ;
  assign w37250 = ~w36671 & w37129 ;
  assign w37251 = w37130 ^ w37250 ;
  assign w37252 = ~w37179 & w37251 ;
  assign w37253 = ( w36663 & w37176 ) | ( w36663 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37254 = ~w37178 & w37253 ;
  assign w37255 = w37252 | w37254 ;
  assign w37256 = ~\pi113 & w37255 ;
  assign w37257 = ~w36678 & w37126 ;
  assign w37258 = w37127 ^ w37257 ;
  assign w37259 = ~w37179 & w37258 ;
  assign w37260 = ( w36670 & w37176 ) | ( w36670 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37261 = ~w37178 & w37260 ;
  assign w37262 = w37259 | w37261 ;
  assign w37263 = ~\pi112 & w37262 ;
  assign w37264 = ~w36685 & w37123 ;
  assign w37265 = w37124 ^ w37264 ;
  assign w37266 = ~w37179 & w37265 ;
  assign w37267 = ( w36677 & w37176 ) | ( w36677 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37268 = ~w37178 & w37267 ;
  assign w37269 = w37266 | w37268 ;
  assign w37270 = ~\pi111 & w37269 ;
  assign w37271 = ~w36692 & w37120 ;
  assign w37272 = w37121 ^ w37271 ;
  assign w37273 = ~w37179 & w37272 ;
  assign w37274 = ( w36684 & w37176 ) | ( w36684 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37275 = ~w37178 & w37274 ;
  assign w37276 = w37273 | w37275 ;
  assign w37277 = ~\pi110 & w37276 ;
  assign w37278 = ~w36699 & w37117 ;
  assign w37279 = w37118 ^ w37278 ;
  assign w37280 = ~w37179 & w37279 ;
  assign w37281 = ( w36691 & w37176 ) | ( w36691 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37282 = ~w37178 & w37281 ;
  assign w37283 = w37280 | w37282 ;
  assign w37284 = ~\pi109 & w37283 ;
  assign w37285 = ~w36706 & w37114 ;
  assign w37286 = w37115 ^ w37285 ;
  assign w37287 = ~w37179 & w37286 ;
  assign w37288 = ( w36698 & w37176 ) | ( w36698 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37289 = ~w37178 & w37288 ;
  assign w37290 = w37287 | w37289 ;
  assign w37291 = ~\pi108 & w37290 ;
  assign w37292 = ~w36713 & w37111 ;
  assign w37293 = w37112 ^ w37292 ;
  assign w37294 = ~w37179 & w37293 ;
  assign w37295 = ( w36705 & w37176 ) | ( w36705 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37296 = ~w37178 & w37295 ;
  assign w37297 = w37294 | w37296 ;
  assign w37298 = ~\pi107 & w37297 ;
  assign w37299 = ~w36720 & w37108 ;
  assign w37300 = w37109 ^ w37299 ;
  assign w37301 = ~w37179 & w37300 ;
  assign w37302 = ( w36712 & w37176 ) | ( w36712 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37303 = ~w37178 & w37302 ;
  assign w37304 = w37301 | w37303 ;
  assign w37305 = ~\pi106 & w37304 ;
  assign w37306 = ~w36727 & w37105 ;
  assign w37307 = w37106 ^ w37306 ;
  assign w37308 = ~w37179 & w37307 ;
  assign w37309 = ( w36719 & w37176 ) | ( w36719 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37310 = ~w37178 & w37309 ;
  assign w37311 = w37308 | w37310 ;
  assign w37312 = ~\pi105 & w37311 ;
  assign w37313 = ~w36734 & w37102 ;
  assign w37314 = w37103 ^ w37313 ;
  assign w37315 = ~w37179 & w37314 ;
  assign w37316 = ( w36726 & w37176 ) | ( w36726 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37317 = ~w37178 & w37316 ;
  assign w37318 = w37315 | w37317 ;
  assign w37319 = ~\pi104 & w37318 ;
  assign w37320 = ~w36741 & w37099 ;
  assign w37321 = w37100 ^ w37320 ;
  assign w37322 = ~w37179 & w37321 ;
  assign w37323 = ( w36733 & w37176 ) | ( w36733 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37324 = ~w37178 & w37323 ;
  assign w37325 = w37322 | w37324 ;
  assign w37326 = ~\pi103 & w37325 ;
  assign w37327 = ~w36748 & w37096 ;
  assign w37328 = w37097 ^ w37327 ;
  assign w37329 = ~w37179 & w37328 ;
  assign w37330 = ( w36740 & w37176 ) | ( w36740 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37331 = ~w37178 & w37330 ;
  assign w37332 = w37329 | w37331 ;
  assign w37333 = ~\pi102 & w37332 ;
  assign w37334 = ~w36755 & w37093 ;
  assign w37335 = w37094 ^ w37334 ;
  assign w37336 = ~w37179 & w37335 ;
  assign w37337 = ( w36747 & w37176 ) | ( w36747 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37338 = ~w37178 & w37337 ;
  assign w37339 = w37336 | w37338 ;
  assign w37340 = ~\pi101 & w37339 ;
  assign w37341 = ~w36762 & w37090 ;
  assign w37342 = w37091 ^ w37341 ;
  assign w37343 = ~w37179 & w37342 ;
  assign w37344 = ( w36754 & w37176 ) | ( w36754 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37345 = ~w37178 & w37344 ;
  assign w37346 = w37343 | w37345 ;
  assign w37347 = ~\pi100 & w37346 ;
  assign w37348 = ~w36769 & w37087 ;
  assign w37349 = w37088 ^ w37348 ;
  assign w37350 = ~w37179 & w37349 ;
  assign w37351 = ( w36761 & w37176 ) | ( w36761 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37352 = ~w37178 & w37351 ;
  assign w37353 = w37350 | w37352 ;
  assign w37354 = ~\pi099 & w37353 ;
  assign w37355 = ~w36776 & w37084 ;
  assign w37356 = w37085 ^ w37355 ;
  assign w37357 = ~w37179 & w37356 ;
  assign w37358 = ( w36768 & w37176 ) | ( w36768 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37359 = ~w37178 & w37358 ;
  assign w37360 = w37357 | w37359 ;
  assign w37361 = ~\pi098 & w37360 ;
  assign w37362 = ~w36783 & w37081 ;
  assign w37363 = w37082 ^ w37362 ;
  assign w37364 = ~w37179 & w37363 ;
  assign w37365 = ( w36775 & w37176 ) | ( w36775 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37366 = ~w37178 & w37365 ;
  assign w37367 = w37364 | w37366 ;
  assign w37368 = ~\pi097 & w37367 ;
  assign w37369 = ~w36790 & w37078 ;
  assign w37370 = w37079 ^ w37369 ;
  assign w37371 = ~w37179 & w37370 ;
  assign w37372 = ( w36782 & w37176 ) | ( w36782 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37373 = ~w37178 & w37372 ;
  assign w37374 = w37371 | w37373 ;
  assign w37375 = ~\pi096 & w37374 ;
  assign w37376 = ~w36797 & w37075 ;
  assign w37377 = w37076 ^ w37376 ;
  assign w37378 = ~w37179 & w37377 ;
  assign w37379 = ( w36789 & w37176 ) | ( w36789 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37380 = ~w37178 & w37379 ;
  assign w37381 = w37378 | w37380 ;
  assign w37382 = ~\pi095 & w37381 ;
  assign w37383 = ~w36804 & w37072 ;
  assign w37384 = w37073 ^ w37383 ;
  assign w37385 = ~w37179 & w37384 ;
  assign w37386 = ( w36796 & w37176 ) | ( w36796 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37387 = ~w37178 & w37386 ;
  assign w37388 = w37385 | w37387 ;
  assign w37389 = ~\pi094 & w37388 ;
  assign w37390 = ~w36811 & w37069 ;
  assign w37391 = w37070 ^ w37390 ;
  assign w37392 = ~w37179 & w37391 ;
  assign w37393 = ( w36803 & w37176 ) | ( w36803 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37394 = ~w37178 & w37393 ;
  assign w37395 = w37392 | w37394 ;
  assign w37396 = ~\pi093 & w37395 ;
  assign w37397 = ~w36818 & w37066 ;
  assign w37398 = w37067 ^ w37397 ;
  assign w37399 = ~w37179 & w37398 ;
  assign w37400 = ( w36810 & w37176 ) | ( w36810 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37401 = ~w37178 & w37400 ;
  assign w37402 = w37399 | w37401 ;
  assign w37403 = ~\pi092 & w37402 ;
  assign w37404 = ~w36825 & w37063 ;
  assign w37405 = w37064 ^ w37404 ;
  assign w37406 = ~w37179 & w37405 ;
  assign w37407 = ( w36817 & w37176 ) | ( w36817 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37408 = ~w37178 & w37407 ;
  assign w37409 = w37406 | w37408 ;
  assign w37410 = ~\pi091 & w37409 ;
  assign w37411 = ~w36832 & w37060 ;
  assign w37412 = w37061 ^ w37411 ;
  assign w37413 = ~w37179 & w37412 ;
  assign w37414 = ( w36824 & w37176 ) | ( w36824 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37415 = ~w37178 & w37414 ;
  assign w37416 = w37413 | w37415 ;
  assign w37417 = ~\pi090 & w37416 ;
  assign w37418 = ~w36839 & w37057 ;
  assign w37419 = w37058 ^ w37418 ;
  assign w37420 = ~w37179 & w37419 ;
  assign w37421 = ( w36831 & w37176 ) | ( w36831 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37422 = ~w37178 & w37421 ;
  assign w37423 = w37420 | w37422 ;
  assign w37424 = ~\pi089 & w37423 ;
  assign w37425 = ~w36846 & w37054 ;
  assign w37426 = w37055 ^ w37425 ;
  assign w37427 = ~w37179 & w37426 ;
  assign w37428 = ( w36838 & w37176 ) | ( w36838 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37429 = ~w37178 & w37428 ;
  assign w37430 = w37427 | w37429 ;
  assign w37431 = ~\pi088 & w37430 ;
  assign w37432 = ~w36853 & w37051 ;
  assign w37433 = w37052 ^ w37432 ;
  assign w37434 = ~w37179 & w37433 ;
  assign w37435 = ( w36845 & w37176 ) | ( w36845 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37436 = ~w37178 & w37435 ;
  assign w37437 = w37434 | w37436 ;
  assign w37438 = ~\pi087 & w37437 ;
  assign w37439 = ~w36860 & w37048 ;
  assign w37440 = w37049 ^ w37439 ;
  assign w37441 = ~w37179 & w37440 ;
  assign w37442 = ( w36852 & w37176 ) | ( w36852 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37443 = ~w37178 & w37442 ;
  assign w37444 = w37441 | w37443 ;
  assign w37445 = ~\pi086 & w37444 ;
  assign w37446 = ~w36867 & w37045 ;
  assign w37447 = w37046 ^ w37446 ;
  assign w37448 = ~w37179 & w37447 ;
  assign w37449 = ( w36859 & w37176 ) | ( w36859 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37450 = ~w37178 & w37449 ;
  assign w37451 = w37448 | w37450 ;
  assign w37452 = ~\pi085 & w37451 ;
  assign w37453 = ~w36874 & w37042 ;
  assign w37454 = w37043 ^ w37453 ;
  assign w37455 = ~w37179 & w37454 ;
  assign w37456 = ( w36866 & w37176 ) | ( w36866 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37457 = ~w37178 & w37456 ;
  assign w37458 = w37455 | w37457 ;
  assign w37459 = ~\pi084 & w37458 ;
  assign w37460 = ~w36881 & w37039 ;
  assign w37461 = w37040 ^ w37460 ;
  assign w37462 = ~w37179 & w37461 ;
  assign w37463 = ( w36873 & w37176 ) | ( w36873 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37464 = ~w37178 & w37463 ;
  assign w37465 = w37462 | w37464 ;
  assign w37466 = ~\pi083 & w37465 ;
  assign w37467 = ~w36888 & w37036 ;
  assign w37468 = w37037 ^ w37467 ;
  assign w37469 = ~w37179 & w37468 ;
  assign w37470 = ( w36880 & w37176 ) | ( w36880 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37471 = ~w37178 & w37470 ;
  assign w37472 = w37469 | w37471 ;
  assign w37473 = ~\pi082 & w37472 ;
  assign w37474 = ~w36895 & w37033 ;
  assign w37475 = w37034 ^ w37474 ;
  assign w37476 = ~w37179 & w37475 ;
  assign w37477 = ( w36887 & w37176 ) | ( w36887 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37478 = ~w37178 & w37477 ;
  assign w37479 = w37476 | w37478 ;
  assign w37480 = ~\pi081 & w37479 ;
  assign w37481 = ~w36902 & w37030 ;
  assign w37482 = w37031 ^ w37481 ;
  assign w37483 = ~w37179 & w37482 ;
  assign w37484 = ( w36894 & w37176 ) | ( w36894 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37485 = ~w37178 & w37484 ;
  assign w37486 = w37483 | w37485 ;
  assign w37487 = ~\pi080 & w37486 ;
  assign w37488 = ~w36909 & w37027 ;
  assign w37489 = w37028 ^ w37488 ;
  assign w37490 = ~w37179 & w37489 ;
  assign w37491 = ( w36901 & w37176 ) | ( w36901 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37492 = ~w37178 & w37491 ;
  assign w37493 = w37490 | w37492 ;
  assign w37494 = ~\pi079 & w37493 ;
  assign w37495 = ~w36916 & w37024 ;
  assign w37496 = w37025 ^ w37495 ;
  assign w37497 = ~w37179 & w37496 ;
  assign w37498 = ( w36908 & w37176 ) | ( w36908 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37499 = ~w37178 & w37498 ;
  assign w37500 = w37497 | w37499 ;
  assign w37501 = ~\pi078 & w37500 ;
  assign w37502 = ~w36923 & w37021 ;
  assign w37503 = w37022 ^ w37502 ;
  assign w37504 = ~w37179 & w37503 ;
  assign w37505 = ( w36915 & w37176 ) | ( w36915 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37506 = ~w37178 & w37505 ;
  assign w37507 = w37504 | w37506 ;
  assign w37508 = ~\pi077 & w37507 ;
  assign w37509 = ~w36930 & w37018 ;
  assign w37510 = w37019 ^ w37509 ;
  assign w37511 = ~w37179 & w37510 ;
  assign w37512 = ( w36922 & w37176 ) | ( w36922 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37513 = ~w37178 & w37512 ;
  assign w37514 = w37511 | w37513 ;
  assign w37515 = ~\pi076 & w37514 ;
  assign w37516 = ~w36937 & w37015 ;
  assign w37517 = w37016 ^ w37516 ;
  assign w37518 = ~w37179 & w37517 ;
  assign w37519 = ( w36929 & w37176 ) | ( w36929 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37520 = ~w37178 & w37519 ;
  assign w37521 = w37518 | w37520 ;
  assign w37522 = ~\pi075 & w37521 ;
  assign w37523 = ~w36944 & w37012 ;
  assign w37524 = w37013 ^ w37523 ;
  assign w37525 = ~w37179 & w37524 ;
  assign w37526 = ( w36936 & w37176 ) | ( w36936 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37527 = ~w37178 & w37526 ;
  assign w37528 = w37525 | w37527 ;
  assign w37529 = ~\pi074 & w37528 ;
  assign w37530 = ~w36951 & w37009 ;
  assign w37531 = w37010 ^ w37530 ;
  assign w37532 = ~w37179 & w37531 ;
  assign w37533 = ( w36943 & w37176 ) | ( w36943 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37534 = ~w37178 & w37533 ;
  assign w37535 = w37532 | w37534 ;
  assign w37536 = ~\pi073 & w37535 ;
  assign w37537 = ~w36958 & w37006 ;
  assign w37538 = w37007 ^ w37537 ;
  assign w37539 = ~w37179 & w37538 ;
  assign w37540 = ( w36950 & w37176 ) | ( w36950 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37541 = ~w37178 & w37540 ;
  assign w37542 = w37539 | w37541 ;
  assign w37543 = ~\pi072 & w37542 ;
  assign w37544 = ~w36965 & w37003 ;
  assign w37545 = w37004 ^ w37544 ;
  assign w37546 = ~w37179 & w37545 ;
  assign w37547 = ( w36957 & w37176 ) | ( w36957 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37548 = ~w37178 & w37547 ;
  assign w37549 = w37546 | w37548 ;
  assign w37550 = ~\pi071 & w37549 ;
  assign w37551 = ~w36972 & w37000 ;
  assign w37552 = w37001 ^ w37551 ;
  assign w37553 = ~w37179 & w37552 ;
  assign w37554 = ( w36964 & w37176 ) | ( w36964 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37555 = ~w37178 & w37554 ;
  assign w37556 = w37553 | w37555 ;
  assign w37557 = ~\pi070 & w37556 ;
  assign w37558 = ~w36978 & w36997 ;
  assign w37559 = w36998 ^ w37558 ;
  assign w37560 = ~w37179 & w37559 ;
  assign w37561 = ( w36971 & w37176 ) | ( w36971 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37562 = ~w37178 & w37561 ;
  assign w37563 = w37560 | w37562 ;
  assign w37564 = ~\pi069 & w37563 ;
  assign w37565 = ~w36986 & w36994 ;
  assign w37566 = w36995 ^ w37565 ;
  assign w37567 = ~w37179 & w37566 ;
  assign w37568 = ( w36977 & w37176 ) | ( w36977 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37569 = ~w37178 & w37568 ;
  assign w37570 = w37567 | w37569 ;
  assign w37571 = ~\pi068 & w37570 ;
  assign w37572 = \pi064 & ~w36587 ;
  assign w37573 = \pi005 ^ w37572 ;
  assign w37574 = ( \pi065 & w18236 ) | ( \pi065 & ~w37573 ) | ( w18236 & ~w37573 ) ;
  assign w37575 = w36990 ^ w37574 ;
  assign w37576 = ~w37179 & w37575 ;
  assign w37577 = ( w36985 & w37176 ) | ( w36985 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37578 = ~w37178 & w37577 ;
  assign w37579 = w37576 | w37578 ;
  assign w37580 = ~\pi067 & w37579 ;
  assign w37581 = \pi004 ^ w36587 ;
  assign w37582 = ( \pi064 & w37179 ) | ( \pi064 & w37581 ) | ( w37179 & w37581 ) ;
  assign w37583 = w18244 ^ w37582 ;
  assign w37584 = ~w37179 & w37583 ;
  assign w37585 = w37179 & w37573 ;
  assign w37586 = w37584 | w37585 ;
  assign w37587 = ~\pi066 & w37586 ;
  assign w37588 = \pi066 ^ w37586 ;
  assign w37589 = ( \pi064 & ~w37179 ) | ( \pi064 & w37588 ) | ( ~w37179 & w37588 ) ;
  assign w37590 = \pi004 ^ w37589 ;
  assign w37591 = ( \pi065 & w18843 ) | ( \pi065 & ~w37590 ) | ( w18843 & ~w37590 ) ;
  assign w37592 = w37588 | w37591 ;
  assign w37593 = \pi067 ^ w37579 ;
  assign w37594 = ( ~w37587 & w37592 ) | ( ~w37587 & w37593 ) | ( w37592 & w37593 ) ;
  assign w37595 = w37593 | w37594 ;
  assign w37596 = \pi068 ^ w37570 ;
  assign w37597 = ( ~w37580 & w37595 ) | ( ~w37580 & w37596 ) | ( w37595 & w37596 ) ;
  assign w37598 = w37596 | w37597 ;
  assign w37599 = \pi069 ^ w37563 ;
  assign w37600 = ( ~w37571 & w37598 ) | ( ~w37571 & w37599 ) | ( w37598 & w37599 ) ;
  assign w37601 = w37599 | w37600 ;
  assign w37602 = \pi070 ^ w37556 ;
  assign w37603 = ( ~w37564 & w37601 ) | ( ~w37564 & w37602 ) | ( w37601 & w37602 ) ;
  assign w37604 = w37602 | w37603 ;
  assign w37605 = \pi071 ^ w37549 ;
  assign w37606 = ( ~w37557 & w37604 ) | ( ~w37557 & w37605 ) | ( w37604 & w37605 ) ;
  assign w37607 = w37605 | w37606 ;
  assign w37608 = \pi072 ^ w37542 ;
  assign w37609 = ( ~w37550 & w37607 ) | ( ~w37550 & w37608 ) | ( w37607 & w37608 ) ;
  assign w37610 = w37608 | w37609 ;
  assign w37611 = \pi073 ^ w37535 ;
  assign w37612 = ( ~w37543 & w37610 ) | ( ~w37543 & w37611 ) | ( w37610 & w37611 ) ;
  assign w37613 = w37611 | w37612 ;
  assign w37614 = \pi074 ^ w37528 ;
  assign w37615 = ( ~w37536 & w37613 ) | ( ~w37536 & w37614 ) | ( w37613 & w37614 ) ;
  assign w37616 = w37614 | w37615 ;
  assign w37617 = \pi075 ^ w37521 ;
  assign w37618 = ( ~w37529 & w37616 ) | ( ~w37529 & w37617 ) | ( w37616 & w37617 ) ;
  assign w37619 = w37617 | w37618 ;
  assign w37620 = \pi076 ^ w37514 ;
  assign w37621 = ( ~w37522 & w37619 ) | ( ~w37522 & w37620 ) | ( w37619 & w37620 ) ;
  assign w37622 = w37620 | w37621 ;
  assign w37623 = \pi077 ^ w37507 ;
  assign w37624 = ( ~w37515 & w37622 ) | ( ~w37515 & w37623 ) | ( w37622 & w37623 ) ;
  assign w37625 = w37623 | w37624 ;
  assign w37626 = \pi078 ^ w37500 ;
  assign w37627 = ( ~w37508 & w37625 ) | ( ~w37508 & w37626 ) | ( w37625 & w37626 ) ;
  assign w37628 = w37626 | w37627 ;
  assign w37629 = \pi079 ^ w37493 ;
  assign w37630 = ( ~w37501 & w37628 ) | ( ~w37501 & w37629 ) | ( w37628 & w37629 ) ;
  assign w37631 = w37629 | w37630 ;
  assign w37632 = \pi080 ^ w37486 ;
  assign w37633 = ( ~w37494 & w37631 ) | ( ~w37494 & w37632 ) | ( w37631 & w37632 ) ;
  assign w37634 = w37632 | w37633 ;
  assign w37635 = \pi081 ^ w37479 ;
  assign w37636 = ( ~w37487 & w37634 ) | ( ~w37487 & w37635 ) | ( w37634 & w37635 ) ;
  assign w37637 = w37635 | w37636 ;
  assign w37638 = \pi082 ^ w37472 ;
  assign w37639 = ( ~w37480 & w37637 ) | ( ~w37480 & w37638 ) | ( w37637 & w37638 ) ;
  assign w37640 = w37638 | w37639 ;
  assign w37641 = \pi083 ^ w37465 ;
  assign w37642 = ( ~w37473 & w37640 ) | ( ~w37473 & w37641 ) | ( w37640 & w37641 ) ;
  assign w37643 = w37641 | w37642 ;
  assign w37644 = \pi084 ^ w37458 ;
  assign w37645 = ( ~w37466 & w37643 ) | ( ~w37466 & w37644 ) | ( w37643 & w37644 ) ;
  assign w37646 = w37644 | w37645 ;
  assign w37647 = \pi085 ^ w37451 ;
  assign w37648 = ( ~w37459 & w37646 ) | ( ~w37459 & w37647 ) | ( w37646 & w37647 ) ;
  assign w37649 = w37647 | w37648 ;
  assign w37650 = \pi086 ^ w37444 ;
  assign w37651 = ( ~w37452 & w37649 ) | ( ~w37452 & w37650 ) | ( w37649 & w37650 ) ;
  assign w37652 = w37650 | w37651 ;
  assign w37653 = \pi087 ^ w37437 ;
  assign w37654 = ( ~w37445 & w37652 ) | ( ~w37445 & w37653 ) | ( w37652 & w37653 ) ;
  assign w37655 = w37653 | w37654 ;
  assign w37656 = \pi088 ^ w37430 ;
  assign w37657 = ( ~w37438 & w37655 ) | ( ~w37438 & w37656 ) | ( w37655 & w37656 ) ;
  assign w37658 = w37656 | w37657 ;
  assign w37659 = \pi089 ^ w37423 ;
  assign w37660 = ( ~w37431 & w37658 ) | ( ~w37431 & w37659 ) | ( w37658 & w37659 ) ;
  assign w37661 = w37659 | w37660 ;
  assign w37662 = \pi090 ^ w37416 ;
  assign w37663 = ( ~w37424 & w37661 ) | ( ~w37424 & w37662 ) | ( w37661 & w37662 ) ;
  assign w37664 = w37662 | w37663 ;
  assign w37665 = \pi091 ^ w37409 ;
  assign w37666 = ( ~w37417 & w37664 ) | ( ~w37417 & w37665 ) | ( w37664 & w37665 ) ;
  assign w37667 = w37665 | w37666 ;
  assign w37668 = \pi092 ^ w37402 ;
  assign w37669 = ( ~w37410 & w37667 ) | ( ~w37410 & w37668 ) | ( w37667 & w37668 ) ;
  assign w37670 = w37668 | w37669 ;
  assign w37671 = \pi093 ^ w37395 ;
  assign w37672 = ( ~w37403 & w37670 ) | ( ~w37403 & w37671 ) | ( w37670 & w37671 ) ;
  assign w37673 = w37671 | w37672 ;
  assign w37674 = \pi094 ^ w37388 ;
  assign w37675 = ( ~w37396 & w37673 ) | ( ~w37396 & w37674 ) | ( w37673 & w37674 ) ;
  assign w37676 = w37674 | w37675 ;
  assign w37677 = \pi095 ^ w37381 ;
  assign w37678 = ( ~w37389 & w37676 ) | ( ~w37389 & w37677 ) | ( w37676 & w37677 ) ;
  assign w37679 = w37677 | w37678 ;
  assign w37680 = \pi096 ^ w37374 ;
  assign w37681 = ( ~w37382 & w37679 ) | ( ~w37382 & w37680 ) | ( w37679 & w37680 ) ;
  assign w37682 = w37680 | w37681 ;
  assign w37683 = \pi097 ^ w37367 ;
  assign w37684 = ( ~w37375 & w37682 ) | ( ~w37375 & w37683 ) | ( w37682 & w37683 ) ;
  assign w37685 = w37683 | w37684 ;
  assign w37686 = \pi098 ^ w37360 ;
  assign w37687 = ( ~w37368 & w37685 ) | ( ~w37368 & w37686 ) | ( w37685 & w37686 ) ;
  assign w37688 = w37686 | w37687 ;
  assign w37689 = \pi099 ^ w37353 ;
  assign w37690 = ( ~w37361 & w37688 ) | ( ~w37361 & w37689 ) | ( w37688 & w37689 ) ;
  assign w37691 = w37689 | w37690 ;
  assign w37692 = \pi100 ^ w37346 ;
  assign w37693 = ( ~w37354 & w37691 ) | ( ~w37354 & w37692 ) | ( w37691 & w37692 ) ;
  assign w37694 = w37692 | w37693 ;
  assign w37695 = \pi101 ^ w37339 ;
  assign w37696 = ( ~w37347 & w37694 ) | ( ~w37347 & w37695 ) | ( w37694 & w37695 ) ;
  assign w37697 = w37695 | w37696 ;
  assign w37698 = \pi102 ^ w37332 ;
  assign w37699 = ( ~w37340 & w37697 ) | ( ~w37340 & w37698 ) | ( w37697 & w37698 ) ;
  assign w37700 = w37698 | w37699 ;
  assign w37701 = \pi103 ^ w37325 ;
  assign w37702 = ( ~w37333 & w37700 ) | ( ~w37333 & w37701 ) | ( w37700 & w37701 ) ;
  assign w37703 = w37701 | w37702 ;
  assign w37704 = \pi104 ^ w37318 ;
  assign w37705 = ( ~w37326 & w37703 ) | ( ~w37326 & w37704 ) | ( w37703 & w37704 ) ;
  assign w37706 = w37704 | w37705 ;
  assign w37707 = \pi105 ^ w37311 ;
  assign w37708 = ( ~w37319 & w37706 ) | ( ~w37319 & w37707 ) | ( w37706 & w37707 ) ;
  assign w37709 = w37707 | w37708 ;
  assign w37710 = \pi106 ^ w37304 ;
  assign w37711 = ( ~w37312 & w37709 ) | ( ~w37312 & w37710 ) | ( w37709 & w37710 ) ;
  assign w37712 = w37710 | w37711 ;
  assign w37713 = \pi107 ^ w37297 ;
  assign w37714 = ( ~w37305 & w37712 ) | ( ~w37305 & w37713 ) | ( w37712 & w37713 ) ;
  assign w37715 = w37713 | w37714 ;
  assign w37716 = \pi108 ^ w37290 ;
  assign w37717 = ( ~w37298 & w37715 ) | ( ~w37298 & w37716 ) | ( w37715 & w37716 ) ;
  assign w37718 = w37716 | w37717 ;
  assign w37719 = \pi109 ^ w37283 ;
  assign w37720 = ( ~w37291 & w37718 ) | ( ~w37291 & w37719 ) | ( w37718 & w37719 ) ;
  assign w37721 = w37719 | w37720 ;
  assign w37722 = \pi110 ^ w37276 ;
  assign w37723 = ( ~w37284 & w37721 ) | ( ~w37284 & w37722 ) | ( w37721 & w37722 ) ;
  assign w37724 = w37722 | w37723 ;
  assign w37725 = \pi111 ^ w37269 ;
  assign w37726 = ( ~w37277 & w37724 ) | ( ~w37277 & w37725 ) | ( w37724 & w37725 ) ;
  assign w37727 = w37725 | w37726 ;
  assign w37728 = \pi112 ^ w37262 ;
  assign w37729 = ( ~w37270 & w37727 ) | ( ~w37270 & w37728 ) | ( w37727 & w37728 ) ;
  assign w37730 = w37728 | w37729 ;
  assign w37731 = \pi113 ^ w37255 ;
  assign w37732 = ( ~w37263 & w37730 ) | ( ~w37263 & w37731 ) | ( w37730 & w37731 ) ;
  assign w37733 = w37731 | w37732 ;
  assign w37734 = \pi114 ^ w37248 ;
  assign w37735 = ( ~w37256 & w37733 ) | ( ~w37256 & w37734 ) | ( w37733 & w37734 ) ;
  assign w37736 = w37734 | w37735 ;
  assign w37737 = \pi115 ^ w37241 ;
  assign w37738 = ( ~w37249 & w37736 ) | ( ~w37249 & w37737 ) | ( w37736 & w37737 ) ;
  assign w37739 = w37737 | w37738 ;
  assign w37740 = \pi116 ^ w37234 ;
  assign w37741 = ( ~w37242 & w37739 ) | ( ~w37242 & w37740 ) | ( w37739 & w37740 ) ;
  assign w37742 = w37740 | w37741 ;
  assign w37743 = \pi117 ^ w37227 ;
  assign w37744 = ( ~w37235 & w37742 ) | ( ~w37235 & w37743 ) | ( w37742 & w37743 ) ;
  assign w37745 = w37743 | w37744 ;
  assign w37746 = \pi118 ^ w37220 ;
  assign w37747 = ( ~w37228 & w37745 ) | ( ~w37228 & w37746 ) | ( w37745 & w37746 ) ;
  assign w37748 = w37746 | w37747 ;
  assign w37749 = \pi119 ^ w37213 ;
  assign w37750 = ( ~w37221 & w37748 ) | ( ~w37221 & w37749 ) | ( w37748 & w37749 ) ;
  assign w37751 = w37749 | w37750 ;
  assign w37752 = \pi120 ^ w37206 ;
  assign w37753 = ( ~w37214 & w37751 ) | ( ~w37214 & w37752 ) | ( w37751 & w37752 ) ;
  assign w37754 = w37752 | w37753 ;
  assign w37755 = \pi121 ^ w37199 ;
  assign w37756 = ( ~w37207 & w37754 ) | ( ~w37207 & w37755 ) | ( w37754 & w37755 ) ;
  assign w37757 = w37755 | w37756 ;
  assign w37758 = \pi122 ^ w37192 ;
  assign w37759 = ( ~w37200 & w37757 ) | ( ~w37200 & w37758 ) | ( w37757 & w37758 ) ;
  assign w37760 = w37758 | w37759 ;
  assign w37761 = \pi123 ^ w37185 ;
  assign w37762 = ( ~w37193 & w37760 ) | ( ~w37193 & w37761 ) | ( w37760 & w37761 ) ;
  assign w37763 = w37761 | w37762 ;
  assign w37764 = ( ~w36594 & w37162 ) | ( ~w36594 & w37179 ) | ( w37162 & w37179 ) ;
  assign w37765 = w37173 ^ w37764 ;
  assign w37766 = ~w37179 & w37765 ;
  assign w37767 = ( w37169 & w37176 ) | ( w37169 & w37178 ) | ( w37176 & w37178 ) ;
  assign w37768 = ~w37178 & w37767 ;
  assign w37769 = w37766 | w37768 ;
  assign w37770 = ~\pi124 & w37769 ;
  assign w37771 = ( \pi124 & ~w37766 ) | ( \pi124 & w37768 ) | ( ~w37766 & w37768 ) ;
  assign w37772 = ~w37768 & w37771 ;
  assign w37773 = w37770 | w37772 ;
  assign w37774 = ( ~w37186 & w37763 ) | ( ~w37186 & w37773 ) | ( w37763 & w37773 ) ;
  assign w37775 = ( w269 & ~w37773 ) | ( w269 & w37774 ) | ( ~w37773 & w37774 ) ;
  assign w37776 = w37773 | w37775 ;
  assign w37777 = ~w147 & w37769 ;
  assign w37778 = w37776 & ~w37777 ;
  assign w37779 = ~w37193 & w37760 ;
  assign w37780 = w37761 ^ w37779 ;
  assign w37781 = ~w37778 & w37780 ;
  assign w37782 = ( w37185 & w37776 ) | ( w37185 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37783 = ~w37777 & w37782 ;
  assign w37784 = w37781 | w37783 ;
  assign w37785 = ~\pi124 & w37784 ;
  assign w37786 = ~w37200 & w37757 ;
  assign w37787 = w37758 ^ w37786 ;
  assign w37788 = ~w37778 & w37787 ;
  assign w37789 = ( w37192 & w37776 ) | ( w37192 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37790 = ~w37777 & w37789 ;
  assign w37791 = w37788 | w37790 ;
  assign w37792 = ~\pi123 & w37791 ;
  assign w37793 = ~w37207 & w37754 ;
  assign w37794 = w37755 ^ w37793 ;
  assign w37795 = ~w37778 & w37794 ;
  assign w37796 = ( w37199 & w37776 ) | ( w37199 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37797 = ~w37777 & w37796 ;
  assign w37798 = w37795 | w37797 ;
  assign w37799 = ~\pi122 & w37798 ;
  assign w37800 = ~w37214 & w37751 ;
  assign w37801 = w37752 ^ w37800 ;
  assign w37802 = ~w37778 & w37801 ;
  assign w37803 = ( w37206 & w37776 ) | ( w37206 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37804 = ~w37777 & w37803 ;
  assign w37805 = w37802 | w37804 ;
  assign w37806 = ~\pi121 & w37805 ;
  assign w37807 = ~w37221 & w37748 ;
  assign w37808 = w37749 ^ w37807 ;
  assign w37809 = ~w37778 & w37808 ;
  assign w37810 = ( w37213 & w37776 ) | ( w37213 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37811 = ~w37777 & w37810 ;
  assign w37812 = w37809 | w37811 ;
  assign w37813 = ~\pi120 & w37812 ;
  assign w37814 = ~w37228 & w37745 ;
  assign w37815 = w37746 ^ w37814 ;
  assign w37816 = ~w37778 & w37815 ;
  assign w37817 = ( w37220 & w37776 ) | ( w37220 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37818 = ~w37777 & w37817 ;
  assign w37819 = w37816 | w37818 ;
  assign w37820 = ~\pi119 & w37819 ;
  assign w37821 = ~w37235 & w37742 ;
  assign w37822 = w37743 ^ w37821 ;
  assign w37823 = ~w37778 & w37822 ;
  assign w37824 = ( w37227 & w37776 ) | ( w37227 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37825 = ~w37777 & w37824 ;
  assign w37826 = w37823 | w37825 ;
  assign w37827 = ~\pi118 & w37826 ;
  assign w37828 = ~w37242 & w37739 ;
  assign w37829 = w37740 ^ w37828 ;
  assign w37830 = ~w37778 & w37829 ;
  assign w37831 = ( w37234 & w37776 ) | ( w37234 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37832 = ~w37777 & w37831 ;
  assign w37833 = w37830 | w37832 ;
  assign w37834 = ~\pi117 & w37833 ;
  assign w37835 = ~w37249 & w37736 ;
  assign w37836 = w37737 ^ w37835 ;
  assign w37837 = ~w37778 & w37836 ;
  assign w37838 = ( w37241 & w37776 ) | ( w37241 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37839 = ~w37777 & w37838 ;
  assign w37840 = w37837 | w37839 ;
  assign w37841 = ~\pi116 & w37840 ;
  assign w37842 = ~w37256 & w37733 ;
  assign w37843 = w37734 ^ w37842 ;
  assign w37844 = ~w37778 & w37843 ;
  assign w37845 = ( w37248 & w37776 ) | ( w37248 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37846 = ~w37777 & w37845 ;
  assign w37847 = w37844 | w37846 ;
  assign w37848 = ~\pi115 & w37847 ;
  assign w37849 = ~w37263 & w37730 ;
  assign w37850 = w37731 ^ w37849 ;
  assign w37851 = ~w37778 & w37850 ;
  assign w37852 = ( w37255 & w37776 ) | ( w37255 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37853 = ~w37777 & w37852 ;
  assign w37854 = w37851 | w37853 ;
  assign w37855 = ~\pi114 & w37854 ;
  assign w37856 = ~w37270 & w37727 ;
  assign w37857 = w37728 ^ w37856 ;
  assign w37858 = ~w37778 & w37857 ;
  assign w37859 = ( w37262 & w37776 ) | ( w37262 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37860 = ~w37777 & w37859 ;
  assign w37861 = w37858 | w37860 ;
  assign w37862 = ~\pi113 & w37861 ;
  assign w37863 = ~w37277 & w37724 ;
  assign w37864 = w37725 ^ w37863 ;
  assign w37865 = ~w37778 & w37864 ;
  assign w37866 = ( w37269 & w37776 ) | ( w37269 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37867 = ~w37777 & w37866 ;
  assign w37868 = w37865 | w37867 ;
  assign w37869 = ~\pi112 & w37868 ;
  assign w37870 = ~w37284 & w37721 ;
  assign w37871 = w37722 ^ w37870 ;
  assign w37872 = ~w37778 & w37871 ;
  assign w37873 = ( w37276 & w37776 ) | ( w37276 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37874 = ~w37777 & w37873 ;
  assign w37875 = w37872 | w37874 ;
  assign w37876 = ~\pi111 & w37875 ;
  assign w37877 = ~w37291 & w37718 ;
  assign w37878 = w37719 ^ w37877 ;
  assign w37879 = ~w37778 & w37878 ;
  assign w37880 = ( w37283 & w37776 ) | ( w37283 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37881 = ~w37777 & w37880 ;
  assign w37882 = w37879 | w37881 ;
  assign w37883 = ~\pi110 & w37882 ;
  assign w37884 = ~w37298 & w37715 ;
  assign w37885 = w37716 ^ w37884 ;
  assign w37886 = ~w37778 & w37885 ;
  assign w37887 = ( w37290 & w37776 ) | ( w37290 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37888 = ~w37777 & w37887 ;
  assign w37889 = w37886 | w37888 ;
  assign w37890 = ~\pi109 & w37889 ;
  assign w37891 = ~w37305 & w37712 ;
  assign w37892 = w37713 ^ w37891 ;
  assign w37893 = ~w37778 & w37892 ;
  assign w37894 = ( w37297 & w37776 ) | ( w37297 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37895 = ~w37777 & w37894 ;
  assign w37896 = w37893 | w37895 ;
  assign w37897 = ~\pi108 & w37896 ;
  assign w37898 = ~w37312 & w37709 ;
  assign w37899 = w37710 ^ w37898 ;
  assign w37900 = ~w37778 & w37899 ;
  assign w37901 = ( w37304 & w37776 ) | ( w37304 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37902 = ~w37777 & w37901 ;
  assign w37903 = w37900 | w37902 ;
  assign w37904 = ~\pi107 & w37903 ;
  assign w37905 = ~w37319 & w37706 ;
  assign w37906 = w37707 ^ w37905 ;
  assign w37907 = ~w37778 & w37906 ;
  assign w37908 = ( w37311 & w37776 ) | ( w37311 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37909 = ~w37777 & w37908 ;
  assign w37910 = w37907 | w37909 ;
  assign w37911 = ~\pi106 & w37910 ;
  assign w37912 = ~w37326 & w37703 ;
  assign w37913 = w37704 ^ w37912 ;
  assign w37914 = ~w37778 & w37913 ;
  assign w37915 = ( w37318 & w37776 ) | ( w37318 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37916 = ~w37777 & w37915 ;
  assign w37917 = w37914 | w37916 ;
  assign w37918 = ~\pi105 & w37917 ;
  assign w37919 = ~w37333 & w37700 ;
  assign w37920 = w37701 ^ w37919 ;
  assign w37921 = ~w37778 & w37920 ;
  assign w37922 = ( w37325 & w37776 ) | ( w37325 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37923 = ~w37777 & w37922 ;
  assign w37924 = w37921 | w37923 ;
  assign w37925 = ~\pi104 & w37924 ;
  assign w37926 = ~w37340 & w37697 ;
  assign w37927 = w37698 ^ w37926 ;
  assign w37928 = ~w37778 & w37927 ;
  assign w37929 = ( w37332 & w37776 ) | ( w37332 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37930 = ~w37777 & w37929 ;
  assign w37931 = w37928 | w37930 ;
  assign w37932 = ~\pi103 & w37931 ;
  assign w37933 = ~w37347 & w37694 ;
  assign w37934 = w37695 ^ w37933 ;
  assign w37935 = ~w37778 & w37934 ;
  assign w37936 = ( w37339 & w37776 ) | ( w37339 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37937 = ~w37777 & w37936 ;
  assign w37938 = w37935 | w37937 ;
  assign w37939 = ~\pi102 & w37938 ;
  assign w37940 = ~w37354 & w37691 ;
  assign w37941 = w37692 ^ w37940 ;
  assign w37942 = ~w37778 & w37941 ;
  assign w37943 = ( w37346 & w37776 ) | ( w37346 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37944 = ~w37777 & w37943 ;
  assign w37945 = w37942 | w37944 ;
  assign w37946 = ~\pi101 & w37945 ;
  assign w37947 = ~w37361 & w37688 ;
  assign w37948 = w37689 ^ w37947 ;
  assign w37949 = ~w37778 & w37948 ;
  assign w37950 = ( w37353 & w37776 ) | ( w37353 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37951 = ~w37777 & w37950 ;
  assign w37952 = w37949 | w37951 ;
  assign w37953 = ~\pi100 & w37952 ;
  assign w37954 = ~w37368 & w37685 ;
  assign w37955 = w37686 ^ w37954 ;
  assign w37956 = ~w37778 & w37955 ;
  assign w37957 = ( w37360 & w37776 ) | ( w37360 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37958 = ~w37777 & w37957 ;
  assign w37959 = w37956 | w37958 ;
  assign w37960 = ~\pi099 & w37959 ;
  assign w37961 = ~w37375 & w37682 ;
  assign w37962 = w37683 ^ w37961 ;
  assign w37963 = ~w37778 & w37962 ;
  assign w37964 = ( w37367 & w37776 ) | ( w37367 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37965 = ~w37777 & w37964 ;
  assign w37966 = w37963 | w37965 ;
  assign w37967 = ~\pi098 & w37966 ;
  assign w37968 = ~w37382 & w37679 ;
  assign w37969 = w37680 ^ w37968 ;
  assign w37970 = ~w37778 & w37969 ;
  assign w37971 = ( w37374 & w37776 ) | ( w37374 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37972 = ~w37777 & w37971 ;
  assign w37973 = w37970 | w37972 ;
  assign w37974 = ~\pi097 & w37973 ;
  assign w37975 = ~w37389 & w37676 ;
  assign w37976 = w37677 ^ w37975 ;
  assign w37977 = ~w37778 & w37976 ;
  assign w37978 = ( w37381 & w37776 ) | ( w37381 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37979 = ~w37777 & w37978 ;
  assign w37980 = w37977 | w37979 ;
  assign w37981 = ~\pi096 & w37980 ;
  assign w37982 = ~w37396 & w37673 ;
  assign w37983 = w37674 ^ w37982 ;
  assign w37984 = ~w37778 & w37983 ;
  assign w37985 = ( w37388 & w37776 ) | ( w37388 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37986 = ~w37777 & w37985 ;
  assign w37987 = w37984 | w37986 ;
  assign w37988 = ~\pi095 & w37987 ;
  assign w37989 = ~w37403 & w37670 ;
  assign w37990 = w37671 ^ w37989 ;
  assign w37991 = ~w37778 & w37990 ;
  assign w37992 = ( w37395 & w37776 ) | ( w37395 & w37777 ) | ( w37776 & w37777 ) ;
  assign w37993 = ~w37777 & w37992 ;
  assign w37994 = w37991 | w37993 ;
  assign w37995 = ~\pi094 & w37994 ;
  assign w37996 = ~w37410 & w37667 ;
  assign w37997 = w37668 ^ w37996 ;
  assign w37998 = ~w37778 & w37997 ;
  assign w37999 = ( w37402 & w37776 ) | ( w37402 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38000 = ~w37777 & w37999 ;
  assign w38001 = w37998 | w38000 ;
  assign w38002 = ~\pi093 & w38001 ;
  assign w38003 = ~w37417 & w37664 ;
  assign w38004 = w37665 ^ w38003 ;
  assign w38005 = ~w37778 & w38004 ;
  assign w38006 = ( w37409 & w37776 ) | ( w37409 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38007 = ~w37777 & w38006 ;
  assign w38008 = w38005 | w38007 ;
  assign w38009 = ~\pi092 & w38008 ;
  assign w38010 = ~w37424 & w37661 ;
  assign w38011 = w37662 ^ w38010 ;
  assign w38012 = ~w37778 & w38011 ;
  assign w38013 = ( w37416 & w37776 ) | ( w37416 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38014 = ~w37777 & w38013 ;
  assign w38015 = w38012 | w38014 ;
  assign w38016 = ~\pi091 & w38015 ;
  assign w38017 = ~w37431 & w37658 ;
  assign w38018 = w37659 ^ w38017 ;
  assign w38019 = ~w37778 & w38018 ;
  assign w38020 = ( w37423 & w37776 ) | ( w37423 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38021 = ~w37777 & w38020 ;
  assign w38022 = w38019 | w38021 ;
  assign w38023 = ~\pi090 & w38022 ;
  assign w38024 = ~w37438 & w37655 ;
  assign w38025 = w37656 ^ w38024 ;
  assign w38026 = ~w37778 & w38025 ;
  assign w38027 = ( w37430 & w37776 ) | ( w37430 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38028 = ~w37777 & w38027 ;
  assign w38029 = w38026 | w38028 ;
  assign w38030 = ~\pi089 & w38029 ;
  assign w38031 = ~w37445 & w37652 ;
  assign w38032 = w37653 ^ w38031 ;
  assign w38033 = ~w37778 & w38032 ;
  assign w38034 = ( w37437 & w37776 ) | ( w37437 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38035 = ~w37777 & w38034 ;
  assign w38036 = w38033 | w38035 ;
  assign w38037 = ~\pi088 & w38036 ;
  assign w38038 = ~w37452 & w37649 ;
  assign w38039 = w37650 ^ w38038 ;
  assign w38040 = ~w37778 & w38039 ;
  assign w38041 = ( w37444 & w37776 ) | ( w37444 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38042 = ~w37777 & w38041 ;
  assign w38043 = w38040 | w38042 ;
  assign w38044 = ~\pi087 & w38043 ;
  assign w38045 = ~w37459 & w37646 ;
  assign w38046 = w37647 ^ w38045 ;
  assign w38047 = ~w37778 & w38046 ;
  assign w38048 = ( w37451 & w37776 ) | ( w37451 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38049 = ~w37777 & w38048 ;
  assign w38050 = w38047 | w38049 ;
  assign w38051 = ~\pi086 & w38050 ;
  assign w38052 = ~w37466 & w37643 ;
  assign w38053 = w37644 ^ w38052 ;
  assign w38054 = ~w37778 & w38053 ;
  assign w38055 = ( w37458 & w37776 ) | ( w37458 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38056 = ~w37777 & w38055 ;
  assign w38057 = w38054 | w38056 ;
  assign w38058 = ~\pi085 & w38057 ;
  assign w38059 = ~w37473 & w37640 ;
  assign w38060 = w37641 ^ w38059 ;
  assign w38061 = ~w37778 & w38060 ;
  assign w38062 = ( w37465 & w37776 ) | ( w37465 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38063 = ~w37777 & w38062 ;
  assign w38064 = w38061 | w38063 ;
  assign w38065 = ~\pi084 & w38064 ;
  assign w38066 = ~w37480 & w37637 ;
  assign w38067 = w37638 ^ w38066 ;
  assign w38068 = ~w37778 & w38067 ;
  assign w38069 = ( w37472 & w37776 ) | ( w37472 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38070 = ~w37777 & w38069 ;
  assign w38071 = w38068 | w38070 ;
  assign w38072 = ~\pi083 & w38071 ;
  assign w38073 = ~w37487 & w37634 ;
  assign w38074 = w37635 ^ w38073 ;
  assign w38075 = ~w37778 & w38074 ;
  assign w38076 = ( w37479 & w37776 ) | ( w37479 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38077 = ~w37777 & w38076 ;
  assign w38078 = w38075 | w38077 ;
  assign w38079 = ~\pi082 & w38078 ;
  assign w38080 = ~w37494 & w37631 ;
  assign w38081 = w37632 ^ w38080 ;
  assign w38082 = ~w37778 & w38081 ;
  assign w38083 = ( w37486 & w37776 ) | ( w37486 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38084 = ~w37777 & w38083 ;
  assign w38085 = w38082 | w38084 ;
  assign w38086 = ~\pi081 & w38085 ;
  assign w38087 = ~w37501 & w37628 ;
  assign w38088 = w37629 ^ w38087 ;
  assign w38089 = ~w37778 & w38088 ;
  assign w38090 = ( w37493 & w37776 ) | ( w37493 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38091 = ~w37777 & w38090 ;
  assign w38092 = w38089 | w38091 ;
  assign w38093 = ~\pi080 & w38092 ;
  assign w38094 = ~w37508 & w37625 ;
  assign w38095 = w37626 ^ w38094 ;
  assign w38096 = ~w37778 & w38095 ;
  assign w38097 = ( w37500 & w37776 ) | ( w37500 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38098 = ~w37777 & w38097 ;
  assign w38099 = w38096 | w38098 ;
  assign w38100 = ~\pi079 & w38099 ;
  assign w38101 = ~w37515 & w37622 ;
  assign w38102 = w37623 ^ w38101 ;
  assign w38103 = ~w37778 & w38102 ;
  assign w38104 = ( w37507 & w37776 ) | ( w37507 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38105 = ~w37777 & w38104 ;
  assign w38106 = w38103 | w38105 ;
  assign w38107 = ~\pi078 & w38106 ;
  assign w38108 = ~w37522 & w37619 ;
  assign w38109 = w37620 ^ w38108 ;
  assign w38110 = ~w37778 & w38109 ;
  assign w38111 = ( w37514 & w37776 ) | ( w37514 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38112 = ~w37777 & w38111 ;
  assign w38113 = w38110 | w38112 ;
  assign w38114 = ~\pi077 & w38113 ;
  assign w38115 = ~w37529 & w37616 ;
  assign w38116 = w37617 ^ w38115 ;
  assign w38117 = ~w37778 & w38116 ;
  assign w38118 = ( w37521 & w37776 ) | ( w37521 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38119 = ~w37777 & w38118 ;
  assign w38120 = w38117 | w38119 ;
  assign w38121 = ~\pi076 & w38120 ;
  assign w38122 = ~w37536 & w37613 ;
  assign w38123 = w37614 ^ w38122 ;
  assign w38124 = ~w37778 & w38123 ;
  assign w38125 = ( w37528 & w37776 ) | ( w37528 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38126 = ~w37777 & w38125 ;
  assign w38127 = w38124 | w38126 ;
  assign w38128 = ~\pi075 & w38127 ;
  assign w38129 = ~w37543 & w37610 ;
  assign w38130 = w37611 ^ w38129 ;
  assign w38131 = ~w37778 & w38130 ;
  assign w38132 = ( w37535 & w37776 ) | ( w37535 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38133 = ~w37777 & w38132 ;
  assign w38134 = w38131 | w38133 ;
  assign w38135 = ~\pi074 & w38134 ;
  assign w38136 = ~w37550 & w37607 ;
  assign w38137 = w37608 ^ w38136 ;
  assign w38138 = ~w37778 & w38137 ;
  assign w38139 = ( w37542 & w37776 ) | ( w37542 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38140 = ~w37777 & w38139 ;
  assign w38141 = w38138 | w38140 ;
  assign w38142 = ~\pi073 & w38141 ;
  assign w38143 = ~w37557 & w37604 ;
  assign w38144 = w37605 ^ w38143 ;
  assign w38145 = ~w37778 & w38144 ;
  assign w38146 = ( w37549 & w37776 ) | ( w37549 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38147 = ~w37777 & w38146 ;
  assign w38148 = w38145 | w38147 ;
  assign w38149 = ~\pi072 & w38148 ;
  assign w38150 = ~w37564 & w37601 ;
  assign w38151 = w37602 ^ w38150 ;
  assign w38152 = ~w37778 & w38151 ;
  assign w38153 = ( w37556 & w37776 ) | ( w37556 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38154 = ~w37777 & w38153 ;
  assign w38155 = w38152 | w38154 ;
  assign w38156 = ~\pi071 & w38155 ;
  assign w38157 = ~w37571 & w37598 ;
  assign w38158 = w37599 ^ w38157 ;
  assign w38159 = ~w37778 & w38158 ;
  assign w38160 = ( w37563 & w37776 ) | ( w37563 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38161 = ~w37777 & w38160 ;
  assign w38162 = w38159 | w38161 ;
  assign w38163 = ~\pi070 & w38162 ;
  assign w38164 = ~w37580 & w37595 ;
  assign w38165 = w37596 ^ w38164 ;
  assign w38166 = ~w37778 & w38165 ;
  assign w38167 = ( w37570 & w37776 ) | ( w37570 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38168 = ~w37777 & w38167 ;
  assign w38169 = w38166 | w38168 ;
  assign w38170 = ~\pi069 & w38169 ;
  assign w38171 = ~w37587 & w37592 ;
  assign w38172 = w37593 ^ w38171 ;
  assign w38173 = ~w37778 & w38172 ;
  assign w38174 = ( w37579 & w37776 ) | ( w37579 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38175 = ~w37777 & w38174 ;
  assign w38176 = w38173 | w38175 ;
  assign w38177 = ~\pi068 & w38176 ;
  assign w38178 = \pi064 & ~w37179 ;
  assign w38179 = \pi004 ^ w38178 ;
  assign w38180 = ( \pi065 & w18843 ) | ( \pi065 & ~w38179 ) | ( w18843 & ~w38179 ) ;
  assign w38181 = w37588 ^ w38180 ;
  assign w38182 = ~w37778 & w38181 ;
  assign w38183 = ( w37586 & w37776 ) | ( w37586 & w37777 ) | ( w37776 & w37777 ) ;
  assign w38184 = ~w37777 & w38183 ;
  assign w38185 = w38182 | w38184 ;
  assign w38186 = ~\pi067 & w38185 ;
  assign w38187 = \pi003 ^ w37179 ;
  assign w38188 = ( \pi064 & w37778 ) | ( \pi064 & w38187 ) | ( w37778 & w38187 ) ;
  assign w38189 = w18851 ^ w38188 ;
  assign w38190 = ~w37778 & w38189 ;
  assign w38191 = w37778 & w38179 ;
  assign w38192 = w38190 | w38191 ;
  assign w38193 = ~\pi066 & w38192 ;
  assign w38194 = \pi066 ^ w38192 ;
  assign w38195 = ( \pi064 & ~w37778 ) | ( \pi064 & w38194 ) | ( ~w37778 & w38194 ) ;
  assign w38196 = \pi003 ^ w38195 ;
  assign w38197 = ( \pi065 & w19461 ) | ( \pi065 & ~w38196 ) | ( w19461 & ~w38196 ) ;
  assign w38198 = w38194 | w38197 ;
  assign w38199 = \pi067 ^ w38185 ;
  assign w38200 = ( ~w38193 & w38198 ) | ( ~w38193 & w38199 ) | ( w38198 & w38199 ) ;
  assign w38201 = w38199 | w38200 ;
  assign w38202 = \pi068 ^ w38176 ;
  assign w38203 = ( ~w38186 & w38201 ) | ( ~w38186 & w38202 ) | ( w38201 & w38202 ) ;
  assign w38204 = w38202 | w38203 ;
  assign w38205 = \pi069 ^ w38169 ;
  assign w38206 = ( ~w38177 & w38204 ) | ( ~w38177 & w38205 ) | ( w38204 & w38205 ) ;
  assign w38207 = w38205 | w38206 ;
  assign w38208 = \pi070 ^ w38162 ;
  assign w38209 = ( ~w38170 & w38207 ) | ( ~w38170 & w38208 ) | ( w38207 & w38208 ) ;
  assign w38210 = w38208 | w38209 ;
  assign w38211 = \pi071 ^ w38155 ;
  assign w38212 = ( ~w38163 & w38210 ) | ( ~w38163 & w38211 ) | ( w38210 & w38211 ) ;
  assign w38213 = w38211 | w38212 ;
  assign w38214 = \pi072 ^ w38148 ;
  assign w38215 = ( ~w38156 & w38213 ) | ( ~w38156 & w38214 ) | ( w38213 & w38214 ) ;
  assign w38216 = w38214 | w38215 ;
  assign w38217 = \pi073 ^ w38141 ;
  assign w38218 = ( ~w38149 & w38216 ) | ( ~w38149 & w38217 ) | ( w38216 & w38217 ) ;
  assign w38219 = w38217 | w38218 ;
  assign w38220 = \pi074 ^ w38134 ;
  assign w38221 = ( ~w38142 & w38219 ) | ( ~w38142 & w38220 ) | ( w38219 & w38220 ) ;
  assign w38222 = w38220 | w38221 ;
  assign w38223 = \pi075 ^ w38127 ;
  assign w38224 = ( ~w38135 & w38222 ) | ( ~w38135 & w38223 ) | ( w38222 & w38223 ) ;
  assign w38225 = w38223 | w38224 ;
  assign w38226 = \pi076 ^ w38120 ;
  assign w38227 = ( ~w38128 & w38225 ) | ( ~w38128 & w38226 ) | ( w38225 & w38226 ) ;
  assign w38228 = w38226 | w38227 ;
  assign w38229 = \pi077 ^ w38113 ;
  assign w38230 = ( ~w38121 & w38228 ) | ( ~w38121 & w38229 ) | ( w38228 & w38229 ) ;
  assign w38231 = w38229 | w38230 ;
  assign w38232 = \pi078 ^ w38106 ;
  assign w38233 = ( ~w38114 & w38231 ) | ( ~w38114 & w38232 ) | ( w38231 & w38232 ) ;
  assign w38234 = w38232 | w38233 ;
  assign w38235 = \pi079 ^ w38099 ;
  assign w38236 = ( ~w38107 & w38234 ) | ( ~w38107 & w38235 ) | ( w38234 & w38235 ) ;
  assign w38237 = w38235 | w38236 ;
  assign w38238 = \pi080 ^ w38092 ;
  assign w38239 = ( ~w38100 & w38237 ) | ( ~w38100 & w38238 ) | ( w38237 & w38238 ) ;
  assign w38240 = w38238 | w38239 ;
  assign w38241 = \pi081 ^ w38085 ;
  assign w38242 = ( ~w38093 & w38240 ) | ( ~w38093 & w38241 ) | ( w38240 & w38241 ) ;
  assign w38243 = w38241 | w38242 ;
  assign w38244 = \pi082 ^ w38078 ;
  assign w38245 = ( ~w38086 & w38243 ) | ( ~w38086 & w38244 ) | ( w38243 & w38244 ) ;
  assign w38246 = w38244 | w38245 ;
  assign w38247 = \pi083 ^ w38071 ;
  assign w38248 = ( ~w38079 & w38246 ) | ( ~w38079 & w38247 ) | ( w38246 & w38247 ) ;
  assign w38249 = w38247 | w38248 ;
  assign w38250 = \pi084 ^ w38064 ;
  assign w38251 = ( ~w38072 & w38249 ) | ( ~w38072 & w38250 ) | ( w38249 & w38250 ) ;
  assign w38252 = w38250 | w38251 ;
  assign w38253 = \pi085 ^ w38057 ;
  assign w38254 = ( ~w38065 & w38252 ) | ( ~w38065 & w38253 ) | ( w38252 & w38253 ) ;
  assign w38255 = w38253 | w38254 ;
  assign w38256 = \pi086 ^ w38050 ;
  assign w38257 = ( ~w38058 & w38255 ) | ( ~w38058 & w38256 ) | ( w38255 & w38256 ) ;
  assign w38258 = w38256 | w38257 ;
  assign w38259 = \pi087 ^ w38043 ;
  assign w38260 = ( ~w38051 & w38258 ) | ( ~w38051 & w38259 ) | ( w38258 & w38259 ) ;
  assign w38261 = w38259 | w38260 ;
  assign w38262 = \pi088 ^ w38036 ;
  assign w38263 = ( ~w38044 & w38261 ) | ( ~w38044 & w38262 ) | ( w38261 & w38262 ) ;
  assign w38264 = w38262 | w38263 ;
  assign w38265 = \pi089 ^ w38029 ;
  assign w38266 = ( ~w38037 & w38264 ) | ( ~w38037 & w38265 ) | ( w38264 & w38265 ) ;
  assign w38267 = w38265 | w38266 ;
  assign w38268 = \pi090 ^ w38022 ;
  assign w38269 = ( ~w38030 & w38267 ) | ( ~w38030 & w38268 ) | ( w38267 & w38268 ) ;
  assign w38270 = w38268 | w38269 ;
  assign w38271 = \pi091 ^ w38015 ;
  assign w38272 = ( ~w38023 & w38270 ) | ( ~w38023 & w38271 ) | ( w38270 & w38271 ) ;
  assign w38273 = w38271 | w38272 ;
  assign w38274 = \pi092 ^ w38008 ;
  assign w38275 = ( ~w38016 & w38273 ) | ( ~w38016 & w38274 ) | ( w38273 & w38274 ) ;
  assign w38276 = w38274 | w38275 ;
  assign w38277 = \pi093 ^ w38001 ;
  assign w38278 = ( ~w38009 & w38276 ) | ( ~w38009 & w38277 ) | ( w38276 & w38277 ) ;
  assign w38279 = w38277 | w38278 ;
  assign w38280 = \pi094 ^ w37994 ;
  assign w38281 = ( ~w38002 & w38279 ) | ( ~w38002 & w38280 ) | ( w38279 & w38280 ) ;
  assign w38282 = w38280 | w38281 ;
  assign w38283 = \pi095 ^ w37987 ;
  assign w38284 = ( ~w37995 & w38282 ) | ( ~w37995 & w38283 ) | ( w38282 & w38283 ) ;
  assign w38285 = w38283 | w38284 ;
  assign w38286 = \pi096 ^ w37980 ;
  assign w38287 = ( ~w37988 & w38285 ) | ( ~w37988 & w38286 ) | ( w38285 & w38286 ) ;
  assign w38288 = w38286 | w38287 ;
  assign w38289 = \pi097 ^ w37973 ;
  assign w38290 = ( ~w37981 & w38288 ) | ( ~w37981 & w38289 ) | ( w38288 & w38289 ) ;
  assign w38291 = w38289 | w38290 ;
  assign w38292 = \pi098 ^ w37966 ;
  assign w38293 = ( ~w37974 & w38291 ) | ( ~w37974 & w38292 ) | ( w38291 & w38292 ) ;
  assign w38294 = w38292 | w38293 ;
  assign w38295 = \pi099 ^ w37959 ;
  assign w38296 = ( ~w37967 & w38294 ) | ( ~w37967 & w38295 ) | ( w38294 & w38295 ) ;
  assign w38297 = w38295 | w38296 ;
  assign w38298 = \pi100 ^ w37952 ;
  assign w38299 = ( ~w37960 & w38297 ) | ( ~w37960 & w38298 ) | ( w38297 & w38298 ) ;
  assign w38300 = w38298 | w38299 ;
  assign w38301 = \pi101 ^ w37945 ;
  assign w38302 = ( ~w37953 & w38300 ) | ( ~w37953 & w38301 ) | ( w38300 & w38301 ) ;
  assign w38303 = w38301 | w38302 ;
  assign w38304 = \pi102 ^ w37938 ;
  assign w38305 = ( ~w37946 & w38303 ) | ( ~w37946 & w38304 ) | ( w38303 & w38304 ) ;
  assign w38306 = w38304 | w38305 ;
  assign w38307 = \pi103 ^ w37931 ;
  assign w38308 = ( ~w37939 & w38306 ) | ( ~w37939 & w38307 ) | ( w38306 & w38307 ) ;
  assign w38309 = w38307 | w38308 ;
  assign w38310 = \pi104 ^ w37924 ;
  assign w38311 = ( ~w37932 & w38309 ) | ( ~w37932 & w38310 ) | ( w38309 & w38310 ) ;
  assign w38312 = w38310 | w38311 ;
  assign w38313 = \pi105 ^ w37917 ;
  assign w38314 = ( ~w37925 & w38312 ) | ( ~w37925 & w38313 ) | ( w38312 & w38313 ) ;
  assign w38315 = w38313 | w38314 ;
  assign w38316 = \pi106 ^ w37910 ;
  assign w38317 = ( ~w37918 & w38315 ) | ( ~w37918 & w38316 ) | ( w38315 & w38316 ) ;
  assign w38318 = w38316 | w38317 ;
  assign w38319 = \pi107 ^ w37903 ;
  assign w38320 = ( ~w37911 & w38318 ) | ( ~w37911 & w38319 ) | ( w38318 & w38319 ) ;
  assign w38321 = w38319 | w38320 ;
  assign w38322 = \pi108 ^ w37896 ;
  assign w38323 = ( ~w37904 & w38321 ) | ( ~w37904 & w38322 ) | ( w38321 & w38322 ) ;
  assign w38324 = w38322 | w38323 ;
  assign w38325 = \pi109 ^ w37889 ;
  assign w38326 = ( ~w37897 & w38324 ) | ( ~w37897 & w38325 ) | ( w38324 & w38325 ) ;
  assign w38327 = w38325 | w38326 ;
  assign w38328 = \pi110 ^ w37882 ;
  assign w38329 = ( ~w37890 & w38327 ) | ( ~w37890 & w38328 ) | ( w38327 & w38328 ) ;
  assign w38330 = w38328 | w38329 ;
  assign w38331 = \pi111 ^ w37875 ;
  assign w38332 = ( ~w37883 & w38330 ) | ( ~w37883 & w38331 ) | ( w38330 & w38331 ) ;
  assign w38333 = w38331 | w38332 ;
  assign w38334 = \pi112 ^ w37868 ;
  assign w38335 = ( ~w37876 & w38333 ) | ( ~w37876 & w38334 ) | ( w38333 & w38334 ) ;
  assign w38336 = w38334 | w38335 ;
  assign w38337 = \pi113 ^ w37861 ;
  assign w38338 = ( ~w37869 & w38336 ) | ( ~w37869 & w38337 ) | ( w38336 & w38337 ) ;
  assign w38339 = w38337 | w38338 ;
  assign w38340 = \pi114 ^ w37854 ;
  assign w38341 = ( ~w37862 & w38339 ) | ( ~w37862 & w38340 ) | ( w38339 & w38340 ) ;
  assign w38342 = w38340 | w38341 ;
  assign w38343 = \pi115 ^ w37847 ;
  assign w38344 = ( ~w37855 & w38342 ) | ( ~w37855 & w38343 ) | ( w38342 & w38343 ) ;
  assign w38345 = w38343 | w38344 ;
  assign w38346 = \pi116 ^ w37840 ;
  assign w38347 = ( ~w37848 & w38345 ) | ( ~w37848 & w38346 ) | ( w38345 & w38346 ) ;
  assign w38348 = w38346 | w38347 ;
  assign w38349 = \pi117 ^ w37833 ;
  assign w38350 = ( ~w37841 & w38348 ) | ( ~w37841 & w38349 ) | ( w38348 & w38349 ) ;
  assign w38351 = w38349 | w38350 ;
  assign w38352 = \pi118 ^ w37826 ;
  assign w38353 = ( ~w37834 & w38351 ) | ( ~w37834 & w38352 ) | ( w38351 & w38352 ) ;
  assign w38354 = w38352 | w38353 ;
  assign w38355 = \pi119 ^ w37819 ;
  assign w38356 = ( ~w37827 & w38354 ) | ( ~w37827 & w38355 ) | ( w38354 & w38355 ) ;
  assign w38357 = w38355 | w38356 ;
  assign w38358 = \pi120 ^ w37812 ;
  assign w38359 = ( ~w37820 & w38357 ) | ( ~w37820 & w38358 ) | ( w38357 & w38358 ) ;
  assign w38360 = w38358 | w38359 ;
  assign w38361 = \pi121 ^ w37805 ;
  assign w38362 = ( ~w37813 & w38360 ) | ( ~w37813 & w38361 ) | ( w38360 & w38361 ) ;
  assign w38363 = w38361 | w38362 ;
  assign w38364 = \pi122 ^ w37798 ;
  assign w38365 = ( ~w37806 & w38363 ) | ( ~w37806 & w38364 ) | ( w38363 & w38364 ) ;
  assign w38366 = w38364 | w38365 ;
  assign w38367 = \pi123 ^ w37791 ;
  assign w38368 = ( ~w37799 & w38366 ) | ( ~w37799 & w38367 ) | ( w38366 & w38367 ) ;
  assign w38369 = w38367 | w38368 ;
  assign w38370 = \pi124 ^ w37784 ;
  assign w38371 = ( ~w37792 & w38369 ) | ( ~w37792 & w38370 ) | ( w38369 & w38370 ) ;
  assign w38372 = w38370 | w38371 ;
  assign w38373 = ( ~w37186 & w37763 ) | ( ~w37186 & w37778 ) | ( w37763 & w37778 ) ;
  assign w38374 = w37773 ^ w38373 ;
  assign w38375 = ~w37778 & w38374 ;
  assign w38376 = ( w147 & ~w37769 ) | ( w147 & w37776 ) | ( ~w37769 & w37776 ) ;
  assign w38377 = w37769 & w38376 ;
  assign w38378 = w38375 | w38377 ;
  assign w38379 = ~\pi125 & w38378 ;
  assign w38380 = ( \pi125 & ~w38375 ) | ( \pi125 & w38377 ) | ( ~w38375 & w38377 ) ;
  assign w38381 = ~w38377 & w38380 ;
  assign w38382 = ( ~w37785 & w38372 ) | ( ~w37785 & w38379 ) | ( w38372 & w38379 ) ;
  assign w38383 = ( \pi127 & w38379 ) | ( \pi127 & ~w38382 ) | ( w38379 & ~w38382 ) ;
  assign w38384 = ( \pi126 & w38381 ) | ( \pi126 & ~w38382 ) | ( w38381 & ~w38382 ) ;
  assign w38385 = ( w38382 & ~w38383 ) | ( w38382 & w38384 ) | ( ~w38383 & w38384 ) ;
  assign w38386 = w38383 | w38385 ;
  assign w38387 = ~w269 & w38378 ;
  assign w38388 = w38386 & ~w38387 ;
  assign w38389 = ~w37792 & w38369 ;
  assign w38390 = w38370 ^ w38389 ;
  assign w38391 = ~w38388 & w38390 ;
  assign w38392 = ( w37784 & w38386 ) | ( w37784 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38393 = ~w38387 & w38392 ;
  assign w38394 = w38391 | w38393 ;
  assign w38395 = ~\pi125 & w38394 ;
  assign w38396 = ~w37799 & w38366 ;
  assign w38397 = w38367 ^ w38396 ;
  assign w38398 = ~w38388 & w38397 ;
  assign w38399 = ( w37791 & w38386 ) | ( w37791 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38400 = ~w38387 & w38399 ;
  assign w38401 = w38398 | w38400 ;
  assign w38402 = ~\pi124 & w38401 ;
  assign w38403 = ~w37806 & w38363 ;
  assign w38404 = w38364 ^ w38403 ;
  assign w38405 = ~w38388 & w38404 ;
  assign w38406 = ( w37798 & w38386 ) | ( w37798 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38407 = ~w38387 & w38406 ;
  assign w38408 = w38405 | w38407 ;
  assign w38409 = ~\pi123 & w38408 ;
  assign w38410 = ~w37813 & w38360 ;
  assign w38411 = w38361 ^ w38410 ;
  assign w38412 = ~w38388 & w38411 ;
  assign w38413 = ( w37805 & w38386 ) | ( w37805 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38414 = ~w38387 & w38413 ;
  assign w38415 = w38412 | w38414 ;
  assign w38416 = ~\pi122 & w38415 ;
  assign w38417 = ~w37820 & w38357 ;
  assign w38418 = w38358 ^ w38417 ;
  assign w38419 = ~w38388 & w38418 ;
  assign w38420 = ( w37812 & w38386 ) | ( w37812 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38421 = ~w38387 & w38420 ;
  assign w38422 = w38419 | w38421 ;
  assign w38423 = ~\pi121 & w38422 ;
  assign w38424 = ~w37827 & w38354 ;
  assign w38425 = w38355 ^ w38424 ;
  assign w38426 = ~w38388 & w38425 ;
  assign w38427 = ( w37819 & w38386 ) | ( w37819 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38428 = ~w38387 & w38427 ;
  assign w38429 = w38426 | w38428 ;
  assign w38430 = ~\pi120 & w38429 ;
  assign w38431 = ~w37834 & w38351 ;
  assign w38432 = w38352 ^ w38431 ;
  assign w38433 = ~w38388 & w38432 ;
  assign w38434 = ( w37826 & w38386 ) | ( w37826 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38435 = ~w38387 & w38434 ;
  assign w38436 = w38433 | w38435 ;
  assign w38437 = ~\pi119 & w38436 ;
  assign w38438 = ~w37841 & w38348 ;
  assign w38439 = w38349 ^ w38438 ;
  assign w38440 = ~w38388 & w38439 ;
  assign w38441 = ( w37833 & w38386 ) | ( w37833 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38442 = ~w38387 & w38441 ;
  assign w38443 = w38440 | w38442 ;
  assign w38444 = ~\pi118 & w38443 ;
  assign w38445 = ~w37848 & w38345 ;
  assign w38446 = w38346 ^ w38445 ;
  assign w38447 = ~w38388 & w38446 ;
  assign w38448 = ( w37840 & w38386 ) | ( w37840 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38449 = ~w38387 & w38448 ;
  assign w38450 = w38447 | w38449 ;
  assign w38451 = ~\pi117 & w38450 ;
  assign w38452 = ~w37855 & w38342 ;
  assign w38453 = w38343 ^ w38452 ;
  assign w38454 = ~w38388 & w38453 ;
  assign w38455 = ( w37847 & w38386 ) | ( w37847 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38456 = ~w38387 & w38455 ;
  assign w38457 = w38454 | w38456 ;
  assign w38458 = ~\pi116 & w38457 ;
  assign w38459 = ~w37862 & w38339 ;
  assign w38460 = w38340 ^ w38459 ;
  assign w38461 = ~w38388 & w38460 ;
  assign w38462 = ( w37854 & w38386 ) | ( w37854 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38463 = ~w38387 & w38462 ;
  assign w38464 = w38461 | w38463 ;
  assign w38465 = ~\pi115 & w38464 ;
  assign w38466 = ~w37869 & w38336 ;
  assign w38467 = w38337 ^ w38466 ;
  assign w38468 = ~w38388 & w38467 ;
  assign w38469 = ( w37861 & w38386 ) | ( w37861 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38470 = ~w38387 & w38469 ;
  assign w38471 = w38468 | w38470 ;
  assign w38472 = ~\pi114 & w38471 ;
  assign w38473 = ~w37876 & w38333 ;
  assign w38474 = w38334 ^ w38473 ;
  assign w38475 = ~w38388 & w38474 ;
  assign w38476 = ( w37868 & w38386 ) | ( w37868 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38477 = ~w38387 & w38476 ;
  assign w38478 = w38475 | w38477 ;
  assign w38479 = ~\pi113 & w38478 ;
  assign w38480 = ~w37883 & w38330 ;
  assign w38481 = w38331 ^ w38480 ;
  assign w38482 = ~w38388 & w38481 ;
  assign w38483 = ( w37875 & w38386 ) | ( w37875 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38484 = ~w38387 & w38483 ;
  assign w38485 = w38482 | w38484 ;
  assign w38486 = ~\pi112 & w38485 ;
  assign w38487 = ~w37890 & w38327 ;
  assign w38488 = w38328 ^ w38487 ;
  assign w38489 = ~w38388 & w38488 ;
  assign w38490 = ( w37882 & w38386 ) | ( w37882 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38491 = ~w38387 & w38490 ;
  assign w38492 = w38489 | w38491 ;
  assign w38493 = ~\pi111 & w38492 ;
  assign w38494 = ~w37897 & w38324 ;
  assign w38495 = w38325 ^ w38494 ;
  assign w38496 = ~w38388 & w38495 ;
  assign w38497 = ( w37889 & w38386 ) | ( w37889 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38498 = ~w38387 & w38497 ;
  assign w38499 = w38496 | w38498 ;
  assign w38500 = ~\pi110 & w38499 ;
  assign w38501 = ~w37904 & w38321 ;
  assign w38502 = w38322 ^ w38501 ;
  assign w38503 = ~w38388 & w38502 ;
  assign w38504 = ( w37896 & w38386 ) | ( w37896 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38505 = ~w38387 & w38504 ;
  assign w38506 = w38503 | w38505 ;
  assign w38507 = ~\pi109 & w38506 ;
  assign w38508 = ~w37911 & w38318 ;
  assign w38509 = w38319 ^ w38508 ;
  assign w38510 = ~w38388 & w38509 ;
  assign w38511 = ( w37903 & w38386 ) | ( w37903 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38512 = ~w38387 & w38511 ;
  assign w38513 = w38510 | w38512 ;
  assign w38514 = ~\pi108 & w38513 ;
  assign w38515 = ~w37918 & w38315 ;
  assign w38516 = w38316 ^ w38515 ;
  assign w38517 = ~w38388 & w38516 ;
  assign w38518 = ( w37910 & w38386 ) | ( w37910 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38519 = ~w38387 & w38518 ;
  assign w38520 = w38517 | w38519 ;
  assign w38521 = ~\pi107 & w38520 ;
  assign w38522 = ~w37925 & w38312 ;
  assign w38523 = w38313 ^ w38522 ;
  assign w38524 = ~w38388 & w38523 ;
  assign w38525 = ( w37917 & w38386 ) | ( w37917 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38526 = ~w38387 & w38525 ;
  assign w38527 = w38524 | w38526 ;
  assign w38528 = ~\pi106 & w38527 ;
  assign w38529 = ~w37932 & w38309 ;
  assign w38530 = w38310 ^ w38529 ;
  assign w38531 = ~w38388 & w38530 ;
  assign w38532 = ( w37924 & w38386 ) | ( w37924 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38533 = ~w38387 & w38532 ;
  assign w38534 = w38531 | w38533 ;
  assign w38535 = ~\pi105 & w38534 ;
  assign w38536 = ~w37939 & w38306 ;
  assign w38537 = w38307 ^ w38536 ;
  assign w38538 = ~w38388 & w38537 ;
  assign w38539 = ( w37931 & w38386 ) | ( w37931 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38540 = ~w38387 & w38539 ;
  assign w38541 = w38538 | w38540 ;
  assign w38542 = ~\pi104 & w38541 ;
  assign w38543 = ~w37946 & w38303 ;
  assign w38544 = w38304 ^ w38543 ;
  assign w38545 = ~w38388 & w38544 ;
  assign w38546 = ( w37938 & w38386 ) | ( w37938 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38547 = ~w38387 & w38546 ;
  assign w38548 = w38545 | w38547 ;
  assign w38549 = ~\pi103 & w38548 ;
  assign w38550 = ~w37953 & w38300 ;
  assign w38551 = w38301 ^ w38550 ;
  assign w38552 = ~w38388 & w38551 ;
  assign w38553 = ( w37945 & w38386 ) | ( w37945 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38554 = ~w38387 & w38553 ;
  assign w38555 = w38552 | w38554 ;
  assign w38556 = ~\pi102 & w38555 ;
  assign w38557 = ~w37960 & w38297 ;
  assign w38558 = w38298 ^ w38557 ;
  assign w38559 = ~w38388 & w38558 ;
  assign w38560 = ( w37952 & w38386 ) | ( w37952 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38561 = ~w38387 & w38560 ;
  assign w38562 = w38559 | w38561 ;
  assign w38563 = ~\pi101 & w38562 ;
  assign w38564 = ~w37967 & w38294 ;
  assign w38565 = w38295 ^ w38564 ;
  assign w38566 = ~w38388 & w38565 ;
  assign w38567 = ( w37959 & w38386 ) | ( w37959 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38568 = ~w38387 & w38567 ;
  assign w38569 = w38566 | w38568 ;
  assign w38570 = ~\pi100 & w38569 ;
  assign w38571 = ~w37974 & w38291 ;
  assign w38572 = w38292 ^ w38571 ;
  assign w38573 = ~w38388 & w38572 ;
  assign w38574 = ( w37966 & w38386 ) | ( w37966 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38575 = ~w38387 & w38574 ;
  assign w38576 = w38573 | w38575 ;
  assign w38577 = ~\pi099 & w38576 ;
  assign w38578 = ~w37981 & w38288 ;
  assign w38579 = w38289 ^ w38578 ;
  assign w38580 = ~w38388 & w38579 ;
  assign w38581 = ( w37973 & w38386 ) | ( w37973 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38582 = ~w38387 & w38581 ;
  assign w38583 = w38580 | w38582 ;
  assign w38584 = ~\pi098 & w38583 ;
  assign w38585 = ~w37988 & w38285 ;
  assign w38586 = w38286 ^ w38585 ;
  assign w38587 = ~w38388 & w38586 ;
  assign w38588 = ( w37980 & w38386 ) | ( w37980 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38589 = ~w38387 & w38588 ;
  assign w38590 = w38587 | w38589 ;
  assign w38591 = ~\pi097 & w38590 ;
  assign w38592 = ~w37995 & w38282 ;
  assign w38593 = w38283 ^ w38592 ;
  assign w38594 = ~w38388 & w38593 ;
  assign w38595 = ( w37987 & w38386 ) | ( w37987 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38596 = ~w38387 & w38595 ;
  assign w38597 = w38594 | w38596 ;
  assign w38598 = ~\pi096 & w38597 ;
  assign w38599 = ~w38002 & w38279 ;
  assign w38600 = w38280 ^ w38599 ;
  assign w38601 = ~w38388 & w38600 ;
  assign w38602 = ( w37994 & w38386 ) | ( w37994 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38603 = ~w38387 & w38602 ;
  assign w38604 = w38601 | w38603 ;
  assign w38605 = ~\pi095 & w38604 ;
  assign w38606 = ~w38009 & w38276 ;
  assign w38607 = w38277 ^ w38606 ;
  assign w38608 = ~w38388 & w38607 ;
  assign w38609 = ( w38001 & w38386 ) | ( w38001 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38610 = ~w38387 & w38609 ;
  assign w38611 = w38608 | w38610 ;
  assign w38612 = ~\pi094 & w38611 ;
  assign w38613 = ~w38016 & w38273 ;
  assign w38614 = w38274 ^ w38613 ;
  assign w38615 = ~w38388 & w38614 ;
  assign w38616 = ( w38008 & w38386 ) | ( w38008 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38617 = ~w38387 & w38616 ;
  assign w38618 = w38615 | w38617 ;
  assign w38619 = ~\pi093 & w38618 ;
  assign w38620 = ~w38023 & w38270 ;
  assign w38621 = w38271 ^ w38620 ;
  assign w38622 = ~w38388 & w38621 ;
  assign w38623 = ( w38015 & w38386 ) | ( w38015 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38624 = ~w38387 & w38623 ;
  assign w38625 = w38622 | w38624 ;
  assign w38626 = ~\pi092 & w38625 ;
  assign w38627 = ~w38030 & w38267 ;
  assign w38628 = w38268 ^ w38627 ;
  assign w38629 = ~w38388 & w38628 ;
  assign w38630 = ( w38022 & w38386 ) | ( w38022 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38631 = ~w38387 & w38630 ;
  assign w38632 = w38629 | w38631 ;
  assign w38633 = ~\pi091 & w38632 ;
  assign w38634 = ~w38037 & w38264 ;
  assign w38635 = w38265 ^ w38634 ;
  assign w38636 = ~w38388 & w38635 ;
  assign w38637 = ( w38029 & w38386 ) | ( w38029 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38638 = ~w38387 & w38637 ;
  assign w38639 = w38636 | w38638 ;
  assign w38640 = ~\pi090 & w38639 ;
  assign w38641 = ~w38044 & w38261 ;
  assign w38642 = w38262 ^ w38641 ;
  assign w38643 = ~w38388 & w38642 ;
  assign w38644 = ( w38036 & w38386 ) | ( w38036 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38645 = ~w38387 & w38644 ;
  assign w38646 = w38643 | w38645 ;
  assign w38647 = ~\pi089 & w38646 ;
  assign w38648 = ~w38051 & w38258 ;
  assign w38649 = w38259 ^ w38648 ;
  assign w38650 = ~w38388 & w38649 ;
  assign w38651 = ( w38043 & w38386 ) | ( w38043 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38652 = ~w38387 & w38651 ;
  assign w38653 = w38650 | w38652 ;
  assign w38654 = ~\pi088 & w38653 ;
  assign w38655 = ~w38058 & w38255 ;
  assign w38656 = w38256 ^ w38655 ;
  assign w38657 = ~w38388 & w38656 ;
  assign w38658 = ( w38050 & w38386 ) | ( w38050 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38659 = ~w38387 & w38658 ;
  assign w38660 = w38657 | w38659 ;
  assign w38661 = ~\pi087 & w38660 ;
  assign w38662 = ~w38065 & w38252 ;
  assign w38663 = w38253 ^ w38662 ;
  assign w38664 = ~w38388 & w38663 ;
  assign w38665 = ( w38057 & w38386 ) | ( w38057 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38666 = ~w38387 & w38665 ;
  assign w38667 = w38664 | w38666 ;
  assign w38668 = ~\pi086 & w38667 ;
  assign w38669 = ~w38072 & w38249 ;
  assign w38670 = w38250 ^ w38669 ;
  assign w38671 = ~w38388 & w38670 ;
  assign w38672 = ( w38064 & w38386 ) | ( w38064 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38673 = ~w38387 & w38672 ;
  assign w38674 = w38671 | w38673 ;
  assign w38675 = ~\pi085 & w38674 ;
  assign w38676 = ~w38079 & w38246 ;
  assign w38677 = w38247 ^ w38676 ;
  assign w38678 = ~w38388 & w38677 ;
  assign w38679 = ( w38071 & w38386 ) | ( w38071 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38680 = ~w38387 & w38679 ;
  assign w38681 = w38678 | w38680 ;
  assign w38682 = ~\pi084 & w38681 ;
  assign w38683 = ~w38086 & w38243 ;
  assign w38684 = w38244 ^ w38683 ;
  assign w38685 = ~w38388 & w38684 ;
  assign w38686 = ( w38078 & w38386 ) | ( w38078 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38687 = ~w38387 & w38686 ;
  assign w38688 = w38685 | w38687 ;
  assign w38689 = ~\pi083 & w38688 ;
  assign w38690 = ~w38093 & w38240 ;
  assign w38691 = w38241 ^ w38690 ;
  assign w38692 = ~w38388 & w38691 ;
  assign w38693 = ( w38085 & w38386 ) | ( w38085 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38694 = ~w38387 & w38693 ;
  assign w38695 = w38692 | w38694 ;
  assign w38696 = ~\pi082 & w38695 ;
  assign w38697 = ~w38100 & w38237 ;
  assign w38698 = w38238 ^ w38697 ;
  assign w38699 = ~w38388 & w38698 ;
  assign w38700 = ( w38092 & w38386 ) | ( w38092 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38701 = ~w38387 & w38700 ;
  assign w38702 = w38699 | w38701 ;
  assign w38703 = ~\pi081 & w38702 ;
  assign w38704 = ~w38107 & w38234 ;
  assign w38705 = w38235 ^ w38704 ;
  assign w38706 = ~w38388 & w38705 ;
  assign w38707 = ( w38099 & w38386 ) | ( w38099 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38708 = ~w38387 & w38707 ;
  assign w38709 = w38706 | w38708 ;
  assign w38710 = ~\pi080 & w38709 ;
  assign w38711 = ~w38114 & w38231 ;
  assign w38712 = w38232 ^ w38711 ;
  assign w38713 = ~w38388 & w38712 ;
  assign w38714 = ( w38106 & w38386 ) | ( w38106 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38715 = ~w38387 & w38714 ;
  assign w38716 = w38713 | w38715 ;
  assign w38717 = ~\pi079 & w38716 ;
  assign w38718 = ~w38121 & w38228 ;
  assign w38719 = w38229 ^ w38718 ;
  assign w38720 = ~w38388 & w38719 ;
  assign w38721 = ( w38113 & w38386 ) | ( w38113 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38722 = ~w38387 & w38721 ;
  assign w38723 = w38720 | w38722 ;
  assign w38724 = ~\pi078 & w38723 ;
  assign w38725 = ~w38128 & w38225 ;
  assign w38726 = w38226 ^ w38725 ;
  assign w38727 = ~w38388 & w38726 ;
  assign w38728 = ( w38120 & w38386 ) | ( w38120 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38729 = ~w38387 & w38728 ;
  assign w38730 = w38727 | w38729 ;
  assign w38731 = ~\pi077 & w38730 ;
  assign w38732 = ~w38135 & w38222 ;
  assign w38733 = w38223 ^ w38732 ;
  assign w38734 = ~w38388 & w38733 ;
  assign w38735 = ( w38127 & w38386 ) | ( w38127 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38736 = ~w38387 & w38735 ;
  assign w38737 = w38734 | w38736 ;
  assign w38738 = ~\pi076 & w38737 ;
  assign w38739 = ~w38142 & w38219 ;
  assign w38740 = w38220 ^ w38739 ;
  assign w38741 = ~w38388 & w38740 ;
  assign w38742 = ( w38134 & w38386 ) | ( w38134 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38743 = ~w38387 & w38742 ;
  assign w38744 = w38741 | w38743 ;
  assign w38745 = ~\pi075 & w38744 ;
  assign w38746 = ~w38149 & w38216 ;
  assign w38747 = w38217 ^ w38746 ;
  assign w38748 = ~w38388 & w38747 ;
  assign w38749 = ( w38141 & w38386 ) | ( w38141 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38750 = ~w38387 & w38749 ;
  assign w38751 = w38748 | w38750 ;
  assign w38752 = ~\pi074 & w38751 ;
  assign w38753 = ~w38156 & w38213 ;
  assign w38754 = w38214 ^ w38753 ;
  assign w38755 = ~w38388 & w38754 ;
  assign w38756 = ( w38148 & w38386 ) | ( w38148 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38757 = ~w38387 & w38756 ;
  assign w38758 = w38755 | w38757 ;
  assign w38759 = ~\pi073 & w38758 ;
  assign w38760 = ~w38163 & w38210 ;
  assign w38761 = w38211 ^ w38760 ;
  assign w38762 = ~w38388 & w38761 ;
  assign w38763 = ( w38155 & w38386 ) | ( w38155 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38764 = ~w38387 & w38763 ;
  assign w38765 = w38762 | w38764 ;
  assign w38766 = ~\pi072 & w38765 ;
  assign w38767 = ~w38170 & w38207 ;
  assign w38768 = w38208 ^ w38767 ;
  assign w38769 = ~w38388 & w38768 ;
  assign w38770 = ( w38162 & w38386 ) | ( w38162 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38771 = ~w38387 & w38770 ;
  assign w38772 = w38769 | w38771 ;
  assign w38773 = ~\pi071 & w38772 ;
  assign w38774 = ~w38177 & w38204 ;
  assign w38775 = w38205 ^ w38774 ;
  assign w38776 = ~w38388 & w38775 ;
  assign w38777 = ( w38169 & w38386 ) | ( w38169 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38778 = ~w38387 & w38777 ;
  assign w38779 = w38776 | w38778 ;
  assign w38780 = ~\pi070 & w38779 ;
  assign w38781 = ~w38186 & w38201 ;
  assign w38782 = w38202 ^ w38781 ;
  assign w38783 = ~w38388 & w38782 ;
  assign w38784 = ( w38176 & w38386 ) | ( w38176 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38785 = ~w38387 & w38784 ;
  assign w38786 = w38783 | w38785 ;
  assign w38787 = ~\pi069 & w38786 ;
  assign w38788 = ~w38193 & w38198 ;
  assign w38789 = w38199 ^ w38788 ;
  assign w38790 = ~w38388 & w38789 ;
  assign w38791 = ( w38185 & w38386 ) | ( w38185 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38792 = ~w38387 & w38791 ;
  assign w38793 = w38790 | w38792 ;
  assign w38794 = ~\pi068 & w38793 ;
  assign w38795 = \pi064 & ~w37778 ;
  assign w38796 = \pi003 ^ w38795 ;
  assign w38797 = ( \pi065 & w19461 ) | ( \pi065 & ~w38796 ) | ( w19461 & ~w38796 ) ;
  assign w38798 = w38194 ^ w38797 ;
  assign w38799 = ~w38388 & w38798 ;
  assign w38800 = ( w38192 & w38386 ) | ( w38192 & w38387 ) | ( w38386 & w38387 ) ;
  assign w38801 = ~w38387 & w38800 ;
  assign w38802 = w38799 | w38801 ;
  assign w38803 = ~\pi067 & w38802 ;
  assign w38804 = \pi002 ^ w37778 ;
  assign w38805 = ( \pi064 & w38388 ) | ( \pi064 & w38804 ) | ( w38388 & w38804 ) ;
  assign w38806 = w19469 ^ w38805 ;
  assign w38807 = ~w38388 & w38806 ;
  assign w38808 = w38388 & w38796 ;
  assign w38809 = w38807 | w38808 ;
  assign w38810 = ~\pi066 & w38809 ;
  assign w38811 = \pi066 ^ w38809 ;
  assign w38812 = ( \pi064 & ~w38388 ) | ( \pi064 & w38811 ) | ( ~w38388 & w38811 ) ;
  assign w38813 = \pi002 ^ w38812 ;
  assign w38814 = ( \pi065 & w19790 ) | ( \pi065 & ~w38813 ) | ( w19790 & ~w38813 ) ;
  assign w38815 = w38811 | w38814 ;
  assign w38816 = \pi067 ^ w38802 ;
  assign w38817 = ( ~w38810 & w38815 ) | ( ~w38810 & w38816 ) | ( w38815 & w38816 ) ;
  assign w38818 = w38816 | w38817 ;
  assign w38819 = \pi068 ^ w38793 ;
  assign w38820 = ( ~w38803 & w38818 ) | ( ~w38803 & w38819 ) | ( w38818 & w38819 ) ;
  assign w38821 = w38819 | w38820 ;
  assign w38822 = \pi069 ^ w38786 ;
  assign w38823 = ( ~w38794 & w38821 ) | ( ~w38794 & w38822 ) | ( w38821 & w38822 ) ;
  assign w38824 = w38822 | w38823 ;
  assign w38825 = \pi070 ^ w38779 ;
  assign w38826 = ( ~w38787 & w38824 ) | ( ~w38787 & w38825 ) | ( w38824 & w38825 ) ;
  assign w38827 = w38825 | w38826 ;
  assign w38828 = \pi071 ^ w38772 ;
  assign w38829 = ( ~w38780 & w38827 ) | ( ~w38780 & w38828 ) | ( w38827 & w38828 ) ;
  assign w38830 = w38828 | w38829 ;
  assign w38831 = \pi072 ^ w38765 ;
  assign w38832 = ( ~w38773 & w38830 ) | ( ~w38773 & w38831 ) | ( w38830 & w38831 ) ;
  assign w38833 = w38831 | w38832 ;
  assign w38834 = \pi073 ^ w38758 ;
  assign w38835 = ( ~w38766 & w38833 ) | ( ~w38766 & w38834 ) | ( w38833 & w38834 ) ;
  assign w38836 = w38834 | w38835 ;
  assign w38837 = \pi074 ^ w38751 ;
  assign w38838 = ( ~w38759 & w38836 ) | ( ~w38759 & w38837 ) | ( w38836 & w38837 ) ;
  assign w38839 = w38837 | w38838 ;
  assign w38840 = \pi075 ^ w38744 ;
  assign w38841 = ( ~w38752 & w38839 ) | ( ~w38752 & w38840 ) | ( w38839 & w38840 ) ;
  assign w38842 = w38840 | w38841 ;
  assign w38843 = \pi076 ^ w38737 ;
  assign w38844 = ( ~w38745 & w38842 ) | ( ~w38745 & w38843 ) | ( w38842 & w38843 ) ;
  assign w38845 = w38843 | w38844 ;
  assign w38846 = \pi077 ^ w38730 ;
  assign w38847 = ( ~w38738 & w38845 ) | ( ~w38738 & w38846 ) | ( w38845 & w38846 ) ;
  assign w38848 = w38846 | w38847 ;
  assign w38849 = \pi078 ^ w38723 ;
  assign w38850 = ( ~w38731 & w38848 ) | ( ~w38731 & w38849 ) | ( w38848 & w38849 ) ;
  assign w38851 = w38849 | w38850 ;
  assign w38852 = \pi079 ^ w38716 ;
  assign w38853 = ( ~w38724 & w38851 ) | ( ~w38724 & w38852 ) | ( w38851 & w38852 ) ;
  assign w38854 = w38852 | w38853 ;
  assign w38855 = \pi080 ^ w38709 ;
  assign w38856 = ( ~w38717 & w38854 ) | ( ~w38717 & w38855 ) | ( w38854 & w38855 ) ;
  assign w38857 = w38855 | w38856 ;
  assign w38858 = \pi081 ^ w38702 ;
  assign w38859 = ( ~w38710 & w38857 ) | ( ~w38710 & w38858 ) | ( w38857 & w38858 ) ;
  assign w38860 = w38858 | w38859 ;
  assign w38861 = \pi082 ^ w38695 ;
  assign w38862 = ( ~w38703 & w38860 ) | ( ~w38703 & w38861 ) | ( w38860 & w38861 ) ;
  assign w38863 = w38861 | w38862 ;
  assign w38864 = \pi083 ^ w38688 ;
  assign w38865 = ( ~w38696 & w38863 ) | ( ~w38696 & w38864 ) | ( w38863 & w38864 ) ;
  assign w38866 = w38864 | w38865 ;
  assign w38867 = \pi084 ^ w38681 ;
  assign w38868 = ( ~w38689 & w38866 ) | ( ~w38689 & w38867 ) | ( w38866 & w38867 ) ;
  assign w38869 = w38867 | w38868 ;
  assign w38870 = \pi085 ^ w38674 ;
  assign w38871 = ( ~w38682 & w38869 ) | ( ~w38682 & w38870 ) | ( w38869 & w38870 ) ;
  assign w38872 = w38870 | w38871 ;
  assign w38873 = \pi086 ^ w38667 ;
  assign w38874 = ( ~w38675 & w38872 ) | ( ~w38675 & w38873 ) | ( w38872 & w38873 ) ;
  assign w38875 = w38873 | w38874 ;
  assign w38876 = \pi087 ^ w38660 ;
  assign w38877 = ( ~w38668 & w38875 ) | ( ~w38668 & w38876 ) | ( w38875 & w38876 ) ;
  assign w38878 = w38876 | w38877 ;
  assign w38879 = \pi088 ^ w38653 ;
  assign w38880 = ( ~w38661 & w38878 ) | ( ~w38661 & w38879 ) | ( w38878 & w38879 ) ;
  assign w38881 = w38879 | w38880 ;
  assign w38882 = \pi089 ^ w38646 ;
  assign w38883 = ( ~w38654 & w38881 ) | ( ~w38654 & w38882 ) | ( w38881 & w38882 ) ;
  assign w38884 = w38882 | w38883 ;
  assign w38885 = \pi090 ^ w38639 ;
  assign w38886 = ( ~w38647 & w38884 ) | ( ~w38647 & w38885 ) | ( w38884 & w38885 ) ;
  assign w38887 = w38885 | w38886 ;
  assign w38888 = \pi091 ^ w38632 ;
  assign w38889 = ( ~w38640 & w38887 ) | ( ~w38640 & w38888 ) | ( w38887 & w38888 ) ;
  assign w38890 = w38888 | w38889 ;
  assign w38891 = \pi092 ^ w38625 ;
  assign w38892 = ( ~w38633 & w38890 ) | ( ~w38633 & w38891 ) | ( w38890 & w38891 ) ;
  assign w38893 = w38891 | w38892 ;
  assign w38894 = \pi093 ^ w38618 ;
  assign w38895 = ( ~w38626 & w38893 ) | ( ~w38626 & w38894 ) | ( w38893 & w38894 ) ;
  assign w38896 = w38894 | w38895 ;
  assign w38897 = \pi094 ^ w38611 ;
  assign w38898 = ( ~w38619 & w38896 ) | ( ~w38619 & w38897 ) | ( w38896 & w38897 ) ;
  assign w38899 = w38897 | w38898 ;
  assign w38900 = \pi095 ^ w38604 ;
  assign w38901 = ( ~w38612 & w38899 ) | ( ~w38612 & w38900 ) | ( w38899 & w38900 ) ;
  assign w38902 = w38900 | w38901 ;
  assign w38903 = \pi096 ^ w38597 ;
  assign w38904 = ( ~w38605 & w38902 ) | ( ~w38605 & w38903 ) | ( w38902 & w38903 ) ;
  assign w38905 = w38903 | w38904 ;
  assign w38906 = \pi097 ^ w38590 ;
  assign w38907 = ( ~w38598 & w38905 ) | ( ~w38598 & w38906 ) | ( w38905 & w38906 ) ;
  assign w38908 = w38906 | w38907 ;
  assign w38909 = \pi098 ^ w38583 ;
  assign w38910 = ( ~w38591 & w38908 ) | ( ~w38591 & w38909 ) | ( w38908 & w38909 ) ;
  assign w38911 = w38909 | w38910 ;
  assign w38912 = \pi099 ^ w38576 ;
  assign w38913 = ( ~w38584 & w38911 ) | ( ~w38584 & w38912 ) | ( w38911 & w38912 ) ;
  assign w38914 = w38912 | w38913 ;
  assign w38915 = \pi100 ^ w38569 ;
  assign w38916 = ( ~w38577 & w38914 ) | ( ~w38577 & w38915 ) | ( w38914 & w38915 ) ;
  assign w38917 = w38915 | w38916 ;
  assign w38918 = \pi101 ^ w38562 ;
  assign w38919 = ( ~w38570 & w38917 ) | ( ~w38570 & w38918 ) | ( w38917 & w38918 ) ;
  assign w38920 = w38918 | w38919 ;
  assign w38921 = \pi102 ^ w38555 ;
  assign w38922 = ( ~w38563 & w38920 ) | ( ~w38563 & w38921 ) | ( w38920 & w38921 ) ;
  assign w38923 = w38921 | w38922 ;
  assign w38924 = \pi103 ^ w38548 ;
  assign w38925 = ( ~w38556 & w38923 ) | ( ~w38556 & w38924 ) | ( w38923 & w38924 ) ;
  assign w38926 = w38924 | w38925 ;
  assign w38927 = \pi104 ^ w38541 ;
  assign w38928 = ( ~w38549 & w38926 ) | ( ~w38549 & w38927 ) | ( w38926 & w38927 ) ;
  assign w38929 = w38927 | w38928 ;
  assign w38930 = \pi105 ^ w38534 ;
  assign w38931 = ( ~w38542 & w38929 ) | ( ~w38542 & w38930 ) | ( w38929 & w38930 ) ;
  assign w38932 = w38930 | w38931 ;
  assign w38933 = \pi106 ^ w38527 ;
  assign w38934 = ( ~w38535 & w38932 ) | ( ~w38535 & w38933 ) | ( w38932 & w38933 ) ;
  assign w38935 = w38933 | w38934 ;
  assign w38936 = \pi107 ^ w38520 ;
  assign w38937 = ( ~w38528 & w38935 ) | ( ~w38528 & w38936 ) | ( w38935 & w38936 ) ;
  assign w38938 = w38936 | w38937 ;
  assign w38939 = \pi108 ^ w38513 ;
  assign w38940 = ( ~w38521 & w38938 ) | ( ~w38521 & w38939 ) | ( w38938 & w38939 ) ;
  assign w38941 = w38939 | w38940 ;
  assign w38942 = \pi109 ^ w38506 ;
  assign w38943 = ( ~w38514 & w38941 ) | ( ~w38514 & w38942 ) | ( w38941 & w38942 ) ;
  assign w38944 = w38942 | w38943 ;
  assign w38945 = \pi110 ^ w38499 ;
  assign w38946 = ( ~w38507 & w38944 ) | ( ~w38507 & w38945 ) | ( w38944 & w38945 ) ;
  assign w38947 = w38945 | w38946 ;
  assign w38948 = \pi111 ^ w38492 ;
  assign w38949 = ( ~w38500 & w38947 ) | ( ~w38500 & w38948 ) | ( w38947 & w38948 ) ;
  assign w38950 = w38948 | w38949 ;
  assign w38951 = \pi112 ^ w38485 ;
  assign w38952 = ( ~w38493 & w38950 ) | ( ~w38493 & w38951 ) | ( w38950 & w38951 ) ;
  assign w38953 = w38951 | w38952 ;
  assign w38954 = \pi113 ^ w38478 ;
  assign w38955 = ( ~w38486 & w38953 ) | ( ~w38486 & w38954 ) | ( w38953 & w38954 ) ;
  assign w38956 = w38954 | w38955 ;
  assign w38957 = \pi114 ^ w38471 ;
  assign w38958 = ( ~w38479 & w38956 ) | ( ~w38479 & w38957 ) | ( w38956 & w38957 ) ;
  assign w38959 = w38957 | w38958 ;
  assign w38960 = \pi115 ^ w38464 ;
  assign w38961 = ( ~w38472 & w38959 ) | ( ~w38472 & w38960 ) | ( w38959 & w38960 ) ;
  assign w38962 = w38960 | w38961 ;
  assign w38963 = \pi116 ^ w38457 ;
  assign w38964 = ( ~w38465 & w38962 ) | ( ~w38465 & w38963 ) | ( w38962 & w38963 ) ;
  assign w38965 = w38963 | w38964 ;
  assign w38966 = \pi117 ^ w38450 ;
  assign w38967 = ( ~w38458 & w38965 ) | ( ~w38458 & w38966 ) | ( w38965 & w38966 ) ;
  assign w38968 = w38966 | w38967 ;
  assign w38969 = \pi118 ^ w38443 ;
  assign w38970 = ( ~w38451 & w38968 ) | ( ~w38451 & w38969 ) | ( w38968 & w38969 ) ;
  assign w38971 = w38969 | w38970 ;
  assign w38972 = \pi119 ^ w38436 ;
  assign w38973 = ( ~w38444 & w38971 ) | ( ~w38444 & w38972 ) | ( w38971 & w38972 ) ;
  assign w38974 = w38972 | w38973 ;
  assign w38975 = \pi120 ^ w38429 ;
  assign w38976 = ( ~w38437 & w38974 ) | ( ~w38437 & w38975 ) | ( w38974 & w38975 ) ;
  assign w38977 = w38975 | w38976 ;
  assign w38978 = \pi121 ^ w38422 ;
  assign w38979 = ( ~w38430 & w38977 ) | ( ~w38430 & w38978 ) | ( w38977 & w38978 ) ;
  assign w38980 = w38978 | w38979 ;
  assign w38981 = \pi122 ^ w38415 ;
  assign w38982 = ( ~w38423 & w38980 ) | ( ~w38423 & w38981 ) | ( w38980 & w38981 ) ;
  assign w38983 = w38981 | w38982 ;
  assign w38984 = \pi123 ^ w38408 ;
  assign w38985 = ( ~w38416 & w38983 ) | ( ~w38416 & w38984 ) | ( w38983 & w38984 ) ;
  assign w38986 = w38984 | w38985 ;
  assign w38987 = \pi124 ^ w38401 ;
  assign w38988 = ( ~w38409 & w38986 ) | ( ~w38409 & w38987 ) | ( w38986 & w38987 ) ;
  assign w38989 = w38987 | w38988 ;
  assign w38990 = \pi125 ^ w38394 ;
  assign w38991 = ( ~w38402 & w38989 ) | ( ~w38402 & w38990 ) | ( w38989 & w38990 ) ;
  assign w38992 = w38990 | w38991 ;
  assign w38993 = w38379 | w38381 ;
  assign w38994 = ( ~w37785 & w38372 ) | ( ~w37785 & w38388 ) | ( w38372 & w38388 ) ;
  assign w38995 = w38993 ^ w38994 ;
  assign w38996 = ~w38388 & w38995 ;
  assign w38997 = ( w269 & ~w38378 ) | ( w269 & w38386 ) | ( ~w38378 & w38386 ) ;
  assign w38998 = w38378 & w38997 ;
  assign w38999 = w38996 | w38998 ;
  assign w39000 = ~\pi126 & w38999 ;
  assign w39001 = ( \pi126 & ~w38996 ) | ( \pi126 & w38998 ) | ( ~w38996 & w38998 ) ;
  assign w39002 = ~w38998 & w39001 ;
  assign w39003 = w39000 | w39002 ;
  assign w39004 = ( ~w38395 & w38992 ) | ( ~w38395 & w39003 ) | ( w38992 & w39003 ) ;
  assign w39005 = ( \pi127 & ~w39003 ) | ( \pi127 & w39004 ) | ( ~w39003 & w39004 ) ;
  assign w39006 = w39003 | w39005 ;
  assign w39007 = ( \pi126 & ~\pi127 ) | ( \pi126 & w38999 ) | ( ~\pi127 & w38999 ) ;
  assign w39008 = ~\pi126 & w39007 ;
  assign w39009 = w39006 & ~w39008 ;
  assign w39010 = ( ~w38395 & w38992 ) | ( ~w38395 & w39009 ) | ( w38992 & w39009 ) ;
  assign w39011 = w39003 ^ w39010 ;
  assign w39012 = ~w39009 & w39011 ;
  assign w39013 = ( w38999 & w39006 ) | ( w38999 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39014 = ~w39008 & w39013 ;
  assign w39015 = w39012 | w39014 ;
  assign w39016 = ~\pi127 & w39015 ;
  assign w39017 = ~w38402 & w38989 ;
  assign w39018 = w38990 ^ w39017 ;
  assign w39019 = ~w39009 & w39018 ;
  assign w39020 = ( w38394 & w39006 ) | ( w38394 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39021 = ~w39008 & w39020 ;
  assign w39022 = w39019 | w39021 ;
  assign w39023 = ~\pi126 & w39022 ;
  assign w39024 = ~w38409 & w38986 ;
  assign w39025 = w38987 ^ w39024 ;
  assign w39026 = ~w39009 & w39025 ;
  assign w39027 = ( w38401 & w39006 ) | ( w38401 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39028 = ~w39008 & w39027 ;
  assign w39029 = w39026 | w39028 ;
  assign w39030 = ~\pi125 & w39029 ;
  assign w39031 = ~w38416 & w38983 ;
  assign w39032 = w38984 ^ w39031 ;
  assign w39033 = ~w39009 & w39032 ;
  assign w39034 = ( w38408 & w39006 ) | ( w38408 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39035 = ~w39008 & w39034 ;
  assign w39036 = w39033 | w39035 ;
  assign w39037 = ~\pi124 & w39036 ;
  assign w39038 = ~w38423 & w38980 ;
  assign w39039 = w38981 ^ w39038 ;
  assign w39040 = ~w39009 & w39039 ;
  assign w39041 = ( w38415 & w39006 ) | ( w38415 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39042 = ~w39008 & w39041 ;
  assign w39043 = w39040 | w39042 ;
  assign w39044 = ~\pi123 & w39043 ;
  assign w39045 = ~w38430 & w38977 ;
  assign w39046 = w38978 ^ w39045 ;
  assign w39047 = ~w39009 & w39046 ;
  assign w39048 = ( w38422 & w39006 ) | ( w38422 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39049 = ~w39008 & w39048 ;
  assign w39050 = w39047 | w39049 ;
  assign w39051 = ~\pi122 & w39050 ;
  assign w39052 = ~w38437 & w38974 ;
  assign w39053 = w38975 ^ w39052 ;
  assign w39054 = ~w39009 & w39053 ;
  assign w39055 = ( w38429 & w39006 ) | ( w38429 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39056 = ~w39008 & w39055 ;
  assign w39057 = w39054 | w39056 ;
  assign w39058 = ~\pi121 & w39057 ;
  assign w39059 = ~w38444 & w38971 ;
  assign w39060 = w38972 ^ w39059 ;
  assign w39061 = ~w39009 & w39060 ;
  assign w39062 = ( w38436 & w39006 ) | ( w38436 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39063 = ~w39008 & w39062 ;
  assign w39064 = w39061 | w39063 ;
  assign w39065 = ~\pi120 & w39064 ;
  assign w39066 = ~w38451 & w38968 ;
  assign w39067 = w38969 ^ w39066 ;
  assign w39068 = ~w39009 & w39067 ;
  assign w39069 = ( w38443 & w39006 ) | ( w38443 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39070 = ~w39008 & w39069 ;
  assign w39071 = w39068 | w39070 ;
  assign w39072 = ~\pi119 & w39071 ;
  assign w39073 = ~w38458 & w38965 ;
  assign w39074 = w38966 ^ w39073 ;
  assign w39075 = ~w39009 & w39074 ;
  assign w39076 = ( w38450 & w39006 ) | ( w38450 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39077 = ~w39008 & w39076 ;
  assign w39078 = w39075 | w39077 ;
  assign w39079 = ~\pi118 & w39078 ;
  assign w39080 = ~w38465 & w38962 ;
  assign w39081 = w38963 ^ w39080 ;
  assign w39082 = ~w39009 & w39081 ;
  assign w39083 = ( w38457 & w39006 ) | ( w38457 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39084 = ~w39008 & w39083 ;
  assign w39085 = w39082 | w39084 ;
  assign w39086 = ~\pi117 & w39085 ;
  assign w39087 = ~w38472 & w38959 ;
  assign w39088 = w38960 ^ w39087 ;
  assign w39089 = ~w39009 & w39088 ;
  assign w39090 = ( w38464 & w39006 ) | ( w38464 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39091 = ~w39008 & w39090 ;
  assign w39092 = w39089 | w39091 ;
  assign w39093 = ~\pi116 & w39092 ;
  assign w39094 = ~w38479 & w38956 ;
  assign w39095 = w38957 ^ w39094 ;
  assign w39096 = ~w39009 & w39095 ;
  assign w39097 = ( w38471 & w39006 ) | ( w38471 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39098 = ~w39008 & w39097 ;
  assign w39099 = w39096 | w39098 ;
  assign w39100 = ~\pi115 & w39099 ;
  assign w39101 = ~w38486 & w38953 ;
  assign w39102 = w38954 ^ w39101 ;
  assign w39103 = ~w39009 & w39102 ;
  assign w39104 = ( w38478 & w39006 ) | ( w38478 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39105 = ~w39008 & w39104 ;
  assign w39106 = w39103 | w39105 ;
  assign w39107 = ~\pi114 & w39106 ;
  assign w39108 = ~w38493 & w38950 ;
  assign w39109 = w38951 ^ w39108 ;
  assign w39110 = ~w39009 & w39109 ;
  assign w39111 = ( w38485 & w39006 ) | ( w38485 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39112 = ~w39008 & w39111 ;
  assign w39113 = w39110 | w39112 ;
  assign w39114 = ~\pi113 & w39113 ;
  assign w39115 = ~w38500 & w38947 ;
  assign w39116 = w38948 ^ w39115 ;
  assign w39117 = ~w39009 & w39116 ;
  assign w39118 = ( w38492 & w39006 ) | ( w38492 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39119 = ~w39008 & w39118 ;
  assign w39120 = w39117 | w39119 ;
  assign w39121 = ~\pi112 & w39120 ;
  assign w39122 = ~w38507 & w38944 ;
  assign w39123 = w38945 ^ w39122 ;
  assign w39124 = ~w39009 & w39123 ;
  assign w39125 = ( w38499 & w39006 ) | ( w38499 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39126 = ~w39008 & w39125 ;
  assign w39127 = w39124 | w39126 ;
  assign w39128 = ~\pi111 & w39127 ;
  assign w39129 = ~w38514 & w38941 ;
  assign w39130 = w38942 ^ w39129 ;
  assign w39131 = ~w39009 & w39130 ;
  assign w39132 = ( w38506 & w39006 ) | ( w38506 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39133 = ~w39008 & w39132 ;
  assign w39134 = w39131 | w39133 ;
  assign w39135 = ~\pi110 & w39134 ;
  assign w39136 = ~w38521 & w38938 ;
  assign w39137 = w38939 ^ w39136 ;
  assign w39138 = ~w39009 & w39137 ;
  assign w39139 = ( w38513 & w39006 ) | ( w38513 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39140 = ~w39008 & w39139 ;
  assign w39141 = w39138 | w39140 ;
  assign w39142 = ~\pi109 & w39141 ;
  assign w39143 = ~w38528 & w38935 ;
  assign w39144 = w38936 ^ w39143 ;
  assign w39145 = ~w39009 & w39144 ;
  assign w39146 = ( w38520 & w39006 ) | ( w38520 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39147 = ~w39008 & w39146 ;
  assign w39148 = w39145 | w39147 ;
  assign w39149 = ~\pi108 & w39148 ;
  assign w39150 = ~w38535 & w38932 ;
  assign w39151 = w38933 ^ w39150 ;
  assign w39152 = ~w39009 & w39151 ;
  assign w39153 = ( w38527 & w39006 ) | ( w38527 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39154 = ~w39008 & w39153 ;
  assign w39155 = w39152 | w39154 ;
  assign w39156 = ~\pi107 & w39155 ;
  assign w39157 = ~w38542 & w38929 ;
  assign w39158 = w38930 ^ w39157 ;
  assign w39159 = ~w39009 & w39158 ;
  assign w39160 = ( w38534 & w39006 ) | ( w38534 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39161 = ~w39008 & w39160 ;
  assign w39162 = w39159 | w39161 ;
  assign w39163 = ~\pi106 & w39162 ;
  assign w39164 = ~w38549 & w38926 ;
  assign w39165 = w38927 ^ w39164 ;
  assign w39166 = ~w39009 & w39165 ;
  assign w39167 = ( w38541 & w39006 ) | ( w38541 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39168 = ~w39008 & w39167 ;
  assign w39169 = w39166 | w39168 ;
  assign w39170 = ~\pi105 & w39169 ;
  assign w39171 = ~w38556 & w38923 ;
  assign w39172 = w38924 ^ w39171 ;
  assign w39173 = ~w39009 & w39172 ;
  assign w39174 = ( w38548 & w39006 ) | ( w38548 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39175 = ~w39008 & w39174 ;
  assign w39176 = w39173 | w39175 ;
  assign w39177 = ~\pi104 & w39176 ;
  assign w39178 = ~w38563 & w38920 ;
  assign w39179 = w38921 ^ w39178 ;
  assign w39180 = ~w39009 & w39179 ;
  assign w39181 = ( w38555 & w39006 ) | ( w38555 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39182 = ~w39008 & w39181 ;
  assign w39183 = w39180 | w39182 ;
  assign w39184 = ~\pi103 & w39183 ;
  assign w39185 = ~w38570 & w38917 ;
  assign w39186 = w38918 ^ w39185 ;
  assign w39187 = ~w39009 & w39186 ;
  assign w39188 = ( w38562 & w39006 ) | ( w38562 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39189 = ~w39008 & w39188 ;
  assign w39190 = w39187 | w39189 ;
  assign w39191 = ~\pi102 & w39190 ;
  assign w39192 = ~w38577 & w38914 ;
  assign w39193 = w38915 ^ w39192 ;
  assign w39194 = ~w39009 & w39193 ;
  assign w39195 = ( w38569 & w39006 ) | ( w38569 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39196 = ~w39008 & w39195 ;
  assign w39197 = w39194 | w39196 ;
  assign w39198 = ~\pi101 & w39197 ;
  assign w39199 = ~w38584 & w38911 ;
  assign w39200 = w38912 ^ w39199 ;
  assign w39201 = ~w39009 & w39200 ;
  assign w39202 = ( w38576 & w39006 ) | ( w38576 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39203 = ~w39008 & w39202 ;
  assign w39204 = w39201 | w39203 ;
  assign w39205 = ~\pi100 & w39204 ;
  assign w39206 = ~w38591 & w38908 ;
  assign w39207 = w38909 ^ w39206 ;
  assign w39208 = ~w39009 & w39207 ;
  assign w39209 = ( w38583 & w39006 ) | ( w38583 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39210 = ~w39008 & w39209 ;
  assign w39211 = w39208 | w39210 ;
  assign w39212 = ~\pi099 & w39211 ;
  assign w39213 = ~w38598 & w38905 ;
  assign w39214 = w38906 ^ w39213 ;
  assign w39215 = ~w39009 & w39214 ;
  assign w39216 = ( w38590 & w39006 ) | ( w38590 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39217 = ~w39008 & w39216 ;
  assign w39218 = w39215 | w39217 ;
  assign w39219 = ~\pi098 & w39218 ;
  assign w39220 = ~w38605 & w38902 ;
  assign w39221 = w38903 ^ w39220 ;
  assign w39222 = ~w39009 & w39221 ;
  assign w39223 = ( w38597 & w39006 ) | ( w38597 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39224 = ~w39008 & w39223 ;
  assign w39225 = w39222 | w39224 ;
  assign w39226 = ~\pi097 & w39225 ;
  assign w39227 = ~w38612 & w38899 ;
  assign w39228 = w38900 ^ w39227 ;
  assign w39229 = ~w39009 & w39228 ;
  assign w39230 = ( w38604 & w39006 ) | ( w38604 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39231 = ~w39008 & w39230 ;
  assign w39232 = w39229 | w39231 ;
  assign w39233 = ~\pi096 & w39232 ;
  assign w39234 = ~w38619 & w38896 ;
  assign w39235 = w38897 ^ w39234 ;
  assign w39236 = ~w39009 & w39235 ;
  assign w39237 = ( w38611 & w39006 ) | ( w38611 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39238 = ~w39008 & w39237 ;
  assign w39239 = w39236 | w39238 ;
  assign w39240 = ~\pi095 & w39239 ;
  assign w39241 = ~w38626 & w38893 ;
  assign w39242 = w38894 ^ w39241 ;
  assign w39243 = ~w39009 & w39242 ;
  assign w39244 = ( w38618 & w39006 ) | ( w38618 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39245 = ~w39008 & w39244 ;
  assign w39246 = w39243 | w39245 ;
  assign w39247 = ~\pi094 & w39246 ;
  assign w39248 = ~w38633 & w38890 ;
  assign w39249 = w38891 ^ w39248 ;
  assign w39250 = ~w39009 & w39249 ;
  assign w39251 = ( w38625 & w39006 ) | ( w38625 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39252 = ~w39008 & w39251 ;
  assign w39253 = w39250 | w39252 ;
  assign w39254 = ~\pi093 & w39253 ;
  assign w39255 = ~w38640 & w38887 ;
  assign w39256 = w38888 ^ w39255 ;
  assign w39257 = ~w39009 & w39256 ;
  assign w39258 = ( w38632 & w39006 ) | ( w38632 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39259 = ~w39008 & w39258 ;
  assign w39260 = w39257 | w39259 ;
  assign w39261 = ~\pi092 & w39260 ;
  assign w39262 = ~w38647 & w38884 ;
  assign w39263 = w38885 ^ w39262 ;
  assign w39264 = ~w39009 & w39263 ;
  assign w39265 = ( w38639 & w39006 ) | ( w38639 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39266 = ~w39008 & w39265 ;
  assign w39267 = w39264 | w39266 ;
  assign w39268 = ~\pi091 & w39267 ;
  assign w39269 = ~w38654 & w38881 ;
  assign w39270 = w38882 ^ w39269 ;
  assign w39271 = ~w39009 & w39270 ;
  assign w39272 = ( w38646 & w39006 ) | ( w38646 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39273 = ~w39008 & w39272 ;
  assign w39274 = w39271 | w39273 ;
  assign w39275 = ~\pi090 & w39274 ;
  assign w39276 = ~w38661 & w38878 ;
  assign w39277 = w38879 ^ w39276 ;
  assign w39278 = ~w39009 & w39277 ;
  assign w39279 = ( w38653 & w39006 ) | ( w38653 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39280 = ~w39008 & w39279 ;
  assign w39281 = w39278 | w39280 ;
  assign w39282 = ~\pi089 & w39281 ;
  assign w39283 = ~w38668 & w38875 ;
  assign w39284 = w38876 ^ w39283 ;
  assign w39285 = ~w39009 & w39284 ;
  assign w39286 = ( w38660 & w39006 ) | ( w38660 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39287 = ~w39008 & w39286 ;
  assign w39288 = w39285 | w39287 ;
  assign w39289 = ~\pi088 & w39288 ;
  assign w39290 = ~w38675 & w38872 ;
  assign w39291 = w38873 ^ w39290 ;
  assign w39292 = ~w39009 & w39291 ;
  assign w39293 = ( w38667 & w39006 ) | ( w38667 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39294 = ~w39008 & w39293 ;
  assign w39295 = w39292 | w39294 ;
  assign w39296 = ~\pi087 & w39295 ;
  assign w39297 = ~w38682 & w38869 ;
  assign w39298 = w38870 ^ w39297 ;
  assign w39299 = ~w39009 & w39298 ;
  assign w39300 = ( w38674 & w39006 ) | ( w38674 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39301 = ~w39008 & w39300 ;
  assign w39302 = w39299 | w39301 ;
  assign w39303 = ~\pi086 & w39302 ;
  assign w39304 = ~w38689 & w38866 ;
  assign w39305 = w38867 ^ w39304 ;
  assign w39306 = ~w39009 & w39305 ;
  assign w39307 = ( w38681 & w39006 ) | ( w38681 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39308 = ~w39008 & w39307 ;
  assign w39309 = w39306 | w39308 ;
  assign w39310 = ~\pi085 & w39309 ;
  assign w39311 = ~w38696 & w38863 ;
  assign w39312 = w38864 ^ w39311 ;
  assign w39313 = ~w39009 & w39312 ;
  assign w39314 = ( w38688 & w39006 ) | ( w38688 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39315 = ~w39008 & w39314 ;
  assign w39316 = w39313 | w39315 ;
  assign w39317 = ~\pi084 & w39316 ;
  assign w39318 = ~w38703 & w38860 ;
  assign w39319 = w38861 ^ w39318 ;
  assign w39320 = ~w39009 & w39319 ;
  assign w39321 = ( w38695 & w39006 ) | ( w38695 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39322 = ~w39008 & w39321 ;
  assign w39323 = w39320 | w39322 ;
  assign w39324 = ~\pi083 & w39323 ;
  assign w39325 = ~w38710 & w38857 ;
  assign w39326 = w38858 ^ w39325 ;
  assign w39327 = ~w39009 & w39326 ;
  assign w39328 = ( w38702 & w39006 ) | ( w38702 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39329 = ~w39008 & w39328 ;
  assign w39330 = w39327 | w39329 ;
  assign w39331 = ~\pi082 & w39330 ;
  assign w39332 = ~w38717 & w38854 ;
  assign w39333 = w38855 ^ w39332 ;
  assign w39334 = ~w39009 & w39333 ;
  assign w39335 = ( w38709 & w39006 ) | ( w38709 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39336 = ~w39008 & w39335 ;
  assign w39337 = w39334 | w39336 ;
  assign w39338 = ~\pi081 & w39337 ;
  assign w39339 = ~w38724 & w38851 ;
  assign w39340 = w38852 ^ w39339 ;
  assign w39341 = ~w39009 & w39340 ;
  assign w39342 = ( w38716 & w39006 ) | ( w38716 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39343 = ~w39008 & w39342 ;
  assign w39344 = w39341 | w39343 ;
  assign w39345 = ~\pi080 & w39344 ;
  assign w39346 = ~w38731 & w38848 ;
  assign w39347 = w38849 ^ w39346 ;
  assign w39348 = ~w39009 & w39347 ;
  assign w39349 = ( w38723 & w39006 ) | ( w38723 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39350 = ~w39008 & w39349 ;
  assign w39351 = w39348 | w39350 ;
  assign w39352 = ~\pi079 & w39351 ;
  assign w39353 = ~w38738 & w38845 ;
  assign w39354 = w38846 ^ w39353 ;
  assign w39355 = ~w39009 & w39354 ;
  assign w39356 = ( w38730 & w39006 ) | ( w38730 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39357 = ~w39008 & w39356 ;
  assign w39358 = w39355 | w39357 ;
  assign w39359 = ~\pi078 & w39358 ;
  assign w39360 = ~w38745 & w38842 ;
  assign w39361 = w38843 ^ w39360 ;
  assign w39362 = ~w39009 & w39361 ;
  assign w39363 = ( w38737 & w39006 ) | ( w38737 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39364 = ~w39008 & w39363 ;
  assign w39365 = w39362 | w39364 ;
  assign w39366 = ~\pi077 & w39365 ;
  assign w39367 = ~w38752 & w38839 ;
  assign w39368 = w38840 ^ w39367 ;
  assign w39369 = ~w39009 & w39368 ;
  assign w39370 = ( w38744 & w39006 ) | ( w38744 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39371 = ~w39008 & w39370 ;
  assign w39372 = w39369 | w39371 ;
  assign w39373 = ~\pi076 & w39372 ;
  assign w39374 = ~w38759 & w38836 ;
  assign w39375 = w38837 ^ w39374 ;
  assign w39376 = ~w39009 & w39375 ;
  assign w39377 = ( w38751 & w39006 ) | ( w38751 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39378 = ~w39008 & w39377 ;
  assign w39379 = w39376 | w39378 ;
  assign w39380 = ~\pi075 & w39379 ;
  assign w39381 = ~w38766 & w38833 ;
  assign w39382 = w38834 ^ w39381 ;
  assign w39383 = ~w39009 & w39382 ;
  assign w39384 = ( w38758 & w39006 ) | ( w38758 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39385 = ~w39008 & w39384 ;
  assign w39386 = w39383 | w39385 ;
  assign w39387 = ~\pi074 & w39386 ;
  assign w39388 = ~w38773 & w38830 ;
  assign w39389 = w38831 ^ w39388 ;
  assign w39390 = ~w39009 & w39389 ;
  assign w39391 = ( w38765 & w39006 ) | ( w38765 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39392 = ~w39008 & w39391 ;
  assign w39393 = w39390 | w39392 ;
  assign w39394 = ~\pi073 & w39393 ;
  assign w39395 = ~w38780 & w38827 ;
  assign w39396 = w38828 ^ w39395 ;
  assign w39397 = ~w39009 & w39396 ;
  assign w39398 = ( w38772 & w39006 ) | ( w38772 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39399 = ~w39008 & w39398 ;
  assign w39400 = w39397 | w39399 ;
  assign w39401 = ~\pi072 & w39400 ;
  assign w39402 = ~w38787 & w38824 ;
  assign w39403 = w38825 ^ w39402 ;
  assign w39404 = ~w39009 & w39403 ;
  assign w39405 = ( w38779 & w39006 ) | ( w38779 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39406 = ~w39008 & w39405 ;
  assign w39407 = w39404 | w39406 ;
  assign w39408 = ~\pi071 & w39407 ;
  assign w39409 = ~w38794 & w38821 ;
  assign w39410 = w38822 ^ w39409 ;
  assign w39411 = ~w39009 & w39410 ;
  assign w39412 = ( w38786 & w39006 ) | ( w38786 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39413 = ~w39008 & w39412 ;
  assign w39414 = w39411 | w39413 ;
  assign w39415 = ~\pi070 & w39414 ;
  assign w39416 = ~w38803 & w38818 ;
  assign w39417 = w38819 ^ w39416 ;
  assign w39418 = ~w39009 & w39417 ;
  assign w39419 = ( w38793 & w39006 ) | ( w38793 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39420 = ~w39008 & w39419 ;
  assign w39421 = w39418 | w39420 ;
  assign w39422 = ~\pi069 & w39421 ;
  assign w39423 = ~w38810 & w38815 ;
  assign w39424 = w38816 ^ w39423 ;
  assign w39425 = ~w39009 & w39424 ;
  assign w39426 = ( w38802 & w39006 ) | ( w38802 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39427 = ~w39008 & w39426 ;
  assign w39428 = w39425 | w39427 ;
  assign w39429 = ~\pi068 & w39428 ;
  assign w39430 = \pi064 & ~w38388 ;
  assign w39431 = \pi002 ^ w39430 ;
  assign w39432 = ( \pi065 & w19790 ) | ( \pi065 & ~w39431 ) | ( w19790 & ~w39431 ) ;
  assign w39433 = w38811 ^ w39432 ;
  assign w39434 = ~w39009 & w39433 ;
  assign w39435 = ( w38809 & w39006 ) | ( w38809 & w39008 ) | ( w39006 & w39008 ) ;
  assign w39436 = ~w39008 & w39435 ;
  assign w39437 = w39434 | w39436 ;
  assign w39438 = ~\pi067 & w39437 ;
  assign w39439 = \pi001 ^ w38388 ;
  assign w39440 = ( \pi064 & w39009 ) | ( \pi064 & w39439 ) | ( w39009 & w39439 ) ;
  assign w39441 = w19795 ^ w39440 ;
  assign w39442 = ~w39009 & w39441 ;
  assign w39443 = w39009 & w39431 ;
  assign w39444 = w39442 | w39443 ;
  assign w39445 = ~\pi066 & w39444 ;
  assign w39446 = \pi066 ^ w39444 ;
  assign w39447 = ( \pi064 & ~w39009 ) | ( \pi064 & w39446 ) | ( ~w39009 & w39446 ) ;
  assign w39448 = \pi001 ^ w39447 ;
  assign w39449 = ( \pi065 & w19805 ) | ( \pi065 & ~w39448 ) | ( w19805 & ~w39448 ) ;
  assign w39450 = w39446 | w39449 ;
  assign w39451 = \pi067 ^ w39437 ;
  assign w39452 = ( ~w39445 & w39450 ) | ( ~w39445 & w39451 ) | ( w39450 & w39451 ) ;
  assign w39453 = w39451 | w39452 ;
  assign w39454 = \pi068 ^ w39428 ;
  assign w39455 = ( ~w39438 & w39453 ) | ( ~w39438 & w39454 ) | ( w39453 & w39454 ) ;
  assign w39456 = w39454 | w39455 ;
  assign w39457 = \pi069 ^ w39421 ;
  assign w39458 = ( ~w39429 & w39456 ) | ( ~w39429 & w39457 ) | ( w39456 & w39457 ) ;
  assign w39459 = w39457 | w39458 ;
  assign w39460 = \pi070 ^ w39414 ;
  assign w39461 = ( ~w39422 & w39459 ) | ( ~w39422 & w39460 ) | ( w39459 & w39460 ) ;
  assign w39462 = w39460 | w39461 ;
  assign w39463 = \pi071 ^ w39407 ;
  assign w39464 = ( ~w39415 & w39462 ) | ( ~w39415 & w39463 ) | ( w39462 & w39463 ) ;
  assign w39465 = w39463 | w39464 ;
  assign w39466 = \pi072 ^ w39400 ;
  assign w39467 = ( ~w39408 & w39465 ) | ( ~w39408 & w39466 ) | ( w39465 & w39466 ) ;
  assign w39468 = w39466 | w39467 ;
  assign w39469 = \pi073 ^ w39393 ;
  assign w39470 = ( ~w39401 & w39468 ) | ( ~w39401 & w39469 ) | ( w39468 & w39469 ) ;
  assign w39471 = w39469 | w39470 ;
  assign w39472 = \pi074 ^ w39386 ;
  assign w39473 = ( ~w39394 & w39471 ) | ( ~w39394 & w39472 ) | ( w39471 & w39472 ) ;
  assign w39474 = w39472 | w39473 ;
  assign w39475 = \pi075 ^ w39379 ;
  assign w39476 = ( ~w39387 & w39474 ) | ( ~w39387 & w39475 ) | ( w39474 & w39475 ) ;
  assign w39477 = w39475 | w39476 ;
  assign w39478 = \pi076 ^ w39372 ;
  assign w39479 = ( ~w39380 & w39477 ) | ( ~w39380 & w39478 ) | ( w39477 & w39478 ) ;
  assign w39480 = w39478 | w39479 ;
  assign w39481 = \pi077 ^ w39365 ;
  assign w39482 = ( ~w39373 & w39480 ) | ( ~w39373 & w39481 ) | ( w39480 & w39481 ) ;
  assign w39483 = w39481 | w39482 ;
  assign w39484 = \pi078 ^ w39358 ;
  assign w39485 = ( ~w39366 & w39483 ) | ( ~w39366 & w39484 ) | ( w39483 & w39484 ) ;
  assign w39486 = w39484 | w39485 ;
  assign w39487 = \pi079 ^ w39351 ;
  assign w39488 = ( ~w39359 & w39486 ) | ( ~w39359 & w39487 ) | ( w39486 & w39487 ) ;
  assign w39489 = w39487 | w39488 ;
  assign w39490 = \pi080 ^ w39344 ;
  assign w39491 = ( ~w39352 & w39489 ) | ( ~w39352 & w39490 ) | ( w39489 & w39490 ) ;
  assign w39492 = w39490 | w39491 ;
  assign w39493 = \pi081 ^ w39337 ;
  assign w39494 = ( ~w39345 & w39492 ) | ( ~w39345 & w39493 ) | ( w39492 & w39493 ) ;
  assign w39495 = w39493 | w39494 ;
  assign w39496 = \pi082 ^ w39330 ;
  assign w39497 = ( ~w39338 & w39495 ) | ( ~w39338 & w39496 ) | ( w39495 & w39496 ) ;
  assign w39498 = w39496 | w39497 ;
  assign w39499 = \pi083 ^ w39323 ;
  assign w39500 = ( ~w39331 & w39498 ) | ( ~w39331 & w39499 ) | ( w39498 & w39499 ) ;
  assign w39501 = w39499 | w39500 ;
  assign w39502 = \pi084 ^ w39316 ;
  assign w39503 = ( ~w39324 & w39501 ) | ( ~w39324 & w39502 ) | ( w39501 & w39502 ) ;
  assign w39504 = w39502 | w39503 ;
  assign w39505 = \pi085 ^ w39309 ;
  assign w39506 = ( ~w39317 & w39504 ) | ( ~w39317 & w39505 ) | ( w39504 & w39505 ) ;
  assign w39507 = w39505 | w39506 ;
  assign w39508 = \pi086 ^ w39302 ;
  assign w39509 = ( ~w39310 & w39507 ) | ( ~w39310 & w39508 ) | ( w39507 & w39508 ) ;
  assign w39510 = w39508 | w39509 ;
  assign w39511 = \pi087 ^ w39295 ;
  assign w39512 = ( ~w39303 & w39510 ) | ( ~w39303 & w39511 ) | ( w39510 & w39511 ) ;
  assign w39513 = w39511 | w39512 ;
  assign w39514 = \pi088 ^ w39288 ;
  assign w39515 = ( ~w39296 & w39513 ) | ( ~w39296 & w39514 ) | ( w39513 & w39514 ) ;
  assign w39516 = w39514 | w39515 ;
  assign w39517 = \pi089 ^ w39281 ;
  assign w39518 = ( ~w39289 & w39516 ) | ( ~w39289 & w39517 ) | ( w39516 & w39517 ) ;
  assign w39519 = w39517 | w39518 ;
  assign w39520 = \pi090 ^ w39274 ;
  assign w39521 = ( ~w39282 & w39519 ) | ( ~w39282 & w39520 ) | ( w39519 & w39520 ) ;
  assign w39522 = w39520 | w39521 ;
  assign w39523 = \pi091 ^ w39267 ;
  assign w39524 = ( ~w39275 & w39522 ) | ( ~w39275 & w39523 ) | ( w39522 & w39523 ) ;
  assign w39525 = w39523 | w39524 ;
  assign w39526 = \pi092 ^ w39260 ;
  assign w39527 = ( ~w39268 & w39525 ) | ( ~w39268 & w39526 ) | ( w39525 & w39526 ) ;
  assign w39528 = w39526 | w39527 ;
  assign w39529 = \pi093 ^ w39253 ;
  assign w39530 = ( ~w39261 & w39528 ) | ( ~w39261 & w39529 ) | ( w39528 & w39529 ) ;
  assign w39531 = w39529 | w39530 ;
  assign w39532 = \pi094 ^ w39246 ;
  assign w39533 = ( ~w39254 & w39531 ) | ( ~w39254 & w39532 ) | ( w39531 & w39532 ) ;
  assign w39534 = w39532 | w39533 ;
  assign w39535 = \pi095 ^ w39239 ;
  assign w39536 = ( ~w39247 & w39534 ) | ( ~w39247 & w39535 ) | ( w39534 & w39535 ) ;
  assign w39537 = w39535 | w39536 ;
  assign w39538 = \pi096 ^ w39232 ;
  assign w39539 = ( ~w39240 & w39537 ) | ( ~w39240 & w39538 ) | ( w39537 & w39538 ) ;
  assign w39540 = w39538 | w39539 ;
  assign w39541 = \pi097 ^ w39225 ;
  assign w39542 = ( ~w39233 & w39540 ) | ( ~w39233 & w39541 ) | ( w39540 & w39541 ) ;
  assign w39543 = w39541 | w39542 ;
  assign w39544 = \pi098 ^ w39218 ;
  assign w39545 = ( ~w39226 & w39543 ) | ( ~w39226 & w39544 ) | ( w39543 & w39544 ) ;
  assign w39546 = w39544 | w39545 ;
  assign w39547 = \pi099 ^ w39211 ;
  assign w39548 = ( ~w39219 & w39546 ) | ( ~w39219 & w39547 ) | ( w39546 & w39547 ) ;
  assign w39549 = w39547 | w39548 ;
  assign w39550 = \pi100 ^ w39204 ;
  assign w39551 = ( ~w39212 & w39549 ) | ( ~w39212 & w39550 ) | ( w39549 & w39550 ) ;
  assign w39552 = w39550 | w39551 ;
  assign w39553 = \pi101 ^ w39197 ;
  assign w39554 = ( ~w39205 & w39552 ) | ( ~w39205 & w39553 ) | ( w39552 & w39553 ) ;
  assign w39555 = w39553 | w39554 ;
  assign w39556 = \pi102 ^ w39190 ;
  assign w39557 = ( ~w39198 & w39555 ) | ( ~w39198 & w39556 ) | ( w39555 & w39556 ) ;
  assign w39558 = w39556 | w39557 ;
  assign w39559 = \pi103 ^ w39183 ;
  assign w39560 = ( ~w39191 & w39558 ) | ( ~w39191 & w39559 ) | ( w39558 & w39559 ) ;
  assign w39561 = w39559 | w39560 ;
  assign w39562 = \pi104 ^ w39176 ;
  assign w39563 = ( ~w39184 & w39561 ) | ( ~w39184 & w39562 ) | ( w39561 & w39562 ) ;
  assign w39564 = w39562 | w39563 ;
  assign w39565 = \pi105 ^ w39169 ;
  assign w39566 = ( ~w39177 & w39564 ) | ( ~w39177 & w39565 ) | ( w39564 & w39565 ) ;
  assign w39567 = w39565 | w39566 ;
  assign w39568 = \pi106 ^ w39162 ;
  assign w39569 = ( ~w39170 & w39567 ) | ( ~w39170 & w39568 ) | ( w39567 & w39568 ) ;
  assign w39570 = w39568 | w39569 ;
  assign w39571 = \pi107 ^ w39155 ;
  assign w39572 = ( ~w39163 & w39570 ) | ( ~w39163 & w39571 ) | ( w39570 & w39571 ) ;
  assign w39573 = w39571 | w39572 ;
  assign w39574 = \pi108 ^ w39148 ;
  assign w39575 = ( ~w39156 & w39573 ) | ( ~w39156 & w39574 ) | ( w39573 & w39574 ) ;
  assign w39576 = w39574 | w39575 ;
  assign w39577 = \pi109 ^ w39141 ;
  assign w39578 = ( ~w39149 & w39576 ) | ( ~w39149 & w39577 ) | ( w39576 & w39577 ) ;
  assign w39579 = w39577 | w39578 ;
  assign w39580 = \pi110 ^ w39134 ;
  assign w39581 = ( ~w39142 & w39579 ) | ( ~w39142 & w39580 ) | ( w39579 & w39580 ) ;
  assign w39582 = w39580 | w39581 ;
  assign w39583 = \pi111 ^ w39127 ;
  assign w39584 = ( ~w39135 & w39582 ) | ( ~w39135 & w39583 ) | ( w39582 & w39583 ) ;
  assign w39585 = w39583 | w39584 ;
  assign w39586 = \pi112 ^ w39120 ;
  assign w39587 = ( ~w39128 & w39585 ) | ( ~w39128 & w39586 ) | ( w39585 & w39586 ) ;
  assign w39588 = w39586 | w39587 ;
  assign w39589 = \pi113 ^ w39113 ;
  assign w39590 = ( ~w39121 & w39588 ) | ( ~w39121 & w39589 ) | ( w39588 & w39589 ) ;
  assign w39591 = w39589 | w39590 ;
  assign w39592 = \pi114 ^ w39106 ;
  assign w39593 = ( ~w39114 & w39591 ) | ( ~w39114 & w39592 ) | ( w39591 & w39592 ) ;
  assign w39594 = w39592 | w39593 ;
  assign w39595 = \pi115 ^ w39099 ;
  assign w39596 = ( ~w39107 & w39594 ) | ( ~w39107 & w39595 ) | ( w39594 & w39595 ) ;
  assign w39597 = w39595 | w39596 ;
  assign w39598 = \pi116 ^ w39092 ;
  assign w39599 = ( ~w39100 & w39597 ) | ( ~w39100 & w39598 ) | ( w39597 & w39598 ) ;
  assign w39600 = w39598 | w39599 ;
  assign w39601 = \pi117 ^ w39085 ;
  assign w39602 = ( ~w39093 & w39600 ) | ( ~w39093 & w39601 ) | ( w39600 & w39601 ) ;
  assign w39603 = w39601 | w39602 ;
  assign w39604 = \pi118 ^ w39078 ;
  assign w39605 = ( ~w39086 & w39603 ) | ( ~w39086 & w39604 ) | ( w39603 & w39604 ) ;
  assign w39606 = w39604 | w39605 ;
  assign w39607 = \pi119 ^ w39071 ;
  assign w39608 = ( ~w39079 & w39606 ) | ( ~w39079 & w39607 ) | ( w39606 & w39607 ) ;
  assign w39609 = w39607 | w39608 ;
  assign w39610 = \pi120 ^ w39064 ;
  assign w39611 = ( ~w39072 & w39609 ) | ( ~w39072 & w39610 ) | ( w39609 & w39610 ) ;
  assign w39612 = w39610 | w39611 ;
  assign w39613 = \pi121 ^ w39057 ;
  assign w39614 = ( ~w39065 & w39612 ) | ( ~w39065 & w39613 ) | ( w39612 & w39613 ) ;
  assign w39615 = w39613 | w39614 ;
  assign w39616 = \pi122 ^ w39050 ;
  assign w39617 = ( ~w39058 & w39615 ) | ( ~w39058 & w39616 ) | ( w39615 & w39616 ) ;
  assign w39618 = w39616 | w39617 ;
  assign w39619 = \pi123 ^ w39043 ;
  assign w39620 = ( ~w39051 & w39618 ) | ( ~w39051 & w39619 ) | ( w39618 & w39619 ) ;
  assign w39621 = w39619 | w39620 ;
  assign w39622 = \pi124 ^ w39036 ;
  assign w39623 = ( ~w39044 & w39621 ) | ( ~w39044 & w39622 ) | ( w39621 & w39622 ) ;
  assign w39624 = w39622 | w39623 ;
  assign w39625 = \pi125 ^ w39029 ;
  assign w39626 = ( ~w39037 & w39624 ) | ( ~w39037 & w39625 ) | ( w39624 & w39625 ) ;
  assign w39627 = w39625 | w39626 ;
  assign w39628 = \pi126 ^ w39022 ;
  assign w39629 = ( ~w39030 & w39627 ) | ( ~w39030 & w39628 ) | ( w39627 & w39628 ) ;
  assign w39630 = w39628 | w39629 ;
  assign w39631 = \pi127 ^ w39015 ;
  assign w39632 = ( ~w39023 & w39630 ) | ( ~w39023 & w39631 ) | ( w39630 & w39631 ) ;
  assign w39633 = w39631 | w39632 ;
  assign w39634 = w39016 & w39633 ;
  assign w39635 = ( \pi064 & ~w39633 ) | ( \pi064 & w39634 ) | ( ~w39633 & w39634 ) ;
  assign w39636 = \pi000 ^ w39635 ;
  assign w39637 = \pi001 ^ \pi065 ;
  assign w39638 = \pi000 ^ w39009 ;
  assign w39639 = \pi064 & w39638 ;
  assign w39640 = w39637 ^ w39639 ;
  assign w39641 = ( ~\pi064 & w39009 ) | ( ~\pi064 & w39633 ) | ( w39009 & w39633 ) ;
  assign w39642 = \pi001 ^ w39641 ;
  assign w39643 = ~w39016 & w39633 ;
  assign w39644 = w39642 ^ w39643 ;
  assign w39645 = ( w39640 & ~w39642 ) | ( w39640 & w39644 ) | ( ~w39642 & w39644 ) ;
  assign w39646 = \pi064 & ~w39009 ;
  assign w39647 = \pi001 ^ w39646 ;
  assign w39648 = ( \pi065 & w19805 ) | ( \pi065 & ~w39647 ) | ( w19805 & ~w39647 ) ;
  assign w39649 = w39446 ^ w39648 ;
  assign w39650 = w39643 ^ w39649 ;
  assign w39651 = ( w39444 & w39649 ) | ( w39444 & w39650 ) | ( w39649 & w39650 ) ;
  assign w39652 = ~w39445 & w39450 ;
  assign w39653 = w39451 ^ w39652 ;
  assign w39654 = w39437 ^ w39643 ;
  assign w39655 = ( w39437 & w39653 ) | ( w39437 & ~w39654 ) | ( w39653 & ~w39654 ) ;
  assign w39656 = ~w39438 & w39453 ;
  assign w39657 = w39454 ^ w39656 ;
  assign w39658 = w39428 ^ w39643 ;
  assign w39659 = ( w39428 & w39657 ) | ( w39428 & ~w39658 ) | ( w39657 & ~w39658 ) ;
  assign w39660 = ~w39429 & w39456 ;
  assign w39661 = w39457 ^ w39660 ;
  assign w39662 = w39421 ^ w39643 ;
  assign w39663 = ( w39421 & w39661 ) | ( w39421 & ~w39662 ) | ( w39661 & ~w39662 ) ;
  assign w39664 = ~w39422 & w39459 ;
  assign w39665 = w39460 ^ w39664 ;
  assign w39666 = w39414 ^ w39643 ;
  assign w39667 = ( w39414 & w39665 ) | ( w39414 & ~w39666 ) | ( w39665 & ~w39666 ) ;
  assign w39668 = ~w39415 & w39462 ;
  assign w39669 = w39463 ^ w39668 ;
  assign w39670 = w39407 ^ w39643 ;
  assign w39671 = ( w39407 & w39669 ) | ( w39407 & ~w39670 ) | ( w39669 & ~w39670 ) ;
  assign w39672 = ~w39408 & w39465 ;
  assign w39673 = w39466 ^ w39672 ;
  assign w39674 = w39400 ^ w39643 ;
  assign w39675 = ( w39400 & w39673 ) | ( w39400 & ~w39674 ) | ( w39673 & ~w39674 ) ;
  assign w39676 = ~w39401 & w39468 ;
  assign w39677 = w39469 ^ w39676 ;
  assign w39678 = w39393 ^ w39643 ;
  assign w39679 = ( w39393 & w39677 ) | ( w39393 & ~w39678 ) | ( w39677 & ~w39678 ) ;
  assign w39680 = ~w39394 & w39471 ;
  assign w39681 = w39472 ^ w39680 ;
  assign w39682 = w39386 ^ w39643 ;
  assign w39683 = ( w39386 & w39681 ) | ( w39386 & ~w39682 ) | ( w39681 & ~w39682 ) ;
  assign w39684 = ~w39387 & w39474 ;
  assign w39685 = w39475 ^ w39684 ;
  assign w39686 = w39379 ^ w39643 ;
  assign w39687 = ( w39379 & w39685 ) | ( w39379 & ~w39686 ) | ( w39685 & ~w39686 ) ;
  assign w39688 = ~w39380 & w39477 ;
  assign w39689 = w39478 ^ w39688 ;
  assign w39690 = w39372 ^ w39643 ;
  assign w39691 = ( w39372 & w39689 ) | ( w39372 & ~w39690 ) | ( w39689 & ~w39690 ) ;
  assign w39692 = ~w39373 & w39480 ;
  assign w39693 = w39481 ^ w39692 ;
  assign w39694 = w39365 ^ w39643 ;
  assign w39695 = ( w39365 & w39693 ) | ( w39365 & ~w39694 ) | ( w39693 & ~w39694 ) ;
  assign w39696 = ~w39366 & w39483 ;
  assign w39697 = w39484 ^ w39696 ;
  assign w39698 = w39358 ^ w39643 ;
  assign w39699 = ( w39358 & w39697 ) | ( w39358 & ~w39698 ) | ( w39697 & ~w39698 ) ;
  assign w39700 = ~w39359 & w39486 ;
  assign w39701 = w39487 ^ w39700 ;
  assign w39702 = w39351 ^ w39643 ;
  assign w39703 = ( w39351 & w39701 ) | ( w39351 & ~w39702 ) | ( w39701 & ~w39702 ) ;
  assign w39704 = ~w39352 & w39489 ;
  assign w39705 = w39490 ^ w39704 ;
  assign w39706 = w39344 ^ w39643 ;
  assign w39707 = ( w39344 & w39705 ) | ( w39344 & ~w39706 ) | ( w39705 & ~w39706 ) ;
  assign w39708 = ~w39345 & w39492 ;
  assign w39709 = w39493 ^ w39708 ;
  assign w39710 = w39337 ^ w39643 ;
  assign w39711 = ( w39337 & w39709 ) | ( w39337 & ~w39710 ) | ( w39709 & ~w39710 ) ;
  assign w39712 = ~w39338 & w39495 ;
  assign w39713 = w39496 ^ w39712 ;
  assign w39714 = w39330 ^ w39643 ;
  assign w39715 = ( w39330 & w39713 ) | ( w39330 & ~w39714 ) | ( w39713 & ~w39714 ) ;
  assign w39716 = ~w39331 & w39498 ;
  assign w39717 = w39499 ^ w39716 ;
  assign w39718 = w39323 ^ w39643 ;
  assign w39719 = ( w39323 & w39717 ) | ( w39323 & ~w39718 ) | ( w39717 & ~w39718 ) ;
  assign w39720 = ~w39324 & w39501 ;
  assign w39721 = w39502 ^ w39720 ;
  assign w39722 = w39316 ^ w39643 ;
  assign w39723 = ( w39316 & w39721 ) | ( w39316 & ~w39722 ) | ( w39721 & ~w39722 ) ;
  assign w39724 = ~w39317 & w39504 ;
  assign w39725 = w39505 ^ w39724 ;
  assign w39726 = w39309 ^ w39643 ;
  assign w39727 = ( w39309 & w39725 ) | ( w39309 & ~w39726 ) | ( w39725 & ~w39726 ) ;
  assign w39728 = ~w39310 & w39507 ;
  assign w39729 = w39508 ^ w39728 ;
  assign w39730 = w39302 ^ w39643 ;
  assign w39731 = ( w39302 & w39729 ) | ( w39302 & ~w39730 ) | ( w39729 & ~w39730 ) ;
  assign w39732 = ~w39303 & w39510 ;
  assign w39733 = w39511 ^ w39732 ;
  assign w39734 = w39295 ^ w39643 ;
  assign w39735 = ( w39295 & w39733 ) | ( w39295 & ~w39734 ) | ( w39733 & ~w39734 ) ;
  assign w39736 = ~w39296 & w39513 ;
  assign w39737 = w39514 ^ w39736 ;
  assign w39738 = w39288 ^ w39643 ;
  assign w39739 = ( w39288 & w39737 ) | ( w39288 & ~w39738 ) | ( w39737 & ~w39738 ) ;
  assign w39740 = ~w39289 & w39516 ;
  assign w39741 = w39517 ^ w39740 ;
  assign w39742 = w39281 ^ w39643 ;
  assign w39743 = ( w39281 & w39741 ) | ( w39281 & ~w39742 ) | ( w39741 & ~w39742 ) ;
  assign w39744 = ~w39282 & w39519 ;
  assign w39745 = w39520 ^ w39744 ;
  assign w39746 = w39274 ^ w39643 ;
  assign w39747 = ( w39274 & w39745 ) | ( w39274 & ~w39746 ) | ( w39745 & ~w39746 ) ;
  assign w39748 = ~w39275 & w39522 ;
  assign w39749 = w39523 ^ w39748 ;
  assign w39750 = w39267 ^ w39643 ;
  assign w39751 = ( w39267 & w39749 ) | ( w39267 & ~w39750 ) | ( w39749 & ~w39750 ) ;
  assign w39752 = ~w39268 & w39525 ;
  assign w39753 = w39526 ^ w39752 ;
  assign w39754 = w39260 ^ w39643 ;
  assign w39755 = ( w39260 & w39753 ) | ( w39260 & ~w39754 ) | ( w39753 & ~w39754 ) ;
  assign w39756 = ~w39261 & w39528 ;
  assign w39757 = w39529 ^ w39756 ;
  assign w39758 = w39253 ^ w39643 ;
  assign w39759 = ( w39253 & w39757 ) | ( w39253 & ~w39758 ) | ( w39757 & ~w39758 ) ;
  assign w39760 = ~w39254 & w39531 ;
  assign w39761 = w39532 ^ w39760 ;
  assign w39762 = w39246 ^ w39643 ;
  assign w39763 = ( w39246 & w39761 ) | ( w39246 & ~w39762 ) | ( w39761 & ~w39762 ) ;
  assign w39764 = ~w39247 & w39534 ;
  assign w39765 = w39535 ^ w39764 ;
  assign w39766 = w39239 ^ w39643 ;
  assign w39767 = ( w39239 & w39765 ) | ( w39239 & ~w39766 ) | ( w39765 & ~w39766 ) ;
  assign w39768 = ~w39240 & w39537 ;
  assign w39769 = w39538 ^ w39768 ;
  assign w39770 = w39232 ^ w39643 ;
  assign w39771 = ( w39232 & w39769 ) | ( w39232 & ~w39770 ) | ( w39769 & ~w39770 ) ;
  assign w39772 = ~w39233 & w39540 ;
  assign w39773 = w39541 ^ w39772 ;
  assign w39774 = w39225 ^ w39643 ;
  assign w39775 = ( w39225 & w39773 ) | ( w39225 & ~w39774 ) | ( w39773 & ~w39774 ) ;
  assign w39776 = ~w39226 & w39543 ;
  assign w39777 = w39544 ^ w39776 ;
  assign w39778 = w39218 ^ w39643 ;
  assign w39779 = ( w39218 & w39777 ) | ( w39218 & ~w39778 ) | ( w39777 & ~w39778 ) ;
  assign w39780 = ~w39219 & w39546 ;
  assign w39781 = w39547 ^ w39780 ;
  assign w39782 = w39211 ^ w39643 ;
  assign w39783 = ( w39211 & w39781 ) | ( w39211 & ~w39782 ) | ( w39781 & ~w39782 ) ;
  assign w39784 = ~w39212 & w39549 ;
  assign w39785 = w39550 ^ w39784 ;
  assign w39786 = w39204 ^ w39643 ;
  assign w39787 = ( w39204 & w39785 ) | ( w39204 & ~w39786 ) | ( w39785 & ~w39786 ) ;
  assign w39788 = ~w39205 & w39552 ;
  assign w39789 = w39553 ^ w39788 ;
  assign w39790 = w39197 ^ w39643 ;
  assign w39791 = ( w39197 & w39789 ) | ( w39197 & ~w39790 ) | ( w39789 & ~w39790 ) ;
  assign w39792 = ~w39198 & w39555 ;
  assign w39793 = w39556 ^ w39792 ;
  assign w39794 = w39190 ^ w39643 ;
  assign w39795 = ( w39190 & w39793 ) | ( w39190 & ~w39794 ) | ( w39793 & ~w39794 ) ;
  assign w39796 = ~w39191 & w39558 ;
  assign w39797 = w39559 ^ w39796 ;
  assign w39798 = w39183 ^ w39643 ;
  assign w39799 = ( w39183 & w39797 ) | ( w39183 & ~w39798 ) | ( w39797 & ~w39798 ) ;
  assign w39800 = ~w39184 & w39561 ;
  assign w39801 = w39562 ^ w39800 ;
  assign w39802 = w39176 ^ w39643 ;
  assign w39803 = ( w39176 & w39801 ) | ( w39176 & ~w39802 ) | ( w39801 & ~w39802 ) ;
  assign w39804 = ~w39177 & w39564 ;
  assign w39805 = w39565 ^ w39804 ;
  assign w39806 = w39169 ^ w39643 ;
  assign w39807 = ( w39169 & w39805 ) | ( w39169 & ~w39806 ) | ( w39805 & ~w39806 ) ;
  assign w39808 = ~w39170 & w39567 ;
  assign w39809 = w39568 ^ w39808 ;
  assign w39810 = w39162 ^ w39643 ;
  assign w39811 = ( w39162 & w39809 ) | ( w39162 & ~w39810 ) | ( w39809 & ~w39810 ) ;
  assign w39812 = ~w39163 & w39570 ;
  assign w39813 = w39571 ^ w39812 ;
  assign w39814 = w39155 ^ w39643 ;
  assign w39815 = ( w39155 & w39813 ) | ( w39155 & ~w39814 ) | ( w39813 & ~w39814 ) ;
  assign w39816 = ~w39156 & w39573 ;
  assign w39817 = w39574 ^ w39816 ;
  assign w39818 = w39148 ^ w39643 ;
  assign w39819 = ( w39148 & w39817 ) | ( w39148 & ~w39818 ) | ( w39817 & ~w39818 ) ;
  assign w39820 = ~w39149 & w39576 ;
  assign w39821 = w39577 ^ w39820 ;
  assign w39822 = w39141 ^ w39643 ;
  assign w39823 = ( w39141 & w39821 ) | ( w39141 & ~w39822 ) | ( w39821 & ~w39822 ) ;
  assign w39824 = ~w39142 & w39579 ;
  assign w39825 = w39580 ^ w39824 ;
  assign w39826 = w39134 ^ w39643 ;
  assign w39827 = ( w39134 & w39825 ) | ( w39134 & ~w39826 ) | ( w39825 & ~w39826 ) ;
  assign w39828 = ~w39135 & w39582 ;
  assign w39829 = w39583 ^ w39828 ;
  assign w39830 = w39127 ^ w39643 ;
  assign w39831 = ( w39127 & w39829 ) | ( w39127 & ~w39830 ) | ( w39829 & ~w39830 ) ;
  assign w39832 = ~w39128 & w39585 ;
  assign w39833 = w39586 ^ w39832 ;
  assign w39834 = w39120 ^ w39643 ;
  assign w39835 = ( w39120 & w39833 ) | ( w39120 & ~w39834 ) | ( w39833 & ~w39834 ) ;
  assign w39836 = ~w39121 & w39588 ;
  assign w39837 = w39589 ^ w39836 ;
  assign w39838 = w39113 ^ w39643 ;
  assign w39839 = ( w39113 & w39837 ) | ( w39113 & ~w39838 ) | ( w39837 & ~w39838 ) ;
  assign w39840 = ~w39114 & w39591 ;
  assign w39841 = w39592 ^ w39840 ;
  assign w39842 = w39106 ^ w39643 ;
  assign w39843 = ( w39106 & w39841 ) | ( w39106 & ~w39842 ) | ( w39841 & ~w39842 ) ;
  assign w39844 = ~w39107 & w39594 ;
  assign w39845 = w39595 ^ w39844 ;
  assign w39846 = w39099 ^ w39643 ;
  assign w39847 = ( w39099 & w39845 ) | ( w39099 & ~w39846 ) | ( w39845 & ~w39846 ) ;
  assign w39848 = ~w39100 & w39597 ;
  assign w39849 = w39598 ^ w39848 ;
  assign w39850 = w39092 ^ w39643 ;
  assign w39851 = ( w39092 & w39849 ) | ( w39092 & ~w39850 ) | ( w39849 & ~w39850 ) ;
  assign w39852 = ~w39093 & w39600 ;
  assign w39853 = w39601 ^ w39852 ;
  assign w39854 = w39085 ^ w39643 ;
  assign w39855 = ( w39085 & w39853 ) | ( w39085 & ~w39854 ) | ( w39853 & ~w39854 ) ;
  assign w39856 = ~w39086 & w39603 ;
  assign w39857 = w39604 ^ w39856 ;
  assign w39858 = w39078 ^ w39643 ;
  assign w39859 = ( w39078 & w39857 ) | ( w39078 & ~w39858 ) | ( w39857 & ~w39858 ) ;
  assign w39860 = ~w39079 & w39606 ;
  assign w39861 = w39607 ^ w39860 ;
  assign w39862 = w39071 ^ w39643 ;
  assign w39863 = ( w39071 & w39861 ) | ( w39071 & ~w39862 ) | ( w39861 & ~w39862 ) ;
  assign w39864 = ~w39072 & w39609 ;
  assign w39865 = w39610 ^ w39864 ;
  assign w39866 = w39064 ^ w39643 ;
  assign w39867 = ( w39064 & w39865 ) | ( w39064 & ~w39866 ) | ( w39865 & ~w39866 ) ;
  assign w39868 = ~w39065 & w39612 ;
  assign w39869 = w39613 ^ w39868 ;
  assign w39870 = w39057 ^ w39643 ;
  assign w39871 = ( w39057 & w39869 ) | ( w39057 & ~w39870 ) | ( w39869 & ~w39870 ) ;
  assign w39872 = ~w39058 & w39615 ;
  assign w39873 = w39616 ^ w39872 ;
  assign w39874 = w39050 ^ w39643 ;
  assign w39875 = ( w39050 & w39873 ) | ( w39050 & ~w39874 ) | ( w39873 & ~w39874 ) ;
  assign w39876 = ~w39051 & w39618 ;
  assign w39877 = w39619 ^ w39876 ;
  assign w39878 = w39043 ^ w39643 ;
  assign w39879 = ( w39043 & w39877 ) | ( w39043 & ~w39878 ) | ( w39877 & ~w39878 ) ;
  assign w39880 = ~w39044 & w39621 ;
  assign w39881 = w39622 ^ w39880 ;
  assign w39882 = w39036 ^ w39643 ;
  assign w39883 = ( w39036 & w39881 ) | ( w39036 & ~w39882 ) | ( w39881 & ~w39882 ) ;
  assign w39884 = ~w39037 & w39624 ;
  assign w39885 = w39625 ^ w39884 ;
  assign w39886 = w39029 ^ w39643 ;
  assign w39887 = ( w39029 & w39885 ) | ( w39029 & ~w39886 ) | ( w39885 & ~w39886 ) ;
  assign w39888 = ~w39030 & w39627 ;
  assign w39889 = w39628 ^ w39888 ;
  assign w39890 = w39022 ^ w39643 ;
  assign w39891 = ( w39022 & w39889 ) | ( w39022 & ~w39890 ) | ( w39889 & ~w39890 ) ;
  assign w39892 = ~w39023 & w39630 ;
  assign w39893 = ( ~w39015 & w39631 ) | ( ~w39015 & w39892 ) | ( w39631 & w39892 ) ;
  assign w39894 = ( \pi127 & w39015 ) | ( \pi127 & ~w39892 ) | ( w39015 & ~w39892 ) ;
  assign w39895 = w39631 & w39894 ;
  assign w39896 = ( w39892 & ~w39893 ) | ( w39892 & w39895 ) | ( ~w39893 & w39895 ) ;
  assign \po000 = ~w20150 ;
  assign \po001 = ~w19673 ;
  assign \po002 = ~w19054 ;
  assign \po003 = ~w18443 ;
  assign \po004 = ~w17843 ;
  assign \po005 = ~w17250 ;
  assign \po006 = ~w16708 ;
  assign \po007 = ~w16139 ;
  assign \po008 = ~w15578 ;
  assign \po009 = ~w15064 ;
  assign \po010 = ~w14524 ;
  assign \po011 = ~w13994 ;
  assign \po012 = ~w13509 ;
  assign \po013 = ~w13002 ;
  assign \po014 = ~w12502 ;
  assign \po015 = ~w12039 ;
  assign \po016 = ~w11562 ;
  assign \po017 = ~w11093 ;
  assign \po018 = ~w10651 ;
  assign \po019 = ~w10200 ;
  assign \po020 = ~w9756 ;
  assign \po021 = ~w9352 ;
  assign \po022 = ~w8931 ;
  assign \po023 = ~w8544 ;
  assign \po024 = ~w8170 ;
  assign \po025 = ~w7783 ;
  assign \po026 = ~w7420 ;
  assign \po027 = ~w7066 ;
  assign \po028 = ~w6710 ;
  assign \po029 = ~w6380 ;
  assign \po030 = ~w6048 ;
  assign \po031 = ~w5716 ;
  assign \po032 = ~w5416 ;
  assign \po033 = ~w5118 ;
  assign \po034 = ~w4816 ;
  assign \po035 = ~w4536 ;
  assign \po036 = ~w4267 ;
  assign \po037 = ~w3999 ;
  assign \po038 = ~w3744 ;
  assign \po039 = ~w3495 ;
  assign \po040 = ~w3255 ;
  assign \po041 = ~w3026 ;
  assign \po042 = ~w2800 ;
  assign \po043 = ~w2587 ;
  assign \po044 = ~w2390 ;
  assign \po045 = ~w2198 ;
  assign \po046 = ~w2017 ;
  assign \po047 = ~w1842 ;
  assign \po048 = ~w1683 ;
  assign \po049 = ~w1534 ;
  assign \po050 = ~w1385 ;
  assign \po051 = ~w1246 ;
  assign \po052 = ~w1124 ;
  assign \po053 = ~w1008 ;
  assign \po054 = ~w890 ;
  assign \po055 = ~w795 ;
  assign \po056 = ~w704 ;
  assign \po057 = ~w613 ;
  assign \po058 = ~w551 ;
  assign \po059 = ~w20151 ;
  assign \po060 = ~w373 ;
  assign \po061 = ~w310 ;
  assign \po062 = ~w20153 ;
  assign \po063 = ~w20159 ;
  assign \po064 = w39636 ;
  assign \po065 = w39645 ;
  assign \po066 = w39651 ;
  assign \po067 = w39655 ;
  assign \po068 = w39659 ;
  assign \po069 = w39663 ;
  assign \po070 = w39667 ;
  assign \po071 = w39671 ;
  assign \po072 = w39675 ;
  assign \po073 = w39679 ;
  assign \po074 = w39683 ;
  assign \po075 = w39687 ;
  assign \po076 = w39691 ;
  assign \po077 = w39695 ;
  assign \po078 = w39699 ;
  assign \po079 = w39703 ;
  assign \po080 = w39707 ;
  assign \po081 = w39711 ;
  assign \po082 = w39715 ;
  assign \po083 = w39719 ;
  assign \po084 = w39723 ;
  assign \po085 = w39727 ;
  assign \po086 = w39731 ;
  assign \po087 = w39735 ;
  assign \po088 = w39739 ;
  assign \po089 = w39743 ;
  assign \po090 = w39747 ;
  assign \po091 = w39751 ;
  assign \po092 = w39755 ;
  assign \po093 = w39759 ;
  assign \po094 = w39763 ;
  assign \po095 = w39767 ;
  assign \po096 = w39771 ;
  assign \po097 = w39775 ;
  assign \po098 = w39779 ;
  assign \po099 = w39783 ;
  assign \po100 = w39787 ;
  assign \po101 = w39791 ;
  assign \po102 = w39795 ;
  assign \po103 = w39799 ;
  assign \po104 = w39803 ;
  assign \po105 = w39807 ;
  assign \po106 = w39811 ;
  assign \po107 = w39815 ;
  assign \po108 = w39819 ;
  assign \po109 = w39823 ;
  assign \po110 = w39827 ;
  assign \po111 = w39831 ;
  assign \po112 = w39835 ;
  assign \po113 = w39839 ;
  assign \po114 = w39843 ;
  assign \po115 = w39847 ;
  assign \po116 = w39851 ;
  assign \po117 = w39855 ;
  assign \po118 = w39859 ;
  assign \po119 = w39863 ;
  assign \po120 = w39867 ;
  assign \po121 = w39871 ;
  assign \po122 = w39875 ;
  assign \po123 = w39879 ;
  assign \po124 = w39883 ;
  assign \po125 = w39887 ;
  assign \po126 = w39891 ;
  assign \po127 = w39896 ;
endmodule
