module log2( \pi00 , \pi01 , \pi02 , \pi03 , \pi04 , \pi05 , \pi06 , \pi07 , \pi08 , \pi09 , \pi10 , \pi11 , \pi12 , \pi13 , \pi14 , \pi15 , \pi16 , \pi17 , \pi18 , \pi19 , \pi20 , \pi21 , \pi22 , \pi23 , \pi24 , \pi25 , \pi26 , \pi27 , \pi28 , \pi29 , \pi30 , \pi31 , \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po23 , \po24 , \po25 , \po26 , \po27 , \po28 , \po29 , \po30 , \po31 );
  input \pi00 , \pi01 , \pi02 , \pi03 , \pi04 , \pi05 , \pi06 , \pi07 , \pi08 , \pi09 , \pi10 , \pi11 , \pi12 , \pi13 , \pi14 , \pi15 , \pi16 , \pi17 , \pi18 , \pi19 , \pi20 , \pi21 , \pi22 , \pi23 , \pi24 , \pi25 , \pi26 , \pi27 , \pi28 , \pi29 , \pi30 , \pi31 ;
  output \po00 , \po01 , \po02 , \po03 , \po04 , \po05 , \po06 , \po07 , \po08 , \po09 , \po10 , \po11 , \po12 , \po13 , \po14 , \po15 , \po16 , \po17 , \po18 , \po19 , \po20 , \po21 , \po22 , \po23 , \po24 , \po25 , \po26 , \po27 , \po28 , \po29 , \po30 , \po31 ;
  wire zero , w33 , w34 , w35 , w36 , w37 , w38 , w39 , w40 , w41 , w42 , w43 , w44 , w45 , w46 , w47 , w48 , w49 , w50 , w51 , w52 , w53 , w54 , w55 , w56 , w57 , w58 , w59 , w60 , w61 , w62 , w63 , w64 , w65 , w66 , w67 , w68 , w69 , w70 , w71 , w72 , w73 , w74 , w75 , w76 , w77 , w78 , w79 , w80 , w81 , w82 , w83 , w84 , w85 , w86 , w87 , w88 , w89 , w90 , w91 , w92 , w93 , w94 , w95 , w96 , w97 , w98 , w99 , w100 , w101 , w102 , w103 , w104 , w105 , w106 , w107 , w108 , w109 , w110 , w111 , w112 , w113 , w114 , w115 , w116 , w117 , w118 , w119 , w120 , w121 , w122 , w123 , w124 , w125 , w126 , w127 , w128 , w129 , w130 , w131 , w132 , w133 , w134 , w135 , w136 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w146 , w147 , w148 , w149 , w150 , w151 , w152 , w153 , w154 , w155 , w156 , w157 , w158 , w159 , w160 , w161 , w162 , w163 , w164 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w174 , w175 , w176 , w177 , w178 , w179 , w180 , w181 , w182 , w183 , w184 , w185 , w186 , w187 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w203 , w204 , w205 , w206 , w207 , w208 , w209 , w210 , w211 , w212 , w213 , w214 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w224 , w225 , w226 , w227 , w228 , w229 , w230 , w231 , w232 , w233 , w234 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w250 , w251 , w252 , w253 , w254 , w255 , w256 , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 , w2495 , w2496 , w2497 , w2498 , w2499 , w2500 , w2501 , w2502 , w2503 , w2504 , w2505 , w2506 , w2507 , w2508 , w2509 , w2510 , w2511 , w2512 , w2513 , w2514 , w2515 , w2516 , w2517 , w2518 , w2519 , w2520 , w2521 , w2522 , w2523 , w2524 , w2525 , w2526 , w2527 , w2528 , w2529 , w2530 , w2531 , w2532 , w2533 , w2534 , w2535 , w2536 , w2537 , w2538 , w2539 , w2540 , w2541 , w2542 , w2543 , w2544 , w2545 , w2546 , w2547 , w2548 , w2549 , w2550 , w2551 , w2552 , w2553 , w2554 , w2555 , w2556 , w2557 , w2558 , w2559 , w2560 , w2561 , w2562 , w2563 , w2564 , w2565 , w2566 , w2567 , w2568 , w2569 , w2570 , w2571 , w2572 , w2573 , w2574 , w2575 , w2576 , w2577 , w2578 , w2579 , w2580 , w2581 , w2582 , w2583 , w2584 , w2585 , w2586 , w2587 , w2588 , w2589 , w2590 , w2591 , w2592 , w2593 , w2594 , w2595 , w2596 , w2597 , w2598 , w2599 , w2600 , w2601 , w2602 , w2603 , w2604 , w2605 , w2606 , w2607 , w2608 , w2609 , w2610 , w2611 , w2612 , w2613 , w2614 , w2615 , w2616 , w2617 , w2618 , w2619 , w2620 , w2621 , w2622 , w2623 , w2624 , w2625 , w2626 , w2627 , w2628 , w2629 , w2630 , w2631 , w2632 , w2633 , w2634 , w2635 , w2636 , w2637 , w2638 , w2639 , w2640 , w2641 , w2642 , w2643 , w2644 , w2645 , w2646 , w2647 , w2648 , w2649 , w2650 , w2651 , w2652 , w2653 , w2654 , w2655 , w2656 , w2657 , w2658 , w2659 , w2660 , w2661 , w2662 , w2663 , w2664 , w2665 , w2666 , w2667 , w2668 , w2669 , w2670 , w2671 , w2672 , w2673 , w2674 , w2675 , w2676 , w2677 , w2678 , w2679 , w2680 , w2681 , w2682 , w2683 , w2684 , w2685 , w2686 , w2687 , w2688 , w2689 , w2690 , w2691 , w2692 , w2693 , w2694 , w2695 , w2696 , w2697 , w2698 , w2699 , w2700 , w2701 , w2702 , w2703 , w2704 , w2705 , w2706 , w2707 , w2708 , w2709 , w2710 , w2711 , w2712 , w2713 , w2714 , w2715 , w2716 , w2717 , w2718 , w2719 , w2720 , w2721 , w2722 , w2723 , w2724 , w2725 , w2726 , w2727 , w2728 , w2729 , w2730 , w2731 , w2732 , w2733 , w2734 , w2735 , w2736 , w2737 , w2738 , w2739 , w2740 , w2741 , w2742 , w2743 , w2744 , w2745 , w2746 , w2747 , w2748 , w2749 , w2750 , w2751 , w2752 , w2753 , w2754 , w2755 , w2756 , w2757 , w2758 , w2759 , w2760 , w2761 , w2762 , w2763 , w2764 , w2765 , w2766 , w2767 , w2768 , w2769 , w2770 , w2771 , w2772 , w2773 , w2774 , w2775 , w2776 , w2777 , w2778 , w2779 , w2780 , w2781 , w2782 , w2783 , w2784 , w2785 , w2786 , w2787 , w2788 , w2789 , w2790 , w2791 , w2792 , w2793 , w2794 , w2795 , w2796 , w2797 , w2798 , w2799 , w2800 , w2801 , w2802 , w2803 , w2804 , w2805 , w2806 , w2807 , w2808 , w2809 , w2810 , w2811 , w2812 , w2813 , w2814 , w2815 , w2816 , w2817 , w2818 , w2819 , w2820 , w2821 , w2822 , w2823 , w2824 , w2825 , w2826 , w2827 , w2828 , w2829 , w2830 , w2831 , w2832 , w2833 , w2834 , w2835 , w2836 , w2837 , w2838 , w2839 , w2840 , w2841 , w2842 , w2843 , w2844 , w2845 , w2846 , w2847 , w2848 , w2849 , w2850 , w2851 , w2852 , w2853 , w2854 , w2855 , w2856 , w2857 , w2858 , w2859 , w2860 , w2861 , w2862 , w2863 , w2864 , w2865 , w2866 , w2867 , w2868 , w2869 , w2870 , w2871 , w2872 , w2873 , w2874 , w2875 , w2876 , w2877 , w2878 , w2879 , w2880 , w2881 , w2882 , w2883 , w2884 , w2885 , w2886 , w2887 , w2888 , w2889 , w2890 , w2891 , w2892 , w2893 , w2894 , w2895 , w2896 , w2897 , w2898 , w2899 , w2900 , w2901 , w2902 , w2903 , w2904 , w2905 , w2906 , w2907 , w2908 , w2909 , w2910 , w2911 , w2912 , w2913 , w2914 , w2915 , w2916 , w2917 , w2918 , w2919 , w2920 , w2921 , w2922 , w2923 , w2924 , w2925 , w2926 , w2927 , w2928 , w2929 , w2930 , w2931 , w2932 , w2933 , w2934 , w2935 , w2936 , w2937 , w2938 , w2939 , w2940 , w2941 , w2942 , w2943 , w2944 , w2945 , w2946 , w2947 , w2948 , w2949 , w2950 , w2951 , w2952 , w2953 , w2954 , w2955 , w2956 , w2957 , w2958 , w2959 , w2960 , w2961 , w2962 , w2963 , w2964 , w2965 , w2966 , w2967 , w2968 , w2969 , w2970 , w2971 , w2972 , w2973 , w2974 , w2975 , w2976 , w2977 , w2978 , w2979 , w2980 , w2981 , w2982 , w2983 , w2984 , w2985 , w2986 , w2987 , w2988 , w2989 , w2990 , w2991 , w2992 , w2993 , w2994 , w2995 , w2996 , w2997 , w2998 , w2999 , w3000 , w3001 , w3002 , w3003 , w3004 , w3005 , w3006 , w3007 , w3008 , w3009 , w3010 , w3011 , w3012 , w3013 , w3014 , w3015 , w3016 , w3017 , w3018 , w3019 , w3020 , w3021 , w3022 , w3023 , w3024 , w3025 , w3026 , w3027 , w3028 , w3029 , w3030 , w3031 , w3032 , w3033 , w3034 , w3035 , w3036 , w3037 , w3038 , w3039 , w3040 , w3041 , w3042 , w3043 , w3044 , w3045 , w3046 , w3047 , w3048 , w3049 , w3050 , w3051 , w3052 , w3053 , w3054 , w3055 , w3056 , w3057 , w3058 , w3059 , w3060 , w3061 , w3062 , w3063 , w3064 , w3065 , w3066 , w3067 , w3068 , w3069 , w3070 , w3071 , w3072 , w3073 , w3074 , w3075 , w3076 , w3077 , w3078 , w3079 , w3080 , w3081 , w3082 , w3083 , w3084 , w3085 , w3086 , w3087 , w3088 , w3089 , w3090 , w3091 , w3092 , w3093 , w3094 , w3095 , w3096 , w3097 , w3098 , w3099 , w3100 , w3101 , w3102 , w3103 , w3104 , w3105 , w3106 , w3107 , w3108 , w3109 , w3110 , w3111 , w3112 , w3113 , w3114 , w3115 , w3116 , w3117 , w3118 , w3119 , w3120 , w3121 , w3122 , w3123 , w3124 , w3125 , w3126 , w3127 , w3128 , w3129 , w3130 , w3131 , w3132 , w3133 , w3134 , w3135 , w3136 , w3137 , w3138 , w3139 , w3140 , w3141 , w3142 , w3143 , w3144 , w3145 , w3146 , w3147 , w3148 , w3149 , w3150 , w3151 , w3152 , w3153 , w3154 , w3155 , w3156 , w3157 , w3158 , w3159 , w3160 , w3161 , w3162 , w3163 , w3164 , w3165 , w3166 , w3167 , w3168 , w3169 , w3170 , w3171 , w3172 , w3173 , w3174 , w3175 , w3176 , w3177 , w3178 , w3179 , w3180 , w3181 , w3182 , w3183 , w3184 , w3185 , w3186 , w3187 , w3188 , w3189 , w3190 , w3191 , w3192 , w3193 , w3194 , w3195 , w3196 , w3197 , w3198 , w3199 , w3200 , w3201 , w3202 , w3203 , w3204 , w3205 , w3206 , w3207 , w3208 , w3209 , w3210 , w3211 , w3212 , w3213 , w3214 , w3215 , w3216 , w3217 , w3218 , w3219 , w3220 , w3221 , w3222 , w3223 , w3224 , w3225 , w3226 , w3227 , w3228 , w3229 , w3230 , w3231 , w3232 , w3233 , w3234 , w3235 , w3236 , w3237 , w3238 , w3239 , w3240 , w3241 , w3242 , w3243 , w3244 , w3245 , w3246 , w3247 , w3248 , w3249 , w3250 , w3251 , w3252 , w3253 , w3254 , w3255 , w3256 , w3257 , w3258 , w3259 , w3260 , w3261 , w3262 , w3263 , w3264 , w3265 , w3266 , w3267 , w3268 , w3269 , w3270 , w3271 , w3272 , w3273 , w3274 , w3275 , w3276 , w3277 , w3278 , w3279 , w3280 , w3281 , w3282 , w3283 , w3284 , w3285 , w3286 , w3287 , w3288 , w3289 , w3290 , w3291 , w3292 , w3293 , w3294 , w3295 , w3296 , w3297 , w3298 , w3299 , w3300 , w3301 , w3302 , w3303 , w3304 , w3305 , w3306 , w3307 , w3308 , w3309 , w3310 , w3311 , w3312 , w3313 , w3314 , w3315 , w3316 , w3317 , w3318 , w3319 , w3320 , w3321 , w3322 , w3323 , w3324 , w3325 , w3326 , w3327 , w3328 , w3329 , w3330 , w3331 , w3332 , w3333 , w3334 , w3335 , w3336 , w3337 , w3338 , w3339 , w3340 , w3341 , w3342 , w3343 , w3344 , w3345 , w3346 , w3347 , w3348 , w3349 , w3350 , w3351 , w3352 , w3353 , w3354 , w3355 , w3356 , w3357 , w3358 , w3359 , w3360 , w3361 , w3362 , w3363 , w3364 , w3365 , w3366 , w3367 , w3368 , w3369 , w3370 , w3371 , w3372 , w3373 , w3374 , w3375 , w3376 , w3377 , w3378 , w3379 , w3380 , w3381 , w3382 , w3383 , w3384 , w3385 , w3386 , w3387 , w3388 , w3389 , w3390 , w3391 , w3392 , w3393 , w3394 , w3395 , w3396 , w3397 , w3398 , w3399 , w3400 , w3401 , w3402 , w3403 , w3404 , w3405 , w3406 , w3407 , w3408 , w3409 , w3410 , w3411 , w3412 , w3413 , w3414 , w3415 , w3416 , w3417 , w3418 , w3419 , w3420 , w3421 , w3422 , w3423 , w3424 , w3425 , w3426 , w3427 , w3428 , w3429 , w3430 , w3431 , w3432 , w3433 , w3434 , w3435 , w3436 , w3437 , w3438 , w3439 , w3440 , w3441 , w3442 , w3443 , w3444 , w3445 , w3446 , w3447 , w3448 , w3449 , w3450 , w3451 , w3452 , w3453 , w3454 , w3455 , w3456 , w3457 , w3458 , w3459 , w3460 , w3461 , w3462 , w3463 , w3464 , w3465 , w3466 , w3467 , w3468 , w3469 , w3470 , w3471 , w3472 , w3473 , w3474 , w3475 , w3476 , w3477 , w3478 , w3479 , w3480 , w3481 , w3482 , w3483 , w3484 , w3485 , w3486 , w3487 , w3488 , w3489 , w3490 , w3491 , w3492 , w3493 , w3494 , w3495 , w3496 , w3497 , w3498 , w3499 , w3500 , w3501 , w3502 , w3503 , w3504 , w3505 , w3506 , w3507 , w3508 , w3509 , w3510 , w3511 , w3512 , w3513 , w3514 , w3515 , w3516 , w3517 , w3518 , w3519 , w3520 , w3521 , w3522 , w3523 , w3524 , w3525 , w3526 , w3527 , w3528 , w3529 , w3530 , w3531 , w3532 , w3533 , w3534 , w3535 , w3536 , w3537 , w3538 , w3539 , w3540 , w3541 , w3542 , w3543 , w3544 , w3545 , w3546 , w3547 , w3548 , w3549 , w3550 , w3551 , w3552 , w3553 , w3554 , w3555 , w3556 , w3557 , w3558 , w3559 , w3560 , w3561 , w3562 , w3563 , w3564 , w3565 , w3566 , w3567 , w3568 , w3569 , w3570 , w3571 , w3572 , w3573 , w3574 , w3575 , w3576 , w3577 , w3578 , w3579 , w3580 , w3581 , w3582 , w3583 , w3584 , w3585 , w3586 , w3587 , w3588 , w3589 , w3590 , w3591 , w3592 , w3593 , w3594 , w3595 , w3596 , w3597 , w3598 , w3599 , w3600 , w3601 , w3602 , w3603 , w3604 , w3605 , w3606 , w3607 , w3608 , w3609 , w3610 , w3611 , w3612 , w3613 , w3614 , w3615 , w3616 , w3617 , w3618 , w3619 , w3620 , w3621 , w3622 , w3623 , w3624 , w3625 , w3626 , w3627 , w3628 , w3629 , w3630 , w3631 , w3632 , w3633 , w3634 , w3635 , w3636 , w3637 , w3638 , w3639 , w3640 , w3641 , w3642 , w3643 , w3644 , w3645 , w3646 , w3647 , w3648 , w3649 , w3650 , w3651 , w3652 , w3653 , w3654 , w3655 , w3656 , w3657 , w3658 , w3659 , w3660 , w3661 , w3662 , w3663 , w3664 , w3665 , w3666 , w3667 , w3668 , w3669 , w3670 , w3671 , w3672 , w3673 , w3674 , w3675 , w3676 , w3677 , w3678 , w3679 , w3680 , w3681 , w3682 , w3683 , w3684 , w3685 , w3686 , w3687 , w3688 , w3689 , w3690 , w3691 , w3692 , w3693 , w3694 , w3695 , w3696 , w3697 , w3698 , w3699 , w3700 , w3701 , w3702 , w3703 , w3704 , w3705 , w3706 , w3707 , w3708 , w3709 , w3710 , w3711 , w3712 , w3713 , w3714 , w3715 , w3716 , w3717 , w3718 , w3719 , w3720 , w3721 , w3722 , w3723 , w3724 , w3725 , w3726 , w3727 , w3728 , w3729 , w3730 , w3731 , w3732 , w3733 , w3734 , w3735 , w3736 , w3737 , w3738 , w3739 , w3740 , w3741 , w3742 , w3743 , w3744 , w3745 , w3746 , w3747 , w3748 , w3749 , w3750 , w3751 , w3752 , w3753 , w3754 , w3755 , w3756 , w3757 , w3758 , w3759 , w3760 , w3761 , w3762 , w3763 , w3764 , w3765 , w3766 , w3767 , w3768 , w3769 , w3770 , w3771 , w3772 , w3773 , w3774 , w3775 , w3776 , w3777 , w3778 , w3779 , w3780 , w3781 , w3782 , w3783 , w3784 , w3785 , w3786 , w3787 , w3788 , w3789 , w3790 , w3791 , w3792 , w3793 , w3794 , w3795 , w3796 , w3797 , w3798 , w3799 , w3800 , w3801 , w3802 , w3803 , w3804 , w3805 , w3806 , w3807 , w3808 , w3809 , w3810 , w3811 , w3812 , w3813 , w3814 , w3815 , w3816 , w3817 , w3818 , w3819 , w3820 , w3821 , w3822 , w3823 , w3824 , w3825 , w3826 , w3827 , w3828 , w3829 , w3830 , w3831 , w3832 , w3833 , w3834 , w3835 , w3836 , w3837 , w3838 , w3839 , w3840 , w3841 , w3842 , w3843 , w3844 , w3845 , w3846 , w3847 , w3848 , w3849 , w3850 , w3851 , w3852 , w3853 , w3854 , w3855 , w3856 , w3857 , w3858 , w3859 , w3860 , w3861 , w3862 , w3863 , w3864 , w3865 , w3866 , w3867 , w3868 , w3869 , w3870 , w3871 , w3872 , w3873 , w3874 , w3875 , w3876 , w3877 , w3878 , w3879 , w3880 , w3881 , w3882 , w3883 , w3884 , w3885 , w3886 , w3887 , w3888 , w3889 , w3890 , w3891 , w3892 , w3893 , w3894 , w3895 , w3896 , w3897 , w3898 , w3899 , w3900 , w3901 , w3902 , w3903 , w3904 , w3905 , w3906 , w3907 , w3908 , w3909 , w3910 , w3911 , w3912 , w3913 , w3914 , w3915 , w3916 , w3917 , w3918 , w3919 , w3920 , w3921 , w3922 , w3923 , w3924 , w3925 , w3926 , w3927 , w3928 , w3929 , w3930 , w3931 , w3932 , w3933 , w3934 , w3935 , w3936 , w3937 , w3938 , w3939 , w3940 , w3941 , w3942 , w3943 , w3944 , w3945 , w3946 , w3947 , w3948 , w3949 , w3950 , w3951 , w3952 , w3953 , w3954 , w3955 , w3956 , w3957 , w3958 , w3959 , w3960 , w3961 , w3962 , w3963 , w3964 , w3965 , w3966 , w3967 , w3968 , w3969 , w3970 , w3971 , w3972 , w3973 , w3974 , w3975 , w3976 , w3977 , w3978 , w3979 , w3980 , w3981 , w3982 , w3983 , w3984 , w3985 , w3986 , w3987 , w3988 , w3989 , w3990 , w3991 , w3992 , w3993 , w3994 , w3995 , w3996 , w3997 , w3998 , w3999 , w4000 , w4001 , w4002 , w4003 , w4004 , w4005 , w4006 , w4007 , w4008 , w4009 , w4010 , w4011 , w4012 , w4013 , w4014 , w4015 , w4016 , w4017 , w4018 , w4019 , w4020 , w4021 , w4022 , w4023 , w4024 , w4025 , w4026 , w4027 , w4028 , w4029 , w4030 , w4031 , w4032 , w4033 , w4034 , w4035 , w4036 , w4037 , w4038 , w4039 , w4040 , w4041 , w4042 , w4043 , w4044 , w4045 , w4046 , w4047 , w4048 , w4049 , w4050 , w4051 , w4052 , w4053 , w4054 , w4055 , w4056 , w4057 , w4058 , w4059 , w4060 , w4061 , w4062 , w4063 , w4064 , w4065 , w4066 , w4067 , w4068 , w4069 , w4070 , w4071 , w4072 , w4073 , w4074 , w4075 , w4076 , w4077 , w4078 , w4079 , w4080 , w4081 , w4082 , w4083 , w4084 , w4085 , w4086 , w4087 , w4088 , w4089 , w4090 , w4091 , w4092 , w4093 , w4094 , w4095 , w4096 , w4097 , w4098 , w4099 , w4100 , w4101 , w4102 , w4103 , w4104 , w4105 , w4106 , w4107 , w4108 , w4109 , w4110 , w4111 , w4112 , w4113 , w4114 , w4115 , w4116 , w4117 , w4118 , w4119 , w4120 , w4121 , w4122 , w4123 , w4124 , w4125 , w4126 , w4127 , w4128 , w4129 , w4130 , w4131 , w4132 , w4133 , w4134 , w4135 , w4136 , w4137 , w4138 , w4139 , w4140 , w4141 , w4142 , w4143 , w4144 , w4145 , w4146 , w4147 , w4148 , w4149 , w4150 , w4151 , w4152 , w4153 , w4154 , w4155 , w4156 , w4157 , w4158 , w4159 , w4160 , w4161 , w4162 , w4163 , w4164 , w4165 , w4166 , w4167 , w4168 , w4169 , w4170 , w4171 , w4172 , w4173 , w4174 , w4175 , w4176 , w4177 , w4178 , w4179 , w4180 , w4181 , w4182 , w4183 , w4184 , w4185 , w4186 , w4187 , w4188 , w4189 , w4190 , w4191 , w4192 , w4193 , w4194 , w4195 , w4196 , w4197 , w4198 , w4199 , w4200 , w4201 , w4202 , w4203 , w4204 , w4205 , w4206 , w4207 , w4208 , w4209 , w4210 , w4211 , w4212 , w4213 , w4214 , w4215 , w4216 , w4217 , w4218 , w4219 , w4220 , w4221 , w4222 , w4223 , w4224 , w4225 , w4226 , w4227 , w4228 , w4229 , w4230 , w4231 , w4232 , w4233 , w4234 , w4235 , w4236 , w4237 , w4238 , w4239 , w4240 , w4241 , w4242 , w4243 , w4244 , w4245 , w4246 , w4247 , w4248 , w4249 , w4250 , w4251 , w4252 , w4253 , w4254 , w4255 , w4256 , w4257 , w4258 , w4259 , w4260 , w4261 , w4262 , w4263 , w4264 , w4265 , w4266 , w4267 , w4268 , w4269 , w4270 , w4271 , w4272 , w4273 , w4274 , w4275 , w4276 , w4277 , w4278 , w4279 , w4280 , w4281 , w4282 , w4283 , w4284 , w4285 , w4286 , w4287 , w4288 , w4289 , w4290 , w4291 , w4292 , w4293 , w4294 , w4295 , w4296 , w4297 , w4298 , w4299 , w4300 , w4301 , w4302 , w4303 , w4304 , w4305 , w4306 , w4307 , w4308 , w4309 , w4310 , w4311 , w4312 , w4313 , w4314 , w4315 , w4316 , w4317 , w4318 , w4319 , w4320 , w4321 , w4322 , w4323 , w4324 , w4325 , w4326 , w4327 , w4328 , w4329 , w4330 , w4331 , w4332 , w4333 , w4334 , w4335 , w4336 , w4337 , w4338 , w4339 , w4340 , w4341 , w4342 , w4343 , w4344 , w4345 , w4346 , w4347 , w4348 , w4349 , w4350 , w4351 , w4352 , w4353 , w4354 , w4355 , w4356 , w4357 , w4358 , w4359 , w4360 , w4361 , w4362 , w4363 , w4364 , w4365 , w4366 , w4367 , w4368 , w4369 , w4370 , w4371 , w4372 , w4373 , w4374 , w4375 , w4376 , w4377 , w4378 , w4379 , w4380 , w4381 , w4382 , w4383 , w4384 , w4385 , w4386 , w4387 , w4388 , w4389 , w4390 , w4391 , w4392 , w4393 , w4394 , w4395 , w4396 , w4397 , w4398 , w4399 , w4400 , w4401 , w4402 , w4403 , w4404 , w4405 , w4406 , w4407 , w4408 , w4409 , w4410 , w4411 , w4412 , w4413 , w4414 , w4415 , w4416 , w4417 , w4418 , w4419 , w4420 , w4421 , w4422 , w4423 , w4424 , w4425 , w4426 , w4427 , w4428 , w4429 , w4430 , w4431 , w4432 , w4433 , w4434 , w4435 , w4436 , w4437 , w4438 , w4439 , w4440 , w4441 , w4442 , w4443 , w4444 , w4445 , w4446 , w4447 , w4448 , w4449 , w4450 , w4451 , w4452 , w4453 , w4454 , w4455 , w4456 , w4457 , w4458 , w4459 , w4460 , w4461 , w4462 , w4463 , w4464 , w4465 , w4466 , w4467 , w4468 , w4469 , w4470 , w4471 , w4472 , w4473 , w4474 , w4475 , w4476 , w4477 , w4478 , w4479 , w4480 , w4481 , w4482 , w4483 , w4484 , w4485 , w4486 , w4487 , w4488 , w4489 , w4490 , w4491 , w4492 , w4493 , w4494 , w4495 , w4496 , w4497 , w4498 , w4499 , w4500 , w4501 , w4502 , w4503 , w4504 , w4505 , w4506 , w4507 , w4508 , w4509 , w4510 , w4511 , w4512 , w4513 , w4514 , w4515 , w4516 , w4517 , w4518 , w4519 , w4520 , w4521 , w4522 , w4523 , w4524 , w4525 , w4526 , w4527 , w4528 , w4529 , w4530 , w4531 , w4532 , w4533 , w4534 , w4535 , w4536 , w4537 , w4538 , w4539 , w4540 , w4541 , w4542 , w4543 , w4544 , w4545 , w4546 , w4547 , w4548 , w4549 , w4550 , w4551 , w4552 , w4553 , w4554 , w4555 , w4556 , w4557 , w4558 , w4559 , w4560 , w4561 , w4562 , w4563 , w4564 , w4565 , w4566 , w4567 , w4568 , w4569 , w4570 , w4571 , w4572 , w4573 , w4574 , w4575 , w4576 , w4577 , w4578 , w4579 , w4580 , w4581 , w4582 , w4583 , w4584 , w4585 , w4586 , w4587 , w4588 , w4589 , w4590 , w4591 , w4592 , w4593 , w4594 , w4595 , w4596 , w4597 , w4598 , w4599 , w4600 , w4601 , w4602 , w4603 , w4604 , w4605 , w4606 , w4607 , w4608 , w4609 , w4610 , w4611 , w4612 , w4613 , w4614 , w4615 , w4616 , w4617 , w4618 , w4619 , w4620 , w4621 , w4622 , w4623 , w4624 , w4625 , w4626 , w4627 , w4628 , w4629 , w4630 , w4631 , w4632 , w4633 , w4634 , w4635 , w4636 , w4637 , w4638 , w4639 , w4640 , w4641 , w4642 , w4643 , w4644 , w4645 , w4646 , w4647 , w4648 , w4649 , w4650 , w4651 , w4652 , w4653 , w4654 , w4655 , w4656 , w4657 , w4658 , w4659 , w4660 , w4661 , w4662 , w4663 , w4664 , w4665 , w4666 , w4667 , w4668 , w4669 , w4670 , w4671 , w4672 , w4673 , w4674 , w4675 , w4676 , w4677 , w4678 , w4679 , w4680 , w4681 , w4682 , w4683 , w4684 , w4685 , w4686 , w4687 , w4688 , w4689 , w4690 , w4691 , w4692 , w4693 , w4694 , w4695 , w4696 , w4697 , w4698 , w4699 , w4700 , w4701 , w4702 , w4703 , w4704 , w4705 , w4706 , w4707 , w4708 , w4709 , w4710 , w4711 , w4712 , w4713 , w4714 , w4715 , w4716 , w4717 , w4718 , w4719 , w4720 , w4721 , w4722 , w4723 , w4724 , w4725 , w4726 , w4727 , w4728 , w4729 , w4730 , w4731 , w4732 , w4733 , w4734 , w4735 , w4736 , w4737 , w4738 , w4739 , w4740 , w4741 , w4742 , w4743 , w4744 , w4745 , w4746 , w4747 , w4748 , w4749 , w4750 , w4751 , w4752 , w4753 , w4754 , w4755 , w4756 , w4757 , w4758 , w4759 , w4760 , w4761 , w4762 , w4763 , w4764 , w4765 , w4766 , w4767 , w4768 , w4769 , w4770 , w4771 , w4772 , w4773 , w4774 , w4775 , w4776 , w4777 , w4778 , w4779 , w4780 , w4781 , w4782 , w4783 , w4784 , w4785 , w4786 , w4787 , w4788 , w4789 , w4790 , w4791 , w4792 , w4793 , w4794 , w4795 , w4796 , w4797 , w4798 , w4799 , w4800 , w4801 , w4802 , w4803 , w4804 , w4805 , w4806 , w4807 , w4808 , w4809 , w4810 , w4811 , w4812 , w4813 , w4814 , w4815 , w4816 , w4817 , w4818 , w4819 , w4820 , w4821 , w4822 , w4823 , w4824 , w4825 , w4826 , w4827 , w4828 , w4829 , w4830 , w4831 , w4832 , w4833 , w4834 , w4835 , w4836 , w4837 , w4838 , w4839 , w4840 , w4841 , w4842 , w4843 , w4844 , w4845 , w4846 , w4847 , w4848 , w4849 , w4850 , w4851 , w4852 , w4853 , w4854 , w4855 , w4856 , w4857 , w4858 , w4859 , w4860 , w4861 , w4862 , w4863 , w4864 , w4865 , w4866 , w4867 , w4868 , w4869 , w4870 , w4871 , w4872 , w4873 , w4874 , w4875 , w4876 , w4877 , w4878 , w4879 , w4880 , w4881 , w4882 , w4883 , w4884 , w4885 , w4886 , w4887 , w4888 , w4889 , w4890 , w4891 , w4892 , w4893 , w4894 , w4895 , w4896 , w4897 , w4898 , w4899 , w4900 , w4901 , w4902 , w4903 , w4904 , w4905 , w4906 , w4907 , w4908 , w4909 , w4910 , w4911 , w4912 , w4913 , w4914 , w4915 , w4916 , w4917 , w4918 , w4919 , w4920 , w4921 , w4922 , w4923 , w4924 , w4925 , w4926 , w4927 , w4928 , w4929 , w4930 , w4931 , w4932 , w4933 , w4934 , w4935 , w4936 , w4937 , w4938 , w4939 , w4940 , w4941 , w4942 , w4943 , w4944 , w4945 , w4946 , w4947 , w4948 , w4949 , w4950 , w4951 , w4952 , w4953 , w4954 , w4955 , w4956 , w4957 , w4958 , w4959 , w4960 , w4961 , w4962 , w4963 , w4964 , w4965 , w4966 , w4967 , w4968 , w4969 , w4970 , w4971 , w4972 , w4973 , w4974 , w4975 , w4976 , w4977 , w4978 , w4979 , w4980 , w4981 , w4982 , w4983 , w4984 , w4985 , w4986 , w4987 , w4988 , w4989 , w4990 , w4991 , w4992 , w4993 , w4994 , w4995 , w4996 , w4997 , w4998 , w4999 , w5000 , w5001 , w5002 , w5003 , w5004 , w5005 , w5006 , w5007 , w5008 , w5009 , w5010 , w5011 , w5012 , w5013 , w5014 , w5015 , w5016 , w5017 , w5018 , w5019 , w5020 , w5021 , w5022 , w5023 , w5024 , w5025 , w5026 , w5027 , w5028 , w5029 , w5030 , w5031 , w5032 , w5033 , w5034 , w5035 , w5036 , w5037 , w5038 , w5039 , w5040 , w5041 , w5042 , w5043 , w5044 , w5045 , w5046 , w5047 , w5048 , w5049 , w5050 , w5051 , w5052 , w5053 , w5054 , w5055 , w5056 , w5057 , w5058 , w5059 , w5060 , w5061 , w5062 , w5063 , w5064 , w5065 , w5066 , w5067 , w5068 , w5069 , w5070 , w5071 , w5072 , w5073 , w5074 , w5075 , w5076 , w5077 , w5078 , w5079 , w5080 , w5081 , w5082 , w5083 , w5084 , w5085 , w5086 , w5087 , w5088 , w5089 , w5090 , w5091 , w5092 , w5093 , w5094 , w5095 , w5096 , w5097 , w5098 , w5099 , w5100 , w5101 , w5102 , w5103 , w5104 , w5105 , w5106 , w5107 , w5108 , w5109 , w5110 , w5111 , w5112 , w5113 , w5114 , w5115 , w5116 , w5117 , w5118 , w5119 , w5120 , w5121 , w5122 , w5123 , w5124 , w5125 , w5126 , w5127 , w5128 , w5129 , w5130 , w5131 , w5132 , w5133 , w5134 , w5135 , w5136 , w5137 , w5138 , w5139 , w5140 , w5141 , w5142 , w5143 , w5144 , w5145 , w5146 , w5147 , w5148 , w5149 , w5150 , w5151 , w5152 , w5153 , w5154 , w5155 , w5156 , w5157 , w5158 , w5159 , w5160 , w5161 , w5162 , w5163 , w5164 , w5165 , w5166 , w5167 , w5168 , w5169 , w5170 , w5171 , w5172 , w5173 , w5174 , w5175 , w5176 , w5177 , w5178 , w5179 , w5180 , w5181 , w5182 , w5183 , w5184 , w5185 , w5186 , w5187 , w5188 , w5189 , w5190 , w5191 , w5192 , w5193 , w5194 , w5195 , w5196 , w5197 , w5198 , w5199 , w5200 , w5201 , w5202 , w5203 , w5204 , w5205 , w5206 , w5207 , w5208 , w5209 , w5210 , w5211 , w5212 , w5213 , w5214 , w5215 , w5216 , w5217 , w5218 , w5219 , w5220 , w5221 , w5222 , w5223 , w5224 , w5225 , w5226 , w5227 , w5228 , w5229 , w5230 , w5231 , w5232 , w5233 , w5234 , w5235 , w5236 , w5237 , w5238 , w5239 , w5240 , w5241 , w5242 , w5243 , w5244 , w5245 , w5246 , w5247 , w5248 , w5249 , w5250 , w5251 , w5252 , w5253 , w5254 , w5255 , w5256 , w5257 , w5258 , w5259 , w5260 , w5261 , w5262 , w5263 , w5264 , w5265 , w5266 , w5267 , w5268 , w5269 , w5270 , w5271 , w5272 , w5273 , w5274 , w5275 , w5276 , w5277 , w5278 , w5279 , w5280 , w5281 , w5282 , w5283 , w5284 , w5285 , w5286 , w5287 , w5288 , w5289 , w5290 , w5291 , w5292 , w5293 , w5294 , w5295 , w5296 , w5297 , w5298 , w5299 , w5300 , w5301 , w5302 , w5303 , w5304 , w5305 , w5306 , w5307 , w5308 , w5309 , w5310 , w5311 , w5312 , w5313 , w5314 , w5315 , w5316 , w5317 , w5318 , w5319 , w5320 , w5321 , w5322 , w5323 , w5324 , w5325 , w5326 , w5327 , w5328 , w5329 , w5330 , w5331 , w5332 , w5333 , w5334 , w5335 , w5336 , w5337 , w5338 , w5339 , w5340 , w5341 , w5342 , w5343 , w5344 , w5345 , w5346 , w5347 , w5348 , w5349 , w5350 , w5351 , w5352 , w5353 , w5354 , w5355 , w5356 , w5357 , w5358 , w5359 , w5360 , w5361 , w5362 , w5363 , w5364 , w5365 , w5366 , w5367 , w5368 , w5369 , w5370 , w5371 , w5372 , w5373 , w5374 , w5375 , w5376 , w5377 , w5378 , w5379 , w5380 , w5381 , w5382 , w5383 , w5384 , w5385 , w5386 , w5387 , w5388 , w5389 , w5390 , w5391 , w5392 , w5393 , w5394 , w5395 , w5396 , w5397 , w5398 , w5399 , w5400 , w5401 , w5402 , w5403 , w5404 , w5405 , w5406 , w5407 , w5408 , w5409 , w5410 , w5411 , w5412 , w5413 , w5414 , w5415 , w5416 , w5417 , w5418 , w5419 , w5420 , w5421 , w5422 , w5423 , w5424 , w5425 , w5426 , w5427 , w5428 , w5429 , w5430 , w5431 , w5432 , w5433 , w5434 , w5435 , w5436 , w5437 , w5438 , w5439 , w5440 , w5441 , w5442 , w5443 , w5444 , w5445 , w5446 , w5447 , w5448 , w5449 , w5450 , w5451 , w5452 , w5453 , w5454 , w5455 , w5456 , w5457 , w5458 , w5459 , w5460 , w5461 , w5462 , w5463 , w5464 , w5465 , w5466 , w5467 , w5468 , w5469 , w5470 , w5471 , w5472 , w5473 , w5474 , w5475 , w5476 , w5477 , w5478 , w5479 , w5480 , w5481 , w5482 , w5483 , w5484 , w5485 , w5486 , w5487 , w5488 , w5489 , w5490 , w5491 , w5492 , w5493 , w5494 , w5495 , w5496 , w5497 , w5498 , w5499 , w5500 , w5501 , w5502 , w5503 , w5504 , w5505 , w5506 , w5507 , w5508 , w5509 , w5510 , w5511 , w5512 , w5513 , w5514 , w5515 , w5516 , w5517 , w5518 , w5519 , w5520 , w5521 , w5522 , w5523 , w5524 , w5525 , w5526 , w5527 , w5528 , w5529 , w5530 , w5531 , w5532 , w5533 , w5534 , w5535 , w5536 , w5537 , w5538 , w5539 , w5540 , w5541 , w5542 , w5543 , w5544 , w5545 , w5546 , w5547 , w5548 , w5549 , w5550 , w5551 , w5552 , w5553 , w5554 , w5555 , w5556 , w5557 , w5558 , w5559 , w5560 , w5561 , w5562 , w5563 , w5564 , w5565 , w5566 , w5567 , w5568 , w5569 , w5570 , w5571 , w5572 , w5573 , w5574 , w5575 , w5576 , w5577 , w5578 , w5579 , w5580 , w5581 , w5582 , w5583 , w5584 , w5585 , w5586 , w5587 , w5588 , w5589 , w5590 , w5591 , w5592 , w5593 , w5594 , w5595 , w5596 , w5597 , w5598 , w5599 , w5600 , w5601 , w5602 , w5603 , w5604 , w5605 , w5606 , w5607 , w5608 , w5609 , w5610 , w5611 , w5612 , w5613 , w5614 , w5615 , w5616 , w5617 , w5618 , w5619 , w5620 , w5621 , w5622 , w5623 , w5624 , w5625 , w5626 , w5627 , w5628 , w5629 , w5630 , w5631 , w5632 , w5633 , w5634 , w5635 , w5636 , w5637 , w5638 , w5639 , w5640 , w5641 , w5642 , w5643 , w5644 , w5645 , w5646 , w5647 , w5648 , w5649 , w5650 , w5651 , w5652 , w5653 , w5654 , w5655 , w5656 , w5657 , w5658 , w5659 , w5660 , w5661 , w5662 , w5663 , w5664 , w5665 , w5666 , w5667 , w5668 , w5669 , w5670 , w5671 , w5672 , w5673 , w5674 , w5675 , w5676 , w5677 , w5678 , w5679 , w5680 , w5681 , w5682 , w5683 , w5684 , w5685 , w5686 , w5687 , w5688 , w5689 , w5690 , w5691 , w5692 , w5693 , w5694 , w5695 , w5696 , w5697 , w5698 , w5699 , w5700 , w5701 , w5702 , w5703 , w5704 , w5705 , w5706 , w5707 , w5708 , w5709 , w5710 , w5711 , w5712 , w5713 , w5714 , w5715 , w5716 , w5717 , w5718 , w5719 , w5720 , w5721 , w5722 , w5723 , w5724 , w5725 , w5726 , w5727 , w5728 , w5729 , w5730 , w5731 , w5732 , w5733 , w5734 , w5735 , w5736 , w5737 , w5738 , w5739 , w5740 , w5741 , w5742 , w5743 , w5744 , w5745 , w5746 , w5747 , w5748 , w5749 , w5750 , w5751 , w5752 , w5753 , w5754 , w5755 , w5756 , w5757 , w5758 , w5759 , w5760 , w5761 , w5762 , w5763 , w5764 , w5765 , w5766 , w5767 , w5768 , w5769 , w5770 , w5771 , w5772 , w5773 , w5774 , w5775 , w5776 , w5777 , w5778 , w5779 , w5780 , w5781 , w5782 , w5783 , w5784 , w5785 , w5786 , w5787 , w5788 , w5789 , w5790 , w5791 , w5792 , w5793 , w5794 , w5795 , w5796 , w5797 , w5798 , w5799 , w5800 , w5801 , w5802 , w5803 , w5804 , w5805 , w5806 , w5807 , w5808 , w5809 , w5810 , w5811 , w5812 , w5813 , w5814 , w5815 , w5816 , w5817 , w5818 , w5819 , w5820 , w5821 , w5822 , w5823 , w5824 , w5825 , w5826 , w5827 , w5828 , w5829 , w5830 , w5831 , w5832 , w5833 , w5834 , w5835 , w5836 , w5837 , w5838 , w5839 , w5840 , w5841 , w5842 , w5843 , w5844 , w5845 , w5846 , w5847 , w5848 , w5849 , w5850 , w5851 , w5852 , w5853 , w5854 , w5855 , w5856 , w5857 , w5858 , w5859 , w5860 , w5861 , w5862 , w5863 , w5864 , w5865 , w5866 , w5867 , w5868 , w5869 , w5870 , w5871 , w5872 , w5873 , w5874 , w5875 , w5876 , w5877 , w5878 , w5879 , w5880 , w5881 , w5882 , w5883 , w5884 , w5885 , w5886 , w5887 , w5888 , w5889 , w5890 , w5891 , w5892 , w5893 , w5894 , w5895 , w5896 , w5897 , w5898 , w5899 , w5900 , w5901 , w5902 , w5903 , w5904 , w5905 , w5906 , w5907 , w5908 , w5909 , w5910 , w5911 , w5912 , w5913 , w5914 , w5915 , w5916 , w5917 , w5918 , w5919 , w5920 , w5921 , w5922 , w5923 , w5924 , w5925 , w5926 , w5927 , w5928 , w5929 , w5930 , w5931 , w5932 , w5933 , w5934 , w5935 , w5936 , w5937 , w5938 , w5939 , w5940 , w5941 , w5942 , w5943 , w5944 , w5945 , w5946 , w5947 , w5948 , w5949 , w5950 , w5951 , w5952 , w5953 , w5954 , w5955 , w5956 , w5957 , w5958 , w5959 , w5960 , w5961 , w5962 , w5963 , w5964 , w5965 , w5966 , w5967 , w5968 , w5969 , w5970 , w5971 , w5972 , w5973 , w5974 , w5975 , w5976 , w5977 , w5978 , w5979 , w5980 , w5981 , w5982 , w5983 , w5984 , w5985 , w5986 , w5987 , w5988 , w5989 , w5990 , w5991 , w5992 , w5993 , w5994 , w5995 , w5996 , w5997 , w5998 , w5999 , w6000 , w6001 , w6002 , w6003 , w6004 , w6005 , w6006 , w6007 , w6008 , w6009 , w6010 , w6011 , w6012 , w6013 , w6014 , w6015 , w6016 , w6017 , w6018 , w6019 , w6020 , w6021 , w6022 , w6023 , w6024 , w6025 , w6026 , w6027 , w6028 , w6029 , w6030 , w6031 , w6032 , w6033 , w6034 , w6035 , w6036 , w6037 , w6038 , w6039 , w6040 , w6041 , w6042 , w6043 , w6044 , w6045 , w6046 , w6047 , w6048 , w6049 , w6050 , w6051 , w6052 , w6053 , w6054 , w6055 , w6056 , w6057 , w6058 , w6059 , w6060 , w6061 , w6062 , w6063 , w6064 , w6065 , w6066 , w6067 , w6068 , w6069 , w6070 , w6071 , w6072 , w6073 , w6074 , w6075 , w6076 , w6077 , w6078 , w6079 , w6080 , w6081 , w6082 , w6083 , w6084 , w6085 , w6086 , w6087 , w6088 , w6089 , w6090 , w6091 , w6092 , w6093 , w6094 , w6095 , w6096 , w6097 , w6098 , w6099 , w6100 , w6101 , w6102 , w6103 , w6104 , w6105 , w6106 , w6107 , w6108 , w6109 , w6110 , w6111 , w6112 , w6113 , w6114 , w6115 , w6116 , w6117 , w6118 , w6119 , w6120 , w6121 , w6122 , w6123 , w6124 , w6125 , w6126 , w6127 , w6128 , w6129 , w6130 , w6131 , w6132 , w6133 , w6134 , w6135 , w6136 , w6137 , w6138 , w6139 , w6140 , w6141 , w6142 , w6143 , w6144 , w6145 , w6146 , w6147 , w6148 , w6149 , w6150 , w6151 , w6152 , w6153 , w6154 , w6155 , w6156 , w6157 , w6158 , w6159 , w6160 , w6161 , w6162 , w6163 , w6164 , w6165 , w6166 , w6167 , w6168 , w6169 , w6170 , w6171 , w6172 , w6173 , w6174 , w6175 , w6176 , w6177 , w6178 , w6179 , w6180 , w6181 , w6182 , w6183 , w6184 , w6185 , w6186 , w6187 , w6188 , w6189 , w6190 , w6191 , w6192 , w6193 , w6194 , w6195 , w6196 , w6197 , w6198 , w6199 , w6200 , w6201 , w6202 , w6203 , w6204 , w6205 , w6206 , w6207 , w6208 , w6209 , w6210 , w6211 , w6212 , w6213 , w6214 , w6215 , w6216 , w6217 , w6218 , w6219 , w6220 , w6221 , w6222 , w6223 , w6224 , w6225 , w6226 , w6227 , w6228 , w6229 , w6230 , w6231 , w6232 , w6233 , w6234 , w6235 , w6236 , w6237 , w6238 , w6239 , w6240 , w6241 , w6242 , w6243 , w6244 , w6245 , w6246 , w6247 , w6248 , w6249 , w6250 , w6251 , w6252 , w6253 , w6254 , w6255 , w6256 , w6257 , w6258 , w6259 , w6260 , w6261 , w6262 , w6263 , w6264 , w6265 , w6266 , w6267 , w6268 , w6269 , w6270 , w6271 , w6272 , w6273 , w6274 , w6275 , w6276 , w6277 , w6278 , w6279 , w6280 , w6281 , w6282 , w6283 , w6284 , w6285 , w6286 , w6287 , w6288 , w6289 , w6290 , w6291 , w6292 , w6293 , w6294 , w6295 , w6296 , w6297 , w6298 , w6299 , w6300 , w6301 , w6302 , w6303 , w6304 , w6305 , w6306 , w6307 , w6308 , w6309 , w6310 , w6311 , w6312 , w6313 , w6314 , w6315 , w6316 , w6317 , w6318 , w6319 , w6320 , w6321 , w6322 , w6323 , w6324 , w6325 , w6326 , w6327 , w6328 , w6329 , w6330 , w6331 , w6332 , w6333 , w6334 , w6335 , w6336 , w6337 , w6338 , w6339 , w6340 , w6341 , w6342 , w6343 , w6344 , w6345 , w6346 , w6347 , w6348 , w6349 , w6350 , w6351 , w6352 , w6353 , w6354 , w6355 , w6356 , w6357 , w6358 , w6359 , w6360 , w6361 , w6362 , w6363 , w6364 , w6365 , w6366 , w6367 , w6368 , w6369 , w6370 , w6371 , w6372 , w6373 , w6374 , w6375 , w6376 , w6377 , w6378 , w6379 , w6380 , w6381 , w6382 , w6383 , w6384 , w6385 , w6386 , w6387 , w6388 , w6389 , w6390 , w6391 , w6392 , w6393 , w6394 , w6395 , w6396 , w6397 , w6398 , w6399 , w6400 , w6401 , w6402 , w6403 , w6404 , w6405 , w6406 , w6407 , w6408 , w6409 , w6410 , w6411 , w6412 , w6413 , w6414 , w6415 , w6416 , w6417 , w6418 , w6419 , w6420 , w6421 , w6422 , w6423 , w6424 , w6425 , w6426 , w6427 , w6428 , w6429 , w6430 , w6431 , w6432 , w6433 , w6434 , w6435 , w6436 , w6437 , w6438 , w6439 , w6440 , w6441 , w6442 , w6443 , w6444 , w6445 , w6446 , w6447 , w6448 , w6449 , w6450 , w6451 , w6452 , w6453 , w6454 , w6455 , w6456 , w6457 , w6458 , w6459 , w6460 , w6461 , w6462 , w6463 , w6464 , w6465 , w6466 , w6467 , w6468 , w6469 , w6470 , w6471 , w6472 , w6473 , w6474 , w6475 , w6476 , w6477 , w6478 , w6479 , w6480 , w6481 , w6482 , w6483 , w6484 , w6485 , w6486 , w6487 , w6488 , w6489 , w6490 , w6491 , w6492 , w6493 , w6494 , w6495 , w6496 , w6497 , w6498 , w6499 , w6500 , w6501 , w6502 , w6503 , w6504 , w6505 , w6506 , w6507 , w6508 , w6509 , w6510 , w6511 , w6512 , w6513 , w6514 , w6515 , w6516 , w6517 , w6518 , w6519 , w6520 , w6521 , w6522 , w6523 , w6524 , w6525 , w6526 , w6527 , w6528 , w6529 , w6530 , w6531 , w6532 , w6533 , w6534 , w6535 , w6536 , w6537 , w6538 , w6539 , w6540 , w6541 , w6542 , w6543 , w6544 , w6545 , w6546 , w6547 , w6548 , w6549 , w6550 , w6551 , w6552 , w6553 , w6554 , w6555 , w6556 , w6557 , w6558 , w6559 , w6560 , w6561 , w6562 , w6563 , w6564 , w6565 , w6566 , w6567 , w6568 , w6569 , w6570 , w6571 , w6572 , w6573 , w6574 , w6575 , w6576 , w6577 , w6578 , w6579 , w6580 , w6581 , w6582 , w6583 , w6584 , w6585 , w6586 , w6587 , w6588 , w6589 , w6590 , w6591 , w6592 , w6593 , w6594 , w6595 , w6596 , w6597 , w6598 , w6599 , w6600 , w6601 , w6602 , w6603 , w6604 , w6605 , w6606 , w6607 , w6608 , w6609 , w6610 , w6611 , w6612 , w6613 , w6614 , w6615 , w6616 , w6617 , w6618 , w6619 , w6620 , w6621 , w6622 , w6623 , w6624 , w6625 , w6626 , w6627 , w6628 , w6629 , w6630 , w6631 , w6632 , w6633 , w6634 , w6635 , w6636 , w6637 , w6638 , w6639 , w6640 , w6641 , w6642 , w6643 , w6644 , w6645 , w6646 , w6647 , w6648 , w6649 , w6650 , w6651 , w6652 , w6653 , w6654 , w6655 , w6656 , w6657 , w6658 , w6659 , w6660 , w6661 , w6662 , w6663 , w6664 , w6665 , w6666 , w6667 , w6668 , w6669 , w6670 , w6671 , w6672 , w6673 , w6674 , w6675 , w6676 , w6677 , w6678 , w6679 , w6680 , w6681 , w6682 , w6683 , w6684 , w6685 , w6686 , w6687 , w6688 , w6689 , w6690 , w6691 , w6692 , w6693 , w6694 , w6695 , w6696 , w6697 , w6698 , w6699 , w6700 , w6701 , w6702 , w6703 , w6704 , w6705 , w6706 , w6707 , w6708 , w6709 , w6710 , w6711 , w6712 , w6713 , w6714 , w6715 , w6716 , w6717 , w6718 , w6719 , w6720 , w6721 , w6722 , w6723 , w6724 , w6725 , w6726 , w6727 , w6728 , w6729 , w6730 , w6731 , w6732 , w6733 , w6734 , w6735 , w6736 , w6737 , w6738 , w6739 , w6740 , w6741 , w6742 , w6743 , w6744 , w6745 , w6746 , w6747 , w6748 , w6749 , w6750 , w6751 , w6752 , w6753 , w6754 , w6755 , w6756 , w6757 , w6758 , w6759 , w6760 , w6761 , w6762 , w6763 , w6764 , w6765 , w6766 , w6767 , w6768 , w6769 , w6770 , w6771 , w6772 , w6773 , w6774 , w6775 , w6776 , w6777 , w6778 , w6779 , w6780 , w6781 , w6782 , w6783 , w6784 , w6785 , w6786 , w6787 , w6788 , w6789 , w6790 , w6791 , w6792 , w6793 , w6794 , w6795 , w6796 , w6797 , w6798 , w6799 , w6800 , w6801 , w6802 , w6803 , w6804 , w6805 , w6806 , w6807 , w6808 , w6809 , w6810 , w6811 , w6812 , w6813 , w6814 , w6815 , w6816 , w6817 , w6818 , w6819 , w6820 , w6821 , w6822 , w6823 , w6824 , w6825 , w6826 , w6827 , w6828 , w6829 , w6830 , w6831 , w6832 , w6833 , w6834 , w6835 , w6836 , w6837 , w6838 , w6839 , w6840 , w6841 , w6842 , w6843 , w6844 , w6845 , w6846 , w6847 , w6848 , w6849 , w6850 , w6851 , w6852 , w6853 , w6854 , w6855 , w6856 , w6857 , w6858 , w6859 , w6860 , w6861 , w6862 , w6863 , w6864 , w6865 , w6866 , w6867 , w6868 , w6869 , w6870 , w6871 , w6872 , w6873 , w6874 , w6875 , w6876 , w6877 , w6878 , w6879 , w6880 , w6881 , w6882 , w6883 , w6884 , w6885 , w6886 , w6887 , w6888 , w6889 , w6890 , w6891 , w6892 , w6893 , w6894 , w6895 , w6896 , w6897 , w6898 , w6899 , w6900 , w6901 , w6902 , w6903 , w6904 , w6905 , w6906 , w6907 , w6908 , w6909 , w6910 , w6911 , w6912 , w6913 , w6914 , w6915 , w6916 , w6917 , w6918 , w6919 , w6920 , w6921 , w6922 , w6923 , w6924 , w6925 , w6926 , w6927 , w6928 , w6929 , w6930 , w6931 , w6932 , w6933 , w6934 , w6935 , w6936 , w6937 , w6938 , w6939 , w6940 , w6941 , w6942 , w6943 , w6944 , w6945 , w6946 , w6947 , w6948 , w6949 , w6950 , w6951 , w6952 , w6953 , w6954 , w6955 , w6956 , w6957 , w6958 , w6959 , w6960 , w6961 , w6962 , w6963 , w6964 , w6965 , w6966 , w6967 , w6968 , w6969 , w6970 , w6971 , w6972 , w6973 , w6974 , w6975 , w6976 , w6977 , w6978 , w6979 , w6980 , w6981 , w6982 , w6983 , w6984 , w6985 , w6986 , w6987 , w6988 , w6989 , w6990 , w6991 , w6992 , w6993 , w6994 , w6995 , w6996 , w6997 , w6998 , w6999 , w7000 , w7001 , w7002 , w7003 , w7004 , w7005 , w7006 , w7007 , w7008 , w7009 , w7010 , w7011 , w7012 , w7013 , w7014 , w7015 , w7016 , w7017 , w7018 , w7019 , w7020 , w7021 , w7022 , w7023 , w7024 , w7025 , w7026 , w7027 , w7028 , w7029 , w7030 , w7031 , w7032 , w7033 , w7034 , w7035 , w7036 , w7037 , w7038 , w7039 , w7040 , w7041 , w7042 , w7043 , w7044 , w7045 , w7046 , w7047 , w7048 , w7049 , w7050 , w7051 , w7052 , w7053 , w7054 , w7055 , w7056 , w7057 , w7058 , w7059 , w7060 , w7061 , w7062 , w7063 , w7064 , w7065 , w7066 , w7067 , w7068 , w7069 , w7070 , w7071 , w7072 , w7073 , w7074 , w7075 , w7076 , w7077 , w7078 , w7079 , w7080 , w7081 , w7082 , w7083 , w7084 , w7085 , w7086 , w7087 , w7088 , w7089 , w7090 , w7091 , w7092 , w7093 , w7094 , w7095 , w7096 , w7097 , w7098 , w7099 , w7100 , w7101 , w7102 , w7103 , w7104 , w7105 , w7106 , w7107 , w7108 , w7109 , w7110 , w7111 , w7112 , w7113 , w7114 , w7115 , w7116 , w7117 , w7118 , w7119 , w7120 , w7121 , w7122 , w7123 , w7124 , w7125 , w7126 , w7127 , w7128 , w7129 , w7130 , w7131 , w7132 , w7133 , w7134 , w7135 , w7136 , w7137 , w7138 , w7139 , w7140 , w7141 , w7142 , w7143 , w7144 , w7145 , w7146 , w7147 , w7148 , w7149 , w7150 , w7151 , w7152 , w7153 , w7154 , w7155 , w7156 , w7157 , w7158 , w7159 , w7160 , w7161 , w7162 , w7163 , w7164 , w7165 , w7166 , w7167 , w7168 , w7169 , w7170 , w7171 , w7172 , w7173 , w7174 , w7175 , w7176 , w7177 , w7178 , w7179 , w7180 , w7181 , w7182 , w7183 , w7184 , w7185 , w7186 , w7187 , w7188 , w7189 , w7190 , w7191 , w7192 , w7193 , w7194 , w7195 , w7196 , w7197 , w7198 , w7199 , w7200 , w7201 , w7202 , w7203 , w7204 , w7205 , w7206 , w7207 , w7208 , w7209 , w7210 , w7211 , w7212 , w7213 , w7214 , w7215 , w7216 , w7217 , w7218 , w7219 , w7220 , w7221 , w7222 , w7223 , w7224 , w7225 , w7226 , w7227 , w7228 , w7229 , w7230 , w7231 , w7232 , w7233 , w7234 , w7235 , w7236 , w7237 , w7238 , w7239 , w7240 , w7241 , w7242 , w7243 , w7244 , w7245 , w7246 , w7247 , w7248 , w7249 , w7250 , w7251 , w7252 , w7253 , w7254 , w7255 , w7256 , w7257 , w7258 , w7259 , w7260 , w7261 , w7262 , w7263 , w7264 , w7265 , w7266 , w7267 , w7268 , w7269 , w7270 , w7271 , w7272 , w7273 , w7274 , w7275 , w7276 , w7277 , w7278 , w7279 , w7280 , w7281 , w7282 , w7283 , w7284 , w7285 , w7286 , w7287 , w7288 , w7289 , w7290 , w7291 , w7292 , w7293 , w7294 , w7295 , w7296 , w7297 , w7298 , w7299 , w7300 , w7301 , w7302 , w7303 , w7304 , w7305 , w7306 , w7307 , w7308 , w7309 , w7310 , w7311 , w7312 , w7313 , w7314 , w7315 , w7316 , w7317 , w7318 , w7319 , w7320 , w7321 , w7322 , w7323 , w7324 , w7325 , w7326 , w7327 , w7328 , w7329 , w7330 , w7331 , w7332 , w7333 , w7334 , w7335 , w7336 , w7337 , w7338 , w7339 , w7340 , w7341 , w7342 , w7343 , w7344 , w7345 , w7346 , w7347 , w7348 , w7349 , w7350 , w7351 , w7352 , w7353 , w7354 , w7355 , w7356 , w7357 , w7358 , w7359 , w7360 , w7361 , w7362 , w7363 , w7364 , w7365 , w7366 , w7367 , w7368 , w7369 , w7370 , w7371 , w7372 , w7373 , w7374 , w7375 , w7376 , w7377 , w7378 , w7379 , w7380 , w7381 , w7382 , w7383 , w7384 , w7385 , w7386 , w7387 , w7388 , w7389 , w7390 , w7391 , w7392 , w7393 , w7394 , w7395 , w7396 , w7397 , w7398 , w7399 , w7400 , w7401 , w7402 , w7403 , w7404 , w7405 , w7406 , w7407 , w7408 , w7409 , w7410 , w7411 , w7412 , w7413 , w7414 , w7415 , w7416 , w7417 , w7418 , w7419 , w7420 , w7421 , w7422 , w7423 , w7424 , w7425 , w7426 , w7427 , w7428 , w7429 , w7430 , w7431 , w7432 , w7433 , w7434 , w7435 , w7436 , w7437 , w7438 , w7439 , w7440 , w7441 , w7442 , w7443 , w7444 , w7445 , w7446 , w7447 , w7448 , w7449 , w7450 , w7451 , w7452 , w7453 , w7454 , w7455 , w7456 , w7457 , w7458 , w7459 , w7460 , w7461 , w7462 , w7463 , w7464 , w7465 , w7466 , w7467 , w7468 , w7469 , w7470 , w7471 , w7472 , w7473 , w7474 , w7475 , w7476 , w7477 , w7478 , w7479 , w7480 , w7481 , w7482 , w7483 , w7484 , w7485 , w7486 , w7487 , w7488 , w7489 , w7490 , w7491 , w7492 , w7493 , w7494 , w7495 , w7496 , w7497 , w7498 , w7499 , w7500 , w7501 , w7502 , w7503 , w7504 , w7505 , w7506 , w7507 , w7508 , w7509 , w7510 , w7511 , w7512 , w7513 , w7514 , w7515 , w7516 , w7517 , w7518 , w7519 , w7520 , w7521 , w7522 , w7523 , w7524 , w7525 , w7526 , w7527 , w7528 , w7529 , w7530 , w7531 , w7532 , w7533 , w7534 , w7535 , w7536 , w7537 , w7538 , w7539 , w7540 , w7541 , w7542 , w7543 , w7544 , w7545 , w7546 , w7547 , w7548 , w7549 , w7550 , w7551 , w7552 , w7553 , w7554 , w7555 , w7556 , w7557 , w7558 , w7559 , w7560 , w7561 , w7562 , w7563 , w7564 , w7565 , w7566 , w7567 , w7568 , w7569 , w7570 , w7571 , w7572 , w7573 , w7574 , w7575 , w7576 , w7577 , w7578 , w7579 , w7580 , w7581 , w7582 , w7583 , w7584 , w7585 , w7586 , w7587 , w7588 , w7589 , w7590 , w7591 , w7592 , w7593 , w7594 , w7595 , w7596 , w7597 , w7598 , w7599 , w7600 , w7601 , w7602 , w7603 , w7604 , w7605 , w7606 , w7607 , w7608 , w7609 , w7610 , w7611 , w7612 , w7613 , w7614 , w7615 , w7616 , w7617 , w7618 , w7619 , w7620 , w7621 , w7622 , w7623 , w7624 , w7625 , w7626 , w7627 , w7628 , w7629 , w7630 , w7631 , w7632 , w7633 , w7634 , w7635 , w7636 , w7637 , w7638 , w7639 , w7640 , w7641 , w7642 , w7643 , w7644 , w7645 , w7646 , w7647 , w7648 , w7649 , w7650 , w7651 , w7652 , w7653 , w7654 , w7655 , w7656 , w7657 , w7658 , w7659 , w7660 , w7661 , w7662 , w7663 , w7664 , w7665 , w7666 , w7667 , w7668 , w7669 , w7670 , w7671 , w7672 , w7673 , w7674 , w7675 , w7676 , w7677 , w7678 , w7679 , w7680 , w7681 , w7682 , w7683 , w7684 , w7685 , w7686 , w7687 , w7688 , w7689 , w7690 , w7691 , w7692 , w7693 , w7694 , w7695 , w7696 , w7697 , w7698 , w7699 , w7700 , w7701 , w7702 , w7703 , w7704 , w7705 , w7706 , w7707 , w7708 , w7709 , w7710 , w7711 , w7712 , w7713 , w7714 , w7715 , w7716 , w7717 , w7718 , w7719 , w7720 , w7721 , w7722 , w7723 , w7724 , w7725 , w7726 , w7727 , w7728 , w7729 , w7730 , w7731 , w7732 , w7733 , w7734 , w7735 , w7736 , w7737 , w7738 , w7739 , w7740 , w7741 , w7742 , w7743 , w7744 , w7745 , w7746 , w7747 , w7748 , w7749 , w7750 , w7751 , w7752 , w7753 , w7754 , w7755 , w7756 , w7757 , w7758 , w7759 , w7760 , w7761 , w7762 , w7763 , w7764 , w7765 , w7766 , w7767 , w7768 , w7769 , w7770 , w7771 , w7772 , w7773 , w7774 , w7775 , w7776 , w7777 , w7778 , w7779 , w7780 , w7781 , w7782 , w7783 , w7784 , w7785 , w7786 , w7787 , w7788 , w7789 , w7790 , w7791 , w7792 , w7793 , w7794 , w7795 , w7796 , w7797 , w7798 , w7799 , w7800 , w7801 , w7802 , w7803 , w7804 , w7805 , w7806 , w7807 , w7808 , w7809 , w7810 , w7811 , w7812 , w7813 , w7814 , w7815 , w7816 , w7817 , w7818 , w7819 , w7820 , w7821 , w7822 , w7823 , w7824 , w7825 , w7826 , w7827 , w7828 , w7829 , w7830 , w7831 , w7832 , w7833 , w7834 , w7835 , w7836 , w7837 , w7838 , w7839 , w7840 , w7841 , w7842 , w7843 , w7844 , w7845 , w7846 , w7847 , w7848 , w7849 , w7850 , w7851 , w7852 , w7853 , w7854 , w7855 , w7856 , w7857 , w7858 , w7859 , w7860 , w7861 , w7862 , w7863 , w7864 , w7865 , w7866 , w7867 , w7868 , w7869 , w7870 , w7871 , w7872 , w7873 , w7874 , w7875 , w7876 , w7877 , w7878 , w7879 , w7880 , w7881 , w7882 , w7883 , w7884 , w7885 , w7886 , w7887 , w7888 , w7889 , w7890 , w7891 , w7892 , w7893 , w7894 , w7895 , w7896 , w7897 , w7898 , w7899 , w7900 , w7901 , w7902 , w7903 , w7904 , w7905 , w7906 , w7907 , w7908 , w7909 , w7910 , w7911 , w7912 , w7913 , w7914 , w7915 , w7916 , w7917 , w7918 , w7919 , w7920 , w7921 , w7922 , w7923 , w7924 , w7925 , w7926 , w7927 , w7928 , w7929 , w7930 , w7931 , w7932 , w7933 , w7934 , w7935 , w7936 , w7937 , w7938 , w7939 , w7940 , w7941 , w7942 , w7943 , w7944 , w7945 , w7946 , w7947 , w7948 , w7949 , w7950 , w7951 , w7952 , w7953 , w7954 , w7955 , w7956 , w7957 , w7958 , w7959 , w7960 , w7961 , w7962 , w7963 , w7964 , w7965 , w7966 , w7967 , w7968 , w7969 , w7970 , w7971 , w7972 , w7973 , w7974 , w7975 , w7976 , w7977 , w7978 , w7979 , w7980 , w7981 , w7982 , w7983 , w7984 , w7985 , w7986 , w7987 , w7988 , w7989 , w7990 , w7991 , w7992 , w7993 , w7994 , w7995 , w7996 , w7997 , w7998 , w7999 , w8000 , w8001 , w8002 , w8003 , w8004 , w8005 , w8006 , w8007 , w8008 , w8009 , w8010 , w8011 , w8012 , w8013 , w8014 , w8015 , w8016 , w8017 , w8018 , w8019 , w8020 , w8021 , w8022 , w8023 , w8024 , w8025 , w8026 , w8027 , w8028 , w8029 , w8030 , w8031 , w8032 , w8033 , w8034 , w8035 , w8036 , w8037 , w8038 , w8039 , w8040 , w8041 , w8042 , w8043 , w8044 , w8045 , w8046 , w8047 , w8048 , w8049 , w8050 , w8051 , w8052 , w8053 , w8054 , w8055 , w8056 , w8057 , w8058 , w8059 , w8060 , w8061 , w8062 , w8063 , w8064 , w8065 , w8066 , w8067 , w8068 , w8069 , w8070 , w8071 , w8072 , w8073 , w8074 , w8075 , w8076 , w8077 , w8078 , w8079 , w8080 , w8081 , w8082 , w8083 , w8084 , w8085 , w8086 , w8087 , w8088 , w8089 , w8090 , w8091 , w8092 , w8093 , w8094 , w8095 , w8096 , w8097 , w8098 , w8099 , w8100 , w8101 , w8102 , w8103 , w8104 , w8105 , w8106 , w8107 , w8108 , w8109 , w8110 , w8111 , w8112 , w8113 , w8114 , w8115 , w8116 , w8117 , w8118 , w8119 , w8120 , w8121 , w8122 , w8123 , w8124 , w8125 , w8126 , w8127 , w8128 , w8129 , w8130 , w8131 , w8132 , w8133 , w8134 , w8135 , w8136 , w8137 , w8138 , w8139 , w8140 , w8141 , w8142 , w8143 , w8144 , w8145 , w8146 , w8147 , w8148 , w8149 , w8150 , w8151 , w8152 , w8153 , w8154 , w8155 , w8156 , w8157 , w8158 , w8159 , w8160 , w8161 , w8162 , w8163 , w8164 , w8165 , w8166 , w8167 , w8168 , w8169 , w8170 , w8171 , w8172 , w8173 , w8174 , w8175 , w8176 , w8177 , w8178 , w8179 , w8180 , w8181 , w8182 , w8183 , w8184 , w8185 , w8186 , w8187 , w8188 , w8189 , w8190 , w8191 , w8192 , w8193 , w8194 , w8195 , w8196 , w8197 , w8198 , w8199 , w8200 , w8201 , w8202 , w8203 , w8204 , w8205 , w8206 , w8207 , w8208 , w8209 , w8210 , w8211 , w8212 , w8213 , w8214 , w8215 , w8216 , w8217 , w8218 , w8219 , w8220 , w8221 , w8222 , w8223 , w8224 , w8225 , w8226 , w8227 , w8228 , w8229 , w8230 , w8231 , w8232 , w8233 , w8234 , w8235 , w8236 , w8237 , w8238 , w8239 , w8240 , w8241 , w8242 , w8243 , w8244 , w8245 , w8246 , w8247 , w8248 , w8249 , w8250 , w8251 , w8252 , w8253 , w8254 , w8255 , w8256 , w8257 , w8258 , w8259 , w8260 , w8261 , w8262 , w8263 , w8264 , w8265 , w8266 , w8267 , w8268 , w8269 , w8270 , w8271 , w8272 , w8273 , w8274 , w8275 , w8276 , w8277 , w8278 , w8279 , w8280 , w8281 , w8282 , w8283 , w8284 , w8285 , w8286 , w8287 , w8288 , w8289 , w8290 , w8291 , w8292 , w8293 , w8294 , w8295 , w8296 , w8297 , w8298 , w8299 , w8300 , w8301 , w8302 , w8303 , w8304 , w8305 , w8306 , w8307 , w8308 , w8309 , w8310 , w8311 , w8312 , w8313 , w8314 , w8315 , w8316 , w8317 , w8318 , w8319 , w8320 , w8321 , w8322 , w8323 , w8324 , w8325 , w8326 , w8327 , w8328 , w8329 , w8330 , w8331 , w8332 , w8333 , w8334 , w8335 , w8336 , w8337 , w8338 , w8339 , w8340 , w8341 , w8342 , w8343 , w8344 , w8345 , w8346 , w8347 , w8348 , w8349 , w8350 , w8351 , w8352 , w8353 , w8354 , w8355 , w8356 , w8357 , w8358 , w8359 , w8360 , w8361 , w8362 , w8363 , w8364 , w8365 , w8366 , w8367 , w8368 , w8369 , w8370 , w8371 , w8372 , w8373 , w8374 , w8375 , w8376 , w8377 , w8378 , w8379 , w8380 , w8381 , w8382 , w8383 , w8384 , w8385 , w8386 , w8387 , w8388 , w8389 , w8390 , w8391 , w8392 , w8393 , w8394 , w8395 , w8396 , w8397 , w8398 , w8399 , w8400 , w8401 , w8402 , w8403 , w8404 , w8405 , w8406 , w8407 , w8408 , w8409 , w8410 , w8411 , w8412 , w8413 , w8414 , w8415 , w8416 , w8417 , w8418 , w8419 , w8420 , w8421 , w8422 , w8423 , w8424 , w8425 , w8426 , w8427 , w8428 , w8429 , w8430 , w8431 , w8432 , w8433 , w8434 , w8435 , w8436 , w8437 , w8438 , w8439 , w8440 , w8441 , w8442 , w8443 , w8444 , w8445 , w8446 , w8447 , w8448 , w8449 , w8450 , w8451 , w8452 , w8453 , w8454 , w8455 , w8456 , w8457 , w8458 , w8459 , w8460 , w8461 , w8462 , w8463 , w8464 , w8465 , w8466 , w8467 , w8468 , w8469 , w8470 , w8471 , w8472 , w8473 , w8474 , w8475 , w8476 , w8477 , w8478 , w8479 , w8480 , w8481 , w8482 , w8483 , w8484 , w8485 , w8486 , w8487 , w8488 , w8489 , w8490 , w8491 , w8492 , w8493 , w8494 , w8495 , w8496 , w8497 , w8498 , w8499 , w8500 , w8501 , w8502 , w8503 , w8504 , w8505 , w8506 , w8507 , w8508 , w8509 , w8510 , w8511 , w8512 , w8513 , w8514 , w8515 , w8516 , w8517 , w8518 , w8519 , w8520 , w8521 , w8522 , w8523 , w8524 , w8525 , w8526 , w8527 , w8528 , w8529 , w8530 , w8531 , w8532 , w8533 , w8534 , w8535 , w8536 , w8537 , w8538 , w8539 , w8540 , w8541 , w8542 , w8543 , w8544 , w8545 , w8546 , w8547 , w8548 , w8549 , w8550 , w8551 , w8552 , w8553 , w8554 , w8555 , w8556 , w8557 , w8558 , w8559 , w8560 , w8561 , w8562 , w8563 , w8564 , w8565 , w8566 , w8567 , w8568 , w8569 , w8570 , w8571 , w8572 , w8573 , w8574 , w8575 , w8576 , w8577 , w8578 , w8579 , w8580 , w8581 , w8582 , w8583 , w8584 , w8585 , w8586 , w8587 , w8588 , w8589 , w8590 , w8591 , w8592 , w8593 , w8594 , w8595 , w8596 , w8597 , w8598 , w8599 , w8600 , w8601 , w8602 , w8603 , w8604 , w8605 , w8606 , w8607 , w8608 , w8609 , w8610 , w8611 , w8612 , w8613 , w8614 , w8615 , w8616 , w8617 , w8618 , w8619 , w8620 , w8621 , w8622 , w8623 , w8624 , w8625 , w8626 , w8627 , w8628 , w8629 , w8630 , w8631 , w8632 , w8633 , w8634 , w8635 , w8636 , w8637 , w8638 , w8639 , w8640 , w8641 , w8642 , w8643 , w8644 , w8645 , w8646 , w8647 , w8648 , w8649 , w8650 , w8651 , w8652 , w8653 , w8654 , w8655 , w8656 , w8657 , w8658 , w8659 , w8660 , w8661 , w8662 , w8663 , w8664 , w8665 , w8666 , w8667 , w8668 , w8669 , w8670 , w8671 , w8672 , w8673 , w8674 , w8675 , w8676 , w8677 , w8678 , w8679 , w8680 , w8681 , w8682 , w8683 , w8684 , w8685 , w8686 , w8687 , w8688 , w8689 , w8690 , w8691 , w8692 , w8693 , w8694 , w8695 , w8696 , w8697 , w8698 , w8699 , w8700 , w8701 , w8702 , w8703 , w8704 , w8705 , w8706 , w8707 , w8708 , w8709 , w8710 , w8711 , w8712 , w8713 , w8714 , w8715 , w8716 , w8717 , w8718 , w8719 , w8720 , w8721 , w8722 , w8723 , w8724 , w8725 , w8726 , w8727 , w8728 , w8729 , w8730 , w8731 , w8732 , w8733 , w8734 , w8735 , w8736 , w8737 , w8738 , w8739 , w8740 , w8741 , w8742 , w8743 , w8744 , w8745 , w8746 , w8747 , w8748 , w8749 , w8750 , w8751 , w8752 , w8753 , w8754 , w8755 , w8756 , w8757 , w8758 , w8759 , w8760 , w8761 , w8762 , w8763 , w8764 , w8765 , w8766 , w8767 , w8768 , w8769 , w8770 , w8771 , w8772 , w8773 , w8774 , w8775 , w8776 , w8777 , w8778 , w8779 , w8780 , w8781 , w8782 , w8783 , w8784 , w8785 , w8786 , w8787 , w8788 , w8789 , w8790 , w8791 , w8792 , w8793 , w8794 , w8795 , w8796 , w8797 , w8798 , w8799 , w8800 , w8801 , w8802 , w8803 , w8804 , w8805 , w8806 , w8807 , w8808 , w8809 , w8810 , w8811 , w8812 , w8813 , w8814 , w8815 , w8816 , w8817 , w8818 , w8819 , w8820 , w8821 , w8822 , w8823 , w8824 , w8825 , w8826 , w8827 , w8828 , w8829 , w8830 , w8831 , w8832 , w8833 , w8834 , w8835 , w8836 , w8837 , w8838 , w8839 , w8840 , w8841 , w8842 , w8843 , w8844 , w8845 , w8846 , w8847 , w8848 , w8849 , w8850 , w8851 , w8852 , w8853 , w8854 , w8855 , w8856 , w8857 , w8858 , w8859 , w8860 , w8861 , w8862 , w8863 , w8864 , w8865 , w8866 , w8867 , w8868 , w8869 , w8870 , w8871 , w8872 , w8873 , w8874 , w8875 , w8876 , w8877 , w8878 , w8879 , w8880 , w8881 , w8882 , w8883 , w8884 , w8885 , w8886 , w8887 , w8888 , w8889 , w8890 , w8891 , w8892 , w8893 , w8894 , w8895 , w8896 , w8897 , w8898 , w8899 , w8900 , w8901 , w8902 , w8903 , w8904 , w8905 , w8906 , w8907 , w8908 , w8909 , w8910 , w8911 , w8912 , w8913 , w8914 , w8915 , w8916 , w8917 , w8918 , w8919 , w8920 , w8921 , w8922 , w8923 , w8924 , w8925 , w8926 , w8927 , w8928 , w8929 , w8930 , w8931 , w8932 , w8933 , w8934 , w8935 , w8936 , w8937 , w8938 , w8939 , w8940 , w8941 , w8942 , w8943 , w8944 , w8945 , w8946 , w8947 , w8948 , w8949 , w8950 , w8951 , w8952 , w8953 , w8954 , w8955 , w8956 , w8957 , w8958 , w8959 , w8960 , w8961 , w8962 , w8963 , w8964 , w8965 , w8966 , w8967 , w8968 , w8969 , w8970 , w8971 , w8972 , w8973 , w8974 , w8975 , w8976 , w8977 , w8978 , w8979 , w8980 , w8981 , w8982 , w8983 , w8984 , w8985 , w8986 , w8987 , w8988 , w8989 , w8990 , w8991 , w8992 , w8993 , w8994 , w8995 , w8996 , w8997 , w8998 , w8999 , w9000 , w9001 , w9002 , w9003 , w9004 , w9005 , w9006 , w9007 , w9008 , w9009 , w9010 , w9011 , w9012 , w9013 , w9014 , w9015 , w9016 , w9017 , w9018 , w9019 , w9020 , w9021 , w9022 , w9023 , w9024 , w9025 , w9026 , w9027 , w9028 , w9029 , w9030 , w9031 , w9032 , w9033 , w9034 , w9035 , w9036 , w9037 , w9038 , w9039 , w9040 , w9041 , w9042 , w9043 , w9044 , w9045 , w9046 , w9047 , w9048 , w9049 , w9050 , w9051 , w9052 , w9053 , w9054 , w9055 , w9056 , w9057 , w9058 , w9059 , w9060 , w9061 , w9062 , w9063 , w9064 , w9065 , w9066 , w9067 , w9068 , w9069 , w9070 , w9071 , w9072 , w9073 , w9074 , w9075 , w9076 , w9077 , w9078 , w9079 , w9080 , w9081 , w9082 , w9083 , w9084 , w9085 , w9086 , w9087 , w9088 , w9089 , w9090 , w9091 , w9092 , w9093 , w9094 , w9095 , w9096 , w9097 , w9098 , w9099 , w9100 , w9101 , w9102 , w9103 , w9104 , w9105 , w9106 , w9107 , w9108 , w9109 , w9110 , w9111 , w9112 , w9113 , w9114 , w9115 , w9116 , w9117 , w9118 , w9119 , w9120 , w9121 , w9122 , w9123 , w9124 , w9125 , w9126 , w9127 , w9128 , w9129 , w9130 , w9131 , w9132 , w9133 , w9134 , w9135 , w9136 , w9137 , w9138 , w9139 , w9140 , w9141 , w9142 , w9143 , w9144 , w9145 , w9146 , w9147 , w9148 , w9149 , w9150 , w9151 , w9152 , w9153 , w9154 , w9155 , w9156 , w9157 , w9158 , w9159 , w9160 , w9161 , w9162 , w9163 , w9164 , w9165 , w9166 , w9167 , w9168 , w9169 , w9170 , w9171 , w9172 , w9173 , w9174 , w9175 , w9176 , w9177 , w9178 , w9179 , w9180 , w9181 , w9182 , w9183 , w9184 , w9185 , w9186 , w9187 , w9188 , w9189 , w9190 , w9191 , w9192 , w9193 , w9194 , w9195 , w9196 , w9197 , w9198 , w9199 , w9200 , w9201 , w9202 , w9203 , w9204 , w9205 , w9206 , w9207 , w9208 , w9209 , w9210 , w9211 , w9212 , w9213 , w9214 , w9215 , w9216 , w9217 , w9218 , w9219 , w9220 , w9221 , w9222 , w9223 , w9224 , w9225 , w9226 , w9227 , w9228 , w9229 , w9230 , w9231 , w9232 , w9233 , w9234 , w9235 , w9236 , w9237 , w9238 , w9239 , w9240 , w9241 , w9242 , w9243 , w9244 , w9245 , w9246 , w9247 , w9248 , w9249 , w9250 , w9251 , w9252 , w9253 , w9254 , w9255 , w9256 , w9257 , w9258 , w9259 , w9260 , w9261 , w9262 , w9263 , w9264 , w9265 , w9266 , w9267 , w9268 , w9269 , w9270 , w9271 , w9272 , w9273 , w9274 , w9275 , w9276 , w9277 , w9278 , w9279 , w9280 , w9281 , w9282 , w9283 , w9284 , w9285 , w9286 , w9287 , w9288 , w9289 , w9290 , w9291 , w9292 , w9293 , w9294 , w9295 , w9296 , w9297 , w9298 , w9299 , w9300 , w9301 , w9302 , w9303 , w9304 , w9305 , w9306 , w9307 , w9308 , w9309 , w9310 , w9311 , w9312 , w9313 , w9314 , w9315 , w9316 , w9317 , w9318 , w9319 , w9320 , w9321 , w9322 , w9323 , w9324 , w9325 , w9326 , w9327 , w9328 , w9329 , w9330 , w9331 , w9332 , w9333 , w9334 , w9335 , w9336 , w9337 , w9338 , w9339 , w9340 , w9341 , w9342 , w9343 , w9344 , w9345 , w9346 , w9347 , w9348 , w9349 , w9350 , w9351 , w9352 , w9353 , w9354 , w9355 , w9356 , w9357 , w9358 , w9359 , w9360 , w9361 , w9362 , w9363 , w9364 , w9365 , w9366 , w9367 , w9368 , w9369 , w9370 , w9371 , w9372 , w9373 , w9374 , w9375 , w9376 , w9377 , w9378 , w9379 , w9380 , w9381 , w9382 , w9383 , w9384 , w9385 , w9386 , w9387 , w9388 , w9389 , w9390 , w9391 , w9392 , w9393 , w9394 , w9395 , w9396 , w9397 , w9398 , w9399 , w9400 , w9401 , w9402 , w9403 , w9404 , w9405 , w9406 , w9407 , w9408 , w9409 , w9410 , w9411 , w9412 , w9413 , w9414 , w9415 , w9416 , w9417 , w9418 , w9419 , w9420 , w9421 , w9422 , w9423 , w9424 , w9425 , w9426 , w9427 , w9428 , w9429 , w9430 , w9431 , w9432 , w9433 , w9434 , w9435 , w9436 , w9437 , w9438 , w9439 , w9440 , w9441 , w9442 , w9443 , w9444 , w9445 , w9446 , w9447 , w9448 , w9449 , w9450 , w9451 , w9452 , w9453 , w9454 , w9455 , w9456 , w9457 , w9458 , w9459 , w9460 , w9461 , w9462 , w9463 , w9464 , w9465 , w9466 , w9467 , w9468 , w9469 , w9470 , w9471 , w9472 , w9473 , w9474 , w9475 , w9476 , w9477 , w9478 , w9479 , w9480 , w9481 , w9482 , w9483 , w9484 , w9485 , w9486 , w9487 , w9488 , w9489 , w9490 , w9491 , w9492 , w9493 , w9494 , w9495 , w9496 , w9497 , w9498 , w9499 , w9500 , w9501 , w9502 , w9503 , w9504 , w9505 , w9506 , w9507 , w9508 , w9509 , w9510 , w9511 , w9512 , w9513 , w9514 , w9515 , w9516 , w9517 , w9518 , w9519 , w9520 , w9521 , w9522 , w9523 , w9524 , w9525 , w9526 , w9527 , w9528 , w9529 , w9530 , w9531 , w9532 , w9533 , w9534 , w9535 , w9536 , w9537 , w9538 , w9539 , w9540 , w9541 , w9542 , w9543 , w9544 , w9545 , w9546 , w9547 , w9548 , w9549 , w9550 , w9551 , w9552 , w9553 , w9554 , w9555 , w9556 , w9557 , w9558 , w9559 , w9560 , w9561 , w9562 , w9563 , w9564 , w9565 , w9566 , w9567 , w9568 , w9569 , w9570 , w9571 , w9572 , w9573 , w9574 , w9575 , w9576 , w9577 , w9578 , w9579 , w9580 , w9581 , w9582 , w9583 , w9584 , w9585 , w9586 , w9587 , w9588 , w9589 , w9590 , w9591 , w9592 , w9593 , w9594 , w9595 , w9596 , w9597 , w9598 , w9599 , w9600 , w9601 , w9602 , w9603 , w9604 , w9605 , w9606 , w9607 , w9608 , w9609 , w9610 , w9611 , w9612 , w9613 , w9614 , w9615 , w9616 , w9617 , w9618 , w9619 , w9620 , w9621 , w9622 , w9623 , w9624 , w9625 , w9626 , w9627 , w9628 , w9629 , w9630 , w9631 , w9632 , w9633 , w9634 , w9635 , w9636 , w9637 , w9638 , w9639 , w9640 , w9641 , w9642 , w9643 , w9644 , w9645 , w9646 , w9647 , w9648 , w9649 , w9650 , w9651 , w9652 , w9653 , w9654 , w9655 , w9656 , w9657 , w9658 , w9659 , w9660 , w9661 , w9662 , w9663 , w9664 , w9665 , w9666 , w9667 , w9668 , w9669 , w9670 , w9671 , w9672 , w9673 , w9674 , w9675 , w9676 , w9677 , w9678 , w9679 , w9680 , w9681 , w9682 , w9683 , w9684 , w9685 , w9686 , w9687 , w9688 , w9689 , w9690 , w9691 , w9692 , w9693 , w9694 , w9695 , w9696 , w9697 , w9698 , w9699 , w9700 , w9701 , w9702 , w9703 , w9704 , w9705 , w9706 , w9707 , w9708 , w9709 , w9710 , w9711 , w9712 , w9713 , w9714 , w9715 , w9716 , w9717 , w9718 , w9719 , w9720 , w9721 , w9722 , w9723 , w9724 , w9725 , w9726 , w9727 , w9728 , w9729 , w9730 , w9731 , w9732 , w9733 , w9734 , w9735 , w9736 , w9737 , w9738 , w9739 , w9740 , w9741 , w9742 , w9743 , w9744 , w9745 , w9746 , w9747 , w9748 , w9749 , w9750 , w9751 , w9752 , w9753 , w9754 , w9755 , w9756 , w9757 , w9758 , w9759 , w9760 , w9761 , w9762 , w9763 , w9764 , w9765 , w9766 , w9767 , w9768 , w9769 , w9770 , w9771 , w9772 , w9773 , w9774 , w9775 , w9776 , w9777 , w9778 , w9779 , w9780 , w9781 , w9782 , w9783 , w9784 , w9785 , w9786 , w9787 , w9788 , w9789 , w9790 , w9791 , w9792 , w9793 , w9794 , w9795 , w9796 , w9797 , w9798 , w9799 , w9800 , w9801 , w9802 , w9803 , w9804 , w9805 , w9806 , w9807 , w9808 , w9809 , w9810 , w9811 , w9812 , w9813 , w9814 , w9815 , w9816 , w9817 , w9818 , w9819 , w9820 , w9821 , w9822 , w9823 , w9824 , w9825 , w9826 , w9827 , w9828 , w9829 , w9830 , w9831 , w9832 , w9833 , w9834 , w9835 , w9836 , w9837 , w9838 , w9839 , w9840 , w9841 , w9842 , w9843 , w9844 , w9845 , w9846 , w9847 , w9848 , w9849 , w9850 , w9851 , w9852 , w9853 , w9854 , w9855 , w9856 , w9857 , w9858 , w9859 , w9860 , w9861 , w9862 , w9863 , w9864 , w9865 , w9866 , w9867 , w9868 , w9869 , w9870 , w9871 , w9872 , w9873 , w9874 , w9875 , w9876 , w9877 , w9878 , w9879 , w9880 , w9881 , w9882 , w9883 , w9884 , w9885 , w9886 , w9887 , w9888 , w9889 , w9890 , w9891 , w9892 , w9893 , w9894 , w9895 , w9896 , w9897 , w9898 , w9899 , w9900 , w9901 , w9902 , w9903 , w9904 , w9905 , w9906 , w9907 , w9908 , w9909 , w9910 , w9911 , w9912 , w9913 , w9914 , w9915 , w9916 , w9917 , w9918 , w9919 , w9920 , w9921 , w9922 , w9923 , w9924 , w9925 , w9926 , w9927 , w9928 , w9929 , w9930 , w9931 , w9932 , w9933 , w9934 , w9935 , w9936 , w9937 , w9938 , w9939 , w9940 , w9941 , w9942 , w9943 , w9944 , w9945 , w9946 , w9947 , w9948 , w9949 , w9950 , w9951 , w9952 , w9953 , w9954 , w9955 , w9956 , w9957 , w9958 , w9959 , w9960 , w9961 , w9962 , w9963 , w9964 , w9965 , w9966 , w9967 , w9968 , w9969 , w9970 , w9971 , w9972 , w9973 , w9974 , w9975 , w9976 , w9977 , w9978 , w9979 , w9980 , w9981 , w9982 , w9983 , w9984 , w9985 , w9986 , w9987 , w9988 , w9989 , w9990 , w9991 , w9992 , w9993 , w9994 , w9995 , w9996 , w9997 , w9998 , w9999 , w10000 , w10001 , w10002 , w10003 , w10004 , w10005 , w10006 , w10007 , w10008 , w10009 , w10010 , w10011 , w10012 , w10013 , w10014 , w10015 , w10016 , w10017 , w10018 , w10019 , w10020 , w10021 , w10022 , w10023 , w10024 , w10025 , w10026 , w10027 , w10028 , w10029 , w10030 , w10031 , w10032 , w10033 , w10034 , w10035 , w10036 , w10037 , w10038 , w10039 , w10040 , w10041 , w10042 , w10043 , w10044 , w10045 , w10046 , w10047 , w10048 , w10049 , w10050 , w10051 , w10052 , w10053 , w10054 , w10055 , w10056 , w10057 , w10058 , w10059 , w10060 , w10061 , w10062 , w10063 , w10064 , w10065 , w10066 , w10067 , w10068 , w10069 , w10070 , w10071 , w10072 , w10073 , w10074 , w10075 , w10076 , w10077 , w10078 , w10079 , w10080 , w10081 , w10082 , w10083 , w10084 , w10085 , w10086 , w10087 , w10088 , w10089 , w10090 , w10091 , w10092 , w10093 , w10094 , w10095 , w10096 , w10097 , w10098 , w10099 , w10100 , w10101 , w10102 , w10103 , w10104 , w10105 , w10106 , w10107 , w10108 , w10109 , w10110 , w10111 , w10112 , w10113 , w10114 , w10115 , w10116 , w10117 , w10118 , w10119 , w10120 , w10121 , w10122 , w10123 , w10124 , w10125 , w10126 , w10127 , w10128 , w10129 , w10130 , w10131 , w10132 , w10133 , w10134 , w10135 , w10136 , w10137 , w10138 , w10139 , w10140 , w10141 , w10142 , w10143 , w10144 , w10145 , w10146 , w10147 , w10148 , w10149 , w10150 , w10151 , w10152 , w10153 , w10154 , w10155 , w10156 , w10157 , w10158 , w10159 , w10160 , w10161 , w10162 , w10163 , w10164 , w10165 , w10166 , w10167 , w10168 , w10169 , w10170 , w10171 , w10172 , w10173 , w10174 , w10175 , w10176 , w10177 , w10178 , w10179 , w10180 , w10181 , w10182 , w10183 , w10184 , w10185 , w10186 , w10187 , w10188 , w10189 , w10190 , w10191 , w10192 , w10193 , w10194 , w10195 , w10196 , w10197 , w10198 , w10199 , w10200 , w10201 , w10202 , w10203 , w10204 , w10205 , w10206 , w10207 , w10208 , w10209 , w10210 , w10211 , w10212 , w10213 , w10214 , w10215 , w10216 , w10217 , w10218 , w10219 , w10220 , w10221 , w10222 , w10223 , w10224 , w10225 , w10226 , w10227 , w10228 , w10229 , w10230 , w10231 , w10232 , w10233 , w10234 , w10235 , w10236 , w10237 , w10238 , w10239 , w10240 , w10241 , w10242 , w10243 , w10244 , w10245 , w10246 , w10247 , w10248 , w10249 , w10250 , w10251 , w10252 , w10253 , w10254 , w10255 , w10256 , w10257 , w10258 , w10259 , w10260 , w10261 , w10262 , w10263 , w10264 , w10265 , w10266 , w10267 , w10268 , w10269 , w10270 , w10271 , w10272 , w10273 , w10274 , w10275 , w10276 , w10277 , w10278 , w10279 , w10280 , w10281 , w10282 , w10283 , w10284 , w10285 , w10286 , w10287 , w10288 , w10289 , w10290 , w10291 , w10292 , w10293 , w10294 , w10295 , w10296 , w10297 , w10298 , w10299 , w10300 , w10301 , w10302 , w10303 , w10304 , w10305 , w10306 , w10307 , w10308 , w10309 , w10310 , w10311 , w10312 , w10313 , w10314 , w10315 , w10316 , w10317 , w10318 , w10319 , w10320 , w10321 , w10322 , w10323 , w10324 , w10325 , w10326 , w10327 , w10328 , w10329 , w10330 , w10331 , w10332 , w10333 , w10334 , w10335 , w10336 , w10337 , w10338 , w10339 , w10340 , w10341 , w10342 , w10343 , w10344 , w10345 , w10346 , w10347 , w10348 , w10349 , w10350 , w10351 , w10352 , w10353 , w10354 , w10355 , w10356 , w10357 , w10358 , w10359 , w10360 , w10361 , w10362 , w10363 , w10364 , w10365 , w10366 , w10367 , w10368 , w10369 , w10370 , w10371 , w10372 , w10373 , w10374 , w10375 , w10376 , w10377 , w10378 , w10379 , w10380 , w10381 , w10382 , w10383 , w10384 , w10385 , w10386 , w10387 , w10388 , w10389 , w10390 , w10391 , w10392 , w10393 , w10394 , w10395 , w10396 , w10397 , w10398 , w10399 , w10400 , w10401 , w10402 , w10403 , w10404 , w10405 , w10406 , w10407 , w10408 , w10409 , w10410 , w10411 , w10412 , w10413 , w10414 , w10415 , w10416 , w10417 , w10418 , w10419 , w10420 , w10421 , w10422 , w10423 , w10424 , w10425 , w10426 , w10427 , w10428 , w10429 , w10430 , w10431 , w10432 , w10433 , w10434 , w10435 , w10436 , w10437 , w10438 , w10439 , w10440 , w10441 , w10442 , w10443 , w10444 , w10445 , w10446 , w10447 , w10448 , w10449 , w10450 , w10451 , w10452 , w10453 , w10454 , w10455 , w10456 , w10457 , w10458 , w10459 , w10460 , w10461 , w10462 , w10463 , w10464 , w10465 , w10466 , w10467 , w10468 , w10469 , w10470 , w10471 , w10472 , w10473 , w10474 , w10475 , w10476 , w10477 , w10478 , w10479 , w10480 , w10481 , w10482 , w10483 , w10484 , w10485 , w10486 , w10487 , w10488 , w10489 , w10490 , w10491 , w10492 , w10493 , w10494 , w10495 , w10496 , w10497 , w10498 , w10499 , w10500 , w10501 , w10502 , w10503 , w10504 , w10505 , w10506 , w10507 , w10508 , w10509 , w10510 , w10511 , w10512 , w10513 , w10514 , w10515 , w10516 , w10517 , w10518 , w10519 , w10520 , w10521 , w10522 , w10523 , w10524 , w10525 , w10526 , w10527 , w10528 , w10529 , w10530 , w10531 , w10532 , w10533 , w10534 , w10535 , w10536 , w10537 , w10538 , w10539 , w10540 , w10541 , w10542 , w10543 , w10544 , w10545 , w10546 , w10547 , w10548 , w10549 , w10550 , w10551 , w10552 , w10553 , w10554 , w10555 , w10556 , w10557 , w10558 , w10559 , w10560 , w10561 , w10562 , w10563 , w10564 , w10565 , w10566 , w10567 , w10568 , w10569 , w10570 , w10571 , w10572 , w10573 , w10574 , w10575 , w10576 , w10577 , w10578 , w10579 , w10580 , w10581 , w10582 , w10583 , w10584 , w10585 , w10586 , w10587 , w10588 , w10589 , w10590 , w10591 , w10592 , w10593 , w10594 , w10595 , w10596 , w10597 , w10598 , w10599 , w10600 , w10601 , w10602 , w10603 , w10604 , w10605 , w10606 , w10607 , w10608 , w10609 , w10610 , w10611 , w10612 , w10613 , w10614 , w10615 , w10616 , w10617 , w10618 , w10619 , w10620 , w10621 , w10622 , w10623 , w10624 , w10625 , w10626 , w10627 , w10628 , w10629 , w10630 , w10631 , w10632 , w10633 , w10634 , w10635 , w10636 , w10637 , w10638 , w10639 , w10640 , w10641 , w10642 , w10643 , w10644 , w10645 , w10646 , w10647 , w10648 , w10649 , w10650 , w10651 , w10652 , w10653 , w10654 , w10655 , w10656 , w10657 , w10658 , w10659 , w10660 , w10661 , w10662 , w10663 , w10664 , w10665 , w10666 , w10667 , w10668 , w10669 , w10670 , w10671 , w10672 , w10673 , w10674 , w10675 , w10676 , w10677 , w10678 , w10679 , w10680 , w10681 , w10682 , w10683 , w10684 , w10685 , w10686 , w10687 , w10688 , w10689 , w10690 , w10691 , w10692 , w10693 , w10694 , w10695 , w10696 , w10697 , w10698 , w10699 , w10700 , w10701 , w10702 , w10703 , w10704 , w10705 , w10706 , w10707 , w10708 , w10709 , w10710 , w10711 , w10712 , w10713 , w10714 , w10715 , w10716 , w10717 , w10718 , w10719 , w10720 , w10721 , w10722 , w10723 , w10724 , w10725 , w10726 , w10727 , w10728 , w10729 , w10730 , w10731 , w10732 , w10733 , w10734 , w10735 , w10736 , w10737 , w10738 , w10739 , w10740 , w10741 , w10742 , w10743 , w10744 , w10745 , w10746 , w10747 , w10748 , w10749 , w10750 , w10751 , w10752 , w10753 , w10754 , w10755 , w10756 , w10757 , w10758 , w10759 , w10760 , w10761 , w10762 , w10763 , w10764 , w10765 , w10766 , w10767 , w10768 , w10769 , w10770 , w10771 , w10772 , w10773 , w10774 , w10775 , w10776 , w10777 , w10778 , w10779 , w10780 , w10781 , w10782 , w10783 , w10784 , w10785 , w10786 , w10787 , w10788 , w10789 , w10790 , w10791 , w10792 , w10793 , w10794 , w10795 , w10796 , w10797 , w10798 , w10799 , w10800 , w10801 , w10802 , w10803 , w10804 , w10805 , w10806 , w10807 , w10808 , w10809 , w10810 , w10811 , w10812 , w10813 , w10814 , w10815 , w10816 , w10817 , w10818 , w10819 , w10820 , w10821 , w10822 , w10823 , w10824 , w10825 , w10826 , w10827 , w10828 , w10829 , w10830 , w10831 , w10832 , w10833 , w10834 , w10835 , w10836 , w10837 , w10838 , w10839 , w10840 , w10841 , w10842 , w10843 , w10844 , w10845 , w10846 , w10847 , w10848 , w10849 , w10850 , w10851 , w10852 , w10853 , w10854 , w10855 , w10856 , w10857 , w10858 , w10859 , w10860 , w10861 , w10862 , w10863 , w10864 , w10865 , w10866 , w10867 , w10868 , w10869 , w10870 , w10871 , w10872 , w10873 , w10874 , w10875 , w10876 , w10877 , w10878 , w10879 , w10880 , w10881 , w10882 , w10883 , w10884 , w10885 , w10886 , w10887 , w10888 , w10889 , w10890 , w10891 , w10892 , w10893 , w10894 , w10895 , w10896 , w10897 , w10898 , w10899 , w10900 , w10901 , w10902 , w10903 , w10904 , w10905 , w10906 , w10907 , w10908 , w10909 , w10910 , w10911 , w10912 , w10913 , w10914 , w10915 , w10916 , w10917 , w10918 , w10919 , w10920 , w10921 , w10922 , w10923 , w10924 , w10925 , w10926 , w10927 , w10928 , w10929 , w10930 , w10931 , w10932 , w10933 , w10934 , w10935 , w10936 , w10937 , w10938 , w10939 , w10940 , w10941 , w10942 , w10943 , w10944 , w10945 , w10946 , w10947 , w10948 , w10949 , w10950 , w10951 , w10952 , w10953 , w10954 , w10955 , w10956 , w10957 , w10958 , w10959 , w10960 , w10961 , w10962 , w10963 , w10964 , w10965 , w10966 , w10967 , w10968 , w10969 , w10970 , w10971 , w10972 , w10973 , w10974 , w10975 , w10976 , w10977 , w10978 , w10979 , w10980 , w10981 , w10982 , w10983 , w10984 , w10985 , w10986 , w10987 , w10988 , w10989 , w10990 , w10991 , w10992 , w10993 , w10994 , w10995 , w10996 , w10997 , w10998 , w10999 , w11000 , w11001 , w11002 , w11003 , w11004 , w11005 , w11006 , w11007 , w11008 , w11009 , w11010 , w11011 , w11012 , w11013 , w11014 , w11015 , w11016 , w11017 , w11018 , w11019 , w11020 , w11021 , w11022 , w11023 , w11024 , w11025 , w11026 , w11027 , w11028 , w11029 , w11030 , w11031 , w11032 , w11033 , w11034 , w11035 , w11036 , w11037 , w11038 , w11039 , w11040 , w11041 , w11042 , w11043 , w11044 , w11045 , w11046 , w11047 , w11048 , w11049 , w11050 , w11051 , w11052 , w11053 , w11054 , w11055 , w11056 , w11057 , w11058 , w11059 , w11060 , w11061 , w11062 , w11063 , w11064 , w11065 , w11066 , w11067 , w11068 , w11069 , w11070 , w11071 , w11072 , w11073 , w11074 , w11075 , w11076 , w11077 , w11078 , w11079 , w11080 , w11081 , w11082 , w11083 , w11084 , w11085 , w11086 , w11087 , w11088 , w11089 , w11090 , w11091 , w11092 , w11093 , w11094 , w11095 , w11096 , w11097 , w11098 , w11099 , w11100 , w11101 , w11102 , w11103 , w11104 , w11105 , w11106 , w11107 , w11108 , w11109 , w11110 , w11111 , w11112 , w11113 , w11114 , w11115 , w11116 , w11117 , w11118 , w11119 , w11120 , w11121 , w11122 , w11123 , w11124 , w11125 , w11126 , w11127 , w11128 , w11129 , w11130 , w11131 , w11132 , w11133 , w11134 , w11135 , w11136 , w11137 , w11138 , w11139 , w11140 , w11141 , w11142 , w11143 , w11144 , w11145 , w11146 , w11147 , w11148 , w11149 , w11150 , w11151 , w11152 , w11153 , w11154 , w11155 , w11156 , w11157 , w11158 , w11159 , w11160 , w11161 , w11162 , w11163 , w11164 , w11165 , w11166 , w11167 , w11168 , w11169 , w11170 , w11171 , w11172 , w11173 , w11174 , w11175 , w11176 , w11177 , w11178 , w11179 , w11180 , w11181 , w11182 , w11183 , w11184 , w11185 , w11186 , w11187 , w11188 , w11189 , w11190 , w11191 , w11192 , w11193 , w11194 , w11195 , w11196 , w11197 , w11198 , w11199 , w11200 , w11201 , w11202 , w11203 , w11204 , w11205 , w11206 , w11207 , w11208 , w11209 , w11210 , w11211 , w11212 , w11213 , w11214 , w11215 , w11216 , w11217 , w11218 , w11219 , w11220 , w11221 , w11222 , w11223 , w11224 , w11225 , w11226 , w11227 , w11228 , w11229 , w11230 , w11231 , w11232 , w11233 , w11234 , w11235 , w11236 , w11237 , w11238 , w11239 , w11240 , w11241 , w11242 , w11243 , w11244 , w11245 , w11246 , w11247 , w11248 , w11249 , w11250 , w11251 , w11252 , w11253 , w11254 , w11255 , w11256 , w11257 , w11258 , w11259 , w11260 , w11261 , w11262 , w11263 , w11264 , w11265 , w11266 , w11267 , w11268 , w11269 , w11270 , w11271 , w11272 , w11273 , w11274 , w11275 , w11276 , w11277 , w11278 , w11279 , w11280 , w11281 , w11282 , w11283 , w11284 , w11285 , w11286 , w11287 , w11288 , w11289 , w11290 , w11291 , w11292 , w11293 , w11294 , w11295 , w11296 , w11297 , w11298 , w11299 , w11300 , w11301 , w11302 , w11303 , w11304 , w11305 , w11306 , w11307 , w11308 , w11309 , w11310 , w11311 , w11312 , w11313 , w11314 , w11315 , w11316 , w11317 , w11318 , w11319 , w11320 , w11321 , w11322 , w11323 , w11324 , w11325 , w11326 , w11327 , w11328 , w11329 , w11330 , w11331 , w11332 , w11333 , w11334 , w11335 , w11336 , w11337 , w11338 , w11339 , w11340 , w11341 , w11342 , w11343 , w11344 , w11345 , w11346 , w11347 , w11348 , w11349 , w11350 , w11351 , w11352 , w11353 , w11354 , w11355 , w11356 , w11357 , w11358 , w11359 , w11360 , w11361 , w11362 , w11363 , w11364 , w11365 , w11366 , w11367 , w11368 , w11369 , w11370 , w11371 , w11372 , w11373 , w11374 , w11375 , w11376 , w11377 , w11378 , w11379 , w11380 , w11381 , w11382 , w11383 , w11384 , w11385 , w11386 , w11387 , w11388 , w11389 , w11390 , w11391 , w11392 , w11393 , w11394 , w11395 , w11396 , w11397 , w11398 , w11399 , w11400 , w11401 , w11402 , w11403 , w11404 , w11405 , w11406 , w11407 , w11408 , w11409 , w11410 , w11411 , w11412 , w11413 , w11414 , w11415 , w11416 , w11417 , w11418 , w11419 , w11420 , w11421 , w11422 , w11423 , w11424 , w11425 , w11426 , w11427 , w11428 , w11429 , w11430 , w11431 , w11432 , w11433 , w11434 , w11435 , w11436 , w11437 , w11438 , w11439 , w11440 , w11441 , w11442 , w11443 , w11444 , w11445 , w11446 , w11447 , w11448 , w11449 , w11450 , w11451 , w11452 , w11453 , w11454 , w11455 , w11456 , w11457 , w11458 , w11459 , w11460 , w11461 , w11462 , w11463 , w11464 , w11465 , w11466 , w11467 , w11468 , w11469 , w11470 , w11471 , w11472 , w11473 , w11474 , w11475 , w11476 , w11477 , w11478 , w11479 , w11480 , w11481 , w11482 , w11483 , w11484 , w11485 , w11486 , w11487 , w11488 , w11489 , w11490 , w11491 , w11492 , w11493 , w11494 , w11495 , w11496 , w11497 , w11498 , w11499 , w11500 , w11501 , w11502 , w11503 , w11504 , w11505 , w11506 , w11507 , w11508 , w11509 , w11510 , w11511 , w11512 , w11513 , w11514 , w11515 , w11516 , w11517 , w11518 , w11519 , w11520 , w11521 , w11522 , w11523 , w11524 , w11525 , w11526 , w11527 , w11528 , w11529 , w11530 , w11531 , w11532 , w11533 , w11534 , w11535 , w11536 , w11537 , w11538 , w11539 , w11540 , w11541 , w11542 , w11543 , w11544 , w11545 , w11546 , w11547 , w11548 , w11549 , w11550 , w11551 , w11552 , w11553 , w11554 , w11555 , w11556 , w11557 , w11558 , w11559 , w11560 , w11561 , w11562 , w11563 , w11564 , w11565 , w11566 , w11567 , w11568 , w11569 , w11570 , w11571 , w11572 , w11573 , w11574 , w11575 , w11576 , w11577 , w11578 , w11579 , w11580 , w11581 , w11582 , w11583 , w11584 , w11585 , w11586 , w11587 , w11588 , w11589 , w11590 , w11591 , w11592 , w11593 , w11594 , w11595 , w11596 , w11597 , w11598 , w11599 , w11600 , w11601 , w11602 , w11603 , w11604 , w11605 , w11606 , w11607 , w11608 , w11609 , w11610 , w11611 , w11612 , w11613 , w11614 , w11615 , w11616 , w11617 , w11618 , w11619 , w11620 , w11621 , w11622 , w11623 , w11624 , w11625 , w11626 , w11627 , w11628 , w11629 , w11630 , w11631 , w11632 , w11633 , w11634 , w11635 , w11636 , w11637 , w11638 , w11639 , w11640 , w11641 , w11642 , w11643 , w11644 , w11645 , w11646 , w11647 , w11648 , w11649 , w11650 , w11651 , w11652 , w11653 , w11654 , w11655 , w11656 , w11657 , w11658 , w11659 , w11660 , w11661 , w11662 , w11663 , w11664 , w11665 , w11666 , w11667 , w11668 , w11669 , w11670 , w11671 , w11672 , w11673 , w11674 , w11675 , w11676 , w11677 , w11678 , w11679 , w11680 , w11681 , w11682 , w11683 , w11684 , w11685 , w11686 , w11687 , w11688 , w11689 , w11690 , w11691 , w11692 , w11693 , w11694 , w11695 , w11696 , w11697 , w11698 , w11699 , w11700 , w11701 , w11702 , w11703 , w11704 , w11705 , w11706 , w11707 , w11708 , w11709 , w11710 , w11711 , w11712 , w11713 , w11714 , w11715 , w11716 , w11717 , w11718 , w11719 , w11720 , w11721 , w11722 , w11723 , w11724 , w11725 , w11726 , w11727 , w11728 , w11729 , w11730 , w11731 , w11732 , w11733 , w11734 , w11735 , w11736 , w11737 , w11738 , w11739 , w11740 , w11741 , w11742 , w11743 , w11744 , w11745 , w11746 , w11747 , w11748 , w11749 , w11750 , w11751 , w11752 , w11753 , w11754 , w11755 , w11756 , w11757 , w11758 , w11759 , w11760 , w11761 , w11762 , w11763 , w11764 , w11765 , w11766 , w11767 , w11768 , w11769 , w11770 , w11771 , w11772 , w11773 , w11774 , w11775 , w11776 , w11777 , w11778 , w11779 , w11780 , w11781 , w11782 , w11783 , w11784 , w11785 , w11786 , w11787 , w11788 , w11789 , w11790 , w11791 , w11792 , w11793 , w11794 , w11795 , w11796 , w11797 , w11798 , w11799 , w11800 , w11801 , w11802 , w11803 , w11804 , w11805 , w11806 , w11807 , w11808 , w11809 , w11810 , w11811 , w11812 , w11813 , w11814 , w11815 , w11816 , w11817 , w11818 , w11819 , w11820 , w11821 , w11822 , w11823 , w11824 , w11825 , w11826 , w11827 , w11828 , w11829 , w11830 , w11831 , w11832 , w11833 , w11834 , w11835 , w11836 , w11837 , w11838 , w11839 , w11840 , w11841 , w11842 , w11843 , w11844 , w11845 , w11846 , w11847 , w11848 , w11849 , w11850 , w11851 , w11852 , w11853 , w11854 , w11855 , w11856 , w11857 , w11858 , w11859 , w11860 , w11861 , w11862 , w11863 , w11864 , w11865 , w11866 , w11867 , w11868 , w11869 , w11870 , w11871 , w11872 , w11873 , w11874 , w11875 , w11876 , w11877 , w11878 , w11879 , w11880 , w11881 , w11882 , w11883 , w11884 , w11885 , w11886 , w11887 , w11888 , w11889 , w11890 , w11891 , w11892 , w11893 , w11894 , w11895 , w11896 , w11897 , w11898 , w11899 , w11900 , w11901 , w11902 , w11903 , w11904 , w11905 , w11906 , w11907 , w11908 , w11909 , w11910 , w11911 , w11912 , w11913 , w11914 , w11915 , w11916 , w11917 , w11918 , w11919 , w11920 , w11921 , w11922 , w11923 , w11924 , w11925 , w11926 , w11927 , w11928 , w11929 , w11930 , w11931 , w11932 , w11933 , w11934 , w11935 , w11936 , w11937 , w11938 , w11939 , w11940 , w11941 , w11942 , w11943 , w11944 , w11945 , w11946 , w11947 , w11948 , w11949 , w11950 , w11951 , w11952 , w11953 , w11954 , w11955 , w11956 , w11957 , w11958 , w11959 , w11960 , w11961 , w11962 , w11963 , w11964 , w11965 , w11966 , w11967 , w11968 , w11969 , w11970 , w11971 , w11972 , w11973 , w11974 , w11975 , w11976 , w11977 , w11978 , w11979 , w11980 , w11981 , w11982 , w11983 , w11984 , w11985 , w11986 , w11987 , w11988 , w11989 , w11990 , w11991 , w11992 , w11993 , w11994 , w11995 , w11996 , w11997 , w11998 , w11999 , w12000 , w12001 , w12002 , w12003 , w12004 , w12005 , w12006 , w12007 , w12008 , w12009 , w12010 , w12011 , w12012 , w12013 , w12014 , w12015 , w12016 , w12017 , w12018 , w12019 , w12020 , w12021 , w12022 , w12023 , w12024 , w12025 , w12026 , w12027 , w12028 , w12029 , w12030 , w12031 , w12032 , w12033 , w12034 , w12035 , w12036 , w12037 , w12038 , w12039 , w12040 , w12041 , w12042 , w12043 , w12044 , w12045 , w12046 , w12047 , w12048 , w12049 , w12050 , w12051 , w12052 , w12053 , w12054 , w12055 , w12056 , w12057 , w12058 , w12059 , w12060 , w12061 , w12062 , w12063 , w12064 , w12065 , w12066 , w12067 , w12068 , w12069 , w12070 , w12071 , w12072 , w12073 , w12074 , w12075 , w12076 , w12077 , w12078 , w12079 , w12080 , w12081 , w12082 , w12083 , w12084 , w12085 , w12086 , w12087 , w12088 , w12089 , w12090 , w12091 , w12092 , w12093 , w12094 , w12095 , w12096 , w12097 , w12098 , w12099 , w12100 , w12101 , w12102 , w12103 , w12104 , w12105 , w12106 , w12107 , w12108 , w12109 , w12110 , w12111 , w12112 , w12113 , w12114 , w12115 , w12116 , w12117 , w12118 , w12119 , w12120 , w12121 , w12122 , w12123 , w12124 , w12125 , w12126 , w12127 , w12128 , w12129 , w12130 , w12131 , w12132 , w12133 , w12134 , w12135 , w12136 , w12137 , w12138 , w12139 , w12140 , w12141 , w12142 , w12143 , w12144 , w12145 , w12146 , w12147 , w12148 , w12149 , w12150 , w12151 , w12152 , w12153 , w12154 , w12155 , w12156 , w12157 , w12158 , w12159 , w12160 , w12161 , w12162 , w12163 , w12164 , w12165 , w12166 , w12167 , w12168 , w12169 , w12170 , w12171 , w12172 , w12173 , w12174 , w12175 , w12176 , w12177 , w12178 , w12179 , w12180 , w12181 , w12182 , w12183 , w12184 , w12185 , w12186 , w12187 , w12188 , w12189 , w12190 , w12191 , w12192 , w12193 , w12194 , w12195 , w12196 , w12197 , w12198 , w12199 , w12200 , w12201 , w12202 , w12203 , w12204 , w12205 , w12206 , w12207 , w12208 , w12209 , w12210 , w12211 , w12212 , w12213 , w12214 , w12215 , w12216 , w12217 , w12218 , w12219 , w12220 , w12221 , w12222 , w12223 , w12224 , w12225 , w12226 , w12227 , w12228 , w12229 , w12230 , w12231 , w12232 , w12233 , w12234 , w12235 , w12236 , w12237 , w12238 , w12239 , w12240 , w12241 , w12242 , w12243 , w12244 , w12245 , w12246 , w12247 , w12248 , w12249 , w12250 , w12251 , w12252 , w12253 , w12254 , w12255 , w12256 , w12257 , w12258 , w12259 , w12260 , w12261 , w12262 , w12263 , w12264 , w12265 , w12266 , w12267 , w12268 , w12269 , w12270 , w12271 , w12272 , w12273 , w12274 , w12275 , w12276 , w12277 , w12278 , w12279 , w12280 , w12281 , w12282 , w12283 , w12284 , w12285 , w12286 , w12287 , w12288 , w12289 , w12290 , w12291 , w12292 , w12293 , w12294 , w12295 , w12296 , w12297 , w12298 , w12299 , w12300 , w12301 , w12302 , w12303 , w12304 , w12305 , w12306 , w12307 , w12308 , w12309 , w12310 , w12311 , w12312 , w12313 , w12314 , w12315 , w12316 , w12317 , w12318 , w12319 , w12320 , w12321 , w12322 , w12323 , w12324 , w12325 , w12326 , w12327 , w12328 , w12329 , w12330 , w12331 , w12332 , w12333 , w12334 , w12335 , w12336 , w12337 , w12338 , w12339 , w12340 , w12341 , w12342 , w12343 , w12344 , w12345 , w12346 , w12347 , w12348 , w12349 , w12350 , w12351 , w12352 , w12353 , w12354 , w12355 , w12356 , w12357 , w12358 , w12359 , w12360 , w12361 , w12362 , w12363 , w12364 , w12365 , w12366 , w12367 , w12368 , w12369 , w12370 , w12371 , w12372 , w12373 , w12374 , w12375 , w12376 , w12377 , w12378 , w12379 , w12380 , w12381 , w12382 , w12383 , w12384 , w12385 , w12386 , w12387 , w12388 , w12389 , w12390 , w12391 , w12392 , w12393 , w12394 , w12395 , w12396 , w12397 , w12398 , w12399 , w12400 , w12401 , w12402 , w12403 , w12404 , w12405 , w12406 , w12407 , w12408 , w12409 , w12410 , w12411 , w12412 , w12413 , w12414 , w12415 , w12416 , w12417 , w12418 , w12419 , w12420 , w12421 , w12422 , w12423 , w12424 , w12425 , w12426 , w12427 , w12428 , w12429 , w12430 , w12431 , w12432 , w12433 , w12434 , w12435 , w12436 , w12437 , w12438 , w12439 , w12440 , w12441 , w12442 , w12443 , w12444 , w12445 , w12446 , w12447 , w12448 , w12449 , w12450 , w12451 , w12452 , w12453 , w12454 , w12455 , w12456 , w12457 , w12458 , w12459 , w12460 , w12461 , w12462 , w12463 , w12464 , w12465 , w12466 , w12467 , w12468 , w12469 , w12470 , w12471 , w12472 , w12473 , w12474 , w12475 , w12476 , w12477 , w12478 , w12479 , w12480 , w12481 , w12482 , w12483 , w12484 , w12485 , w12486 , w12487 , w12488 , w12489 , w12490 , w12491 , w12492 , w12493 , w12494 , w12495 , w12496 , w12497 , w12498 , w12499 , w12500 , w12501 , w12502 , w12503 , w12504 , w12505 , w12506 , w12507 , w12508 , w12509 , w12510 , w12511 , w12512 , w12513 , w12514 , w12515 , w12516 , w12517 , w12518 , w12519 , w12520 , w12521 , w12522 , w12523 , w12524 , w12525 , w12526 , w12527 , w12528 , w12529 , w12530 , w12531 , w12532 , w12533 , w12534 , w12535 , w12536 , w12537 , w12538 , w12539 , w12540 , w12541 , w12542 , w12543 , w12544 , w12545 , w12546 , w12547 , w12548 , w12549 , w12550 , w12551 , w12552 , w12553 , w12554 , w12555 , w12556 , w12557 , w12558 , w12559 , w12560 , w12561 , w12562 , w12563 , w12564 , w12565 , w12566 , w12567 , w12568 , w12569 , w12570 , w12571 , w12572 , w12573 , w12574 , w12575 , w12576 , w12577 , w12578 , w12579 , w12580 , w12581 , w12582 , w12583 , w12584 , w12585 , w12586 , w12587 , w12588 , w12589 , w12590 , w12591 , w12592 , w12593 , w12594 , w12595 , w12596 , w12597 , w12598 , w12599 , w12600 , w12601 , w12602 , w12603 , w12604 , w12605 , w12606 , w12607 , w12608 , w12609 , w12610 , w12611 , w12612 , w12613 , w12614 , w12615 , w12616 , w12617 , w12618 , w12619 , w12620 , w12621 , w12622 , w12623 , w12624 , w12625 , w12626 , w12627 , w12628 , w12629 , w12630 , w12631 , w12632 , w12633 , w12634 , w12635 , w12636 , w12637 , w12638 , w12639 , w12640 , w12641 , w12642 , w12643 , w12644 , w12645 , w12646 , w12647 , w12648 , w12649 , w12650 , w12651 , w12652 , w12653 , w12654 , w12655 , w12656 , w12657 , w12658 , w12659 , w12660 , w12661 , w12662 , w12663 , w12664 , w12665 , w12666 , w12667 , w12668 , w12669 , w12670 , w12671 , w12672 , w12673 , w12674 , w12675 , w12676 , w12677 , w12678 , w12679 , w12680 , w12681 , w12682 , w12683 , w12684 , w12685 , w12686 , w12687 , w12688 , w12689 , w12690 , w12691 , w12692 , w12693 , w12694 , w12695 , w12696 , w12697 , w12698 , w12699 , w12700 , w12701 , w12702 , w12703 , w12704 , w12705 , w12706 , w12707 , w12708 , w12709 , w12710 , w12711 , w12712 , w12713 , w12714 , w12715 , w12716 , w12717 , w12718 , w12719 , w12720 , w12721 , w12722 , w12723 , w12724 , w12725 , w12726 , w12727 , w12728 , w12729 , w12730 , w12731 , w12732 , w12733 , w12734 , w12735 , w12736 , w12737 , w12738 , w12739 , w12740 , w12741 , w12742 , w12743 , w12744 , w12745 , w12746 , w12747 , w12748 , w12749 , w12750 , w12751 , w12752 , w12753 , w12754 , w12755 , w12756 , w12757 , w12758 , w12759 , w12760 , w12761 , w12762 , w12763 , w12764 , w12765 , w12766 , w12767 , w12768 , w12769 , w12770 , w12771 , w12772 , w12773 , w12774 , w12775 , w12776 , w12777 , w12778 , w12779 , w12780 , w12781 , w12782 , w12783 , w12784 , w12785 , w12786 , w12787 , w12788 , w12789 , w12790 , w12791 , w12792 , w12793 , w12794 , w12795 , w12796 , w12797 , w12798 , w12799 , w12800 , w12801 , w12802 , w12803 , w12804 , w12805 , w12806 , w12807 , w12808 , w12809 , w12810 , w12811 , w12812 , w12813 , w12814 , w12815 , w12816 , w12817 , w12818 , w12819 , w12820 , w12821 , w12822 , w12823 , w12824 , w12825 , w12826 , w12827 , w12828 , w12829 , w12830 , w12831 , w12832 , w12833 , w12834 , w12835 , w12836 , w12837 , w12838 , w12839 , w12840 , w12841 , w12842 , w12843 , w12844 , w12845 , w12846 , w12847 , w12848 , w12849 , w12850 , w12851 , w12852 , w12853 , w12854 , w12855 , w12856 , w12857 , w12858 , w12859 , w12860 , w12861 , w12862 , w12863 , w12864 , w12865 , w12866 , w12867 , w12868 , w12869 , w12870 , w12871 , w12872 , w12873 , w12874 , w12875 , w12876 , w12877 , w12878 , w12879 , w12880 , w12881 , w12882 , w12883 , w12884 , w12885 , w12886 , w12887 , w12888 , w12889 , w12890 , w12891 , w12892 , w12893 , w12894 , w12895 , w12896 , w12897 , w12898 , w12899 , w12900 , w12901 , w12902 , w12903 , w12904 , w12905 , w12906 , w12907 , w12908 , w12909 , w12910 , w12911 , w12912 , w12913 , w12914 , w12915 , w12916 , w12917 , w12918 , w12919 , w12920 , w12921 , w12922 , w12923 , w12924 , w12925 , w12926 , w12927 , w12928 , w12929 , w12930 , w12931 , w12932 , w12933 , w12934 , w12935 , w12936 , w12937 , w12938 , w12939 , w12940 , w12941 , w12942 , w12943 , w12944 , w12945 , w12946 , w12947 , w12948 , w12949 , w12950 , w12951 , w12952 , w12953 , w12954 , w12955 , w12956 , w12957 , w12958 , w12959 , w12960 , w12961 , w12962 , w12963 , w12964 , w12965 , w12966 , w12967 , w12968 , w12969 , w12970 , w12971 , w12972 , w12973 , w12974 , w12975 , w12976 , w12977 , w12978 , w12979 , w12980 , w12981 , w12982 , w12983 , w12984 , w12985 , w12986 , w12987 , w12988 , w12989 , w12990 , w12991 , w12992 , w12993 , w12994 , w12995 , w12996 , w12997 , w12998 , w12999 , w13000 , w13001 , w13002 , w13003 , w13004 , w13005 , w13006 , w13007 , w13008 , w13009 , w13010 , w13011 , w13012 , w13013 , w13014 , w13015 , w13016 , w13017 , w13018 , w13019 , w13020 , w13021 , w13022 , w13023 , w13024 , w13025 , w13026 , w13027 , w13028 , w13029 , w13030 , w13031 , w13032 , w13033 , w13034 , w13035 , w13036 , w13037 , w13038 , w13039 , w13040 , w13041 , w13042 , w13043 , w13044 , w13045 , w13046 , w13047 , w13048 , w13049 , w13050 , w13051 , w13052 , w13053 , w13054 , w13055 , w13056 , w13057 , w13058 , w13059 , w13060 , w13061 , w13062 , w13063 , w13064 , w13065 , w13066 , w13067 , w13068 , w13069 , w13070 , w13071 , w13072 , w13073 , w13074 , w13075 , w13076 , w13077 , w13078 , w13079 , w13080 , w13081 , w13082 , w13083 , w13084 , w13085 , w13086 , w13087 , w13088 , w13089 , w13090 , w13091 , w13092 , w13093 , w13094 , w13095 , w13096 , w13097 , w13098 , w13099 , w13100 , w13101 , w13102 , w13103 , w13104 , w13105 , w13106 , w13107 , w13108 , w13109 , w13110 , w13111 , w13112 , w13113 , w13114 , w13115 , w13116 , w13117 , w13118 , w13119 , w13120 , w13121 , w13122 , w13123 , w13124 , w13125 , w13126 , w13127 , w13128 , w13129 , w13130 , w13131 , w13132 , w13133 , w13134 , w13135 , w13136 , w13137 , w13138 , w13139 , w13140 , w13141 , w13142 , w13143 , w13144 , w13145 , w13146 , w13147 , w13148 , w13149 , w13150 , w13151 , w13152 , w13153 , w13154 , w13155 , w13156 , w13157 , w13158 , w13159 , w13160 , w13161 , w13162 , w13163 , w13164 , w13165 , w13166 , w13167 , w13168 , w13169 , w13170 , w13171 , w13172 , w13173 , w13174 , w13175 , w13176 , w13177 , w13178 , w13179 , w13180 , w13181 , w13182 , w13183 , w13184 , w13185 , w13186 , w13187 , w13188 , w13189 , w13190 , w13191 , w13192 , w13193 , w13194 , w13195 , w13196 , w13197 , w13198 , w13199 , w13200 , w13201 , w13202 , w13203 , w13204 , w13205 , w13206 , w13207 , w13208 , w13209 , w13210 , w13211 , w13212 , w13213 , w13214 , w13215 , w13216 , w13217 , w13218 , w13219 , w13220 , w13221 , w13222 , w13223 , w13224 , w13225 , w13226 , w13227 , w13228 , w13229 , w13230 , w13231 , w13232 , w13233 , w13234 , w13235 , w13236 , w13237 , w13238 , w13239 , w13240 , w13241 , w13242 , w13243 , w13244 , w13245 , w13246 , w13247 , w13248 , w13249 , w13250 , w13251 , w13252 , w13253 , w13254 , w13255 , w13256 , w13257 , w13258 , w13259 , w13260 , w13261 , w13262 , w13263 , w13264 , w13265 , w13266 , w13267 , w13268 , w13269 , w13270 , w13271 , w13272 , w13273 , w13274 , w13275 , w13276 , w13277 , w13278 , w13279 , w13280 , w13281 , w13282 , w13283 , w13284 , w13285 , w13286 , w13287 , w13288 , w13289 , w13290 , w13291 , w13292 , w13293 , w13294 , w13295 , w13296 , w13297 , w13298 , w13299 , w13300 , w13301 , w13302 , w13303 , w13304 , w13305 , w13306 , w13307 , w13308 , w13309 , w13310 , w13311 , w13312 , w13313 , w13314 , w13315 , w13316 , w13317 , w13318 , w13319 , w13320 , w13321 , w13322 , w13323 , w13324 , w13325 , w13326 , w13327 , w13328 , w13329 , w13330 , w13331 , w13332 , w13333 , w13334 , w13335 , w13336 , w13337 , w13338 , w13339 , w13340 , w13341 , w13342 , w13343 , w13344 , w13345 , w13346 , w13347 , w13348 , w13349 , w13350 , w13351 , w13352 , w13353 , w13354 , w13355 , w13356 , w13357 , w13358 , w13359 , w13360 , w13361 , w13362 , w13363 , w13364 , w13365 , w13366 , w13367 , w13368 , w13369 , w13370 , w13371 , w13372 , w13373 , w13374 , w13375 , w13376 , w13377 , w13378 , w13379 , w13380 , w13381 , w13382 , w13383 , w13384 , w13385 , w13386 , w13387 , w13388 , w13389 , w13390 , w13391 , w13392 , w13393 , w13394 , w13395 , w13396 , w13397 , w13398 , w13399 , w13400 , w13401 , w13402 , w13403 , w13404 , w13405 , w13406 , w13407 , w13408 , w13409 , w13410 , w13411 , w13412 , w13413 , w13414 , w13415 , w13416 , w13417 , w13418 , w13419 , w13420 , w13421 , w13422 , w13423 , w13424 , w13425 , w13426 , w13427 , w13428 , w13429 , w13430 , w13431 , w13432 , w13433 , w13434 , w13435 , w13436 , w13437 , w13438 , w13439 , w13440 , w13441 , w13442 , w13443 , w13444 , w13445 , w13446 , w13447 , w13448 , w13449 , w13450 , w13451 , w13452 , w13453 , w13454 , w13455 , w13456 , w13457 , w13458 , w13459 , w13460 , w13461 , w13462 , w13463 , w13464 , w13465 , w13466 , w13467 , w13468 , w13469 , w13470 , w13471 , w13472 , w13473 , w13474 , w13475 , w13476 , w13477 , w13478 , w13479 , w13480 , w13481 , w13482 , w13483 , w13484 , w13485 , w13486 , w13487 , w13488 , w13489 , w13490 , w13491 , w13492 , w13493 , w13494 , w13495 , w13496 , w13497 , w13498 , w13499 , w13500 , w13501 , w13502 , w13503 , w13504 , w13505 , w13506 , w13507 , w13508 , w13509 , w13510 , w13511 , w13512 , w13513 , w13514 , w13515 , w13516 , w13517 , w13518 , w13519 , w13520 , w13521 , w13522 , w13523 , w13524 , w13525 , w13526 , w13527 , w13528 , w13529 , w13530 , w13531 , w13532 , w13533 , w13534 , w13535 , w13536 , w13537 , w13538 , w13539 , w13540 , w13541 , w13542 , w13543 , w13544 , w13545 , w13546 , w13547 , w13548 , w13549 , w13550 , w13551 , w13552 , w13553 , w13554 , w13555 , w13556 , w13557 , w13558 , w13559 , w13560 , w13561 , w13562 , w13563 , w13564 , w13565 , w13566 , w13567 , w13568 , w13569 , w13570 , w13571 , w13572 , w13573 , w13574 , w13575 , w13576 , w13577 , w13578 , w13579 , w13580 , w13581 , w13582 , w13583 , w13584 , w13585 , w13586 , w13587 , w13588 , w13589 , w13590 , w13591 , w13592 , w13593 , w13594 , w13595 , w13596 , w13597 , w13598 , w13599 , w13600 , w13601 , w13602 , w13603 , w13604 , w13605 , w13606 , w13607 , w13608 , w13609 , w13610 , w13611 , w13612 , w13613 , w13614 , w13615 , w13616 , w13617 , w13618 , w13619 , w13620 , w13621 , w13622 , w13623 , w13624 , w13625 , w13626 , w13627 , w13628 , w13629 , w13630 , w13631 , w13632 , w13633 , w13634 , w13635 , w13636 , w13637 , w13638 , w13639 , w13640 , w13641 , w13642 , w13643 , w13644 , w13645 , w13646 , w13647 , w13648 , w13649 , w13650 , w13651 , w13652 , w13653 , w13654 , w13655 , w13656 , w13657 , w13658 , w13659 , w13660 , w13661 , w13662 , w13663 , w13664 , w13665 , w13666 , w13667 , w13668 , w13669 , w13670 , w13671 , w13672 , w13673 , w13674 , w13675 , w13676 , w13677 , w13678 , w13679 , w13680 , w13681 , w13682 , w13683 , w13684 , w13685 , w13686 , w13687 , w13688 , w13689 , w13690 , w13691 , w13692 , w13693 , w13694 , w13695 , w13696 , w13697 , w13698 , w13699 , w13700 , w13701 , w13702 , w13703 , w13704 , w13705 , w13706 , w13707 , w13708 , w13709 , w13710 , w13711 , w13712 , w13713 , w13714 , w13715 , w13716 , w13717 , w13718 , w13719 , w13720 , w13721 , w13722 , w13723 , w13724 , w13725 , w13726 , w13727 , w13728 , w13729 , w13730 , w13731 , w13732 , w13733 , w13734 , w13735 , w13736 , w13737 , w13738 , w13739 , w13740 , w13741 , w13742 , w13743 , w13744 , w13745 , w13746 , w13747 , w13748 , w13749 , w13750 , w13751 , w13752 , w13753 , w13754 , w13755 , w13756 , w13757 , w13758 , w13759 , w13760 , w13761 , w13762 , w13763 , w13764 , w13765 , w13766 , w13767 , w13768 , w13769 , w13770 , w13771 , w13772 , w13773 , w13774 , w13775 , w13776 , w13777 , w13778 , w13779 , w13780 , w13781 , w13782 , w13783 , w13784 , w13785 , w13786 , w13787 , w13788 , w13789 , w13790 , w13791 , w13792 , w13793 , w13794 , w13795 , w13796 , w13797 , w13798 , w13799 , w13800 , w13801 , w13802 , w13803 , w13804 , w13805 , w13806 , w13807 , w13808 , w13809 , w13810 , w13811 , w13812 , w13813 , w13814 , w13815 , w13816 , w13817 , w13818 , w13819 , w13820 , w13821 , w13822 , w13823 , w13824 , w13825 , w13826 , w13827 , w13828 , w13829 , w13830 , w13831 , w13832 , w13833 , w13834 , w13835 , w13836 , w13837 , w13838 , w13839 , w13840 , w13841 , w13842 , w13843 , w13844 , w13845 , w13846 , w13847 , w13848 , w13849 , w13850 , w13851 , w13852 , w13853 , w13854 , w13855 , w13856 , w13857 , w13858 , w13859 , w13860 , w13861 , w13862 , w13863 , w13864 , w13865 , w13866 , w13867 , w13868 , w13869 , w13870 , w13871 , w13872 , w13873 , w13874 , w13875 , w13876 , w13877 , w13878 , w13879 , w13880 , w13881 , w13882 , w13883 , w13884 , w13885 , w13886 , w13887 , w13888 , w13889 , w13890 , w13891 , w13892 , w13893 , w13894 , w13895 , w13896 , w13897 , w13898 , w13899 , w13900 , w13901 , w13902 , w13903 , w13904 , w13905 , w13906 , w13907 , w13908 , w13909 , w13910 , w13911 , w13912 , w13913 , w13914 , w13915 , w13916 , w13917 , w13918 , w13919 , w13920 , w13921 , w13922 , w13923 , w13924 , w13925 , w13926 , w13927 , w13928 , w13929 , w13930 , w13931 , w13932 , w13933 , w13934 , w13935 , w13936 , w13937 , w13938 , w13939 , w13940 , w13941 , w13942 , w13943 , w13944 , w13945 , w13946 , w13947 , w13948 , w13949 , w13950 , w13951 , w13952 , w13953 , w13954 , w13955 , w13956 , w13957 , w13958 , w13959 , w13960 , w13961 , w13962 , w13963 , w13964 , w13965 , w13966 , w13967 , w13968 , w13969 , w13970 , w13971 , w13972 , w13973 , w13974 , w13975 , w13976 , w13977 , w13978 , w13979 , w13980 , w13981 , w13982 , w13983 , w13984 , w13985 , w13986 , w13987 , w13988 , w13989 , w13990 , w13991 , w13992 , w13993 , w13994 , w13995 , w13996 , w13997 , w13998 , w13999 , w14000 , w14001 , w14002 , w14003 , w14004 , w14005 , w14006 , w14007 , w14008 , w14009 , w14010 , w14011 , w14012 , w14013 , w14014 , w14015 , w14016 , w14017 , w14018 , w14019 , w14020 , w14021 , w14022 , w14023 , w14024 , w14025 , w14026 , w14027 , w14028 , w14029 , w14030 , w14031 , w14032 , w14033 , w14034 , w14035 , w14036 , w14037 , w14038 , w14039 , w14040 , w14041 , w14042 , w14043 , w14044 , w14045 , w14046 , w14047 , w14048 , w14049 , w14050 , w14051 , w14052 , w14053 , w14054 , w14055 , w14056 , w14057 , w14058 , w14059 , w14060 , w14061 , w14062 , w14063 , w14064 , w14065 , w14066 , w14067 , w14068 , w14069 , w14070 , w14071 , w14072 , w14073 , w14074 , w14075 , w14076 , w14077 , w14078 , w14079 , w14080 , w14081 , w14082 , w14083 , w14084 , w14085 , w14086 , w14087 , w14088 , w14089 , w14090 , w14091 , w14092 , w14093 , w14094 , w14095 , w14096 , w14097 , w14098 , w14099 , w14100 , w14101 , w14102 , w14103 , w14104 , w14105 , w14106 , w14107 , w14108 , w14109 , w14110 , w14111 , w14112 , w14113 , w14114 , w14115 , w14116 , w14117 , w14118 , w14119 , w14120 , w14121 , w14122 , w14123 , w14124 , w14125 , w14126 , w14127 , w14128 , w14129 , w14130 , w14131 , w14132 , w14133 , w14134 , w14135 , w14136 , w14137 , w14138 , w14139 , w14140 , w14141 , w14142 , w14143 , w14144 , w14145 , w14146 , w14147 , w14148 , w14149 , w14150 , w14151 , w14152 , w14153 , w14154 , w14155 , w14156 , w14157 , w14158 , w14159 , w14160 , w14161 , w14162 , w14163 , w14164 , w14165 , w14166 , w14167 , w14168 , w14169 , w14170 , w14171 , w14172 , w14173 , w14174 , w14175 , w14176 , w14177 , w14178 , w14179 , w14180 , w14181 , w14182 , w14183 , w14184 , w14185 , w14186 , w14187 , w14188 , w14189 , w14190 , w14191 , w14192 , w14193 , w14194 , w14195 , w14196 , w14197 , w14198 , w14199 , w14200 , w14201 , w14202 , w14203 , w14204 , w14205 , w14206 , w14207 , w14208 , w14209 , w14210 , w14211 , w14212 , w14213 , w14214 , w14215 , w14216 , w14217 , w14218 , w14219 , w14220 , w14221 , w14222 , w14223 , w14224 , w14225 , w14226 , w14227 , w14228 , w14229 , w14230 , w14231 , w14232 , w14233 , w14234 , w14235 , w14236 , w14237 , w14238 , w14239 , w14240 , w14241 , w14242 , w14243 , w14244 , w14245 , w14246 , w14247 , w14248 , w14249 , w14250 , w14251 , w14252 , w14253 , w14254 , w14255 , w14256 , w14257 , w14258 , w14259 , w14260 , w14261 , w14262 , w14263 , w14264 , w14265 , w14266 , w14267 , w14268 , w14269 , w14270 , w14271 , w14272 , w14273 , w14274 , w14275 , w14276 , w14277 , w14278 , w14279 , w14280 , w14281 , w14282 , w14283 , w14284 , w14285 , w14286 , w14287 , w14288 , w14289 , w14290 , w14291 , w14292 , w14293 , w14294 , w14295 , w14296 , w14297 , w14298 , w14299 , w14300 , w14301 , w14302 , w14303 , w14304 , w14305 , w14306 , w14307 , w14308 , w14309 , w14310 , w14311 , w14312 , w14313 , w14314 , w14315 , w14316 , w14317 , w14318 , w14319 , w14320 , w14321 , w14322 , w14323 , w14324 , w14325 , w14326 , w14327 , w14328 , w14329 , w14330 , w14331 , w14332 , w14333 , w14334 , w14335 , w14336 , w14337 , w14338 , w14339 , w14340 , w14341 , w14342 , w14343 , w14344 , w14345 , w14346 , w14347 , w14348 , w14349 , w14350 , w14351 , w14352 , w14353 , w14354 , w14355 , w14356 , w14357 , w14358 , w14359 , w14360 , w14361 , w14362 , w14363 , w14364 , w14365 , w14366 , w14367 , w14368 , w14369 , w14370 , w14371 , w14372 , w14373 , w14374 , w14375 , w14376 , w14377 , w14378 , w14379 , w14380 , w14381 , w14382 , w14383 , w14384 , w14385 , w14386 , w14387 , w14388 , w14389 , w14390 , w14391 , w14392 , w14393 , w14394 , w14395 , w14396 , w14397 , w14398 , w14399 , w14400 , w14401 , w14402 , w14403 , w14404 , w14405 , w14406 , w14407 , w14408 , w14409 , w14410 , w14411 , w14412 , w14413 , w14414 , w14415 , w14416 , w14417 , w14418 , w14419 , w14420 , w14421 , w14422 , w14423 , w14424 , w14425 , w14426 , w14427 , w14428 , w14429 , w14430 , w14431 , w14432 , w14433 , w14434 , w14435 , w14436 , w14437 , w14438 , w14439 , w14440 , w14441 , w14442 , w14443 , w14444 , w14445 , w14446 , w14447 , w14448 , w14449 , w14450 , w14451 , w14452 , w14453 , w14454 , w14455 , w14456 , w14457 , w14458 , w14459 , w14460 , w14461 , w14462 , w14463 , w14464 , w14465 , w14466 , w14467 , w14468 , w14469 , w14470 , w14471 , w14472 , w14473 , w14474 , w14475 , w14476 , w14477 , w14478 , w14479 , w14480 , w14481 , w14482 , w14483 , w14484 , w14485 , w14486 , w14487 , w14488 , w14489 , w14490 , w14491 , w14492 , w14493 , w14494 , w14495 , w14496 , w14497 , w14498 , w14499 , w14500 , w14501 , w14502 , w14503 , w14504 , w14505 , w14506 , w14507 , w14508 , w14509 , w14510 , w14511 , w14512 , w14513 , w14514 , w14515 , w14516 , w14517 , w14518 , w14519 , w14520 , w14521 , w14522 , w14523 , w14524 , w14525 , w14526 , w14527 , w14528 , w14529 , w14530 , w14531 , w14532 , w14533 , w14534 , w14535 , w14536 , w14537 , w14538 , w14539 , w14540 , w14541 , w14542 , w14543 , w14544 , w14545 , w14546 , w14547 , w14548 , w14549 , w14550 , w14551 , w14552 , w14553 , w14554 , w14555 , w14556 , w14557 , w14558 , w14559 , w14560 , w14561 , w14562 , w14563 , w14564 , w14565 , w14566 , w14567 , w14568 , w14569 , w14570 , w14571 , w14572 , w14573 , w14574 , w14575 , w14576 , w14577 , w14578 , w14579 , w14580 , w14581 , w14582 , w14583 , w14584 , w14585 , w14586 , w14587 , w14588 , w14589 , w14590 , w14591 , w14592 , w14593 , w14594 , w14595 , w14596 , w14597 , w14598 , w14599 , w14600 , w14601 , w14602 , w14603 , w14604 , w14605 , w14606 , w14607 , w14608 , w14609 , w14610 , w14611 , w14612 , w14613 , w14614 , w14615 , w14616 , w14617 , w14618 , w14619 , w14620 , w14621 , w14622 , w14623 , w14624 , w14625 , w14626 , w14627 , w14628 , w14629 , w14630 , w14631 , w14632 , w14633 , w14634 , w14635 , w14636 , w14637 , w14638 , w14639 , w14640 , w14641 , w14642 , w14643 , w14644 , w14645 , w14646 , w14647 , w14648 , w14649 , w14650 , w14651 , w14652 , w14653 , w14654 , w14655 , w14656 , w14657 , w14658 , w14659 , w14660 , w14661 , w14662 , w14663 , w14664 , w14665 , w14666 , w14667 , w14668 , w14669 , w14670 , w14671 , w14672 , w14673 , w14674 , w14675 , w14676 , w14677 , w14678 , w14679 , w14680 , w14681 , w14682 , w14683 , w14684 , w14685 , w14686 , w14687 , w14688 , w14689 , w14690 , w14691 , w14692 , w14693 , w14694 , w14695 , w14696 , w14697 , w14698 , w14699 , w14700 , w14701 , w14702 , w14703 , w14704 , w14705 , w14706 , w14707 , w14708 , w14709 , w14710 , w14711 , w14712 , w14713 , w14714 , w14715 , w14716 , w14717 , w14718 , w14719 , w14720 , w14721 , w14722 , w14723 , w14724 , w14725 , w14726 , w14727 , w14728 , w14729 , w14730 , w14731 , w14732 , w14733 , w14734 , w14735 , w14736 , w14737 , w14738 , w14739 , w14740 , w14741 , w14742 , w14743 , w14744 , w14745 , w14746 , w14747 , w14748 , w14749 , w14750 , w14751 , w14752 , w14753 , w14754 , w14755 , w14756 , w14757 , w14758 , w14759 , w14760 , w14761 , w14762 , w14763 , w14764 , w14765 , w14766 , w14767 , w14768 , w14769 , w14770 , w14771 , w14772 , w14773 , w14774 , w14775 , w14776 , w14777 , w14778 , w14779 , w14780 , w14781 , w14782 , w14783 , w14784 , w14785 , w14786 , w14787 , w14788 , w14789 , w14790 , w14791 , w14792 , w14793 , w14794 , w14795 , w14796 , w14797 , w14798 , w14799 , w14800 , w14801 , w14802 , w14803 , w14804 , w14805 , w14806 , w14807 , w14808 , w14809 , w14810 , w14811 , w14812 , w14813 , w14814 , w14815 , w14816 , w14817 , w14818 , w14819 , w14820 , w14821 , w14822 , w14823 , w14824 , w14825 , w14826 , w14827 , w14828 , w14829 , w14830 , w14831 , w14832 , w14833 , w14834 , w14835 , w14836 , w14837 , w14838 , w14839 , w14840 , w14841 , w14842 , w14843 , w14844 , w14845 , w14846 , w14847 , w14848 , w14849 , w14850 , w14851 , w14852 , w14853 , w14854 , w14855 , w14856 , w14857 , w14858 , w14859 , w14860 , w14861 , w14862 , w14863 , w14864 , w14865 , w14866 , w14867 , w14868 , w14869 , w14870 , w14871 , w14872 , w14873 , w14874 , w14875 , w14876 , w14877 , w14878 , w14879 , w14880 , w14881 , w14882 , w14883 , w14884 , w14885 , w14886 , w14887 , w14888 , w14889 , w14890 , w14891 , w14892 , w14893 , w14894 , w14895 , w14896 , w14897 , w14898 , w14899 , w14900 , w14901 , w14902 , w14903 , w14904 , w14905 , w14906 , w14907 , w14908 , w14909 , w14910 , w14911 , w14912 , w14913 , w14914 , w14915 , w14916 , w14917 , w14918 , w14919 , w14920 , w14921 , w14922 , w14923 , w14924 , w14925 , w14926 , w14927 , w14928 , w14929 , w14930 , w14931 , w14932 , w14933 , w14934 , w14935 , w14936 , w14937 , w14938 , w14939 , w14940 , w14941 , w14942 , w14943 , w14944 , w14945 , w14946 , w14947 , w14948 , w14949 , w14950 , w14951 , w14952 , w14953 , w14954 , w14955 , w14956 , w14957 , w14958 , w14959 , w14960 , w14961 , w14962 , w14963 , w14964 , w14965 , w14966 , w14967 , w14968 , w14969 , w14970 , w14971 , w14972 , w14973 , w14974 , w14975 , w14976 , w14977 , w14978 , w14979 , w14980 , w14981 , w14982 , w14983 , w14984 , w14985 , w14986 , w14987 , w14988 , w14989 , w14990 , w14991 , w14992 , w14993 , w14994 , w14995 , w14996 , w14997 , w14998 , w14999 , w15000 , w15001 , w15002 , w15003 , w15004 , w15005 , w15006 , w15007 , w15008 , w15009 , w15010 , w15011 , w15012 , w15013 , w15014 , w15015 , w15016 , w15017 , w15018 , w15019 , w15020 , w15021 , w15022 , w15023 , w15024 , w15025 , w15026 , w15027 , w15028 , w15029 , w15030 , w15031 , w15032 , w15033 , w15034 , w15035 , w15036 , w15037 , w15038 , w15039 , w15040 , w15041 , w15042 , w15043 , w15044 , w15045 , w15046 , w15047 , w15048 , w15049 , w15050 , w15051 , w15052 , w15053 , w15054 , w15055 , w15056 , w15057 , w15058 , w15059 , w15060 , w15061 , w15062 , w15063 , w15064 , w15065 , w15066 , w15067 , w15068 , w15069 , w15070 , w15071 , w15072 , w15073 , w15074 , w15075 , w15076 , w15077 , w15078 , w15079 , w15080 , w15081 , w15082 , w15083 , w15084 , w15085 , w15086 , w15087 , w15088 , w15089 , w15090 , w15091 , w15092 , w15093 , w15094 , w15095 , w15096 , w15097 , w15098 , w15099 , w15100 , w15101 , w15102 , w15103 , w15104 , w15105 , w15106 , w15107 , w15108 , w15109 , w15110 , w15111 , w15112 , w15113 , w15114 , w15115 , w15116 , w15117 , w15118 , w15119 , w15120 , w15121 , w15122 , w15123 , w15124 , w15125 , w15126 , w15127 , w15128 , w15129 , w15130 , w15131 , w15132 , w15133 , w15134 , w15135 , w15136 , w15137 , w15138 , w15139 , w15140 , w15141 , w15142 , w15143 , w15144 , w15145 , w15146 , w15147 , w15148 , w15149 , w15150 , w15151 , w15152 , w15153 , w15154 , w15155 , w15156 , w15157 , w15158 , w15159 , w15160 , w15161 , w15162 , w15163 , w15164 , w15165 , w15166 , w15167 , w15168 , w15169 , w15170 , w15171 , w15172 , w15173 , w15174 , w15175 , w15176 , w15177 , w15178 , w15179 , w15180 , w15181 , w15182 , w15183 , w15184 , w15185 , w15186 , w15187 , w15188 , w15189 , w15190 , w15191 , w15192 , w15193 , w15194 , w15195 , w15196 , w15197 , w15198 , w15199 , w15200 , w15201 , w15202 , w15203 , w15204 , w15205 , w15206 , w15207 , w15208 , w15209 , w15210 , w15211 , w15212 , w15213 , w15214 , w15215 , w15216 , w15217 , w15218 , w15219 , w15220 , w15221 , w15222 , w15223 , w15224 , w15225 , w15226 , w15227 , w15228 , w15229 , w15230 , w15231 , w15232 , w15233 , w15234 , w15235 , w15236 , w15237 , w15238 , w15239 , w15240 , w15241 , w15242 , w15243 , w15244 , w15245 , w15246 , w15247 , w15248 , w15249 , w15250 , w15251 , w15252 , w15253 , w15254 , w15255 , w15256 , w15257 , w15258 , w15259 , w15260 , w15261 , w15262 , w15263 , w15264 , w15265 , w15266 , w15267 , w15268 , w15269 , w15270 , w15271 , w15272 , w15273 , w15274 , w15275 , w15276 , w15277 , w15278 , w15279 , w15280 , w15281 , w15282 , w15283 , w15284 , w15285 , w15286 , w15287 , w15288 , w15289 , w15290 , w15291 , w15292 , w15293 , w15294 , w15295 , w15296 , w15297 , w15298 , w15299 , w15300 , w15301 , w15302 , w15303 , w15304 , w15305 , w15306 , w15307 , w15308 , w15309 , w15310 , w15311 , w15312 , w15313 , w15314 , w15315 , w15316 , w15317 , w15318 , w15319 , w15320 , w15321 , w15322 , w15323 , w15324 , w15325 , w15326 , w15327 , w15328 , w15329 , w15330 , w15331 , w15332 , w15333 , w15334 , w15335 , w15336 , w15337 , w15338 , w15339 , w15340 , w15341 , w15342 , w15343 , w15344 , w15345 , w15346 , w15347 , w15348 , w15349 , w15350 , w15351 , w15352 , w15353 , w15354 , w15355 , w15356 , w15357 , w15358 , w15359 , w15360 , w15361 , w15362 , w15363 , w15364 , w15365 , w15366 , w15367 , w15368 , w15369 , w15370 , w15371 , w15372 , w15373 , w15374 , w15375 , w15376 , w15377 , w15378 , w15379 , w15380 , w15381 , w15382 , w15383 , w15384 , w15385 , w15386 , w15387 , w15388 , w15389 , w15390 , w15391 , w15392 , w15393 , w15394 , w15395 , w15396 , w15397 , w15398 , w15399 , w15400 , w15401 , w15402 , w15403 , w15404 , w15405 , w15406 , w15407 , w15408 , w15409 , w15410 , w15411 , w15412 , w15413 , w15414 , w15415 , w15416 , w15417 , w15418 , w15419 , w15420 , w15421 , w15422 , w15423 , w15424 , w15425 , w15426 , w15427 , w15428 , w15429 , w15430 , w15431 , w15432 , w15433 , w15434 , w15435 , w15436 , w15437 , w15438 , w15439 , w15440 , w15441 , w15442 , w15443 , w15444 , w15445 , w15446 , w15447 , w15448 , w15449 , w15450 , w15451 , w15452 , w15453 , w15454 , w15455 , w15456 , w15457 , w15458 , w15459 , w15460 , w15461 , w15462 , w15463 , w15464 , w15465 , w15466 , w15467 , w15468 , w15469 , w15470 , w15471 , w15472 , w15473 , w15474 , w15475 , w15476 , w15477 , w15478 , w15479 , w15480 , w15481 , w15482 , w15483 , w15484 , w15485 , w15486 , w15487 , w15488 , w15489 , w15490 , w15491 , w15492 , w15493 , w15494 , w15495 , w15496 , w15497 , w15498 , w15499 , w15500 , w15501 , w15502 , w15503 , w15504 , w15505 , w15506 , w15507 , w15508 , w15509 , w15510 , w15511 , w15512 , w15513 , w15514 , w15515 , w15516 , w15517 , w15518 , w15519 , w15520 , w15521 , w15522 , w15523 , w15524 , w15525 , w15526 , w15527 , w15528 , w15529 , w15530 , w15531 , w15532 , w15533 , w15534 , w15535 , w15536 , w15537 , w15538 , w15539 , w15540 , w15541 , w15542 , w15543 , w15544 , w15545 , w15546 , w15547 , w15548 , w15549 , w15550 , w15551 , w15552 , w15553 , w15554 , w15555 , w15556 , w15557 , w15558 , w15559 , w15560 , w15561 , w15562 , w15563 , w15564 , w15565 , w15566 , w15567 , w15568 , w15569 , w15570 , w15571 , w15572 , w15573 , w15574 , w15575 , w15576 , w15577 , w15578 , w15579 , w15580 , w15581 , w15582 , w15583 , w15584 , w15585 , w15586 , w15587 , w15588 , w15589 , w15590 , w15591 , w15592 , w15593 , w15594 , w15595 , w15596 , w15597 , w15598 , w15599 , w15600 , w15601 , w15602 , w15603 , w15604 , w15605 , w15606 , w15607 , w15608 , w15609 , w15610 , w15611 , w15612 , w15613 , w15614 , w15615 , w15616 , w15617 , w15618 , w15619 , w15620 , w15621 , w15622 , w15623 , w15624 , w15625 , w15626 , w15627 , w15628 , w15629 , w15630 , w15631 , w15632 , w15633 , w15634 , w15635 , w15636 , w15637 , w15638 , w15639 , w15640 , w15641 , w15642 , w15643 , w15644 , w15645 , w15646 , w15647 , w15648 , w15649 , w15650 , w15651 , w15652 , w15653 , w15654 , w15655 , w15656 , w15657 , w15658 , w15659 , w15660 , w15661 , w15662 , w15663 , w15664 , w15665 , w15666 , w15667 , w15668 , w15669 , w15670 , w15671 , w15672 , w15673 , w15674 , w15675 , w15676 , w15677 , w15678 , w15679 , w15680 , w15681 , w15682 , w15683 , w15684 , w15685 , w15686 , w15687 , w15688 , w15689 , w15690 , w15691 , w15692 , w15693 , w15694 , w15695 , w15696 , w15697 , w15698 , w15699 , w15700 , w15701 , w15702 , w15703 , w15704 , w15705 , w15706 , w15707 , w15708 , w15709 , w15710 , w15711 , w15712 , w15713 , w15714 , w15715 , w15716 , w15717 , w15718 , w15719 , w15720 , w15721 , w15722 , w15723 , w15724 , w15725 , w15726 , w15727 , w15728 , w15729 , w15730 , w15731 , w15732 , w15733 , w15734 , w15735 , w15736 , w15737 , w15738 , w15739 , w15740 , w15741 , w15742 , w15743 , w15744 , w15745 , w15746 , w15747 , w15748 , w15749 , w15750 , w15751 , w15752 , w15753 , w15754 , w15755 , w15756 , w15757 , w15758 , w15759 , w15760 , w15761 , w15762 , w15763 , w15764 , w15765 , w15766 , w15767 , w15768 , w15769 , w15770 , w15771 , w15772 , w15773 , w15774 , w15775 , w15776 , w15777 , w15778 , w15779 , w15780 , w15781 , w15782 , w15783 , w15784 , w15785 , w15786 , w15787 , w15788 , w15789 , w15790 , w15791 , w15792 , w15793 , w15794 , w15795 , w15796 , w15797 , w15798 , w15799 , w15800 , w15801 , w15802 , w15803 , w15804 , w15805 , w15806 , w15807 , w15808 , w15809 , w15810 , w15811 , w15812 , w15813 , w15814 , w15815 , w15816 , w15817 , w15818 , w15819 , w15820 , w15821 , w15822 , w15823 , w15824 , w15825 , w15826 , w15827 , w15828 , w15829 , w15830 , w15831 , w15832 , w15833 , w15834 , w15835 , w15836 , w15837 , w15838 , w15839 , w15840 , w15841 , w15842 , w15843 , w15844 , w15845 , w15846 , w15847 , w15848 , w15849 , w15850 , w15851 , w15852 , w15853 , w15854 , w15855 , w15856 , w15857 , w15858 , w15859 , w15860 , w15861 , w15862 , w15863 , w15864 , w15865 , w15866 , w15867 , w15868 , w15869 , w15870 , w15871 , w15872 , w15873 , w15874 , w15875 , w15876 , w15877 , w15878 , w15879 , w15880 , w15881 , w15882 , w15883 , w15884 , w15885 , w15886 , w15887 , w15888 , w15889 , w15890 , w15891 , w15892 , w15893 , w15894 , w15895 , w15896 , w15897 , w15898 , w15899 , w15900 , w15901 , w15902 , w15903 , w15904 , w15905 , w15906 , w15907 , w15908 , w15909 , w15910 , w15911 , w15912 , w15913 , w15914 , w15915 , w15916 , w15917 , w15918 , w15919 , w15920 , w15921 , w15922 , w15923 , w15924 , w15925 , w15926 , w15927 , w15928 , w15929 , w15930 , w15931 , w15932 , w15933 , w15934 , w15935 , w15936 , w15937 , w15938 , w15939 , w15940 , w15941 , w15942 , w15943 , w15944 , w15945 , w15946 , w15947 , w15948 , w15949 , w15950 , w15951 , w15952 , w15953 , w15954 , w15955 , w15956 , w15957 , w15958 , w15959 , w15960 , w15961 , w15962 , w15963 , w15964 , w15965 , w15966 , w15967 , w15968 , w15969 , w15970 , w15971 , w15972 , w15973 , w15974 , w15975 , w15976 , w15977 , w15978 , w15979 , w15980 , w15981 , w15982 , w15983 , w15984 , w15985 , w15986 , w15987 , w15988 , w15989 , w15990 , w15991 , w15992 , w15993 , w15994 , w15995 , w15996 , w15997 , w15998 , w15999 , w16000 , w16001 , w16002 , w16003 , w16004 , w16005 , w16006 , w16007 , w16008 , w16009 , w16010 , w16011 , w16012 , w16013 , w16014 , w16015 , w16016 , w16017 , w16018 , w16019 , w16020 , w16021 , w16022 , w16023 , w16024 , w16025 , w16026 , w16027 , w16028 , w16029 , w16030 , w16031 , w16032 , w16033 , w16034 , w16035 , w16036 , w16037 , w16038 , w16039 , w16040 , w16041 , w16042 , w16043 , w16044 , w16045 , w16046 , w16047 , w16048 , w16049 , w16050 , w16051 , w16052 , w16053 , w16054 , w16055 , w16056 , w16057 , w16058 , w16059 , w16060 , w16061 , w16062 , w16063 , w16064 , w16065 , w16066 , w16067 , w16068 , w16069 , w16070 , w16071 , w16072 , w16073 , w16074 , w16075 , w16076 , w16077 , w16078 , w16079 , w16080 , w16081 , w16082 , w16083 , w16084 , w16085 , w16086 , w16087 , w16088 , w16089 , w16090 , w16091 , w16092 , w16093 , w16094 , w16095 , w16096 , w16097 , w16098 , w16099 , w16100 , w16101 , w16102 , w16103 , w16104 , w16105 , w16106 , w16107 , w16108 , w16109 , w16110 , w16111 , w16112 , w16113 , w16114 , w16115 , w16116 , w16117 , w16118 , w16119 , w16120 , w16121 , w16122 , w16123 , w16124 , w16125 , w16126 , w16127 , w16128 , w16129 , w16130 , w16131 , w16132 , w16133 , w16134 , w16135 , w16136 , w16137 , w16138 , w16139 , w16140 , w16141 , w16142 , w16143 , w16144 , w16145 , w16146 , w16147 , w16148 , w16149 , w16150 , w16151 , w16152 , w16153 , w16154 , w16155 , w16156 , w16157 , w16158 , w16159 , w16160 , w16161 , w16162 , w16163 , w16164 , w16165 , w16166 , w16167 , w16168 , w16169 , w16170 , w16171 , w16172 , w16173 , w16174 , w16175 , w16176 , w16177 , w16178 , w16179 , w16180 , w16181 , w16182 , w16183 , w16184 , w16185 , w16186 , w16187 , w16188 , w16189 , w16190 , w16191 , w16192 , w16193 , w16194 , w16195 , w16196 , w16197 , w16198 , w16199 , w16200 , w16201 , w16202 , w16203 , w16204 , w16205 , w16206 , w16207 , w16208 , w16209 , w16210 , w16211 , w16212 , w16213 , w16214 , w16215 , w16216 , w16217 , w16218 , w16219 , w16220 , w16221 , w16222 , w16223 , w16224 , w16225 , w16226 , w16227 , w16228 , w16229 , w16230 , w16231 , w16232 , w16233 , w16234 , w16235 , w16236 , w16237 , w16238 , w16239 , w16240 , w16241 , w16242 , w16243 , w16244 , w16245 , w16246 , w16247 , w16248 , w16249 , w16250 , w16251 , w16252 , w16253 , w16254 , w16255 , w16256 , w16257 , w16258 , w16259 , w16260 , w16261 , w16262 , w16263 , w16264 , w16265 , w16266 , w16267 , w16268 , w16269 , w16270 , w16271 , w16272 , w16273 , w16274 , w16275 , w16276 , w16277 , w16278 , w16279 , w16280 , w16281 , w16282 , w16283 , w16284 , w16285 , w16286 , w16287 , w16288 , w16289 , w16290 , w16291 , w16292 , w16293 , w16294 , w16295 , w16296 , w16297 , w16298 , w16299 , w16300 , w16301 , w16302 , w16303 , w16304 , w16305 , w16306 , w16307 , w16308 , w16309 , w16310 , w16311 , w16312 , w16313 , w16314 , w16315 , w16316 , w16317 , w16318 , w16319 , w16320 , w16321 , w16322 , w16323 , w16324 , w16325 , w16326 , w16327 , w16328 , w16329 , w16330 , w16331 , w16332 , w16333 , w16334 , w16335 , w16336 , w16337 , w16338 , w16339 , w16340 , w16341 , w16342 , w16343 , w16344 , w16345 , w16346 , w16347 , w16348 , w16349 , w16350 , w16351 , w16352 , w16353 , w16354 , w16355 , w16356 , w16357 , w16358 , w16359 , w16360 , w16361 , w16362 , w16363 , w16364 , w16365 , w16366 , w16367 , w16368 , w16369 , w16370 , w16371 , w16372 , w16373 , w16374 , w16375 , w16376 , w16377 , w16378 , w16379 , w16380 , w16381 , w16382 , w16383 , w16384 , w16385 , w16386 , w16387 , w16388 , w16389 , w16390 , w16391 , w16392 , w16393 , w16394 , w16395 , w16396 , w16397 , w16398 , w16399 , w16400 , w16401 , w16402 , w16403 , w16404 , w16405 , w16406 , w16407 , w16408 , w16409 , w16410 , w16411 , w16412 , w16413 , w16414 , w16415 , w16416 , w16417 , w16418 , w16419 , w16420 , w16421 , w16422 , w16423 , w16424 , w16425 , w16426 , w16427 , w16428 , w16429 , w16430 , w16431 , w16432 , w16433 , w16434 , w16435 , w16436 , w16437 , w16438 , w16439 , w16440 , w16441 , w16442 , w16443 , w16444 , w16445 , w16446 , w16447 , w16448 , w16449 , w16450 , w16451 , w16452 , w16453 , w16454 , w16455 , w16456 , w16457 , w16458 , w16459 , w16460 , w16461 , w16462 , w16463 , w16464 , w16465 , w16466 , w16467 , w16468 , w16469 , w16470 , w16471 , w16472 , w16473 , w16474 , w16475 , w16476 , w16477 , w16478 , w16479 , w16480 , w16481 , w16482 , w16483 , w16484 , w16485 , w16486 , w16487 , w16488 , w16489 , w16490 , w16491 , w16492 , w16493 , w16494 , w16495 , w16496 , w16497 , w16498 , w16499 , w16500 , w16501 , w16502 , w16503 , w16504 , w16505 , w16506 , w16507 , w16508 , w16509 , w16510 , w16511 , w16512 , w16513 , w16514 , w16515 , w16516 , w16517 , w16518 , w16519 , w16520 , w16521 , w16522 , w16523 , w16524 , w16525 , w16526 , w16527 , w16528 , w16529 , w16530 , w16531 , w16532 , w16533 , w16534 , w16535 , w16536 , w16537 , w16538 , w16539 , w16540 , w16541 , w16542 , w16543 , w16544 , w16545 , w16546 , w16547 , w16548 , w16549 , w16550 , w16551 , w16552 , w16553 , w16554 , w16555 , w16556 , w16557 , w16558 , w16559 , w16560 , w16561 , w16562 , w16563 , w16564 , w16565 , w16566 , w16567 , w16568 , w16569 , w16570 , w16571 , w16572 , w16573 , w16574 , w16575 , w16576 , w16577 , w16578 , w16579 , w16580 , w16581 , w16582 , w16583 , w16584 , w16585 , w16586 , w16587 , w16588 , w16589 , w16590 , w16591 , w16592 , w16593 , w16594 , w16595 , w16596 , w16597 , w16598 , w16599 , w16600 , w16601 , w16602 , w16603 , w16604 , w16605 , w16606 , w16607 , w16608 , w16609 , w16610 , w16611 , w16612 , w16613 , w16614 , w16615 , w16616 , w16617 , w16618 , w16619 , w16620 , w16621 , w16622 , w16623 , w16624 , w16625 , w16626 , w16627 , w16628 , w16629 , w16630 , w16631 , w16632 , w16633 , w16634 , w16635 , w16636 , w16637 , w16638 , w16639 , w16640 , w16641 , w16642 , w16643 , w16644 , w16645 , w16646 , w16647 , w16648 , w16649 , w16650 , w16651 , w16652 , w16653 , w16654 , w16655 , w16656 , w16657 , w16658 , w16659 , w16660 , w16661 , w16662 , w16663 , w16664 , w16665 , w16666 , w16667 , w16668 , w16669 , w16670 , w16671 , w16672 , w16673 , w16674 , w16675 , w16676 , w16677 , w16678 , w16679 , w16680 , w16681 , w16682 , w16683 , w16684 , w16685 , w16686 , w16687 , w16688 , w16689 , w16690 , w16691 , w16692 , w16693 , w16694 , w16695 , w16696 , w16697 , w16698 , w16699 , w16700 , w16701 , w16702 , w16703 , w16704 , w16705 , w16706 , w16707 , w16708 , w16709 , w16710 , w16711 , w16712 , w16713 , w16714 , w16715 , w16716 , w16717 , w16718 , w16719 , w16720 , w16721 , w16722 , w16723 , w16724 , w16725 , w16726 , w16727 , w16728 , w16729 , w16730 , w16731 , w16732 , w16733 , w16734 , w16735 , w16736 , w16737 , w16738 , w16739 , w16740 , w16741 , w16742 , w16743 , w16744 , w16745 , w16746 , w16747 , w16748 , w16749 , w16750 , w16751 , w16752 , w16753 , w16754 , w16755 , w16756 , w16757 , w16758 , w16759 , w16760 , w16761 , w16762 , w16763 , w16764 , w16765 , w16766 , w16767 , w16768 , w16769 , w16770 , w16771 , w16772 , w16773 , w16774 , w16775 , w16776 , w16777 , w16778 , w16779 , w16780 , w16781 , w16782 , w16783 , w16784 , w16785 , w16786 , w16787 , w16788 , w16789 , w16790 , w16791 , w16792 , w16793 , w16794 , w16795 , w16796 , w16797 , w16798 , w16799 , w16800 , w16801 , w16802 , w16803 , w16804 , w16805 , w16806 , w16807 , w16808 , w16809 , w16810 , w16811 , w16812 , w16813 , w16814 , w16815 , w16816 , w16817 , w16818 , w16819 , w16820 , w16821 , w16822 , w16823 , w16824 , w16825 , w16826 , w16827 , w16828 , w16829 , w16830 , w16831 , w16832 , w16833 , w16834 , w16835 , w16836 , w16837 , w16838 , w16839 , w16840 , w16841 , w16842 , w16843 , w16844 , w16845 , w16846 , w16847 , w16848 , w16849 , w16850 , w16851 , w16852 , w16853 , w16854 , w16855 , w16856 , w16857 , w16858 , w16859 , w16860 , w16861 , w16862 , w16863 , w16864 , w16865 , w16866 , w16867 , w16868 , w16869 , w16870 , w16871 , w16872 , w16873 , w16874 , w16875 , w16876 , w16877 , w16878 , w16879 , w16880 , w16881 , w16882 , w16883 , w16884 , w16885 , w16886 , w16887 , w16888 , w16889 , w16890 , w16891 , w16892 , w16893 , w16894 , w16895 , w16896 , w16897 , w16898 , w16899 , w16900 , w16901 , w16902 , w16903 , w16904 , w16905 , w16906 , w16907 , w16908 , w16909 , w16910 , w16911 , w16912 , w16913 , w16914 , w16915 , w16916 , w16917 , w16918 , w16919 , w16920 , w16921 , w16922 , w16923 , w16924 , w16925 , w16926 , w16927 , w16928 , w16929 , w16930 , w16931 , w16932 , w16933 , w16934 , w16935 , w16936 , w16937 , w16938 , w16939 , w16940 , w16941 , w16942 , w16943 , w16944 , w16945 , w16946 , w16947 , w16948 , w16949 , w16950 , w16951 , w16952 , w16953 , w16954 , w16955 , w16956 , w16957 , w16958 , w16959 , w16960 , w16961 , w16962 , w16963 , w16964 , w16965 , w16966 , w16967 , w16968 , w16969 , w16970 , w16971 , w16972 , w16973 , w16974 , w16975 , w16976 , w16977 , w16978 , w16979 , w16980 , w16981 , w16982 , w16983 , w16984 , w16985 , w16986 , w16987 , w16988 , w16989 , w16990 , w16991 , w16992 , w16993 , w16994 , w16995 , w16996 , w16997 , w16998 , w16999 , w17000 , w17001 , w17002 , w17003 , w17004 , w17005 , w17006 , w17007 , w17008 , w17009 , w17010 , w17011 , w17012 , w17013 , w17014 , w17015 , w17016 , w17017 , w17018 , w17019 , w17020 , w17021 , w17022 , w17023 , w17024 , w17025 , w17026 , w17027 , w17028 , w17029 , w17030 , w17031 , w17032 , w17033 , w17034 , w17035 , w17036 , w17037 , w17038 , w17039 , w17040 , w17041 , w17042 , w17043 , w17044 , w17045 , w17046 , w17047 , w17048 , w17049 , w17050 , w17051 , w17052 , w17053 , w17054 , w17055 , w17056 , w17057 , w17058 , w17059 , w17060 , w17061 , w17062 , w17063 , w17064 , w17065 , w17066 , w17067 , w17068 , w17069 , w17070 , w17071 , w17072 , w17073 , w17074 , w17075 , w17076 , w17077 , w17078 , w17079 , w17080 , w17081 , w17082 , w17083 , w17084 , w17085 , w17086 , w17087 , w17088 , w17089 , w17090 , w17091 , w17092 , w17093 , w17094 , w17095 , w17096 , w17097 , w17098 , w17099 , w17100 , w17101 , w17102 , w17103 , w17104 , w17105 , w17106 , w17107 , w17108 , w17109 , w17110 , w17111 , w17112 , w17113 , w17114 , w17115 , w17116 , w17117 , w17118 , w17119 , w17120 , w17121 , w17122 , w17123 , w17124 , w17125 , w17126 , w17127 , w17128 , w17129 , w17130 , w17131 , w17132 , w17133 , w17134 , w17135 , w17136 , w17137 , w17138 , w17139 , w17140 , w17141 , w17142 , w17143 , w17144 , w17145 , w17146 , w17147 , w17148 , w17149 , w17150 , w17151 , w17152 , w17153 , w17154 , w17155 , w17156 , w17157 , w17158 , w17159 , w17160 , w17161 , w17162 , w17163 , w17164 , w17165 , w17166 , w17167 , w17168 , w17169 , w17170 , w17171 , w17172 , w17173 , w17174 , w17175 , w17176 , w17177 , w17178 , w17179 , w17180 , w17181 , w17182 , w17183 , w17184 , w17185 , w17186 , w17187 , w17188 , w17189 , w17190 , w17191 , w17192 , w17193 , w17194 , w17195 , w17196 , w17197 , w17198 , w17199 , w17200 , w17201 , w17202 , w17203 , w17204 , w17205 , w17206 , w17207 , w17208 , w17209 , w17210 , w17211 , w17212 , w17213 , w17214 , w17215 , w17216 , w17217 , w17218 , w17219 , w17220 , w17221 , w17222 , w17223 , w17224 , w17225 , w17226 , w17227 , w17228 , w17229 , w17230 , w17231 , w17232 , w17233 , w17234 , w17235 , w17236 , w17237 , w17238 , w17239 , w17240 , w17241 , w17242 , w17243 , w17244 , w17245 , w17246 , w17247 , w17248 , w17249 , w17250 , w17251 , w17252 , w17253 , w17254 , w17255 , w17256 , w17257 , w17258 , w17259 , w17260 , w17261 , w17262 , w17263 , w17264 , w17265 , w17266 , w17267 , w17268 , w17269 , w17270 , w17271 , w17272 , w17273 , w17274 , w17275 , w17276 , w17277 , w17278 , w17279 , w17280 , w17281 , w17282 , w17283 , w17284 , w17285 , w17286 , w17287 , w17288 , w17289 , w17290 , w17291 , w17292 , w17293 , w17294 , w17295 , w17296 , w17297 , w17298 , w17299 , w17300 , w17301 , w17302 , w17303 , w17304 , w17305 , w17306 , w17307 , w17308 , w17309 , w17310 , w17311 , w17312 , w17313 , w17314 , w17315 , w17316 , w17317 , w17318 , w17319 , w17320 , w17321 , w17322 , w17323 , w17324 , w17325 , w17326 , w17327 , w17328 , w17329 , w17330 , w17331 , w17332 , w17333 , w17334 , w17335 , w17336 , w17337 , w17338 , w17339 , w17340 , w17341 , w17342 , w17343 , w17344 , w17345 , w17346 , w17347 , w17348 , w17349 , w17350 , w17351 , w17352 , w17353 , w17354 , w17355 , w17356 , w17357 , w17358 , w17359 , w17360 , w17361 , w17362 , w17363 , w17364 , w17365 , w17366 , w17367 , w17368 , w17369 , w17370 , w17371 , w17372 , w17373 , w17374 , w17375 , w17376 , w17377 , w17378 , w17379 , w17380 , w17381 , w17382 , w17383 , w17384 , w17385 , w17386 , w17387 , w17388 , w17389 , w17390 , w17391 , w17392 , w17393 , w17394 , w17395 , w17396 , w17397 , w17398 , w17399 , w17400 , w17401 , w17402 , w17403 , w17404 , w17405 , w17406 , w17407 , w17408 , w17409 , w17410 , w17411 , w17412 , w17413 , w17414 , w17415 , w17416 , w17417 , w17418 , w17419 , w17420 , w17421 , w17422 , w17423 , w17424 , w17425 , w17426 , w17427 , w17428 , w17429 , w17430 , w17431 , w17432 , w17433 , w17434 , w17435 , w17436 , w17437 , w17438 , w17439 , w17440 , w17441 , w17442 , w17443 , w17444 , w17445 , w17446 , w17447 , w17448 , w17449 , w17450 , w17451 , w17452 , w17453 , w17454 , w17455 , w17456 , w17457 , w17458 , w17459 , w17460 , w17461 , w17462 , w17463 , w17464 , w17465 , w17466 , w17467 , w17468 , w17469 , w17470 , w17471 , w17472 , w17473 , w17474 , w17475 , w17476 , w17477 , w17478 , w17479 , w17480 , w17481 , w17482 , w17483 , w17484 , w17485 , w17486 , w17487 , w17488 , w17489 , w17490 , w17491 , w17492 , w17493 , w17494 , w17495 , w17496 , w17497 , w17498 , w17499 , w17500 , w17501 , w17502 , w17503 , w17504 , w17505 , w17506 , w17507 , w17508 , w17509 , w17510 , w17511 , w17512 , w17513 , w17514 , w17515 , w17516 , w17517 , w17518 , w17519 , w17520 , w17521 , w17522 , w17523 , w17524 , w17525 , w17526 , w17527 , w17528 , w17529 , w17530 , w17531 , w17532 , w17533 , w17534 , w17535 , w17536 , w17537 , w17538 , w17539 , w17540 , w17541 , w17542 , w17543 , w17544 , w17545 , w17546 , w17547 , w17548 , w17549 , w17550 , w17551 , w17552 , w17553 , w17554 , w17555 , w17556 , w17557 , w17558 , w17559 , w17560 , w17561 , w17562 , w17563 , w17564 , w17565 , w17566 , w17567 , w17568 , w17569 , w17570 , w17571 , w17572 , w17573 , w17574 , w17575 , w17576 , w17577 , w17578 , w17579 , w17580 , w17581 , w17582 , w17583 , w17584 , w17585 , w17586 , w17587 , w17588 , w17589 , w17590 , w17591 , w17592 , w17593 , w17594 , w17595 , w17596 , w17597 , w17598 , w17599 , w17600 , w17601 , w17602 , w17603 , w17604 , w17605 , w17606 , w17607 , w17608 , w17609 , w17610 , w17611 , w17612 , w17613 , w17614 , w17615 , w17616 , w17617 , w17618 , w17619 , w17620 , w17621 , w17622 , w17623 , w17624 , w17625 , w17626 , w17627 , w17628 , w17629 , w17630 , w17631 , w17632 , w17633 , w17634 , w17635 , w17636 , w17637 , w17638 , w17639 , w17640 , w17641 , w17642 , w17643 , w17644 , w17645 , w17646 , w17647 , w17648 , w17649 , w17650 , w17651 , w17652 , w17653 , w17654 , w17655 , w17656 , w17657 , w17658 , w17659 , w17660 , w17661 , w17662 , w17663 , w17664 , w17665 , w17666 , w17667 , w17668 , w17669 , w17670 , w17671 , w17672 , w17673 , w17674 , w17675 , w17676 , w17677 , w17678 , w17679 , w17680 , w17681 , w17682 , w17683 , w17684 , w17685 , w17686 , w17687 , w17688 , w17689 , w17690 , w17691 , w17692 , w17693 , w17694 , w17695 , w17696 , w17697 , w17698 , w17699 , w17700 , w17701 , w17702 , w17703 , w17704 , w17705 , w17706 , w17707 , w17708 , w17709 , w17710 , w17711 , w17712 , w17713 , w17714 , w17715 , w17716 , w17717 , w17718 , w17719 , w17720 , w17721 , w17722 , w17723 , w17724 , w17725 , w17726 , w17727 , w17728 , w17729 , w17730 , w17731 , w17732 , w17733 , w17734 , w17735 , w17736 , w17737 , w17738 , w17739 , w17740 , w17741 , w17742 , w17743 , w17744 , w17745 , w17746 , w17747 , w17748 , w17749 , w17750 , w17751 , w17752 , w17753 , w17754 , w17755 , w17756 , w17757 , w17758 , w17759 , w17760 , w17761 , w17762 , w17763 , w17764 , w17765 , w17766 , w17767 , w17768 , w17769 , w17770 , w17771 , w17772 , w17773 , w17774 , w17775 , w17776 , w17777 , w17778 , w17779 , w17780 , w17781 , w17782 , w17783 , w17784 , w17785 , w17786 , w17787 , w17788 , w17789 , w17790 , w17791 , w17792 , w17793 , w17794 , w17795 , w17796 , w17797 , w17798 , w17799 , w17800 , w17801 , w17802 , w17803 , w17804 , w17805 , w17806 , w17807 , w17808 , w17809 , w17810 , w17811 , w17812 , w17813 , w17814 , w17815 , w17816 , w17817 , w17818 , w17819 , w17820 , w17821 , w17822 , w17823 , w17824 , w17825 , w17826 , w17827 , w17828 , w17829 , w17830 , w17831 , w17832 , w17833 , w17834 , w17835 , w17836 , w17837 , w17838 , w17839 , w17840 , w17841 , w17842 , w17843 , w17844 , w17845 , w17846 , w17847 , w17848 , w17849 , w17850 , w17851 , w17852 , w17853 , w17854 , w17855 , w17856 , w17857 , w17858 , w17859 , w17860 , w17861 , w17862 , w17863 , w17864 , w17865 , w17866 , w17867 , w17868 , w17869 , w17870 , w17871 , w17872 , w17873 , w17874 , w17875 , w17876 , w17877 , w17878 , w17879 , w17880 , w17881 , w17882 , w17883 , w17884 , w17885 , w17886 , w17887 , w17888 , w17889 , w17890 , w17891 , w17892 , w17893 , w17894 , w17895 , w17896 , w17897 , w17898 , w17899 , w17900 , w17901 , w17902 , w17903 , w17904 , w17905 , w17906 , w17907 , w17908 , w17909 , w17910 , w17911 , w17912 , w17913 , w17914 , w17915 , w17916 , w17917 , w17918 , w17919 , w17920 , w17921 , w17922 , w17923 , w17924 , w17925 , w17926 , w17927 , w17928 , w17929 , w17930 , w17931 , w17932 , w17933 , w17934 , w17935 , w17936 , w17937 , w17938 , w17939 , w17940 , w17941 , w17942 , w17943 , w17944 , w17945 , w17946 , w17947 , w17948 , w17949 , w17950 , w17951 , w17952 , w17953 , w17954 , w17955 , w17956 , w17957 , w17958 , w17959 , w17960 , w17961 , w17962 , w17963 , w17964 , w17965 , w17966 , w17967 , w17968 , w17969 , w17970 , w17971 , w17972 , w17973 , w17974 , w17975 , w17976 , w17977 , w17978 , w17979 , w17980 , w17981 , w17982 , w17983 , w17984 , w17985 , w17986 , w17987 , w17988 , w17989 , w17990 , w17991 , w17992 , w17993 , w17994 , w17995 , w17996 , w17997 , w17998 , w17999 , w18000 , w18001 , w18002 , w18003 , w18004 , w18005 , w18006 , w18007 , w18008 , w18009 , w18010 , w18011 , w18012 , w18013 , w18014 , w18015 , w18016 , w18017 , w18018 , w18019 , w18020 , w18021 , w18022 , w18023 , w18024 , w18025 , w18026 , w18027 , w18028 , w18029 , w18030 , w18031 , w18032 , w18033 , w18034 , w18035 , w18036 , w18037 , w18038 , w18039 , w18040 , w18041 , w18042 , w18043 , w18044 , w18045 , w18046 , w18047 , w18048 , w18049 , w18050 , w18051 , w18052 , w18053 , w18054 , w18055 , w18056 , w18057 , w18058 , w18059 , w18060 , w18061 , w18062 , w18063 , w18064 , w18065 , w18066 , w18067 , w18068 , w18069 , w18070 , w18071 , w18072 , w18073 , w18074 , w18075 , w18076 , w18077 , w18078 , w18079 , w18080 , w18081 , w18082 , w18083 , w18084 , w18085 , w18086 , w18087 , w18088 , w18089 , w18090 , w18091 , w18092 , w18093 , w18094 , w18095 , w18096 , w18097 , w18098 , w18099 , w18100 , w18101 , w18102 , w18103 , w18104 , w18105 , w18106 , w18107 , w18108 , w18109 , w18110 , w18111 , w18112 , w18113 , w18114 , w18115 , w18116 , w18117 , w18118 , w18119 , w18120 , w18121 , w18122 , w18123 , w18124 , w18125 , w18126 , w18127 , w18128 , w18129 , w18130 , w18131 , w18132 , w18133 , w18134 , w18135 , w18136 , w18137 , w18138 , w18139 , w18140 , w18141 , w18142 , w18143 , w18144 , w18145 , w18146 , w18147 , w18148 , w18149 , w18150 , w18151 , w18152 , w18153 , w18154 , w18155 , w18156 , w18157 , w18158 , w18159 , w18160 , w18161 , w18162 , w18163 , w18164 , w18165 , w18166 , w18167 , w18168 , w18169 , w18170 , w18171 , w18172 , w18173 , w18174 , w18175 , w18176 , w18177 , w18178 , w18179 , w18180 , w18181 , w18182 , w18183 , w18184 , w18185 , w18186 , w18187 , w18188 , w18189 , w18190 , w18191 , w18192 , w18193 , w18194 , w18195 , w18196 , w18197 , w18198 , w18199 , w18200 , w18201 , w18202 , w18203 , w18204 , w18205 , w18206 , w18207 , w18208 , w18209 , w18210 , w18211 , w18212 , w18213 , w18214 , w18215 , w18216 , w18217 , w18218 , w18219 , w18220 , w18221 , w18222 , w18223 , w18224 , w18225 , w18226 , w18227 , w18228 , w18229 , w18230 , w18231 , w18232 , w18233 , w18234 , w18235 , w18236 , w18237 , w18238 , w18239 , w18240 , w18241 , w18242 , w18243 , w18244 , w18245 , w18246 , w18247 , w18248 , w18249 , w18250 , w18251 , w18252 , w18253 , w18254 , w18255 , w18256 , w18257 , w18258 , w18259 , w18260 , w18261 , w18262 , w18263 , w18264 , w18265 , w18266 , w18267 , w18268 , w18269 , w18270 , w18271 , w18272 , w18273 , w18274 , w18275 , w18276 , w18277 , w18278 , w18279 , w18280 , w18281 , w18282 , w18283 , w18284 , w18285 , w18286 , w18287 , w18288 , w18289 , w18290 , w18291 , w18292 , w18293 , w18294 , w18295 , w18296 , w18297 , w18298 , w18299 , w18300 , w18301 , w18302 , w18303 , w18304 , w18305 , w18306 , w18307 , w18308 , w18309 , w18310 , w18311 , w18312 , w18313 , w18314 , w18315 , w18316 , w18317 , w18318 , w18319 , w18320 , w18321 , w18322 , w18323 , w18324 , w18325 , w18326 , w18327 , w18328 , w18329 , w18330 , w18331 , w18332 , w18333 , w18334 , w18335 , w18336 , w18337 , w18338 , w18339 , w18340 , w18341 , w18342 , w18343 , w18344 , w18345 , w18346 , w18347 , w18348 , w18349 , w18350 , w18351 , w18352 , w18353 , w18354 , w18355 , w18356 , w18357 , w18358 , w18359 , w18360 , w18361 , w18362 , w18363 , w18364 , w18365 , w18366 , w18367 , w18368 , w18369 , w18370 , w18371 , w18372 , w18373 , w18374 , w18375 , w18376 , w18377 , w18378 , w18379 , w18380 , w18381 , w18382 , w18383 , w18384 , w18385 , w18386 , w18387 , w18388 , w18389 , w18390 , w18391 , w18392 , w18393 , w18394 , w18395 , w18396 , w18397 , w18398 , w18399 , w18400 , w18401 , w18402 , w18403 , w18404 , w18405 , w18406 , w18407 , w18408 , w18409 , w18410 , w18411 , w18412 , w18413 , w18414 , w18415 , w18416 , w18417 , w18418 , w18419 , w18420 , w18421 , w18422 , w18423 , w18424 , w18425 , w18426 , w18427 , w18428 , w18429 , w18430 , w18431 , w18432 , w18433 , w18434 , w18435 , w18436 , w18437 , w18438 , w18439 , w18440 , w18441 , w18442 , w18443 , w18444 , w18445 , w18446 , w18447 , w18448 , w18449 , w18450 , w18451 , w18452 , w18453 , w18454 , w18455 , w18456 , w18457 , w18458 , w18459 , w18460 , w18461 , w18462 , w18463 , w18464 , w18465 , w18466 , w18467 , w18468 , w18469 , w18470 , w18471 , w18472 , w18473 , w18474 , w18475 , w18476 , w18477 , w18478 , w18479 , w18480 , w18481 , w18482 , w18483 , w18484 , w18485 , w18486 , w18487 , w18488 , w18489 , w18490 , w18491 , w18492 , w18493 , w18494 , w18495 , w18496 , w18497 , w18498 , w18499 , w18500 , w18501 , w18502 , w18503 , w18504 , w18505 , w18506 , w18507 , w18508 , w18509 , w18510 , w18511 , w18512 , w18513 , w18514 , w18515 , w18516 , w18517 , w18518 , w18519 , w18520 , w18521 , w18522 , w18523 , w18524 , w18525 , w18526 , w18527 , w18528 , w18529 , w18530 , w18531 , w18532 , w18533 , w18534 , w18535 , w18536 , w18537 , w18538 , w18539 , w18540 , w18541 , w18542 , w18543 , w18544 , w18545 , w18546 , w18547 , w18548 , w18549 , w18550 , w18551 , w18552 , w18553 , w18554 , w18555 , w18556 , w18557 , w18558 , w18559 , w18560 , w18561 , w18562 , w18563 , w18564 , w18565 , w18566 , w18567 , w18568 , w18569 , w18570 , w18571 , w18572 , w18573 , w18574 , w18575 , w18576 , w18577 , w18578 , w18579 , w18580 , w18581 , w18582 , w18583 , w18584 , w18585 , w18586 , w18587 , w18588 , w18589 , w18590 , w18591 , w18592 , w18593 , w18594 , w18595 , w18596 , w18597 , w18598 , w18599 , w18600 , w18601 , w18602 , w18603 , w18604 , w18605 , w18606 , w18607 , w18608 , w18609 , w18610 , w18611 , w18612 , w18613 , w18614 , w18615 , w18616 , w18617 , w18618 , w18619 , w18620 , w18621 , w18622 , w18623 , w18624 , w18625 , w18626 , w18627 , w18628 , w18629 , w18630 , w18631 , w18632 , w18633 , w18634 , w18635 , w18636 , w18637 , w18638 , w18639 , w18640 , w18641 , w18642 , w18643 , w18644 , w18645 , w18646 , w18647 , w18648 , w18649 , w18650 , w18651 , w18652 , w18653 , w18654 , w18655 , w18656 , w18657 , w18658 , w18659 , w18660 , w18661 , w18662 , w18663 , w18664 , w18665 , w18666 , w18667 , w18668 , w18669 , w18670 , w18671 , w18672 , w18673 , w18674 , w18675 , w18676 , w18677 , w18678 , w18679 , w18680 , w18681 , w18682 , w18683 , w18684 , w18685 , w18686 , w18687 , w18688 , w18689 , w18690 , w18691 , w18692 , w18693 , w18694 , w18695 , w18696 , w18697 , w18698 , w18699 , w18700 , w18701 , w18702 , w18703 , w18704 , w18705 , w18706 , w18707 , w18708 , w18709 , w18710 , w18711 , w18712 , w18713 , w18714 , w18715 , w18716 , w18717 , w18718 , w18719 , w18720 , w18721 , w18722 , w18723 , w18724 , w18725 , w18726 , w18727 , w18728 , w18729 , w18730 , w18731 , w18732 , w18733 , w18734 , w18735 , w18736 , w18737 , w18738 , w18739 , w18740 , w18741 , w18742 , w18743 , w18744 , w18745 , w18746 , w18747 , w18748 , w18749 , w18750 , w18751 , w18752 , w18753 , w18754 , w18755 , w18756 , w18757 , w18758 , w18759 , w18760 , w18761 , w18762 , w18763 , w18764 , w18765 , w18766 , w18767 , w18768 , w18769 , w18770 , w18771 , w18772 , w18773 , w18774 , w18775 , w18776 , w18777 , w18778 , w18779 , w18780 , w18781 , w18782 , w18783 , w18784 , w18785 , w18786 , w18787 , w18788 , w18789 , w18790 , w18791 , w18792 , w18793 , w18794 , w18795 , w18796 , w18797 , w18798 , w18799 , w18800 , w18801 , w18802 , w18803 , w18804 , w18805 , w18806 , w18807 , w18808 , w18809 , w18810 , w18811 , w18812 , w18813 , w18814 , w18815 , w18816 , w18817 , w18818 , w18819 , w18820 , w18821 , w18822 , w18823 , w18824 , w18825 , w18826 , w18827 , w18828 , w18829 , w18830 , w18831 , w18832 , w18833 , w18834 , w18835 , w18836 , w18837 , w18838 , w18839 , w18840 , w18841 , w18842 , w18843 , w18844 , w18845 , w18846 , w18847 , w18848 , w18849 , w18850 , w18851 , w18852 , w18853 , w18854 , w18855 , w18856 , w18857 , w18858 , w18859 , w18860 , w18861 , w18862 , w18863 , w18864 , w18865 , w18866 , w18867 , w18868 , w18869 , w18870 , w18871 , w18872 , w18873 , w18874 , w18875 , w18876 , w18877 , w18878 , w18879 , w18880 , w18881 , w18882 , w18883 , w18884 , w18885 , w18886 , w18887 , w18888 , w18889 , w18890 , w18891 , w18892 , w18893 , w18894 , w18895 , w18896 , w18897 , w18898 , w18899 , w18900 , w18901 , w18902 , w18903 , w18904 , w18905 , w18906 , w18907 , w18908 , w18909 , w18910 , w18911 , w18912 , w18913 , w18914 , w18915 , w18916 , w18917 , w18918 , w18919 , w18920 , w18921 , w18922 , w18923 , w18924 , w18925 , w18926 , w18927 , w18928 , w18929 , w18930 , w18931 , w18932 , w18933 , w18934 , w18935 , w18936 , w18937 , w18938 , w18939 , w18940 , w18941 , w18942 , w18943 , w18944 , w18945 , w18946 , w18947 , w18948 , w18949 , w18950 , w18951 , w18952 , w18953 , w18954 , w18955 , w18956 , w18957 , w18958 , w18959 , w18960 , w18961 , w18962 , w18963 , w18964 , w18965 , w18966 , w18967 , w18968 , w18969 , w18970 , w18971 , w18972 , w18973 , w18974 , w18975 , w18976 , w18977 , w18978 , w18979 , w18980 , w18981 , w18982 , w18983 , w18984 , w18985 , w18986 , w18987 , w18988 , w18989 , w18990 , w18991 , w18992 , w18993 , w18994 , w18995 , w18996 , w18997 , w18998 , w18999 , w19000 , w19001 , w19002 , w19003 , w19004 , w19005 , w19006 , w19007 , w19008 , w19009 , w19010 , w19011 , w19012 , w19013 , w19014 , w19015 , w19016 , w19017 , w19018 , w19019 , w19020 , w19021 , w19022 , w19023 , w19024 , w19025 , w19026 , w19027 , w19028 , w19029 , w19030 , w19031 , w19032 , w19033 , w19034 , w19035 , w19036 , w19037 , w19038 , w19039 , w19040 , w19041 , w19042 , w19043 , w19044 , w19045 , w19046 , w19047 , w19048 , w19049 , w19050 , w19051 , w19052 , w19053 , w19054 , w19055 , w19056 , w19057 , w19058 , w19059 , w19060 , w19061 , w19062 , w19063 , w19064 , w19065 , w19066 , w19067 , w19068 , w19069 , w19070 , w19071 , w19072 , w19073 , w19074 , w19075 , w19076 , w19077 , w19078 , w19079 , w19080 , w19081 , w19082 , w19083 , w19084 , w19085 , w19086 , w19087 , w19088 , w19089 , w19090 , w19091 , w19092 , w19093 , w19094 , w19095 , w19096 , w19097 , w19098 , w19099 , w19100 , w19101 , w19102 , w19103 , w19104 , w19105 , w19106 , w19107 , w19108 , w19109 , w19110 , w19111 , w19112 , w19113 , w19114 , w19115 , w19116 , w19117 , w19118 , w19119 , w19120 , w19121 , w19122 , w19123 , w19124 , w19125 , w19126 , w19127 , w19128 , w19129 , w19130 , w19131 , w19132 , w19133 , w19134 , w19135 , w19136 , w19137 , w19138 , w19139 , w19140 , w19141 , w19142 , w19143 , w19144 , w19145 , w19146 , w19147 , w19148 , w19149 , w19150 , w19151 , w19152 , w19153 , w19154 , w19155 , w19156 , w19157 , w19158 , w19159 , w19160 , w19161 , w19162 , w19163 , w19164 , w19165 , w19166 , w19167 , w19168 , w19169 , w19170 , w19171 , w19172 , w19173 , w19174 , w19175 , w19176 , w19177 , w19178 , w19179 , w19180 , w19181 , w19182 , w19183 , w19184 , w19185 , w19186 , w19187 , w19188 , w19189 , w19190 , w19191 , w19192 , w19193 , w19194 , w19195 , w19196 , w19197 , w19198 , w19199 , w19200 , w19201 , w19202 , w19203 , w19204 , w19205 , w19206 , w19207 , w19208 , w19209 , w19210 , w19211 , w19212 , w19213 , w19214 , w19215 , w19216 , w19217 , w19218 , w19219 , w19220 , w19221 , w19222 , w19223 , w19224 , w19225 , w19226 , w19227 , w19228 , w19229 , w19230 , w19231 , w19232 , w19233 , w19234 , w19235 , w19236 , w19237 , w19238 , w19239 , w19240 , w19241 , w19242 , w19243 , w19244 , w19245 , w19246 , w19247 , w19248 , w19249 , w19250 , w19251 , w19252 , w19253 , w19254 , w19255 , w19256 , w19257 , w19258 , w19259 , w19260 , w19261 , w19262 , w19263 , w19264 , w19265 , w19266 , w19267 , w19268 , w19269 , w19270 , w19271 , w19272 , w19273 , w19274 , w19275 , w19276 , w19277 , w19278 , w19279 , w19280 , w19281 , w19282 , w19283 , w19284 , w19285 , w19286 , w19287 , w19288 , w19289 , w19290 , w19291 , w19292 , w19293 , w19294 , w19295 , w19296 , w19297 , w19298 , w19299 , w19300 , w19301 , w19302 , w19303 , w19304 , w19305 , w19306 , w19307 , w19308 , w19309 , w19310 , w19311 , w19312 , w19313 , w19314 , w19315 , w19316 , w19317 , w19318 , w19319 , w19320 , w19321 , w19322 , w19323 , w19324 , w19325 , w19326 , w19327 , w19328 , w19329 , w19330 , w19331 , w19332 , w19333 , w19334 , w19335 , w19336 , w19337 , w19338 , w19339 , w19340 , w19341 , w19342 , w19343 , w19344 , w19345 , w19346 , w19347 , w19348 , w19349 , w19350 , w19351 , w19352 , w19353 , w19354 , w19355 , w19356 , w19357 , w19358 , w19359 , w19360 , w19361 , w19362 , w19363 , w19364 , w19365 , w19366 , w19367 , w19368 , w19369 , w19370 , w19371 , w19372 , w19373 , w19374 , w19375 , w19376 , w19377 , w19378 , w19379 , w19380 , w19381 , w19382 , w19383 , w19384 , w19385 , w19386 , w19387 , w19388 , w19389 , w19390 , w19391 , w19392 , w19393 , w19394 , w19395 , w19396 , w19397 , w19398 , w19399 , w19400 , w19401 , w19402 , w19403 , w19404 , w19405 , w19406 , w19407 , w19408 , w19409 , w19410 , w19411 , w19412 , w19413 , w19414 , w19415 , w19416 , w19417 , w19418 , w19419 , w19420 , w19421 , w19422 , w19423 , w19424 , w19425 , w19426 , w19427 , w19428 , w19429 , w19430 , w19431 , w19432 , w19433 , w19434 , w19435 , w19436 , w19437 , w19438 , w19439 , w19440 , w19441 , w19442 , w19443 , w19444 , w19445 , w19446 , w19447 , w19448 , w19449 , w19450 , w19451 , w19452 , w19453 , w19454 , w19455 , w19456 , w19457 , w19458 , w19459 , w19460 , w19461 , w19462 , w19463 , w19464 , w19465 , w19466 , w19467 , w19468 , w19469 , w19470 , w19471 , w19472 , w19473 , w19474 , w19475 , w19476 , w19477 , w19478 , w19479 , w19480 , w19481 , w19482 , w19483 , w19484 , w19485 , w19486 , w19487 , w19488 , w19489 , w19490 , w19491 , w19492 , w19493 , w19494 , w19495 , w19496 , w19497 , w19498 , w19499 , w19500 , w19501 , w19502 , w19503 , w19504 , w19505 , w19506 , w19507 , w19508 , w19509 , w19510 , w19511 , w19512 , w19513 , w19514 , w19515 , w19516 , w19517 , w19518 , w19519 , w19520 , w19521 , w19522 , w19523 , w19524 , w19525 , w19526 , w19527 , w19528 , w19529 , w19530 , w19531 , w19532 , w19533 , w19534 , w19535 , w19536 , w19537 , w19538 , w19539 , w19540 , w19541 , w19542 , w19543 , w19544 , w19545 , w19546 , w19547 , w19548 , w19549 , w19550 , w19551 , w19552 , w19553 , w19554 , w19555 , w19556 , w19557 , w19558 , w19559 , w19560 , w19561 , w19562 , w19563 , w19564 , w19565 , w19566 , w19567 , w19568 , w19569 , w19570 , w19571 , w19572 , w19573 , w19574 , w19575 , w19576 , w19577 , w19578 , w19579 , w19580 , w19581 , w19582 , w19583 , w19584 , w19585 , w19586 , w19587 , w19588 , w19589 , w19590 , w19591 , w19592 , w19593 , w19594 , w19595 , w19596 , w19597 , w19598 , w19599 , w19600 , w19601 , w19602 , w19603 , w19604 , w19605 , w19606 , w19607 , w19608 , w19609 , w19610 , w19611 , w19612 , w19613 , w19614 , w19615 , w19616 , w19617 , w19618 , w19619 , w19620 , w19621 , w19622 , w19623 , w19624 , w19625 , w19626 , w19627 , w19628 , w19629 , w19630 , w19631 , w19632 , w19633 , w19634 , w19635 , w19636 , w19637 , w19638 , w19639 , w19640 , w19641 , w19642 , w19643 , w19644 , w19645 , w19646 , w19647 , w19648 , w19649 , w19650 , w19651 , w19652 , w19653 , w19654 , w19655 , w19656 , w19657 , w19658 , w19659 , w19660 , w19661 , w19662 , w19663 , w19664 , w19665 , w19666 , w19667 , w19668 , w19669 , w19670 , w19671 , w19672 , w19673 , w19674 , w19675 , w19676 , w19677 , w19678 , w19679 , w19680 , w19681 , w19682 , w19683 , w19684 , w19685 , w19686 , w19687 , w19688 , w19689 , w19690 , w19691 , w19692 , w19693 , w19694 , w19695 , w19696 , w19697 , w19698 , w19699 , w19700 , w19701 , w19702 , w19703 , w19704 , w19705 , w19706 , w19707 , w19708 , w19709 , w19710 , w19711 , w19712 , w19713 , w19714 , w19715 , w19716 , w19717 , w19718 , w19719 , w19720 , w19721 , w19722 , w19723 , w19724 , w19725 , w19726 , w19727 , w19728 , w19729 , w19730 , w19731 , w19732 , w19733 , w19734 , w19735 , w19736 , w19737 , w19738 , w19739 , w19740 , w19741 , w19742 , w19743 , w19744 , w19745 , w19746 , w19747 , w19748 , w19749 , w19750 , w19751 , w19752 , w19753 , w19754 , w19755 , w19756 , w19757 , w19758 , w19759 , w19760 , w19761 , w19762 , w19763 , w19764 , w19765 , w19766 , w19767 , w19768 , w19769 , w19770 , w19771 , w19772 , w19773 , w19774 , w19775 , w19776 , w19777 , w19778 , w19779 , w19780 , w19781 , w19782 , w19783 , w19784 , w19785 , w19786 , w19787 , w19788 , w19789 , w19790 , w19791 , w19792 , w19793 , w19794 , w19795 , w19796 , w19797 , w19798 , w19799 , w19800 , w19801 , w19802 , w19803 , w19804 , w19805 , w19806 , w19807 , w19808 , w19809 , w19810 , w19811 , w19812 , w19813 , w19814 , w19815 , w19816 , w19817 , w19818 , w19819 , w19820 , w19821 , w19822 , w19823 , w19824 , w19825 , w19826 , w19827 , w19828 , w19829 , w19830 , w19831 , w19832 , w19833 , w19834 , w19835 , w19836 , w19837 , w19838 , w19839 , w19840 , w19841 , w19842 , w19843 , w19844 , w19845 , w19846 , w19847 , w19848 , w19849 , w19850 , w19851 , w19852 , w19853 , w19854 , w19855 , w19856 , w19857 , w19858 , w19859 , w19860 , w19861 , w19862 , w19863 , w19864 , w19865 , w19866 , w19867 , w19868 , w19869 , w19870 , w19871 , w19872 , w19873 , w19874 , w19875 , w19876 , w19877 , w19878 , w19879 , w19880 , w19881 , w19882 , w19883 , w19884 , w19885 , w19886 , w19887 , w19888 , w19889 , w19890 , w19891 , w19892 , w19893 , w19894 , w19895 , w19896 , w19897 , w19898 , w19899 , w19900 , w19901 , w19902 , w19903 , w19904 , w19905 , w19906 , w19907 , w19908 , w19909 , w19910 , w19911 , w19912 , w19913 , w19914 , w19915 , w19916 , w19917 , w19918 , w19919 , w19920 , w19921 , w19922 , w19923 , w19924 , w19925 , w19926 , w19927 , w19928 , w19929 , w19930 , w19931 , w19932 , w19933 , w19934 , w19935 , w19936 , w19937 , w19938 , w19939 , w19940 , w19941 , w19942 , w19943 , w19944 , w19945 , w19946 , w19947 , w19948 , w19949 , w19950 , w19951 , w19952 , w19953 , w19954 , w19955 , w19956 , w19957 , w19958 , w19959 , w19960 , w19961 , w19962 , w19963 , w19964 , w19965 , w19966 , w19967 , w19968 , w19969 , w19970 , w19971 , w19972 , w19973 , w19974 , w19975 , w19976 , w19977 , w19978 , w19979 , w19980 , w19981 , w19982 , w19983 , w19984 , w19985 , w19986 , w19987 , w19988 , w19989 , w19990 , w19991 , w19992 , w19993 , w19994 , w19995 , w19996 , w19997 , w19998 , w19999 , w20000 , w20001 , w20002 , w20003 , w20004 , w20005 , w20006 , w20007 , w20008 , w20009 , w20010 , w20011 , w20012 , w20013 , w20014 , w20015 , w20016 , w20017 , w20018 , w20019 , w20020 , w20021 , w20022 , w20023 , w20024 , w20025 , w20026 , w20027 , w20028 , w20029 , w20030 , w20031 , w20032 , w20033 , w20034 , w20035 , w20036 , w20037 , w20038 , w20039 , w20040 , w20041 , w20042 , w20043 , w20044 , w20045 , w20046 , w20047 , w20048 , w20049 , w20050 , w20051 , w20052 , w20053 , w20054 , w20055 , w20056 , w20057 , w20058 , w20059 , w20060 , w20061 , w20062 , w20063 , w20064 , w20065 , w20066 , w20067 , w20068 , w20069 , w20070 , w20071 , w20072 , w20073 , w20074 , w20075 , w20076 , w20077 , w20078 , w20079 , w20080 , w20081 , w20082 , w20083 , w20084 , w20085 , w20086 , w20087 , w20088 , w20089 , w20090 , w20091 , w20092 , w20093 , w20094 , w20095 , w20096 , w20097 , w20098 , w20099 , w20100 , w20101 , w20102 , w20103 , w20104 , w20105 , w20106 , w20107 , w20108 , w20109 , w20110 , w20111 , w20112 , w20113 , w20114 , w20115 , w20116 , w20117 , w20118 , w20119 , w20120 , w20121 , w20122 , w20123 , w20124 , w20125 , w20126 , w20127 , w20128 , w20129 , w20130 , w20131 , w20132 , w20133 , w20134 , w20135 , w20136 , w20137 , w20138 , w20139 , w20140 , w20141 , w20142 , w20143 , w20144 , w20145 , w20146 , w20147 , w20148 , w20149 , w20150 , w20151 , w20152 , w20153 , w20154 , w20155 , w20156 , w20157 , w20158 , w20159 , w20160 , w20161 , w20162 , w20163 , w20164 , w20165 , w20166 , w20167 , w20168 , w20169 , w20170 , w20171 , w20172 , w20173 , w20174 , w20175 , w20176 , w20177 , w20178 , w20179 , w20180 , w20181 , w20182 , w20183 , w20184 , w20185 , w20186 , w20187 , w20188 , w20189 , w20190 , w20191 , w20192 , w20193 , w20194 , w20195 , w20196 , w20197 , w20198 , w20199 , w20200 , w20201 , w20202 , w20203 , w20204 , w20205 , w20206 , w20207 , w20208 , w20209 , w20210 , w20211 , w20212 , w20213 , w20214 , w20215 , w20216 , w20217 , w20218 , w20219 , w20220 , w20221 , w20222 , w20223 , w20224 , w20225 , w20226 , w20227 , w20228 , w20229 , w20230 , w20231 , w20232 , w20233 , w20234 , w20235 , w20236 , w20237 , w20238 , w20239 , w20240 , w20241 , w20242 , w20243 , w20244 , w20245 , w20246 , w20247 , w20248 , w20249 , w20250 , w20251 , w20252 , w20253 , w20254 , w20255 , w20256 , w20257 , w20258 , w20259 , w20260 , w20261 , w20262 , w20263 , w20264 , w20265 , w20266 , w20267 , w20268 , w20269 , w20270 , w20271 , w20272 , w20273 , w20274 , w20275 , w20276 , w20277 , w20278 , w20279 , w20280 , w20281 , w20282 , w20283 , w20284 , w20285 , w20286 , w20287 , w20288 , w20289 , w20290 , w20291 , w20292 , w20293 , w20294 , w20295 , w20296 , w20297 , w20298 , w20299 , w20300 , w20301 , w20302 , w20303 , w20304 , w20305 , w20306 , w20307 , w20308 , w20309 , w20310 , w20311 , w20312 , w20313 , w20314 , w20315 , w20316 , w20317 , w20318 , w20319 , w20320 , w20321 , w20322 , w20323 , w20324 , w20325 , w20326 , w20327 , w20328 , w20329 , w20330 , w20331 , w20332 , w20333 , w20334 , w20335 , w20336 , w20337 , w20338 , w20339 , w20340 , w20341 , w20342 , w20343 , w20344 , w20345 , w20346 , w20347 , w20348 , w20349 , w20350 , w20351 , w20352 , w20353 , w20354 , w20355 , w20356 , w20357 , w20358 , w20359 , w20360 , w20361 , w20362 , w20363 , w20364 , w20365 , w20366 , w20367 , w20368 , w20369 , w20370 , w20371 , w20372 , w20373 , w20374 , w20375 , w20376 , w20377 , w20378 , w20379 , w20380 , w20381 , w20382 , w20383 , w20384 , w20385 , w20386 , w20387 , w20388 , w20389 , w20390 , w20391 , w20392 , w20393 , w20394 , w20395 , w20396 , w20397 , w20398 , w20399 , w20400 , w20401 , w20402 , w20403 , w20404 , w20405 , w20406 , w20407 , w20408 , w20409 , w20410 , w20411 , w20412 , w20413 , w20414 , w20415 , w20416 , w20417 , w20418 , w20419 , w20420 , w20421 , w20422 , w20423 , w20424 , w20425 , w20426 , w20427 , w20428 , w20429 , w20430 , w20431 , w20432 , w20433 , w20434 , w20435 , w20436 , w20437 , w20438 , w20439 , w20440 , w20441 , w20442 , w20443 , w20444 , w20445 , w20446 , w20447 , w20448 , w20449 , w20450 , w20451 , w20452 , w20453 , w20454 , w20455 , w20456 , w20457 , w20458 , w20459 , w20460 , w20461 , w20462 , w20463 , w20464 , w20465 , w20466 , w20467 , w20468 , w20469 , w20470 , w20471 , w20472 , w20473 , w20474 , w20475 , w20476 , w20477 , w20478 , w20479 , w20480 , w20481 , w20482 , w20483 , w20484 , w20485 , w20486 , w20487 , w20488 , w20489 , w20490 , w20491 , w20492 , w20493 , w20494 , w20495 , w20496 , w20497 , w20498 , w20499 , w20500 , w20501 , w20502 , w20503 , w20504 , w20505 , w20506 , w20507 , w20508 , w20509 , w20510 , w20511 , w20512 , w20513 , w20514 , w20515 , w20516 , w20517 , w20518 , w20519 , w20520 , w20521 , w20522 , w20523 , w20524 , w20525 , w20526 , w20527 , w20528 , w20529 , w20530 , w20531 , w20532 , w20533 , w20534 , w20535 , w20536 , w20537 , w20538 , w20539 , w20540 , w20541 , w20542 , w20543 , w20544 , w20545 , w20546 , w20547 , w20548 , w20549 , w20550 , w20551 , w20552 , w20553 , w20554 , w20555 , w20556 , w20557 , w20558 , w20559 , w20560 , w20561 , w20562 , w20563 , w20564 , w20565 , w20566 , w20567 , w20568 , w20569 , w20570 , w20571 , w20572 , w20573 , w20574 , w20575 , w20576 , w20577 , w20578 , w20579 , w20580 , w20581 , w20582 , w20583 , w20584 , w20585 , w20586 , w20587 , w20588 , w20589 , w20590 , w20591 , w20592 , w20593 , w20594 , w20595 , w20596 , w20597 , w20598 , w20599 , w20600 , w20601 , w20602 , w20603 , w20604 , w20605 , w20606 , w20607 , w20608 , w20609 , w20610 , w20611 , w20612 , w20613 , w20614 , w20615 , w20616 , w20617 , w20618 , w20619 , w20620 , w20621 , w20622 , w20623 , w20624 , w20625 , w20626 , w20627 , w20628 , w20629 , w20630 , w20631 , w20632 , w20633 , w20634 , w20635 , w20636 , w20637 , w20638 , w20639 , w20640 , w20641 , w20642 , w20643 , w20644 , w20645 , w20646 , w20647 , w20648 , w20649 , w20650 , w20651 , w20652 , w20653 , w20654 , w20655 , w20656 , w20657 , w20658 , w20659 , w20660 , w20661 , w20662 , w20663 , w20664 , w20665 , w20666 , w20667 , w20668 , w20669 , w20670 , w20671 , w20672 , w20673 , w20674 , w20675 , w20676 , w20677 , w20678 , w20679 , w20680 , w20681 , w20682 , w20683 , w20684 , w20685 , w20686 , w20687 , w20688 , w20689 , w20690 , w20691 , w20692 , w20693 , w20694 , w20695 , w20696 , w20697 , w20698 , w20699 , w20700 , w20701 , w20702 , w20703 , w20704 , w20705 , w20706 , w20707 , w20708 , w20709 , w20710 , w20711 , w20712 , w20713 , w20714 , w20715 , w20716 , w20717 , w20718 , w20719 , w20720 , w20721 , w20722 , w20723 , w20724 , w20725 , w20726 , w20727 , w20728 , w20729 , w20730 , w20731 , w20732 , w20733 , w20734 , w20735 , w20736 , w20737 , w20738 , w20739 , w20740 , w20741 , w20742 , w20743 , w20744 , w20745 , w20746 , w20747 , w20748 , w20749 , w20750 , w20751 , w20752 , w20753 , w20754 , w20755 , w20756 , w20757 , w20758 , w20759 , w20760 , w20761 , w20762 , w20763 , w20764 , w20765 , w20766 , w20767 , w20768 , w20769 , w20770 , w20771 , w20772 , w20773 , w20774 , w20775 , w20776 , w20777 , w20778 , w20779 , w20780 , w20781 , w20782 , w20783 , w20784 , w20785 , w20786 , w20787 , w20788 , w20789 , w20790 , w20791 , w20792 , w20793 , w20794 , w20795 , w20796 , w20797 , w20798 , w20799 , w20800 , w20801 , w20802 , w20803 , w20804 , w20805 , w20806 , w20807 , w20808 , w20809 , w20810 , w20811 , w20812 , w20813 , w20814 , w20815 , w20816 , w20817 , w20818 , w20819 , w20820 , w20821 , w20822 , w20823 , w20824 , w20825 , w20826 , w20827 , w20828 , w20829 , w20830 , w20831 , w20832 , w20833 , w20834 , w20835 , w20836 , w20837 , w20838 , w20839 , w20840 , w20841 , w20842 , w20843 , w20844 , w20845 , w20846 , w20847 , w20848 , w20849 , w20850 , w20851 , w20852 , w20853 , w20854 , w20855 , w20856 , w20857 , w20858 , w20859 , w20860 , w20861 , w20862 , w20863 , w20864 , w20865 , w20866 , w20867 , w20868 , w20869 , w20870 , w20871 , w20872 , w20873 , w20874 , w20875 , w20876 , w20877 , w20878 , w20879 , w20880 , w20881 , w20882 , w20883 , w20884 , w20885 , w20886 , w20887 , w20888 , w20889 , w20890 , w20891 , w20892 , w20893 , w20894 , w20895 , w20896 , w20897 , w20898 , w20899 , w20900 , w20901 , w20902 , w20903 , w20904 , w20905 , w20906 , w20907 , w20908 , w20909 , w20910 , w20911 , w20912 , w20913 , w20914 , w20915 , w20916 , w20917 , w20918 , w20919 , w20920 , w20921 , w20922 , w20923 , w20924 , w20925 , w20926 , w20927 , w20928 , w20929 , w20930 , w20931 , w20932 , w20933 , w20934 , w20935 , w20936 , w20937 , w20938 , w20939 , w20940 , w20941 , w20942 , w20943 , w20944 , w20945 , w20946 , w20947 , w20948 , w20949 , w20950 , w20951 , w20952 , w20953 , w20954 , w20955 , w20956 , w20957 , w20958 , w20959 , w20960 , w20961 , w20962 , w20963 , w20964 , w20965 , w20966 , w20967 , w20968 , w20969 , w20970 , w20971 , w20972 , w20973 , w20974 , w20975 , w20976 , w20977 , w20978 , w20979 , w20980 , w20981 , w20982 , w20983 , w20984 , w20985 , w20986 , w20987 , w20988 , w20989 , w20990 , w20991 , w20992 , w20993 , w20994 , w20995 , w20996 , w20997 , w20998 , w20999 , w21000 , w21001 , w21002 , w21003 , w21004 , w21005 , w21006 , w21007 , w21008 , w21009 , w21010 , w21011 , w21012 , w21013 , w21014 , w21015 , w21016 , w21017 , w21018 , w21019 , w21020 , w21021 , w21022 , w21023 , w21024 , w21025 , w21026 , w21027 , w21028 , w21029 , w21030 , w21031 , w21032 , w21033 , w21034 , w21035 , w21036 , w21037 , w21038 , w21039 , w21040 , w21041 , w21042 , w21043 , w21044 , w21045 , w21046 , w21047 , w21048 , w21049 , w21050 , w21051 , w21052 , w21053 , w21054 , w21055 , w21056 , w21057 , w21058 , w21059 , w21060 , w21061 , w21062 , w21063 , w21064 , w21065 , w21066 , w21067 , w21068 , w21069 , w21070 , w21071 , w21072 , w21073 , w21074 , w21075 , w21076 , w21077 , w21078 , w21079 , w21080 , w21081 , w21082 , w21083 , w21084 , w21085 , w21086 , w21087 , w21088 , w21089 , w21090 , w21091 , w21092 , w21093 , w21094 , w21095 , w21096 , w21097 , w21098 , w21099 , w21100 , w21101 , w21102 , w21103 , w21104 , w21105 , w21106 , w21107 , w21108 , w21109 , w21110 , w21111 , w21112 , w21113 , w21114 , w21115 , w21116 , w21117 , w21118 , w21119 , w21120 , w21121 , w21122 , w21123 , w21124 , w21125 , w21126 , w21127 , w21128 , w21129 , w21130 , w21131 , w21132 , w21133 , w21134 , w21135 , w21136 , w21137 , w21138 , w21139 , w21140 , w21141 , w21142 , w21143 , w21144 , w21145 , w21146 , w21147 , w21148 , w21149 , w21150 , w21151 , w21152 , w21153 , w21154 , w21155 , w21156 , w21157 , w21158 , w21159 , w21160 , w21161 , w21162 , w21163 , w21164 , w21165 , w21166 , w21167 , w21168 , w21169 , w21170 , w21171 , w21172 , w21173 , w21174 , w21175 , w21176 , w21177 , w21178 , w21179 , w21180 , w21181 , w21182 , w21183 , w21184 , w21185 , w21186 , w21187 , w21188 , w21189 , w21190 , w21191 , w21192 , w21193 , w21194 , w21195 , w21196 , w21197 , w21198 , w21199 , w21200 , w21201 , w21202 , w21203 , w21204 , w21205 , w21206 , w21207 , w21208 , w21209 , w21210 , w21211 , w21212 , w21213 , w21214 , w21215 , w21216 , w21217 , w21218 , w21219 , w21220 , w21221 , w21222 , w21223 , w21224 , w21225 , w21226 , w21227 , w21228 , w21229 , w21230 , w21231 , w21232 , w21233 , w21234 , w21235 , w21236 , w21237 , w21238 , w21239 , w21240 , w21241 , w21242 , w21243 , w21244 , w21245 , w21246 , w21247 , w21248 , w21249 , w21250 , w21251 , w21252 , w21253 , w21254 , w21255 , w21256 , w21257 , w21258 , w21259 , w21260 , w21261 , w21262 , w21263 , w21264 , w21265 , w21266 , w21267 , w21268 , w21269 , w21270 , w21271 , w21272 , w21273 , w21274 , w21275 , w21276 , w21277 , w21278 , w21279 , w21280 , w21281 , w21282 , w21283 , w21284 , w21285 , w21286 , w21287 , w21288 , w21289 , w21290 , w21291 , w21292 , w21293 , w21294 , w21295 , w21296 , w21297 , w21298 , w21299 , w21300 , w21301 , w21302 , w21303 , w21304 , w21305 , w21306 , w21307 , w21308 , w21309 , w21310 , w21311 , w21312 , w21313 , w21314 , w21315 , w21316 , w21317 , w21318 , w21319 , w21320 , w21321 , w21322 , w21323 , w21324 , w21325 , w21326 , w21327 , w21328 , w21329 , w21330 , w21331 , w21332 , w21333 , w21334 , w21335 , w21336 , w21337 , w21338 , w21339 , w21340 , w21341 , w21342 , w21343 , w21344 , w21345 , w21346 , w21347 , w21348 , w21349 , w21350 , w21351 , w21352 , w21353 , w21354 , w21355 , w21356 , w21357 , w21358 , w21359 , w21360 , w21361 , w21362 , w21363 , w21364 , w21365 , w21366 , w21367 , w21368 , w21369 , w21370 , w21371 , w21372 , w21373 , w21374 , w21375 , w21376 , w21377 , w21378 , w21379 , w21380 , w21381 , w21382 , w21383 , w21384 , w21385 , w21386 , w21387 , w21388 , w21389 , w21390 , w21391 , w21392 , w21393 , w21394 , w21395 , w21396 , w21397 , w21398 , w21399 , w21400 , w21401 , w21402 , w21403 , w21404 , w21405 , w21406 , w21407 , w21408 , w21409 , w21410 , w21411 , w21412 , w21413 , w21414 , w21415 , w21416 , w21417 , w21418 , w21419 , w21420 , w21421 , w21422 , w21423 , w21424 , w21425 , w21426 , w21427 , w21428 , w21429 , w21430 , w21431 , w21432 , w21433 , w21434 , w21435 , w21436 , w21437 , w21438 , w21439 , w21440 , w21441 , w21442 , w21443 , w21444 , w21445 , w21446 , w21447 , w21448 , w21449 , w21450 , w21451 , w21452 , w21453 , w21454 , w21455 , w21456 , w21457 , w21458 , w21459 , w21460 , w21461 , w21462 , w21463 , w21464 , w21465 , w21466 , w21467 , w21468 , w21469 , w21470 , w21471 , w21472 , w21473 , w21474 , w21475 , w21476 , w21477 , w21478 , w21479 , w21480 , w21481 , w21482 , w21483 , w21484 , w21485 , w21486 , w21487 , w21488 , w21489 , w21490 , w21491 , w21492 , w21493 , w21494 , w21495 , w21496 , w21497 , w21498 , w21499 , w21500 , w21501 , w21502 , w21503 , w21504 , w21505 , w21506 , w21507 , w21508 , w21509 , w21510 , w21511 , w21512 , w21513 , w21514 , w21515 , w21516 , w21517 , w21518 , w21519 , w21520 , w21521 , w21522 , w21523 , w21524 , w21525 , w21526 , w21527 , w21528 , w21529 , w21530 , w21531 , w21532 , w21533 , w21534 , w21535 , w21536 , w21537 , w21538 , w21539 , w21540 , w21541 , w21542 , w21543 , w21544 , w21545 , w21546 , w21547 , w21548 , w21549 , w21550 , w21551 , w21552 , w21553 , w21554 , w21555 , w21556 , w21557 , w21558 , w21559 , w21560 , w21561 , w21562 , w21563 , w21564 , w21565 , w21566 , w21567 , w21568 , w21569 , w21570 , w21571 , w21572 , w21573 , w21574 , w21575 , w21576 , w21577 , w21578 , w21579 , w21580 , w21581 , w21582 , w21583 , w21584 , w21585 , w21586 , w21587 , w21588 , w21589 , w21590 , w21591 , w21592 , w21593 , w21594 , w21595 , w21596 , w21597 , w21598 , w21599 , w21600 , w21601 , w21602 , w21603 , w21604 , w21605 , w21606 , w21607 , w21608 , w21609 , w21610 , w21611 , w21612 , w21613 , w21614 , w21615 , w21616 , w21617 , w21618 , w21619 , w21620 , w21621 , w21622 , w21623 , w21624 , w21625 , w21626 , w21627 , w21628 , w21629 , w21630 , w21631 , w21632 , w21633 , w21634 , w21635 , w21636 , w21637 , w21638 , w21639 , w21640 , w21641 , w21642 , w21643 , w21644 , w21645 , w21646 , w21647 , w21648 , w21649 , w21650 , w21651 , w21652 , w21653 , w21654 , w21655 , w21656 , w21657 , w21658 , w21659 , w21660 , w21661 , w21662 , w21663 , w21664 , w21665 , w21666 , w21667 , w21668 , w21669 , w21670 , w21671 , w21672 , w21673 , w21674 , w21675 , w21676 , w21677 , w21678 , w21679 , w21680 , w21681 , w21682 , w21683 , w21684 , w21685 , w21686 , w21687 , w21688 , w21689 , w21690 , w21691 , w21692 , w21693 , w21694 , w21695 , w21696 , w21697 , w21698 , w21699 , w21700 , w21701 , w21702 , w21703 , w21704 , w21705 , w21706 , w21707 , w21708 , w21709 , w21710 , w21711 , w21712 , w21713 , w21714 , w21715 , w21716 , w21717 , w21718 , w21719 , w21720 , w21721 , w21722 , w21723 , w21724 , w21725 , w21726 , w21727 , w21728 , w21729 , w21730 , w21731 , w21732 , w21733 , w21734 , w21735 , w21736 , w21737 , w21738 , w21739 , w21740 , w21741 , w21742 , w21743 , w21744 , w21745 , w21746 , w21747 , w21748 , w21749 , w21750 , w21751 , w21752 , w21753 , w21754 , w21755 , w21756 , w21757 , w21758 , w21759 , w21760 , w21761 , w21762 , w21763 , w21764 , w21765 , w21766 , w21767 , w21768 , w21769 , w21770 , w21771 , w21772 , w21773 , w21774 , w21775 , w21776 , w21777 , w21778 , w21779 , w21780 , w21781 , w21782 , w21783 , w21784 , w21785 , w21786 , w21787 , w21788 , w21789 , w21790 , w21791 , w21792 , w21793 , w21794 , w21795 , w21796 , w21797 , w21798 , w21799 , w21800 , w21801 , w21802 , w21803 , w21804 , w21805 , w21806 , w21807 , w21808 , w21809 , w21810 , w21811 , w21812 , w21813 , w21814 , w21815 , w21816 , w21817 , w21818 , w21819 , w21820 , w21821 , w21822 , w21823 , w21824 , w21825 , w21826 , w21827 , w21828 , w21829 , w21830 , w21831 , w21832 , w21833 , w21834 , w21835 , w21836 , w21837 , w21838 , w21839 , w21840 , w21841 , w21842 , w21843 , w21844 , w21845 , w21846 , w21847 , w21848 , w21849 , w21850 , w21851 , w21852 , w21853 , w21854 , w21855 , w21856 , w21857 , w21858 , w21859 , w21860 , w21861 , w21862 , w21863 , w21864 , w21865 , w21866 , w21867 , w21868 , w21869 , w21870 , w21871 , w21872 , w21873 , w21874 , w21875 , w21876 , w21877 , w21878 , w21879 , w21880 , w21881 , w21882 , w21883 , w21884 , w21885 , w21886 , w21887 , w21888 , w21889 , w21890 , w21891 , w21892 , w21893 , w21894 , w21895 , w21896 , w21897 , w21898 , w21899 , w21900 , w21901 , w21902 , w21903 , w21904 , w21905 , w21906 , w21907 , w21908 , w21909 , w21910 , w21911 , w21912 , w21913 , w21914 , w21915 , w21916 , w21917 , w21918 , w21919 , w21920 , w21921 , w21922 , w21923 , w21924 , w21925 , w21926 , w21927 , w21928 , w21929 , w21930 , w21931 , w21932 , w21933 , w21934 , w21935 , w21936 , w21937 , w21938 , w21939 , w21940 , w21941 , w21942 , w21943 , w21944 , w21945 , w21946 , w21947 , w21948 , w21949 , w21950 , w21951 , w21952 , w21953 , w21954 , w21955 , w21956 , w21957 , w21958 , w21959 , w21960 , w21961 , w21962 , w21963 , w21964 , w21965 , w21966 , w21967 , w21968 , w21969 , w21970 , w21971 , w21972 , w21973 , w21974 , w21975 , w21976 , w21977 , w21978 , w21979 , w21980 , w21981 , w21982 , w21983 , w21984 , w21985 , w21986 , w21987 , w21988 , w21989 , w21990 , w21991 , w21992 , w21993 , w21994 , w21995 , w21996 , w21997 , w21998 , w21999 , w22000 , w22001 , w22002 , w22003 , w22004 , w22005 , w22006 , w22007 , w22008 , w22009 , w22010 , w22011 , w22012 , w22013 , w22014 , w22015 , w22016 , w22017 , w22018 , w22019 , w22020 , w22021 , w22022 , w22023 , w22024 , w22025 , w22026 , w22027 , w22028 , w22029 , w22030 , w22031 , w22032 , w22033 , w22034 , w22035 , w22036 , w22037 , w22038 , w22039 , w22040 , w22041 , w22042 , w22043 , w22044 , w22045 , w22046 , w22047 , w22048 , w22049 , w22050 , w22051 , w22052 , w22053 , w22054 , w22055 , w22056 , w22057 , w22058 , w22059 , w22060 , w22061 , w22062 , w22063 , w22064 , w22065 , w22066 , w22067 , w22068 , w22069 , w22070 , w22071 , w22072 , w22073 , w22074 , w22075 , w22076 , w22077 , w22078 , w22079 , w22080 , w22081 , w22082 , w22083 , w22084 , w22085 , w22086 , w22087 , w22088 , w22089 , w22090 , w22091 , w22092 , w22093 , w22094 , w22095 , w22096 , w22097 , w22098 , w22099 , w22100 , w22101 , w22102 , w22103 , w22104 , w22105 , w22106 , w22107 , w22108 , w22109 , w22110 , w22111 , w22112 , w22113 , w22114 , w22115 , w22116 , w22117 , w22118 , w22119 , w22120 , w22121 , w22122 , w22123 , w22124 , w22125 , w22126 , w22127 , w22128 , w22129 , w22130 , w22131 , w22132 , w22133 , w22134 , w22135 , w22136 , w22137 , w22138 , w22139 , w22140 , w22141 , w22142 , w22143 , w22144 , w22145 , w22146 , w22147 , w22148 , w22149 , w22150 , w22151 , w22152 , w22153 , w22154 , w22155 , w22156 , w22157 , w22158 , w22159 , w22160 , w22161 , w22162 , w22163 , w22164 , w22165 , w22166 , w22167 , w22168 , w22169 , w22170 , w22171 , w22172 , w22173 , w22174 , w22175 , w22176 , w22177 , w22178 , w22179 , w22180 , w22181 , w22182 , w22183 , w22184 , w22185 , w22186 , w22187 , w22188 , w22189 , w22190 , w22191 , w22192 , w22193 , w22194 , w22195 , w22196 , w22197 , w22198 , w22199 , w22200 , w22201 , w22202 , w22203 , w22204 , w22205 , w22206 , w22207 , w22208 , w22209 , w22210 , w22211 , w22212 , w22213 , w22214 , w22215 , w22216 , w22217 , w22218 , w22219 , w22220 , w22221 , w22222 , w22223 , w22224 , w22225 , w22226 , w22227 , w22228 , w22229 , w22230 , w22231 , w22232 , w22233 , w22234 , w22235 , w22236 , w22237 , w22238 , w22239 , w22240 , w22241 , w22242 , w22243 , w22244 , w22245 , w22246 , w22247 , w22248 , w22249 , w22250 , w22251 , w22252 , w22253 , w22254 , w22255 , w22256 , w22257 , w22258 , w22259 , w22260 , w22261 , w22262 , w22263 , w22264 , w22265 , w22266 , w22267 , w22268 , w22269 , w22270 , w22271 , w22272 , w22273 , w22274 , w22275 , w22276 , w22277 , w22278 , w22279 , w22280 , w22281 , w22282 , w22283 , w22284 , w22285 , w22286 , w22287 , w22288 , w22289 , w22290 , w22291 , w22292 , w22293 , w22294 , w22295 , w22296 , w22297 , w22298 , w22299 , w22300 , w22301 , w22302 , w22303 , w22304 , w22305 , w22306 , w22307 , w22308 , w22309 , w22310 , w22311 , w22312 , w22313 , w22314 , w22315 , w22316 , w22317 , w22318 , w22319 , w22320 , w22321 , w22322 , w22323 , w22324 , w22325 , w22326 , w22327 , w22328 , w22329 , w22330 , w22331 , w22332 , w22333 , w22334 , w22335 , w22336 , w22337 , w22338 , w22339 , w22340 , w22341 , w22342 , w22343 , w22344 , w22345 , w22346 , w22347 , w22348 , w22349 , w22350 , w22351 , w22352 , w22353 , w22354 , w22355 , w22356 , w22357 , w22358 , w22359 , w22360 , w22361 , w22362 , w22363 , w22364 , w22365 , w22366 , w22367 , w22368 , w22369 , w22370 , w22371 , w22372 , w22373 , w22374 , w22375 , w22376 , w22377 , w22378 , w22379 , w22380 , w22381 , w22382 , w22383 , w22384 , w22385 , w22386 , w22387 , w22388 , w22389 , w22390 , w22391 , w22392 , w22393 , w22394 , w22395 , w22396 , w22397 , w22398 , w22399 , w22400 , w22401 , w22402 , w22403 , w22404 , w22405 , w22406 , w22407 , w22408 , w22409 , w22410 , w22411 , w22412 , w22413 , w22414 , w22415 , w22416 , w22417 , w22418 , w22419 , w22420 , w22421 , w22422 , w22423 , w22424 , w22425 , w22426 , w22427 , w22428 , w22429 , w22430 , w22431 , w22432 , w22433 , w22434 , w22435 , w22436 , w22437 , w22438 , w22439 , w22440 , w22441 , w22442 , w22443 , w22444 , w22445 , w22446 , w22447 , w22448 , w22449 , w22450 , w22451 , w22452 , w22453 , w22454 , w22455 , w22456 , w22457 , w22458 , w22459 , w22460 , w22461 , w22462 , w22463 , w22464 , w22465 , w22466 , w22467 , w22468 , w22469 , w22470 , w22471 , w22472 , w22473 , w22474 , w22475 , w22476 , w22477 , w22478 , w22479 , w22480 , w22481 , w22482 , w22483 , w22484 , w22485 , w22486 , w22487 , w22488 , w22489 , w22490 , w22491 , w22492 , w22493 , w22494 , w22495 , w22496 , w22497 , w22498 , w22499 , w22500 , w22501 , w22502 , w22503 , w22504 , w22505 , w22506 , w22507 , w22508 , w22509 , w22510 , w22511 , w22512 , w22513 , w22514 , w22515 , w22516 , w22517 , w22518 , w22519 , w22520 , w22521 , w22522 , w22523 , w22524 , w22525 , w22526 , w22527 , w22528 , w22529 , w22530 , w22531 , w22532 , w22533 , w22534 , w22535 , w22536 , w22537 , w22538 , w22539 , w22540 , w22541 , w22542 , w22543 , w22544 , w22545 , w22546 , w22547 , w22548 , w22549 , w22550 , w22551 , w22552 , w22553 , w22554 , w22555 , w22556 , w22557 , w22558 , w22559 , w22560 , w22561 , w22562 , w22563 , w22564 , w22565 , w22566 , w22567 , w22568 , w22569 , w22570 , w22571 , w22572 , w22573 , w22574 , w22575 , w22576 , w22577 , w22578 , w22579 , w22580 , w22581 , w22582 , w22583 , w22584 , w22585 , w22586 , w22587 , w22588 , w22589 , w22590 , w22591 , w22592 , w22593 , w22594 , w22595 , w22596 , w22597 , w22598 , w22599 , w22600 , w22601 , w22602 , w22603 , w22604 , w22605 , w22606 , w22607 , w22608 , w22609 , w22610 , w22611 , w22612 , w22613 , w22614 , w22615 , w22616 , w22617 , w22618 , w22619 , w22620 , w22621 , w22622 , w22623 , w22624 , w22625 , w22626 , w22627 , w22628 , w22629 , w22630 , w22631 , w22632 , w22633 , w22634 , w22635 , w22636 , w22637 , w22638 , w22639 , w22640 , w22641 , w22642 , w22643 , w22644 , w22645 , w22646 , w22647 , w22648 , w22649 , w22650 , w22651 , w22652 , w22653 , w22654 , w22655 , w22656 , w22657 , w22658 , w22659 , w22660 , w22661 , w22662 , w22663 , w22664 , w22665 , w22666 , w22667 , w22668 , w22669 , w22670 , w22671 , w22672 , w22673 , w22674 , w22675 , w22676 , w22677 , w22678 , w22679 , w22680 , w22681 , w22682 , w22683 , w22684 , w22685 , w22686 , w22687 , w22688 , w22689 , w22690 , w22691 , w22692 , w22693 , w22694 , w22695 , w22696 , w22697 , w22698 , w22699 , w22700 , w22701 , w22702 , w22703 , w22704 , w22705 , w22706 , w22707 , w22708 , w22709 , w22710 , w22711 , w22712 , w22713 , w22714 , w22715 , w22716 , w22717 , w22718 , w22719 , w22720 , w22721 , w22722 , w22723 , w22724 , w22725 , w22726 , w22727 , w22728 , w22729 , w22730 , w22731 , w22732 , w22733 , w22734 , w22735 , w22736 , w22737 , w22738 , w22739 , w22740 , w22741 , w22742 , w22743 , w22744 , w22745 , w22746 , w22747 , w22748 , w22749 , w22750 , w22751 , w22752 , w22753 , w22754 , w22755 , w22756 , w22757 , w22758 , w22759 , w22760 , w22761 , w22762 , w22763 , w22764 , w22765 , w22766 , w22767 , w22768 , w22769 , w22770 , w22771 , w22772 , w22773 , w22774 , w22775 , w22776 , w22777 , w22778 , w22779 , w22780 , w22781 , w22782 , w22783 , w22784 , w22785 , w22786 , w22787 , w22788 , w22789 , w22790 , w22791 , w22792 , w22793 , w22794 , w22795 , w22796 , w22797 , w22798 , w22799 , w22800 , w22801 , w22802 , w22803 , w22804 , w22805 , w22806 , w22807 , w22808 , w22809 , w22810 , w22811 , w22812 , w22813 , w22814 , w22815 , w22816 , w22817 , w22818 , w22819 , w22820 , w22821 , w22822 , w22823 , w22824 , w22825 , w22826 , w22827 , w22828 , w22829 , w22830 , w22831 , w22832 , w22833 , w22834 , w22835 , w22836 , w22837 , w22838 , w22839 , w22840 , w22841 , w22842 , w22843 , w22844 , w22845 , w22846 , w22847 , w22848 , w22849 , w22850 , w22851 , w22852 , w22853 , w22854 , w22855 , w22856 , w22857 , w22858 , w22859 , w22860 , w22861 , w22862 , w22863 , w22864 , w22865 , w22866 , w22867 , w22868 , w22869 , w22870 , w22871 , w22872 , w22873 , w22874 , w22875 , w22876 , w22877 , w22878 , w22879 , w22880 , w22881 , w22882 , w22883 , w22884 , w22885 , w22886 , w22887 , w22888 , w22889 , w22890 , w22891 , w22892 , w22893 , w22894 , w22895 , w22896 , w22897 , w22898 , w22899 , w22900 , w22901 , w22902 , w22903 , w22904 , w22905 , w22906 , w22907 , w22908 , w22909 , w22910 , w22911 , w22912 , w22913 , w22914 , w22915 , w22916 , w22917 , w22918 , w22919 , w22920 , w22921 , w22922 , w22923 , w22924 , w22925 , w22926 , w22927 , w22928 , w22929 , w22930 , w22931 , w22932 , w22933 , w22934 , w22935 , w22936 , w22937 , w22938 , w22939 , w22940 , w22941 , w22942 , w22943 , w22944 , w22945 , w22946 , w22947 , w22948 , w22949 , w22950 , w22951 , w22952 , w22953 , w22954 , w22955 , w22956 , w22957 , w22958 , w22959 , w22960 , w22961 , w22962 , w22963 , w22964 , w22965 , w22966 , w22967 , w22968 , w22969 , w22970 , w22971 , w22972 , w22973 , w22974 , w22975 , w22976 , w22977 , w22978 , w22979 , w22980 , w22981 , w22982 , w22983 , w22984 , w22985 , w22986 , w22987 , w22988 , w22989 , w22990 , w22991 , w22992 , w22993 , w22994 , w22995 , w22996 , w22997 , w22998 , w22999 , w23000 , w23001 , w23002 , w23003 , w23004 , w23005 , w23006 , w23007 , w23008 , w23009 , w23010 , w23011 , w23012 , w23013 , w23014 , w23015 , w23016 , w23017 , w23018 , w23019 , w23020 , w23021 , w23022 , w23023 , w23024 , w23025 , w23026 , w23027 , w23028 , w23029 , w23030 , w23031 , w23032 , w23033 , w23034 , w23035 , w23036 , w23037 , w23038 ;
  assign zero = 0;
  assign w33 = \pi04 ^ \pi05 ;
  assign w34 = \pi02 ^ \pi03 ;
  assign w35 = ~w33 & w34 ;
  assign w36 = \pi29 ^ \pi30 ;
  assign w37 = \pi31 & w36 ;
  assign w38 = ~\pi24 & \pi26 ;
  assign w39 = ( \pi23 & ~\pi24 ) | ( \pi23 & \pi25 ) | ( ~\pi24 & \pi25 ) ;
  assign w40 = w38 & ~w39 ;
  assign w41 = \pi28 & ~\pi30 ;
  assign w42 = ( \pi27 & ~\pi28 ) | ( \pi27 & \pi29 ) | ( ~\pi28 & \pi29 ) ;
  assign w43 = w41 & w42 ;
  assign w44 = w40 & w43 ;
  assign w45 = \pi28 | \pi30 ;
  assign w46 = ( ~\pi27 & \pi28 ) | ( ~\pi27 & \pi29 ) | ( \pi28 & \pi29 ) ;
  assign w47 = ~w45 & w46 ;
  assign w48 = \pi25 & \pi26 ;
  assign w49 = ~\pi23 & w48 ;
  assign w50 = ( \pi23 & \pi24 ) | ( \pi23 & w47 ) | ( \pi24 & w47 ) ;
  assign w51 = w49 & w50 ;
  assign w52 = \pi24 | \pi26 ;
  assign w53 = w39 | w52 ;
  assign w54 = \pi28 & \pi30 ;
  assign w55 = w42 & w54 ;
  assign w56 = ~w53 & w55 ;
  assign w57 = ( \pi23 & \pi24 ) | ( \pi23 & \pi25 ) | ( \pi24 & \pi25 ) ;
  assign w58 = ~w52 & w57 ;
  assign w59 = w47 & w58 ;
  assign w60 = \pi24 & ~\pi26 ;
  assign w61 = w39 & w60 ;
  assign w62 = w42 | w45 ;
  assign w63 = w61 & ~w62 ;
  assign w64 = w59 | w63 ;
  assign w65 = \pi25 & ~\pi26 ;
  assign w66 = ~\pi23 & w65 ;
  assign w67 = ( \pi23 & ~\pi24 ) | ( \pi23 & w55 ) | ( ~\pi24 & w55 ) ;
  assign w68 = w66 & w67 ;
  assign w69 = ~\pi28 & \pi30 ;
  assign w70 = ( \pi27 & \pi28 ) | ( \pi27 & \pi29 ) | ( \pi28 & \pi29 ) ;
  assign w71 = w69 & w70 ;
  assign w72 = \pi23 & w48 ;
  assign w73 = ( \pi23 & \pi24 ) | ( \pi23 & ~w71 ) | ( \pi24 & ~w71 ) ;
  assign w74 = w72 & ~w73 ;
  assign w75 = w54 & ~w70 ;
  assign w76 = w61 & w75 ;
  assign w77 = ( ~\pi23 & \pi24 ) | ( ~\pi23 & \pi25 ) | ( \pi24 & \pi25 ) ;
  assign w78 = w60 & ~w77 ;
  assign w79 = ( \pi27 & \pi28 ) | ( \pi27 & ~\pi29 ) | ( \pi28 & ~\pi29 ) ;
  assign w80 = w69 & w79 ;
  assign w81 = w78 & w80 ;
  assign w82 = w76 | w81 ;
  assign w83 = w46 & w69 ;
  assign w84 = w58 & w83 ;
  assign w85 = ( \pi23 & \pi24 ) | ( \pi23 & ~w47 ) | ( \pi24 & ~w47 ) ;
  assign w86 = w72 & ~w85 ;
  assign w87 = w84 | w86 ;
  assign w88 = ~w53 & w83 ;
  assign w89 = ~w57 & w60 ;
  assign w90 = w75 & w89 ;
  assign w91 = w38 & w77 ;
  assign w92 = w47 & w91 ;
  assign w93 = \pi24 & \pi26 ;
  assign w94 = ~w77 & w93 ;
  assign w95 = w47 & w94 ;
  assign w96 = w92 | w95 ;
  assign w97 = w41 & ~w70 ;
  assign w98 = w78 & w97 ;
  assign w99 = ( \pi23 & \pi24 ) | ( \pi23 & ~\pi25 ) | ( \pi24 & ~\pi25 ) ;
  assign w100 = ~w52 & w99 ;
  assign w101 = w97 & w100 ;
  assign w102 = ~w42 & w69 ;
  assign w103 = w78 & w102 ;
  assign w104 = w75 & w94 ;
  assign w105 = w103 | w104 ;
  assign w106 = w98 | w105 ;
  assign w107 = ( w96 & ~w98 ) | ( w96 & w101 ) | ( ~w98 & w101 ) ;
  assign w108 = w106 | w107 ;
  assign w109 = ( ~w88 & w90 ) | ( ~w88 & w108 ) | ( w90 & w108 ) ;
  assign w110 = w88 | w109 ;
  assign w111 = ~w62 & w94 ;
  assign w112 = w41 & ~w46 ;
  assign w113 = w89 & w112 ;
  assign w114 = w40 & w112 ;
  assign w115 = w71 & w94 ;
  assign w116 = w40 & w83 ;
  assign w117 = ~w57 & w93 ;
  assign w118 = w83 & w117 ;
  assign w119 = w80 & w91 ;
  assign w120 = w80 & w89 ;
  assign w121 = ( \pi23 & ~\pi24 ) | ( \pi23 & w102 ) | ( ~\pi24 & w102 ) ;
  assign w122 = w66 & w121 ;
  assign w123 = ~w46 & w54 ;
  assign w124 = w94 & w123 ;
  assign w125 = w83 & w91 ;
  assign w126 = w124 | w125 ;
  assign w127 = w58 & w97 ;
  assign w128 = w47 & w117 ;
  assign w129 = w127 | w128 ;
  assign w130 = w41 & ~w79 ;
  assign w131 = w58 & w130 ;
  assign w132 = w39 & w93 ;
  assign w133 = w97 & w132 ;
  assign w134 = ( \pi23 & \pi24 ) | ( \pi23 & w112 ) | ( \pi24 & w112 ) ;
  assign w135 = w49 & w134 ;
  assign w136 = w91 & w112 ;
  assign w137 = ~w45 & w79 ;
  assign w138 = w91 & w137 ;
  assign w139 = w80 & w94 ;
  assign w140 = ( \pi23 & \pi24 ) | ( \pi23 & w123 ) | ( \pi24 & w123 ) ;
  assign w141 = w49 & w140 ;
  assign w142 = w97 & w117 ;
  assign w143 = w80 & w100 ;
  assign w144 = ~w53 & w112 ;
  assign w145 = w54 & ~w79 ;
  assign w146 = ( \pi23 & \pi24 ) | ( \pi23 & ~w145 ) | ( \pi24 & ~w145 ) ;
  assign w147 = w72 & ~w146 ;
  assign w148 = w60 & ~w99 ;
  assign w149 = w83 & w148 ;
  assign w150 = ( w143 & w144 ) | ( w143 & ~w147 ) | ( w144 & ~w147 ) ;
  assign w151 = w141 | w142 ;
  assign w152 = ( ~w142 & w147 ) | ( ~w142 & w149 ) | ( w147 & w149 ) ;
  assign w153 = w151 | w152 ;
  assign w154 = w150 | w153 ;
  assign w155 = ( w135 & w136 ) | ( w135 & ~w138 ) | ( w136 & ~w138 ) ;
  assign w156 = w133 | w154 ;
  assign w157 = ( ~w133 & w138 ) | ( ~w133 & w139 ) | ( w138 & w139 ) ;
  assign w158 = w156 | w157 ;
  assign w159 = w155 | w158 ;
  assign w160 = w131 | w159 ;
  assign w161 = w43 & w91 ;
  assign w162 = ( \pi23 & \pi24 ) | ( \pi23 & ~w80 ) | ( \pi24 & ~w80 ) ;
  assign w163 = w72 & ~w162 ;
  assign w164 = w89 & w123 ;
  assign w165 = ~w62 & w132 ;
  assign w166 = ( \pi23 & ~\pi24 ) | ( \pi23 & w137 ) | ( ~\pi24 & w137 ) ;
  assign w167 = w66 & w166 ;
  assign w168 = w165 | w167 ;
  assign w169 = w75 & w78 ;
  assign w170 = w164 | w169 ;
  assign w171 = w161 | w170 ;
  assign w172 = ( ~w161 & w163 ) | ( ~w161 & w168 ) | ( w163 & w168 ) ;
  assign w173 = w171 | w172 ;
  assign w174 = ~w45 & w70 ;
  assign w175 = w148 & w174 ;
  assign w176 = w94 & w174 ;
  assign w177 = w175 | w176 ;
  assign w178 = w94 & w145 ;
  assign w179 = w58 & w112 ;
  assign w180 = w55 & w117 ;
  assign w181 = w179 | w180 ;
  assign w182 = w178 | w181 ;
  assign w183 = w173 | w182 ;
  assign w184 = ( w160 & ~w173 ) | ( w160 & w177 ) | ( ~w173 & w177 ) ;
  assign w185 = w183 | w184 ;
  assign w186 = w122 | w126 ;
  assign w187 = ( ~w126 & w129 ) | ( ~w126 & w185 ) | ( w129 & w185 ) ;
  assign w188 = w186 | w187 ;
  assign w189 = ( w116 & w118 ) | ( w116 & ~w119 ) | ( w118 & ~w119 ) ;
  assign w190 = w115 | w188 ;
  assign w191 = ( ~w115 & w119 ) | ( ~w115 & w120 ) | ( w119 & w120 ) ;
  assign w192 = w190 | w191 ;
  assign w193 = w189 | w192 ;
  assign w194 = w111 | w114 ;
  assign w195 = ( ~w111 & w113 ) | ( ~w111 & w193 ) | ( w113 & w193 ) ;
  assign w196 = w194 | w195 ;
  assign w197 = ( \pi23 & \pi24 ) | ( \pi23 & w43 ) | ( \pi24 & w43 ) ;
  assign w198 = w49 & w197 ;
  assign w199 = w83 & w132 ;
  assign w200 = ( \pi23 & \pi24 ) | ( \pi23 & w102 ) | ( \pi24 & w102 ) ;
  assign w201 = w49 & w200 ;
  assign w202 = ~w53 & w174 ;
  assign w203 = w58 & w71 ;
  assign w204 = w202 | w203 ;
  assign w205 = w55 & w89 ;
  assign w206 = w40 & w123 ;
  assign w207 = ( \pi23 & \pi24 ) | ( \pi23 & ~w43 ) | ( \pi24 & ~w43 ) ;
  assign w208 = w72 & ~w207 ;
  assign w209 = w94 & w102 ;
  assign w210 = w40 & w145 ;
  assign w211 = ( w208 & ~w209 ) | ( w208 & w210 ) | ( ~w209 & w210 ) ;
  assign w212 = w209 | w211 ;
  assign w213 = ( \pi23 & \pi24 ) | ( \pi23 & w75 ) | ( \pi24 & w75 ) ;
  assign w214 = w49 & w213 ;
  assign w215 = w117 & w174 ;
  assign w216 = w214 | w215 ;
  assign w217 = ( \pi23 & \pi24 ) | ( \pi23 & w83 ) | ( \pi24 & w83 ) ;
  assign w218 = w49 & w217 ;
  assign w219 = w112 & w117 ;
  assign w220 = w123 & w148 ;
  assign w221 = w112 & w148 ;
  assign w222 = w220 | w221 ;
  assign w223 = ~w62 & w91 ;
  assign w224 = w94 & w137 ;
  assign w225 = w71 & w132 ;
  assign w226 = w43 & w100 ;
  assign w227 = w47 & w100 ;
  assign w228 = ( \pi23 & \pi24 ) | ( \pi23 & ~w174 ) | ( \pi24 & ~w174 ) ;
  assign w229 = w72 & ~w228 ;
  assign w230 = w80 & w148 ;
  assign w231 = ( \pi23 & \pi24 ) | ( \pi23 & ~w102 ) | ( \pi24 & ~w102 ) ;
  assign w232 = w72 & ~w231 ;
  assign w233 = ( w227 & w229 ) | ( w227 & ~w230 ) | ( w229 & ~w230 ) ;
  assign w234 = w225 | w226 ;
  assign w235 = ( ~w226 & w230 ) | ( ~w226 & w232 ) | ( w230 & w232 ) ;
  assign w236 = w234 | w235 ;
  assign w237 = w233 | w236 ;
  assign w238 = ( w218 & w219 ) | ( w218 & ~w223 ) | ( w219 & ~w223 ) ;
  assign w239 = w222 | w237 ;
  assign w240 = ( w223 & w224 ) | ( w223 & ~w237 ) | ( w224 & ~w237 ) ;
  assign w241 = w239 | w240 ;
  assign w242 = w238 | w241 ;
  assign w243 = w205 | w206 ;
  assign w244 = w212 | w243 ;
  assign w245 = ( ~w212 & w216 ) | ( ~w212 & w242 ) | ( w216 & w242 ) ;
  assign w246 = w244 | w245 ;
  assign w247 = w199 | w201 ;
  assign w248 = w204 | w247 ;
  assign w249 = ( w198 & ~w204 ) | ( w198 & w246 ) | ( ~w204 & w246 ) ;
  assign w250 = w248 | w249 ;
  assign w251 = w38 & w99 ;
  assign w252 = w43 & w251 ;
  assign w253 = w47 & ~w53 ;
  assign w254 = w100 & w174 ;
  assign w255 = w94 & w97 ;
  assign w256 = w100 & w112 ;
  assign w257 = w78 & w83 ;
  assign w258 = w75 & w100 ;
  assign w259 = w61 & w130 ;
  assign w260 = w102 & w132 ;
  assign w261 = ( \pi23 & ~\pi24 ) | ( \pi23 & w80 ) | ( ~\pi24 & w80 ) ;
  assign w262 = w66 & w261 ;
  assign w263 = w61 & w102 ;
  assign w264 = w262 | w263 ;
  assign w265 = ~w62 & w100 ;
  assign w266 = w102 & w117 ;
  assign w267 = w265 | w266 ;
  assign w268 = w100 & w137 ;
  assign w269 = w55 & w58 ;
  assign w270 = w268 | w269 ;
  assign w271 = w58 & w102 ;
  assign w272 = w61 & w71 ;
  assign w273 = w271 | w272 ;
  assign w274 = w71 & w100 ;
  assign w275 = w47 & w132 ;
  assign w276 = w274 | w275 ;
  assign w277 = w91 & w130 ;
  assign w278 = w58 & w137 ;
  assign w279 = w277 | w278 ;
  assign w280 = ~w62 & w148 ;
  assign w281 = w83 & w100 ;
  assign w282 = w280 | w281 ;
  assign w283 = w75 & w148 ;
  assign w284 = w55 & w91 ;
  assign w285 = ~w53 & w130 ;
  assign w286 = w71 & w251 ;
  assign w287 = w97 & w251 ;
  assign w288 = ( w285 & ~w286 ) | ( w285 & w287 ) | ( ~w286 & w287 ) ;
  assign w289 = w286 | w288 ;
  assign w290 = ( w282 & ~w283 ) | ( w282 & w289 ) | ( ~w283 & w289 ) ;
  assign w291 = w276 | w279 ;
  assign w292 = ( ~w279 & w283 ) | ( ~w279 & w284 ) | ( w283 & w284 ) ;
  assign w293 = w291 | w292 ;
  assign w294 = w290 | w293 ;
  assign w295 = w267 | w273 ;
  assign w296 = ( ~w267 & w270 ) | ( ~w267 & w294 ) | ( w270 & w294 ) ;
  assign w297 = w295 | w296 ;
  assign w298 = ( w257 & w258 ) | ( w257 & ~w259 ) | ( w258 & ~w259 ) ;
  assign w299 = w264 | w297 ;
  assign w300 = ( w259 & w260 ) | ( w259 & ~w264 ) | ( w260 & ~w264 ) ;
  assign w301 = w299 | w300 ;
  assign w302 = w298 | w301 ;
  assign w303 = ( w253 & w254 ) | ( w253 & ~w255 ) | ( w254 & ~w255 ) ;
  assign w304 = w252 | w302 ;
  assign w305 = ( ~w252 & w255 ) | ( ~w252 & w256 ) | ( w255 & w256 ) ;
  assign w306 = w304 | w305 ;
  assign w307 = w303 | w306 ;
  assign w308 = ( \pi23 & ~\pi24 ) | ( \pi23 & w47 ) | ( ~\pi24 & w47 ) ;
  assign w309 = w66 & w308 ;
  assign w310 = w55 & w132 ;
  assign w311 = w132 & w145 ;
  assign w312 = ~w53 & w80 ;
  assign w313 = w40 & w102 ;
  assign w314 = w58 & w123 ;
  assign w315 = w132 & w137 ;
  assign w316 = w130 & w251 ;
  assign w317 = w145 & w148 ;
  assign w318 = w58 & w80 ;
  assign w319 = ( \pi23 & ~\pi24 ) | ( \pi23 & w43 ) | ( ~\pi24 & w43 ) ;
  assign w320 = w66 & w319 ;
  assign w321 = ( \pi23 & \pi24 ) | ( \pi23 & w174 ) | ( \pi24 & w174 ) ;
  assign w322 = w49 & w321 ;
  assign w323 = ( \pi23 & ~\pi24 ) | ( \pi23 & w145 ) | ( ~\pi24 & w145 ) ;
  assign w324 = w66 & w323 ;
  assign w325 = w78 & w130 ;
  assign w326 = w324 | w325 ;
  assign w327 = w320 | w322 ;
  assign w328 = w317 | w327 ;
  assign w329 = ( ~w317 & w318 ) | ( ~w317 & w326 ) | ( w318 & w326 ) ;
  assign w330 = w328 | w329 ;
  assign w331 = ( w313 & w314 ) | ( w313 & ~w315 ) | ( w314 & ~w315 ) ;
  assign w332 = w312 | w330 ;
  assign w333 = ( ~w312 & w315 ) | ( ~w312 & w316 ) | ( w315 & w316 ) ;
  assign w334 = w332 | w333 ;
  assign w335 = w331 | w334 ;
  assign w336 = w309 | w311 ;
  assign w337 = ( ~w309 & w310 ) | ( ~w309 & w335 ) | ( w310 & w335 ) ;
  assign w338 = w336 | w337 ;
  assign w339 = w89 & w145 ;
  assign w340 = w102 & w148 ;
  assign w341 = w91 & w102 ;
  assign w342 = w102 & w251 ;
  assign w343 = w341 | w342 ;
  assign w344 = w55 & w251 ;
  assign w345 = w47 & w251 ;
  assign w346 = w344 | w345 ;
  assign w347 = w339 | w346 ;
  assign w348 = ( ~w339 & w340 ) | ( ~w339 & w343 ) | ( w340 & w343 ) ;
  assign w349 = w347 | w348 ;
  assign w350 = w43 & w58 ;
  assign w351 = w75 & w132 ;
  assign w352 = w61 & w174 ;
  assign w353 = w71 & w78 ;
  assign w354 = ~w62 & w78 ;
  assign w355 = ( w352 & ~w353 ) | ( w352 & w354 ) | ( ~w353 & w354 ) ;
  assign w356 = w353 | w355 ;
  assign w357 = ( \pi23 & \pi24 ) | ( \pi23 & w130 ) | ( \pi24 & w130 ) ;
  assign w358 = w49 & w357 ;
  assign w359 = w53 | w62 ;
  assign w360 = ~w358 & w359 ;
  assign w361 = w55 & w61 ;
  assign w362 = w40 & w97 ;
  assign w363 = ( w350 & w351 ) | ( w350 & ~w361 ) | ( w351 & ~w361 ) ;
  assign w364 = ~w356 & w360 ;
  assign w365 = ( w360 & w361 ) | ( w360 & w362 ) | ( w361 & w362 ) ;
  assign w366 = w364 & ~w365 ;
  assign w367 = ~w363 & w366 ;
  assign w368 = ( w250 & w338 ) | ( w250 & ~w349 ) | ( w338 & ~w349 ) ;
  assign w369 = w196 | w307 ;
  assign w370 = ( w307 & ~w349 ) | ( w307 & w367 ) | ( ~w349 & w367 ) ;
  assign w371 = ~w369 & w370 ;
  assign w372 = ~w368 & w371 ;
  assign w373 = ( ~w68 & w82 ) | ( ~w68 & w87 ) | ( w82 & w87 ) ;
  assign w374 = ~w110 & w372 ;
  assign w375 = ( w68 & w74 ) | ( w68 & ~w110 ) | ( w74 & ~w110 ) ;
  assign w376 = w374 & ~w375 ;
  assign w377 = ~w373 & w376 ;
  assign w378 = w51 | w56 ;
  assign w379 = w64 | w378 ;
  assign w380 = ( ~w44 & w64 ) | ( ~w44 & w377 ) | ( w64 & w377 ) ;
  assign w381 = ~w379 & w380 ;
  assign w382 = ( \pi23 & \pi24 ) | ( \pi23 & w97 ) | ( \pi24 & w97 ) ;
  assign w383 = w49 & w382 ;
  assign w384 = w91 & w97 ;
  assign w385 = w55 & w78 ;
  assign w386 = w40 & w71 ;
  assign w387 = ( \pi23 & \pi24 ) | ( \pi23 & ~w75 ) | ( \pi24 & ~w75 ) ;
  assign w388 = w72 & ~w387 ;
  assign w389 = w100 & w123 ;
  assign w390 = ~w53 & w71 ;
  assign w391 = ( \pi23 & ~\pi24 ) | ( \pi23 & w71 ) | ( ~\pi24 & w71 ) ;
  assign w392 = w66 & w391 ;
  assign w393 = w71 & w117 ;
  assign w394 = w392 | w393 ;
  assign w395 = w362 | w394 ;
  assign w396 = ( w318 & ~w362 ) | ( w318 & w390 ) | ( ~w362 & w390 ) ;
  assign w397 = w395 | w396 ;
  assign w398 = ( w149 & w311 ) | ( w149 & ~w388 ) | ( w311 & ~w388 ) ;
  assign w399 = w76 | w397 ;
  assign w400 = ( ~w76 & w388 ) | ( ~w76 & w389 ) | ( w388 & w389 ) ;
  assign w401 = w399 | w400 ;
  assign w402 = w398 | w401 ;
  assign w403 = ( w281 & w309 ) | ( w281 & ~w385 ) | ( w309 & ~w385 ) ;
  assign w404 = w275 | w402 ;
  assign w405 = ( ~w275 & w385 ) | ( ~w275 & w386 ) | ( w385 & w386 ) ;
  assign w406 = w404 | w405 ;
  assign w407 = w403 | w406 ;
  assign w408 = w40 & w55 ;
  assign w409 = w83 & w89 ;
  assign w410 = w351 | w409 ;
  assign w411 = w61 & w83 ;
  assign w412 = ( \pi23 & \pi24 ) | ( \pi23 & ~w123 ) | ( \pi24 & ~w123 ) ;
  assign w413 = w72 & ~w412 ;
  assign w414 = w411 | w413 ;
  assign w415 = ~w62 & w117 ;
  assign w416 = w115 | w415 ;
  assign w417 = ( \pi23 & ~\pi24 ) | ( \pi23 & w112 ) | ( ~\pi24 & w112 ) ;
  assign w418 = w66 & w417 ;
  assign w419 = w137 & w251 ;
  assign w420 = w80 & w117 ;
  assign w421 = w75 & w117 ;
  assign w422 = w43 & w148 ;
  assign w423 = w43 & w117 ;
  assign w424 = w117 & w137 ;
  assign w425 = w423 | w424 ;
  assign w426 = w176 | w425 ;
  assign w427 = ( w113 & ~w176 ) | ( w113 & w422 ) | ( ~w176 & w422 ) ;
  assign w428 = w426 | w427 ;
  assign w429 = w83 & w251 ;
  assign w430 = w130 & w148 ;
  assign w431 = ~w53 & w137 ;
  assign w432 = w358 | w431 ;
  assign w433 = ( w169 & w421 ) | ( w169 & ~w429 ) | ( w421 & ~w429 ) ;
  assign w434 = w428 | w432 ;
  assign w435 = ( w429 & w430 ) | ( w429 & ~w432 ) | ( w430 & ~w432 ) ;
  assign w436 = w434 | w435 ;
  assign w437 = w433 | w436 ;
  assign w438 = ( w353 & w418 ) | ( w353 & ~w419 ) | ( w418 & ~w419 ) ;
  assign w439 = w262 | w437 ;
  assign w440 = ( ~w262 & w419 ) | ( ~w262 & w420 ) | ( w419 & w420 ) ;
  assign w441 = w439 | w440 ;
  assign w442 = w438 | w441 ;
  assign w443 = w43 & w89 ;
  assign w444 = w253 | w443 ;
  assign w445 = w174 & w251 ;
  assign w446 = ( \pi23 & \pi24 ) | ( \pi23 & ~w62 ) | ( \pi24 & ~w62 ) ;
  assign w447 = w49 & w446 ;
  assign w448 = ( ~\pi23 & \pi24 ) | ( ~\pi23 & w62 ) | ( \pi24 & w62 ) ;
  assign w449 = w66 & ~w448 ;
  assign w450 = w447 | w449 ;
  assign w451 = ( w268 & w271 ) | ( w268 & ~w274 ) | ( w271 & ~w274 ) ;
  assign w452 = w202 | w450 ;
  assign w453 = ( ~w202 & w274 ) | ( ~w202 & w445 ) | ( w274 & w445 ) ;
  assign w454 = w452 | w453 ;
  assign w455 = w451 | w454 ;
  assign w456 = w71 & w148 ;
  assign w457 = ( \pi23 & \pi24 ) | ( \pi23 & w71 ) | ( \pi24 & w71 ) ;
  assign w458 = w49 & w457 ;
  assign w459 = w117 & w123 ;
  assign w460 = w456 | w459 ;
  assign w461 = ( w265 & ~w456 ) | ( w265 & w458 ) | ( ~w456 & w458 ) ;
  assign w462 = w460 | w461 ;
  assign w463 = w61 & w112 ;
  assign w464 = ( \pi23 & \pi24 ) | ( \pi23 & ~w97 ) | ( \pi24 & ~w97 ) ;
  assign w465 = w72 & ~w464 ;
  assign w466 = w58 & w75 ;
  assign w467 = w58 & w174 ;
  assign w468 = w352 | w467 ;
  assign w469 = ( \pi23 & ~\pi24 ) | ( \pi23 & w130 ) | ( ~\pi24 & w130 ) ;
  assign w470 = w66 & w469 ;
  assign w471 = w466 | w470 ;
  assign w472 = w161 | w471 ;
  assign w473 = ( ~w161 & w465 ) | ( ~w161 & w468 ) | ( w465 & w468 ) ;
  assign w474 = w472 | w473 ;
  assign w475 = ( ~w210 & w444 ) | ( ~w210 & w462 ) | ( w444 & w462 ) ;
  assign w476 = w455 | w474 ;
  assign w477 = ( w210 & w463 ) | ( w210 & ~w474 ) | ( w463 & ~w474 ) ;
  assign w478 = w476 | w477 ;
  assign w479 = w475 | w478 ;
  assign w480 = w414 | w416 ;
  assign w481 = w479 | w480 ;
  assign w482 = ( w129 & w442 ) | ( w129 & ~w479 ) | ( w442 & ~w479 ) ;
  assign w483 = w481 | w482 ;
  assign w484 = w320 | w408 ;
  assign w485 = w410 | w484 ;
  assign w486 = ( w230 & ~w410 ) | ( w230 & w483 ) | ( ~w410 & w483 ) ;
  assign w487 = w485 | w486 ;
  assign w488 = w47 & w148 ;
  assign w489 = ( \pi23 & \pi24 ) | ( \pi23 & ~w55 ) | ( \pi24 & ~w55 ) ;
  assign w490 = w72 & ~w489 ;
  assign w491 = w137 & w148 ;
  assign w492 = w97 & w148 ;
  assign w493 = w138 | w492 ;
  assign w494 = ( \pi23 & \pi24 ) | ( \pi23 & w145 ) | ( \pi24 & w145 ) ;
  assign w495 = w49 & w494 ;
  assign w496 = w40 & w137 ;
  assign w497 = w495 | w496 ;
  assign w498 = w163 | w497 ;
  assign w499 = ( ~w163 & w220 ) | ( ~w163 & w493 ) | ( w220 & w493 ) ;
  assign w500 = w498 | w499 ;
  assign w501 = w208 | w491 ;
  assign w502 = ( ~w208 & w272 ) | ( ~w208 & w500 ) | ( w272 & w500 ) ;
  assign w503 = w501 | w502 ;
  assign w504 = w112 & w132 ;
  assign w505 = w61 & w137 ;
  assign w506 = w61 & w145 ;
  assign w507 = w44 | w506 ;
  assign w508 = ( \pi23 & ~\pi24 ) | ( \pi23 & w123 ) | ( ~\pi24 & w123 ) ;
  assign w509 = w66 & w508 ;
  assign w510 = w103 | w509 ;
  assign w511 = w80 & w251 ;
  assign w512 = w71 & w91 ;
  assign w513 = w145 & w251 ;
  assign w514 = w287 | w344 ;
  assign w515 = w61 & w123 ;
  assign w516 = w89 & w130 ;
  assign w517 = w515 | w516 ;
  assign w518 = w316 | w513 ;
  assign w519 = w517 | w518 ;
  assign w520 = ( w131 & w514 ) | ( w131 & ~w517 ) | ( w514 & ~w517 ) ;
  assign w521 = w519 | w520 ;
  assign w522 = ( ~w256 & w512 ) | ( ~w256 & w521 ) | ( w512 & w521 ) ;
  assign w523 = w256 | w522 ;
  assign w524 = w130 & w132 ;
  assign w525 = w71 & w89 ;
  assign w526 = ( w81 & ~w286 ) | ( w81 & w525 ) | ( ~w286 & w525 ) ;
  assign w527 = w286 | w526 ;
  assign w528 = w95 | w199 ;
  assign w529 = ( \pi23 & ~\pi24 ) | ( \pi23 & w174 ) | ( ~\pi24 & w174 ) ;
  assign w530 = w66 & w529 ;
  assign w531 = w117 & w130 ;
  assign w532 = w325 | w531 ;
  assign w533 = w40 & ~w62 ;
  assign w534 = ~w62 & w89 ;
  assign w535 = ( w354 & ~w533 ) | ( w354 & w534 ) | ( ~w533 & w534 ) ;
  assign w536 = w533 | w535 ;
  assign w537 = ( w280 & w322 ) | ( w280 & ~w345 ) | ( w322 & ~w345 ) ;
  assign w538 = w532 | w536 ;
  assign w539 = ( w345 & w530 ) | ( w345 & ~w536 ) | ( w530 & ~w536 ) ;
  assign w540 = w538 | w539 ;
  assign w541 = w537 | w540 ;
  assign w542 = ( ~w254 & w527 ) | ( ~w254 & w528 ) | ( w527 & w528 ) ;
  assign w543 = w523 | w541 ;
  assign w544 = ( w254 & w524 ) | ( w254 & ~w541 ) | ( w524 & ~w541 ) ;
  assign w545 = w543 | w544 ;
  assign w546 = w542 | w545 ;
  assign w547 = w510 | w511 ;
  assign w548 = ( w225 & ~w510 ) | ( w225 & w546 ) | ( ~w510 & w546 ) ;
  assign w549 = w547 | w548 ;
  assign w550 = ( w68 & w74 ) | ( w68 & ~w257 ) | ( w74 & ~w257 ) ;
  assign w551 = w507 | w549 ;
  assign w552 = ( w257 & w317 ) | ( w257 & ~w507 ) | ( w317 & ~w507 ) ;
  assign w553 = w551 | w552 ;
  assign w554 = w550 | w553 ;
  assign w555 = ( w141 & w223 ) | ( w141 & ~w504 ) | ( w223 & ~w504 ) ;
  assign w556 = w116 | w554 ;
  assign w557 = ( ~w116 & w504 ) | ( ~w116 & w505 ) | ( w504 & w505 ) ;
  assign w558 = w556 | w557 ;
  assign w559 = w555 | w558 ;
  assign w560 = ~w53 & w102 ;
  assign w561 = ~w53 & w75 ;
  assign w562 = w259 | w561 ;
  assign w563 = ( w203 & ~w259 ) | ( w203 & w560 ) | ( ~w259 & w560 ) ;
  assign w564 = w562 | w563 ;
  assign w565 = w43 & w132 ;
  assign w566 = ( \pi23 & \pi24 ) | ( \pi23 & w137 ) | ( \pi24 & w137 ) ;
  assign w567 = w49 & w566 ;
  assign w568 = w40 & w130 ;
  assign w569 = ~w62 & w251 ;
  assign w570 = w89 & w137 ;
  assign w571 = w47 & w89 ;
  assign w572 = w570 | w571 ;
  assign w573 = ~w53 & w145 ;
  assign w574 = ( ~w569 & w572 ) | ( ~w569 & w573 ) | ( w572 & w573 ) ;
  assign w575 = w569 | w574 ;
  assign w576 = w567 | w568 ;
  assign w577 = w564 | w576 ;
  assign w578 = ( ~w564 & w565 ) | ( ~w564 & w575 ) | ( w565 & w575 ) ;
  assign w579 = w577 | w578 ;
  assign w580 = ( ~w488 & w503 ) | ( ~w488 & w579 ) | ( w503 & w579 ) ;
  assign w581 = w487 | w559 ;
  assign w582 = ( ~w487 & w488 ) | ( ~w487 & w490 ) | ( w488 & w490 ) ;
  assign w583 = w581 | w582 ;
  assign w584 = w580 | w583 ;
  assign w585 = ( w122 & w168 ) | ( w122 & ~w221 ) | ( w168 & ~w221 ) ;
  assign w586 = w407 | w584 ;
  assign w587 = ( w221 & w284 ) | ( w221 & ~w407 ) | ( w284 & ~w407 ) ;
  assign w588 = w586 | w587 ;
  assign w589 = w585 | w588 ;
  assign w590 = w226 | w384 ;
  assign w591 = ( ~w226 & w383 ) | ( ~w226 & w589 ) | ( w383 & w589 ) ;
  assign w592 = w590 | w591 ;
  assign w593 = w61 & w97 ;
  assign w594 = w161 | w198 ;
  assign w595 = w91 & w174 ;
  assign w596 = w83 & w94 ;
  assign w597 = ( w179 & w205 ) | ( w179 & ~w595 ) | ( w205 & ~w595 ) ;
  assign w598 = w104 | w149 ;
  assign w599 = ( ~w149 & w595 ) | ( ~w149 & w596 ) | ( w595 & w596 ) ;
  assign w600 = w598 | w599 ;
  assign w601 = w597 | w600 ;
  assign w602 = ( ~w86 & w384 ) | ( ~w86 & w601 ) | ( w384 & w601 ) ;
  assign w603 = w86 | w602 ;
  assign w604 = ( \pi23 & \pi24 ) | ( \pi23 & ~w112 ) | ( \pi24 & ~w112 ) ;
  assign w605 = w72 & ~w604 ;
  assign w606 = w80 & w132 ;
  assign w607 = ( \pi23 & ~\pi24 ) | ( \pi23 & w97 ) | ( ~\pi24 & w97 ) ;
  assign w608 = w66 & w607 ;
  assign w609 = w492 | w608 ;
  assign w610 = w345 | w606 ;
  assign w611 = w281 | w610 ;
  assign w612 = ( ~w281 & w344 ) | ( ~w281 & w609 ) | ( w344 & w609 ) ;
  assign w613 = w611 | w612 ;
  assign w614 = ( w221 & w383 ) | ( w221 & ~w467 ) | ( w383 & ~w467 ) ;
  assign w615 = w74 | w613 ;
  assign w616 = ( ~w74 & w467 ) | ( ~w74 & w605 ) | ( w467 & w605 ) ;
  assign w617 = w615 | w616 ;
  assign w618 = w614 | w617 ;
  assign w619 = ( ~w254 & w325 ) | ( ~w254 & w618 ) | ( w325 & w618 ) ;
  assign w620 = w254 | w619 ;
  assign w621 = ( w206 & ~w361 ) | ( w206 & w362 ) | ( ~w361 & w362 ) ;
  assign w622 = w361 | w621 ;
  assign w623 = w75 & w251 ;
  assign w624 = w143 | w623 ;
  assign w625 = w91 & w145 ;
  assign w626 = w100 & w102 ;
  assign w627 = w625 | w626 ;
  assign w628 = w132 & w174 ;
  assign w629 = ( w122 & w135 ) | ( w122 & ~w225 ) | ( w135 & ~w225 ) ;
  assign w630 = w103 | w119 ;
  assign w631 = ( ~w119 & w225 ) | ( ~w119 & w318 ) | ( w225 & w318 ) ;
  assign w632 = w630 | w631 ;
  assign w633 = w629 | w632 ;
  assign w634 = w51 | w628 ;
  assign w635 = ( ~w51 & w531 ) | ( ~w51 & w633 ) | ( w531 & w633 ) ;
  assign w636 = w634 | w635 ;
  assign w637 = w43 & w94 ;
  assign w638 = w418 | w637 ;
  assign w639 = ( \pi23 & ~\pi24 ) | ( \pi23 & w83 ) | ( ~\pi24 & w83 ) ;
  assign w640 = w66 & w639 ;
  assign w641 = w55 & w94 ;
  assign w642 = w40 & w80 ;
  assign w643 = ( w573 & w640 ) | ( w573 & ~w641 ) | ( w640 & ~w641 ) ;
  assign w644 = w491 | w505 ;
  assign w645 = ( ~w505 & w641 ) | ( ~w505 & w642 ) | ( w641 & w642 ) ;
  assign w646 = w644 | w645 ;
  assign w647 = w643 | w646 ;
  assign w648 = w390 | w647 ;
  assign w649 = ( w124 & w638 ) | ( w124 & ~w647 ) | ( w638 & ~w647 ) ;
  assign w650 = w648 | w649 ;
  assign w651 = w220 | w650 ;
  assign w652 = ( w68 & w636 ) | ( w68 & ~w650 ) | ( w636 & ~w650 ) ;
  assign w653 = w651 | w652 ;
  assign w654 = w524 | w627 ;
  assign w655 = ( w147 & ~w627 ) | ( w147 & w653 ) | ( ~w627 & w653 ) ;
  assign w656 = w654 | w655 ;
  assign w657 = w199 | w389 ;
  assign w658 = w624 | w657 ;
  assign w659 = ( w118 & ~w624 ) | ( w118 & w656 ) | ( ~w624 & w656 ) ;
  assign w660 = w658 | w659 ;
  assign w661 = w90 | w92 ;
  assign w662 = w43 & w78 ;
  assign w663 = w58 & w145 ;
  assign w664 = w78 & w174 ;
  assign w665 = ( w421 & w447 ) | ( w421 & ~w663 ) | ( w447 & ~w663 ) ;
  assign w666 = w340 | w420 ;
  assign w667 = ( ~w420 & w663 ) | ( ~w420 & w664 ) | ( w663 & w664 ) ;
  assign w668 = w666 | w667 ;
  assign w669 = w665 | w668 ;
  assign w670 = ( ~w274 & w662 ) | ( ~w274 & w669 ) | ( w662 & w669 ) ;
  assign w671 = w274 | w670 ;
  assign w672 = w265 | w569 ;
  assign w673 = w47 & w61 ;
  assign w674 = w123 & w132 ;
  assign w675 = w673 | w674 ;
  assign w676 = w424 | w675 ;
  assign w677 = ( w263 & ~w424 ) | ( w263 & w516 ) | ( ~w424 & w516 ) ;
  assign w678 = w676 | w677 ;
  assign w679 = ( \pi23 & \pi24 ) | ( \pi23 & ~w130 ) | ( \pi24 & ~w130 ) ;
  assign w680 = w72 & ~w679 ;
  assign w681 = w112 & w251 ;
  assign w682 = ( w113 & w570 ) | ( w113 & ~w680 ) | ( w570 & ~w680 ) ;
  assign w683 = w672 | w678 ;
  assign w684 = ( ~w678 & w680 ) | ( ~w678 & w681 ) | ( w680 & w681 ) ;
  assign w685 = w683 | w684 ;
  assign w686 = w682 | w685 ;
  assign w687 = w661 | w686 ;
  assign w688 = ( w444 & w671 ) | ( w444 & ~w686 ) | ( w671 & ~w686 ) ;
  assign w689 = w687 | w688 ;
  assign w690 = ( w411 & w415 ) | ( w411 & ~w458 ) | ( w415 & ~w458 ) ;
  assign w691 = w314 | w689 ;
  assign w692 = ( ~w314 & w458 ) | ( ~w314 & w525 ) | ( w458 & w525 ) ;
  assign w693 = w691 | w692 ;
  assign w694 = w690 | w693 ;
  assign w695 = ( ~w142 & w565 ) | ( ~w142 & w694 ) | ( w565 & w694 ) ;
  assign w696 = w142 | w695 ;
  assign w697 = w78 & w112 ;
  assign w698 = w313 | w324 ;
  assign w699 = ( w230 & w413 ) | ( w230 & ~w465 ) | ( w413 & ~w465 ) ;
  assign w700 = w114 | w698 ;
  assign w701 = ( ~w114 & w465 ) | ( ~w114 & w533 ) | ( w465 & w533 ) ;
  assign w702 = w700 | w701 ;
  assign w703 = w699 | w702 ;
  assign w704 = ( ~w164 & w622 ) | ( ~w164 & w703 ) | ( w622 & w703 ) ;
  assign w705 = w660 | w696 ;
  assign w706 = ( w164 & ~w696 ) | ( w164 & w697 ) | ( ~w696 & w697 ) ;
  assign w707 = w705 | w706 ;
  assign w708 = w704 | w707 ;
  assign w709 = w315 | w316 ;
  assign w710 = w120 | w709 ;
  assign w711 = ( ~w120 & w311 ) | ( ~w120 & w708 ) | ( w311 & w708 ) ;
  assign w712 = w710 | w711 ;
  assign w713 = ( ~w169 & w177 ) | ( ~w169 & w603 ) | ( w177 & w603 ) ;
  assign w714 = w620 | w712 ;
  assign w715 = ( w169 & w490 ) | ( w169 & ~w620 ) | ( w490 & ~w620 ) ;
  assign w716 = w714 | w715 ;
  assign w717 = w713 | w716 ;
  assign w718 = w513 | w593 ;
  assign w719 = w594 | w718 ;
  assign w720 = ( w310 & ~w594 ) | ( w310 & w717 ) | ( ~w594 & w717 ) ;
  assign w721 = w719 | w720 ;
  assign w722 = w40 & w174 ;
  assign w723 = w89 & w102 ;
  assign w724 = w94 & w112 ;
  assign w725 = w55 & w100 ;
  assign w726 = w78 & w137 ;
  assign w727 = w459 | w726 ;
  assign w728 = w104 | w727 ;
  assign w729 = ( w103 & ~w104 ) | ( w103 & w353 ) | ( ~w104 & w353 ) ;
  assign w730 = w728 | w729 ;
  assign w731 = w135 | w227 ;
  assign w732 = ( w342 & w361 ) | ( w342 & ~w456 ) | ( w361 & ~w456 ) ;
  assign w733 = w116 | w125 ;
  assign w734 = ( ~w125 & w456 ) | ( ~w125 & w466 ) | ( w456 & w466 ) ;
  assign w735 = w733 | w734 ;
  assign w736 = w732 | w735 ;
  assign w737 = ( w268 & w322 ) | ( w268 & ~w383 ) | ( w322 & ~w383 ) ;
  assign w738 = w115 | w736 ;
  assign w739 = ( ~w115 & w383 ) | ( ~w115 & w569 ) | ( w383 & w569 ) ;
  assign w740 = w738 | w739 ;
  assign w741 = w737 | w740 ;
  assign w742 = w114 | w573 ;
  assign w743 = w533 | w663 ;
  assign w744 = w144 | w743 ;
  assign w745 = ( w128 & ~w144 ) | ( w128 & w516 ) | ( ~w144 & w516 ) ;
  assign w746 = w744 | w745 ;
  assign w747 = ( w271 & w286 ) | ( w271 & ~w358 ) | ( w286 & ~w358 ) ;
  assign w748 = w220 | w746 ;
  assign w749 = ( ~w220 & w358 ) | ( ~w220 & w470 ) | ( w358 & w470 ) ;
  assign w750 = w748 | w749 ;
  assign w751 = w747 | w750 ;
  assign w752 = ( w225 & w350 ) | ( w225 & ~w384 ) | ( w350 & ~w384 ) ;
  assign w753 = w59 | w751 ;
  assign w754 = ( ~w59 & w384 ) | ( ~w59 & w449 ) | ( w384 & w449 ) ;
  assign w755 = w753 | w754 ;
  assign w756 = w752 | w755 ;
  assign w757 = ( \pi23 & ~\pi24 ) | ( \pi23 & w75 ) | ( ~\pi24 & w75 ) ;
  assign w758 = w66 & w757 ;
  assign w759 = w180 | w284 ;
  assign w760 = w595 | w758 ;
  assign w761 = w63 | w760 ;
  assign w762 = ( ~w63 & w419 ) | ( ~w63 & w759 ) | ( w419 & w759 ) ;
  assign w763 = w761 | w762 ;
  assign w764 = w91 & w123 ;
  assign w765 = w215 | w490 ;
  assign w766 = ( w168 & ~w215 ) | ( w168 & w285 ) | ( ~w215 & w285 ) ;
  assign w767 = w765 | w766 ;
  assign w768 = ( w124 & ~w567 ) | ( w124 & w767 ) | ( ~w567 & w767 ) ;
  assign w769 = w756 | w763 ;
  assign w770 = ( w567 & ~w763 ) | ( w567 & w764 ) | ( ~w763 & w764 ) ;
  assign w771 = w769 | w770 ;
  assign w772 = w768 | w771 ;
  assign w773 = ( w204 & w730 ) | ( w204 & ~w731 ) | ( w730 & ~w731 ) ;
  assign w774 = w741 | w772 ;
  assign w775 = ( w731 & ~w741 ) | ( w731 & w742 ) | ( ~w741 & w742 ) ;
  assign w776 = w774 | w775 ;
  assign w777 = w773 | w776 ;
  assign w778 = ( w178 & w423 ) | ( w178 & ~w724 ) | ( w423 & ~w724 ) ;
  assign w779 = w136 | w777 ;
  assign w780 = ( ~w136 & w724 ) | ( ~w136 & w725 ) | ( w724 & w725 ) ;
  assign w781 = w779 | w780 ;
  assign w782 = w778 | w781 ;
  assign w783 = w43 & ~w53 ;
  assign w784 = w164 | w219 ;
  assign w785 = w345 | w392 ;
  assign w786 = ( \pi23 & \pi24 ) | ( \pi23 & w55 ) | ( \pi24 & w55 ) ;
  assign w787 = w49 & w786 ;
  assign w788 = ( w320 & w351 ) | ( w320 & ~w421 ) | ( w351 & ~w421 ) ;
  assign w789 = w260 | w312 ;
  assign w790 = ( ~w312 & w421 ) | ( ~w312 & w787 ) | ( w421 & w787 ) ;
  assign w791 = w789 | w790 ;
  assign w792 = w788 | w791 ;
  assign w793 = w272 | w785 ;
  assign w794 = ( w784 & ~w785 ) | ( w784 & w792 ) | ( ~w785 & w792 ) ;
  assign w795 = w793 | w794 ;
  assign w796 = w359 & ~w408 ;
  assign w797 = ~w253 & w796 ;
  assign w798 = ( ~w253 & w344 ) | ( ~w253 & w795 ) | ( w344 & w795 ) ;
  assign w799 = w797 & ~w798 ;
  assign w800 = w393 | w512 ;
  assign w801 = ( \pi23 & \pi24 ) | ( \pi23 & w62 ) | ( \pi24 & w62 ) ;
  assign w802 = w72 & ~w801 ;
  assign w803 = w223 | w802 ;
  assign w804 = w131 | w803 ;
  assign w805 = ( ~w131 & w139 ) | ( ~w131 & w800 ) | ( w139 & w800 ) ;
  assign w806 = w804 | w805 ;
  assign w807 = ( w149 & w467 ) | ( w149 & ~w524 ) | ( w467 & ~w524 ) ;
  assign w808 = w147 | w806 ;
  assign w809 = ( ~w147 & w524 ) | ( ~w147 & w674 ) | ( w524 & w674 ) ;
  assign w810 = w808 | w809 ;
  assign w811 = w807 | w810 ;
  assign w812 = ( w259 & w386 ) | ( w259 & ~w443 ) | ( w386 & ~w443 ) ;
  assign w813 = w51 | w811 ;
  assign w814 = ( ~w51 & w443 ) | ( ~w51 & w492 ) | ( w443 & w492 ) ;
  assign w815 = w813 | w814 ;
  assign w816 = w812 | w815 ;
  assign w817 = w61 & w80 ;
  assign w818 = w362 | w491 ;
  assign w819 = ( w278 & ~w362 ) | ( w278 & w415 ) | ( ~w362 & w415 ) ;
  assign w820 = w818 | w819 ;
  assign w821 = w78 & w145 ;
  assign w822 = w424 | w821 ;
  assign w823 = ( w628 & w642 ) | ( w628 & ~w673 ) | ( w642 & ~w673 ) ;
  assign w824 = w141 | w626 ;
  assign w825 = ( ~w626 & w673 ) | ( ~w626 & w680 ) | ( w673 & w680 ) ;
  assign w826 = w824 | w825 ;
  assign w827 = w823 | w826 ;
  assign w828 = ( w118 & w119 ) | ( w118 & ~w266 ) | ( w119 & ~w266 ) ;
  assign w829 = w822 | w827 ;
  assign w830 = ( w266 & w409 ) | ( w266 & ~w827 ) | ( w409 & ~w827 ) ;
  assign w831 = w829 | w830 ;
  assign w832 = w828 | w831 ;
  assign w833 = w352 | w565 ;
  assign w834 = w205 | w833 ;
  assign w835 = ( ~w205 & w221 ) | ( ~w205 & w832 ) | ( w221 & w832 ) ;
  assign w836 = w834 | w835 ;
  assign w837 = w55 & w148 ;
  assign w838 = w277 | w568 ;
  assign w839 = w413 | w837 ;
  assign w840 = w88 | w839 ;
  assign w841 = ( ~w88 & w224 ) | ( ~w88 & w838 ) | ( w224 & w838 ) ;
  assign w842 = w840 | w841 ;
  assign w843 = ( w252 & w463 ) | ( w252 & ~w504 ) | ( w463 & ~w504 ) ;
  assign w844 = w210 | w842 ;
  assign w845 = ( ~w210 & w504 ) | ( ~w210 & w515 ) | ( w504 & w515 ) ;
  assign w846 = w844 | w845 ;
  assign w847 = w843 | w846 ;
  assign w848 = w495 | w513 ;
  assign w849 = w847 | w848 ;
  assign w850 = ( w820 & w836 ) | ( w820 & ~w847 ) | ( w836 & ~w847 ) ;
  assign w851 = w849 | w850 ;
  assign w852 = ( w310 & w509 ) | ( w310 & ~w511 ) | ( w509 & ~w511 ) ;
  assign w853 = w230 | w851 ;
  assign w854 = ( ~w230 & w511 ) | ( ~w230 & w560 ) | ( w511 & w560 ) ;
  assign w855 = w853 | w854 ;
  assign w856 = w852 | w855 ;
  assign w857 = w262 | w817 ;
  assign w858 = ( ~w262 & w531 ) | ( ~w262 & w856 ) | ( w531 & w856 ) ;
  assign w859 = w857 | w858 ;
  assign w860 = ~w53 & w123 ;
  assign w861 = w623 | w860 ;
  assign w862 = w340 | w861 ;
  assign w863 = ( w199 & ~w340 ) | ( w199 & w561 ) | ( ~w340 & w561 ) ;
  assign w864 = w862 | w863 ;
  assign w865 = ( w87 & w661 ) | ( w87 & ~w864 ) | ( w661 & ~w864 ) ;
  assign w866 = w816 | w859 ;
  assign w867 = ( w163 & ~w816 ) | ( w163 & w864 ) | ( ~w816 & w864 ) ;
  assign w868 = w866 | w867 ;
  assign w869 = w865 | w868 ;
  assign w870 = ( ~w445 & w723 ) | ( ~w445 & w799 ) | ( w723 & w799 ) ;
  assign w871 = w782 | w869 ;
  assign w872 = ( w723 & ~w782 ) | ( w723 & w783 ) | ( ~w782 & w783 ) ;
  assign w873 = w871 | w872 ;
  assign w874 = w870 & ~w873 ;
  assign w875 = ( w120 & w281 ) | ( w120 & ~w496 ) | ( w281 & ~w496 ) ;
  assign w876 = ~w111 & w874 ;
  assign w877 = ( ~w111 & w496 ) | ( ~w111 & w641 ) | ( w496 & w641 ) ;
  assign w878 = w876 & ~w877 ;
  assign w879 = ~w875 & w878 ;
  assign w880 = w488 | w722 ;
  assign w881 = w161 | w880 ;
  assign w882 = ( w161 & ~w465 ) | ( w161 & w879 ) | ( ~w465 & w879 ) ;
  assign w883 = ~w881 & w882 ;
  assign w884 = w230 | w787 ;
  assign w885 = ( w125 & ~w230 ) | ( w125 & w285 ) | ( ~w230 & w285 ) ;
  assign w886 = w884 | w885 ;
  assign w887 = w113 | w723 ;
  assign w888 = w214 | w254 ;
  assign w889 = w43 & w61 ;
  assign w890 = w314 | w725 ;
  assign w891 = w512 | w606 ;
  assign w892 = w179 | w891 ;
  assign w893 = ( ~w179 & w283 ) | ( ~w179 & w890 ) | ( w283 & w890 ) ;
  assign w894 = w892 | w893 ;
  assign w895 = ( ~w309 & w889 ) | ( ~w309 & w894 ) | ( w889 & w894 ) ;
  assign w896 = w309 | w895 ;
  assign w897 = w40 & w47 ;
  assign w898 = ( \pi23 & \pi24 ) | ( \pi23 & ~w83 ) | ( \pi24 & ~w83 ) ;
  assign w899 = w72 & ~w898 ;
  assign w900 = w51 | w278 ;
  assign w901 = w47 & w78 ;
  assign w902 = ( w496 & w565 ) | ( w496 & ~w596 ) | ( w565 & ~w596 ) ;
  assign w903 = w310 | w420 ;
  assign w904 = ( ~w420 & w596 ) | ( ~w420 & w640 ) | ( w596 & w640 ) ;
  assign w905 = w903 | w904 ;
  assign w906 = w902 | w905 ;
  assign w907 = w423 | w901 ;
  assign w908 = w409 | w907 ;
  assign w909 = ( ~w409 & w411 ) | ( ~w409 & w906 ) | ( w411 & w906 ) ;
  assign w910 = w908 | w909 ;
  assign w911 = w419 | w488 ;
  assign w912 = ( w322 & w341 ) | ( w322 & ~w383 ) | ( w341 & ~w383 ) ;
  assign w913 = w730 | w864 ;
  assign w914 = ( w383 & w421 ) | ( w383 & ~w864 ) | ( w421 & ~w864 ) ;
  assign w915 = w913 | w914 ;
  assign w916 = w912 | w915 ;
  assign w917 = ( ~w311 & w536 ) | ( ~w311 & w911 ) | ( w536 & w911 ) ;
  assign w918 = w96 | w916 ;
  assign w919 = ( ~w96 & w311 ) | ( ~w96 & w389 ) | ( w311 & w389 ) ;
  assign w920 = w918 | w919 ;
  assign w921 = w917 | w920 ;
  assign w922 = w900 | w910 ;
  assign w923 = ( w507 & ~w910 ) | ( w507 & w921 ) | ( ~w910 & w921 ) ;
  assign w924 = w922 | w923 ;
  assign w925 = ( w206 & w573 ) | ( w206 & ~w625 ) | ( w573 & ~w625 ) ;
  assign w926 = w572 | w924 ;
  assign w927 = ( ~w572 & w625 ) | ( ~w572 & w899 ) | ( w625 & w899 ) ;
  assign w928 = w926 | w927 ;
  assign w929 = w925 | w928 ;
  assign w930 = w837 | w897 ;
  assign w931 = w315 | w930 ;
  assign w932 = ( ~w315 & w422 ) | ( ~w315 & w929 ) | ( w422 & w929 ) ;
  assign w933 = w931 | w932 ;
  assign w934 = w169 | w637 ;
  assign w935 = ( w98 & ~w169 ) | ( w98 & w593 ) | ( ~w169 & w593 ) ;
  assign w936 = w934 | w935 ;
  assign w937 = w144 | w149 ;
  assign w938 = ( ~w144 & w147 ) | ( ~w144 & w936 ) | ( w147 & w936 ) ;
  assign w939 = w937 | w938 ;
  assign w940 = w318 | w783 ;
  assign w941 = w220 | w940 ;
  assign w942 = ( ~w220 & w232 ) | ( ~w220 & w939 ) | ( w232 & w939 ) ;
  assign w943 = w941 | w942 ;
  assign w944 = ( w312 & w385 ) | ( w312 & ~w458 ) | ( w385 & ~w458 ) ;
  assign w945 = w163 | w943 ;
  assign w946 = ( ~w163 & w458 ) | ( ~w163 & w821 ) | ( w458 & w821 ) ;
  assign w947 = w945 | w946 ;
  assign w948 = w944 | w947 ;
  assign w949 = ( ~w114 & w227 ) | ( ~w114 & w948 ) | ( w227 & w948 ) ;
  assign w950 = w114 | w949 ;
  assign w951 = ~w53 & w97 ;
  assign w952 = w430 | w951 ;
  assign w953 = w111 | w450 ;
  assign w954 = ( w212 & ~w450 ) | ( w212 & w952 ) | ( ~w450 & w952 ) ;
  assign w955 = w953 | w954 ;
  assign w956 = w86 | w431 ;
  assign w957 = w263 | w628 ;
  assign w958 = ( ~w263 & w339 ) | ( ~w263 & w956 ) | ( w339 & w956 ) ;
  assign w959 = w957 | w958 ;
  assign w960 = ( w116 & w161 ) | ( w116 & ~w277 ) | ( w161 & ~w277 ) ;
  assign w961 = w955 | w959 ;
  assign w962 = ( w277 & w470 ) | ( w277 & ~w959 ) | ( w470 & ~w959 ) ;
  assign w963 = w961 | w962 ;
  assign w964 = w960 | w963 ;
  assign w965 = ( ~w887 & w896 ) | ( ~w887 & w964 ) | ( w896 & w964 ) ;
  assign w966 = w933 | w950 ;
  assign w967 = ( w887 & w888 ) | ( w887 & ~w950 ) | ( w888 & ~w950 ) ;
  assign w968 = w966 | w967 ;
  assign w969 = w965 | w968 ;
  assign w970 = ( w201 & ~w221 ) | ( w201 & w886 ) | ( ~w221 & w886 ) ;
  assign w971 = w416 | w969 ;
  assign w972 = ( w221 & ~w416 ) | ( w221 & w758 ) | ( ~w416 & w758 ) ;
  assign w973 = w971 | w972 ;
  assign w974 = w970 | w973 ;
  assign w975 = ( w342 & w361 ) | ( w342 & ~w390 ) | ( w361 & ~w390 ) ;
  assign w976 = w128 | w974 ;
  assign w977 = ( ~w128 & w390 ) | ( ~w128 & w491 ) | ( w390 & w491 ) ;
  assign w978 = w976 | w977 ;
  assign w979 = w975 | w978 ;
  assign w980 = w58 & ~w62 ;
  assign w981 = ( w339 & w388 ) | ( w339 & ~w899 ) | ( w388 & ~w899 ) ;
  assign w982 = w76 | w230 ;
  assign w983 = ( ~w230 & w899 ) | ( ~w230 & w980 ) | ( w899 & w980 ) ;
  assign w984 = w982 | w983 ;
  assign w985 = w981 | w984 ;
  assign w986 = ( ~w68 & w219 ) | ( ~w68 & w985 ) | ( w219 & w985 ) ;
  assign w987 = w68 | w986 ;
  assign w988 = w44 | w320 ;
  assign w989 = w281 | w512 ;
  assign w990 = w136 | w989 ;
  assign w991 = ( ~w136 & w258 ) | ( ~w136 & w988 ) | ( w258 & w988 ) ;
  assign w992 = w990 | w991 ;
  assign w993 = w802 | w897 ;
  assign w994 = w488 | w993 ;
  assign w995 = ( ~w488 & w530 ) | ( ~w488 & w992 ) | ( w530 & w992 ) ;
  assign w996 = w994 | w995 ;
  assign w997 = w384 | w423 ;
  assign w998 = w310 | w641 ;
  assign w999 = w340 | w626 ;
  assign w1000 = ( \pi23 & \pi24 ) | ( \pi23 & ~w137 ) | ( \pi24 & ~w137 ) ;
  assign w1001 = w72 & ~w1000 ;
  assign w1002 = ( w178 & w268 ) | ( w178 & ~w324 ) | ( w268 & ~w324 ) ;
  assign w1003 = w84 | w514 ;
  assign w1004 = ( ~w84 & w324 ) | ( ~w84 & w352 ) | ( w324 & w352 ) ;
  assign w1005 = w1003 | w1004 ;
  assign w1006 = w1002 | w1005 ;
  assign w1007 = w144 | w1001 ;
  assign w1008 = ( ~w144 & w167 ) | ( ~w144 & w1006 ) | ( w167 & w1006 ) ;
  assign w1009 = w1007 | w1008 ;
  assign w1010 = w430 | w593 ;
  assign w1011 = ( w463 & w492 ) | ( w463 & ~w623 ) | ( w492 & ~w623 ) ;
  assign w1012 = w118 | w1010 ;
  assign w1013 = ( ~w118 & w623 ) | ( ~w118 & w837 ) | ( w623 & w837 ) ;
  assign w1014 = w1012 | w1013 ;
  assign w1015 = w1011 | w1014 ;
  assign w1016 = ( w216 & w276 ) | ( w216 & ~w510 ) | ( w276 & ~w510 ) ;
  assign w1017 = w1009 | w1015 ;
  assign w1018 = ( w510 & w999 ) | ( w510 & ~w1015 ) | ( w999 & ~w1015 ) ;
  assign w1019 = w1017 | w1018 ;
  assign w1020 = w1016 | w1019 ;
  assign w1021 = w758 | w998 ;
  assign w1022 = w204 | w1021 ;
  assign w1023 = ( ~w204 & w410 ) | ( ~w204 & w1020 ) | ( w410 & w1020 ) ;
  assign w1024 = w1022 | w1023 ;
  assign w1025 = ( w135 & w149 ) | ( w135 & ~w322 ) | ( w149 & ~w322 ) ;
  assign w1026 = w92 | w1024 ;
  assign w1027 = ( ~w92 & w322 ) | ( ~w92 & w697 ) | ( w322 & w697 ) ;
  assign w1028 = w1026 | w1027 ;
  assign w1029 = w1025 | w1028 ;
  assign w1030 = w100 & w130 ;
  assign w1031 = w78 & w123 ;
  assign w1032 = ( w429 & w680 ) | ( w429 & ~w951 ) | ( w680 & ~w951 ) ;
  assign w1033 = w390 | w421 ;
  assign w1034 = ( ~w421 & w951 ) | ( ~w421 & w1031 ) | ( w951 & w1031 ) ;
  assign w1035 = w1033 | w1034 ;
  assign w1036 = w1032 | w1035 ;
  assign w1037 = w628 | w1030 ;
  assign w1038 = w98 | w1037 ;
  assign w1039 = ( ~w98 & w568 ) | ( ~w98 & w1036 ) | ( w568 & w1036 ) ;
  assign w1040 = w1038 | w1039 ;
  assign w1041 = w226 | w490 ;
  assign w1042 = w201 | w1041 ;
  assign w1043 = ( w164 & ~w201 ) | ( w164 & w210 ) | ( ~w201 & w210 ) ;
  assign w1044 = w1042 | w1043 ;
  assign w1045 = ( w255 & w362 ) | ( w255 & ~w392 ) | ( w362 & ~w392 ) ;
  assign w1046 = w124 | w1044 ;
  assign w1047 = ( ~w124 & w392 ) | ( ~w124 & w393 ) | ( w392 & w393 ) ;
  assign w1048 = w1046 | w1047 ;
  assign w1049 = w1045 | w1048 ;
  assign w1050 = ( w113 & ~w424 ) | ( w113 & w817 ) | ( ~w424 & w817 ) ;
  assign w1051 = w424 | w1050 ;
  assign w1052 = w1049 | w1051 ;
  assign w1053 = ( w222 & w1040 ) | ( w222 & ~w1049 ) | ( w1040 & ~w1049 ) ;
  assign w1054 = w1052 | w1053 ;
  assign w1055 = w119 | w229 ;
  assign w1056 = w759 | w1055 ;
  assign w1057 = ( w90 & ~w759 ) | ( w90 & w1054 ) | ( ~w759 & w1054 ) ;
  assign w1058 = w1056 | w1057 ;
  assign w1059 = ( w227 & w408 ) | ( w227 & ~w415 ) | ( w408 & ~w415 ) ;
  assign w1060 = w111 | w1058 ;
  assign w1061 = ( ~w111 & w415 ) | ( ~w111 & w420 ) | ( w415 & w420 ) ;
  assign w1062 = w1060 | w1061 ;
  assign w1063 = w1059 | w1062 ;
  assign w1064 = w285 | w560 ;
  assign w1065 = w143 | w860 ;
  assign w1066 = w1064 | w1065 ;
  assign w1067 = ( w122 & w572 ) | ( w122 & ~w1064 ) | ( w572 & ~w1064 ) ;
  assign w1068 = w1066 | w1067 ;
  assign w1069 = w138 | w224 ;
  assign w1070 = ( ~w104 & w264 ) | ( ~w104 & w1069 ) | ( w264 & w1069 ) ;
  assign w1071 = w1063 | w1068 ;
  assign w1072 = ( w104 & w133 ) | ( w104 & ~w1068 ) | ( w133 & ~w1068 ) ;
  assign w1073 = w1071 | w1072 ;
  assign w1074 = w1070 | w1073 ;
  assign w1075 = w147 | w524 ;
  assign w1076 = w1074 | w1075 ;
  assign w1077 = ( w997 & w1029 ) | ( w997 & ~w1074 ) | ( w1029 & ~w1074 ) ;
  assign w1078 = w1076 | w1077 ;
  assign w1079 = w606 | w900 ;
  assign w1080 = w996 | w1079 ;
  assign w1081 = ( w987 & ~w996 ) | ( w987 & w1078 ) | ( ~w996 & w1078 ) ;
  assign w1082 = w1080 | w1081 ;
  assign w1083 = w127 | w506 ;
  assign w1084 = ( ~w127 & w419 ) | ( ~w127 & w1082 ) | ( w419 & w1082 ) ;
  assign w1085 = w1083 | w1084 ;
  assign w1086 = w100 & w145 ;
  assign w1087 = w149 | w408 ;
  assign w1088 = w411 | w1031 ;
  assign w1089 = ( w320 & w389 ) | ( w320 & ~w390 ) | ( w389 & ~w390 ) ;
  assign w1090 = w138 | w1088 ;
  assign w1091 = ( ~w138 & w390 ) | ( ~w138 & w889 ) | ( w390 & w889 ) ;
  assign w1092 = w1090 | w1091 ;
  assign w1093 = w1089 | w1092 ;
  assign w1094 = w75 & w91 ;
  assign w1095 = w125 | w1094 ;
  assign w1096 = w229 | w509 ;
  assign w1097 = w136 | w1096 ;
  assign w1098 = ( ~w136 & w215 ) | ( ~w136 & w1095 ) | ( w215 & w1095 ) ;
  assign w1099 = w1097 | w1098 ;
  assign w1100 = ( w118 & w144 ) | ( w118 & ~w283 ) | ( w144 & ~w283 ) ;
  assign w1101 = w74 | w1099 ;
  assign w1102 = ( ~w74 & w283 ) | ( ~w74 & w642 ) | ( w283 & w642 ) ;
  assign w1103 = w1101 | w1102 ;
  assign w1104 = w1100 | w1103 ;
  assign w1105 = w445 | w534 ;
  assign w1106 = w278 | w1105 ;
  assign w1107 = ( w163 & ~w278 ) | ( w163 & w415 ) | ( ~w278 & w415 ) ;
  assign w1108 = w1106 | w1107 ;
  assign w1109 = ( w230 & w232 ) | ( w230 & ~w256 ) | ( w232 & ~w256 ) ;
  assign w1110 = w1104 | w1108 ;
  assign w1111 = ( w256 & w530 ) | ( w256 & ~w1108 ) | ( w530 & ~w1108 ) ;
  assign w1112 = w1110 | w1111 ;
  assign w1113 = w1109 | w1112 ;
  assign w1114 = w1087 | w1093 ;
  assign w1115 = ( w129 & ~w1093 ) | ( w129 & w1113 ) | ( ~w1093 & w1113 ) ;
  assign w1116 = w1114 | w1115 ;
  assign w1117 = ( w81 & w280 ) | ( w81 & ~w593 ) | ( w280 & ~w593 ) ;
  assign w1118 = w572 | w1116 ;
  assign w1119 = ( ~w572 & w593 ) | ( ~w572 & w1086 ) | ( w593 & w1086 ) ;
  assign w1120 = w1118 | w1119 ;
  assign w1121 = w1117 | w1120 ;
  assign w1122 = w352 | w358 ;
  assign w1123 = w253 | w1122 ;
  assign w1124 = ( ~w253 & w325 ) | ( ~w253 & w1121 ) | ( w325 & w1121 ) ;
  assign w1125 = w1123 | w1124 ;
  assign w1126 = w117 & w145 ;
  assign w1127 = ( \pi23 & \pi24 ) | ( \pi23 & w80 ) | ( \pi24 & w80 ) ;
  assign w1128 = w49 & w1127 ;
  assign w1129 = w463 | w1128 ;
  assign w1130 = w89 & w174 ;
  assign w1131 = w516 | w1130 ;
  assign w1132 = ( w608 & w722 ) | ( w608 & ~w764 ) | ( w722 & ~w764 ) ;
  assign w1133 = w143 | w1131 ;
  assign w1134 = ( ~w143 & w764 ) | ( ~w143 & w783 ) | ( w764 & w783 ) ;
  assign w1135 = w1133 | w1134 ;
  assign w1136 = w1132 | w1135 ;
  assign w1137 = w388 | w459 ;
  assign w1138 = w1129 | w1137 ;
  assign w1139 = ( w104 & ~w1129 ) | ( w104 & w1136 ) | ( ~w1129 & w1136 ) ;
  assign w1140 = w1138 | w1139 ;
  assign w1141 = ( w385 & w429 ) | ( w385 & ~w860 ) | ( w429 & ~w860 ) ;
  assign w1142 = w95 | w1140 ;
  assign w1143 = ( ~w95 & w860 ) | ( ~w95 & w1126 ) | ( w860 & w1126 ) ;
  assign w1144 = w1142 | w1143 ;
  assign w1145 = w1141 | w1144 ;
  assign w1146 = ( w218 & ~w224 ) | ( w218 & w255 ) | ( ~w224 & w255 ) ;
  assign w1147 = w224 | w1146 ;
  assign w1148 = ( w176 & w316 ) | ( w176 & ~w392 ) | ( w316 & ~w392 ) ;
  assign w1149 = w113 | w1147 ;
  assign w1150 = ( ~w113 & w392 ) | ( ~w113 & w726 ) | ( w392 & w726 ) ;
  assign w1151 = w1149 | w1150 ;
  assign w1152 = w1148 | w1151 ;
  assign w1153 = w94 & w130 ;
  assign w1154 = w897 | w1153 ;
  assign w1155 = w422 | w466 ;
  assign w1156 = ( w120 & ~w506 ) | ( w120 & w560 ) | ( ~w506 & w560 ) ;
  assign w1157 = w506 | w1156 ;
  assign w1158 = w418 | w817 ;
  assign w1159 = w258 | w673 ;
  assign w1160 = ( w88 & ~w258 ) | ( w88 & w490 ) | ( ~w258 & w490 ) ;
  assign w1161 = w1159 | w1160 ;
  assign w1162 = w384 | w681 ;
  assign w1163 = ( w281 & ~w384 ) | ( w281 & w420 ) | ( ~w384 & w420 ) ;
  assign w1164 = w1162 | w1163 ;
  assign w1165 = w179 | w274 ;
  assign w1166 = w252 | w322 ;
  assign w1167 = ( w133 & ~w257 ) | ( w133 & w1166 ) | ( ~w257 & w1166 ) ;
  assign w1168 = w1164 | w1165 ;
  assign w1169 = ( w257 & w568 ) | ( w257 & ~w1165 ) | ( w568 & ~w1165 ) ;
  assign w1170 = w1168 | w1169 ;
  assign w1171 = w1167 | w1170 ;
  assign w1172 = ( w1155 & w1157 ) | ( w1155 & ~w1158 ) | ( w1157 & ~w1158 ) ;
  assign w1173 = w955 | w1171 ;
  assign w1174 = ( w1158 & w1161 ) | ( w1158 & ~w1171 ) | ( w1161 & ~w1171 ) ;
  assign w1175 = w1173 | w1174 ;
  assign w1176 = w1172 | w1175 ;
  assign w1177 = w353 | w640 ;
  assign w1178 = w661 | w1177 ;
  assign w1179 = ( ~w661 & w1154 ) | ( ~w661 & w1176 ) | ( w1154 & w1176 ) ;
  assign w1180 = w1178 | w1179 ;
  assign w1181 = w285 | w1030 ;
  assign w1182 = w662 | w999 ;
  assign w1183 = ( w101 & w784 ) | ( w101 & ~w999 ) | ( w784 & ~w999 ) ;
  assign w1184 = w1182 | w1183 ;
  assign w1185 = w165 | w465 ;
  assign w1186 = ( w263 & w275 ) | ( w263 & ~w286 ) | ( w275 & ~w286 ) ;
  assign w1187 = w63 | w1185 ;
  assign w1188 = ( ~w63 & w286 ) | ( ~w63 & w724 ) | ( w286 & w724 ) ;
  assign w1189 = w1187 | w1188 ;
  assign w1190 = w1186 | w1189 ;
  assign w1191 = ( ~w260 & w1181 ) | ( ~w260 & w1190 ) | ( w1181 & w1190 ) ;
  assign w1192 = w1180 | w1184 ;
  assign w1193 = ( w260 & w312 ) | ( w260 & ~w1184 ) | ( w312 & ~w1184 ) ;
  assign w1194 = w1192 | w1193 ;
  assign w1195 = w1191 | w1194 ;
  assign w1196 = ( ~w672 & w1145 ) | ( ~w672 & w1152 ) | ( w1145 & w1152 ) ;
  assign w1197 = w1125 | w1195 ;
  assign w1198 = ( w672 & w911 ) | ( w672 & ~w1195 ) | ( w911 & ~w1195 ) ;
  assign w1199 = w1197 | w1198 ;
  assign w1200 = w1196 | w1199 ;
  assign w1201 = ( w456 & w495 ) | ( w456 & ~w565 ) | ( w495 & ~w565 ) ;
  assign w1202 = w956 | w1200 ;
  assign w1203 = ( w565 & w623 ) | ( w565 & ~w956 ) | ( w623 & ~w956 ) ;
  assign w1204 = w1202 | w1203 ;
  assign w1205 = w1201 | w1204 ;
  assign w1206 = w103 | w664 ;
  assign w1207 = w44 | w313 ;
  assign w1208 = w411 | w429 ;
  assign w1209 = w169 | w570 ;
  assign w1210 = w956 | w1209 ;
  assign w1211 = ( w113 & w216 ) | ( w113 & ~w956 ) | ( w216 & ~w956 ) ;
  assign w1212 = w1210 | w1211 ;
  assign w1213 = w1181 | w1208 ;
  assign w1214 = w763 | w1213 ;
  assign w1215 = ( w763 & w799 ) | ( w763 & ~w1212 ) | ( w799 & ~w1212 ) ;
  assign w1216 = ~w1214 & w1215 ;
  assign w1217 = w104 | w283 ;
  assign w1218 = w1207 | w1217 ;
  assign w1219 = ( ~w76 & w1207 ) | ( ~w76 & w1216 ) | ( w1207 & w1216 ) ;
  assign w1220 = ~w1218 & w1219 ;
  assign w1221 = ( w144 & w201 ) | ( w144 & ~w341 ) | ( w201 & ~w341 ) ;
  assign w1222 = ~w135 & w1220 ;
  assign w1223 = ( ~w135 & w341 ) | ( ~w135 & w899 ) | ( w341 & w899 ) ;
  assign w1224 = w1222 & ~w1223 ;
  assign w1225 = ~w1221 & w1224 ;
  assign w1226 = w533 | w662 ;
  assign w1227 = ( w533 & ~w608 ) | ( w533 & w1225 ) | ( ~w608 & w1225 ) ;
  assign w1228 = ~w1226 & w1227 ;
  assign w1229 = w89 & w97 ;
  assign w1230 = ( w525 & w571 ) | ( w525 & ~w889 ) | ( w571 & ~w889 ) ;
  assign w1231 = w311 | w325 ;
  assign w1232 = ( ~w325 & w889 ) | ( ~w325 & w1001 ) | ( w889 & w1001 ) ;
  assign w1233 = w1231 | w1232 ;
  assign w1234 = w1230 | w1233 ;
  assign w1235 = w205 | w1229 ;
  assign w1236 = ( ~w205 & w309 ) | ( ~w205 & w1234 ) | ( w309 & w1234 ) ;
  assign w1237 = w1235 | w1236 ;
  assign w1238 = ( w230 & w315 ) | ( w230 & ~w390 ) | ( w315 & ~w390 ) ;
  assign w1239 = w68 | w124 ;
  assign w1240 = ( ~w124 & w390 ) | ( ~w124 & w593 ) | ( w390 & w593 ) ;
  assign w1241 = w1239 | w1240 ;
  assign w1242 = w1238 | w1241 ;
  assign w1243 = w227 | w567 ;
  assign w1244 = ( w138 & ~w227 ) | ( w138 & w287 ) | ( ~w227 & w287 ) ;
  assign w1245 = w1243 | w1244 ;
  assign w1246 = ( w198 & ~w415 ) | ( w198 & w663 ) | ( ~w415 & w663 ) ;
  assign w1247 = w415 | w1246 ;
  assign w1248 = w268 | w352 ;
  assign w1249 = w1247 | w1248 ;
  assign w1250 = ( w178 & w1245 ) | ( w178 & ~w1247 ) | ( w1245 & ~w1247 ) ;
  assign w1251 = w1249 | w1250 ;
  assign w1252 = ( w1180 & w1237 ) | ( w1180 & ~w1251 ) | ( w1237 & ~w1251 ) ;
  assign w1253 = ~w816 & w1228 ;
  assign w1254 = ( ~w816 & w1242 ) | ( ~w816 & w1251 ) | ( w1242 & w1251 ) ;
  assign w1255 = w1253 & ~w1254 ;
  assign w1256 = ~w1252 & w1255 ;
  assign w1257 = w505 | w515 ;
  assign w1258 = w1206 | w1257 ;
  assign w1259 = ( ~w122 & w1206 ) | ( ~w122 & w1256 ) | ( w1206 & w1256 ) ;
  assign w1260 = ~w1258 & w1259 ;
  assign w1261 = w361 | w605 ;
  assign w1262 = w175 | w1261 ;
  assign w1263 = ( w175 & ~w277 ) | ( w175 & w1260 ) | ( ~w277 & w1260 ) ;
  assign w1264 = ~w1262 & w1263 ;
  assign w1265 = w201 | w388 ;
  assign w1266 = w286 | w409 ;
  assign w1267 = ( w119 & ~w286 ) | ( w119 & w361 ) | ( ~w286 & w361 ) ;
  assign w1268 = w1266 | w1267 ;
  assign w1269 = ( w259 & w392 ) | ( w259 & ~w418 ) | ( w392 & ~w418 ) ;
  assign w1270 = w594 | w1268 ;
  assign w1271 = ( w418 & w496 ) | ( w418 & ~w1268 ) | ( w496 & ~w1268 ) ;
  assign w1272 = w1270 | w1271 ;
  assign w1273 = w1269 | w1272 ;
  assign w1274 = w123 & w251 ;
  assign w1275 = w256 | w466 ;
  assign w1276 = w339 | w1126 ;
  assign w1277 = w284 | w681 ;
  assign w1278 = w227 | w1277 ;
  assign w1279 = ( w167 & ~w227 ) | ( w167 & w283 ) | ( ~w227 & w283 ) ;
  assign w1280 = w1278 | w1279 ;
  assign w1281 = w358 | w504 ;
  assign w1282 = w354 | w783 ;
  assign w1283 = w232 | w565 ;
  assign w1284 = w642 | w673 ;
  assign w1285 = w226 | w1284 ;
  assign w1286 = ( w63 & ~w226 ) | ( w63 & w628 ) | ( ~w226 & w628 ) ;
  assign w1287 = w1285 | w1286 ;
  assign w1288 = ( w128 & ~w144 ) | ( w128 & w1287 ) | ( ~w144 & w1287 ) ;
  assign w1289 = w1282 | w1283 ;
  assign w1290 = ( w144 & w516 ) | ( w144 & ~w1283 ) | ( w516 & ~w1283 ) ;
  assign w1291 = w1289 | w1290 ;
  assign w1292 = w1288 | w1291 ;
  assign w1293 = ( w278 & w495 ) | ( w278 & ~w569 ) | ( w495 & ~w569 ) ;
  assign w1294 = w1281 | w1292 ;
  assign w1295 = ( w569 & w980 ) | ( w569 & ~w1281 ) | ( w980 & ~w1281 ) ;
  assign w1296 = w1294 | w1295 ;
  assign w1297 = w1293 | w1296 ;
  assign w1298 = w534 | w1001 ;
  assign w1299 = w51 | w1298 ;
  assign w1300 = ( ~w51 & w142 ) | ( ~w51 & w222 ) | ( w142 & w222 ) ;
  assign w1301 = w1299 | w1300 ;
  assign w1302 = w421 | w443 ;
  assign w1303 = w513 | w623 ;
  assign w1304 = w124 | w1303 ;
  assign w1305 = ( ~w124 & w389 ) | ( ~w124 & w532 ) | ( w389 & w532 ) ;
  assign w1306 = w1304 | w1305 ;
  assign w1307 = w313 | w899 ;
  assign w1308 = w1129 | w1307 ;
  assign w1309 = ( ~w1129 & w1302 ) | ( ~w1129 & w1306 ) | ( w1302 & w1306 ) ;
  assign w1310 = w1308 | w1309 ;
  assign w1311 = ( w212 & ~w267 ) | ( w212 & w1301 ) | ( ~w267 & w1301 ) ;
  assign w1312 = w1297 | w1310 ;
  assign w1313 = ( w267 & w1280 ) | ( w267 & ~w1310 ) | ( w1280 & ~w1310 ) ;
  assign w1314 = w1312 | w1313 ;
  assign w1315 = w1311 | w1314 ;
  assign w1316 = w420 | w1274 ;
  assign w1317 = w1275 | w1316 ;
  assign w1318 = ( ~w1275 & w1276 ) | ( ~w1275 & w1315 ) | ( w1276 & w1315 ) ;
  assign w1319 = w1317 | w1318 ;
  assign w1320 = ( w269 & w456 ) | ( w269 & ~w571 ) | ( w456 & ~w571 ) ;
  assign w1321 = w163 | w1319 ;
  assign w1322 = ( ~w163 & w571 ) | ( ~w163 & w951 ) | ( w571 & w951 ) ;
  assign w1323 = w1321 | w1322 ;
  assign w1324 = w1320 | w1323 ;
  assign w1325 = w641 | w663 ;
  assign w1326 = w362 | w1325 ;
  assign w1327 = ( w255 & ~w362 ) | ( w255 & w533 ) | ( ~w362 & w533 ) ;
  assign w1328 = w1326 | w1327 ;
  assign w1329 = ( w344 & w345 ) | ( w344 & ~w458 ) | ( w345 & ~w458 ) ;
  assign w1330 = w164 | w1328 ;
  assign w1331 = ( ~w164 & w458 ) | ( ~w164 & w509 ) | ( w458 & w509 ) ;
  assign w1332 = w1330 | w1331 ;
  assign w1333 = w1329 | w1332 ;
  assign w1334 = w430 | w605 ;
  assign w1335 = w92 | w1334 ;
  assign w1336 = ( ~w92 & w165 ) | ( ~w92 & w1333 ) | ( w165 & w1333 ) ;
  assign w1337 = w1335 | w1336 ;
  assign w1338 = ( ~w44 & w637 ) | ( ~w44 & w1337 ) | ( w637 & w1337 ) ;
  assign w1339 = w44 | w1338 ;
  assign w1340 = w40 & w75 ;
  assign w1341 = ( w449 & w625 ) | ( w449 & ~w697 ) | ( w625 & ~w697 ) ;
  assign w1342 = w272 | w385 ;
  assign w1343 = ( ~w385 & w697 ) | ( ~w385 & w1340 ) | ( w697 & w1340 ) ;
  assign w1344 = w1342 | w1343 ;
  assign w1345 = w1341 | w1344 ;
  assign w1346 = ( ~w252 & w315 ) | ( ~w252 & w1345 ) | ( w315 & w1345 ) ;
  assign w1347 = w252 | w1346 ;
  assign w1348 = ( w324 & w384 ) | ( w324 & ~w386 ) | ( w384 & ~w386 ) ;
  assign w1349 = w314 | w1165 ;
  assign w1350 = ( ~w314 & w386 ) | ( ~w314 & w445 ) | ( w386 & w445 ) ;
  assign w1351 = w1349 | w1350 ;
  assign w1352 = w1348 | w1351 ;
  assign w1353 = ( w285 & w320 ) | ( w285 & ~w491 ) | ( w320 & ~w491 ) ;
  assign w1354 = w115 | w1352 ;
  assign w1355 = ( ~w115 & w491 ) | ( ~w115 & w724 ) | ( w491 & w724 ) ;
  assign w1356 = w1354 | w1355 ;
  assign w1357 = w1353 | w1356 ;
  assign w1358 = ( w467 & w515 ) | ( w467 & ~w570 ) | ( w515 & ~w570 ) ;
  assign w1359 = w127 | w422 ;
  assign w1360 = ( ~w422 & w570 ) | ( ~w422 & w664 ) | ( w570 & w664 ) ;
  assign w1361 = w1359 | w1360 ;
  assign w1362 = w1358 | w1361 ;
  assign w1363 = w860 | w901 ;
  assign w1364 = w215 | w281 ;
  assign w1365 = w131 | w1364 ;
  assign w1366 = ( ~w131 & w175 ) | ( ~w131 & w1363 ) | ( w175 & w1363 ) ;
  assign w1367 = w1365 | w1366 ;
  assign w1368 = ( ~w118 & w742 ) | ( ~w118 & w1362 ) | ( w742 & w1362 ) ;
  assign w1369 = w1357 | w1367 ;
  assign w1370 = ( w118 & w606 ) | ( w118 & ~w1367 ) | ( w606 & ~w1367 ) ;
  assign w1371 = w1369 | w1370 ;
  assign w1372 = w1368 | w1371 ;
  assign w1373 = ( w81 & w263 ) | ( w81 & ~w318 ) | ( w263 & ~w318 ) ;
  assign w1374 = w1347 | w1372 ;
  assign w1375 = ( w318 & w758 ) | ( w318 & ~w1347 ) | ( w758 & ~w1347 ) ;
  assign w1376 = w1374 | w1375 ;
  assign w1377 = w1373 | w1376 ;
  assign w1378 = ( ~w203 & w218 ) | ( ~w203 & w1377 ) | ( w218 & w1377 ) ;
  assign w1379 = w203 | w1378 ;
  assign w1380 = ( w84 & w341 ) | ( w84 & ~w353 ) | ( w341 & ~w353 ) ;
  assign w1381 = w842 | w1379 ;
  assign w1382 = ( w353 & w390 ) | ( w353 & ~w842 ) | ( w390 & ~w842 ) ;
  assign w1383 = w1381 | w1382 ;
  assign w1384 = w1380 | w1383 ;
  assign w1385 = ( ~w561 & w1273 ) | ( ~w561 & w1339 ) | ( w1273 & w1339 ) ;
  assign w1386 = w1324 | w1384 ;
  assign w1387 = ( w561 & w817 ) | ( w561 & ~w1324 ) | ( w817 & ~w1324 ) ;
  assign w1388 = w1386 | w1387 ;
  assign w1389 = w1385 | w1388 ;
  assign w1390 = ( w147 & ~w169 ) | ( w147 & w1265 ) | ( ~w169 & w1265 ) ;
  assign w1391 = w956 | w1389 ;
  assign w1392 = ( w169 & w312 ) | ( w169 & ~w956 ) | ( w312 & ~w956 ) ;
  assign w1393 = w1391 | w1392 ;
  assign w1394 = w1390 | w1393 ;
  assign w1395 = ( w415 & w465 ) | ( w415 & ~w530 ) | ( w465 & ~w530 ) ;
  assign w1396 = w352 | w1394 ;
  assign w1397 = ( ~w352 & w530 ) | ( ~w352 & w640 ) | ( w530 & w640 ) ;
  assign w1398 = w1396 | w1397 ;
  assign w1399 = w1395 | w1398 ;
  assign w1400 = w202 | w605 ;
  assign w1401 = w142 | w255 ;
  assign w1402 = w286 | w722 ;
  assign w1403 = ( w224 & ~w286 ) | ( w224 & w506 ) | ( ~w286 & w506 ) ;
  assign w1404 = w1402 | w1403 ;
  assign w1405 = ( w76 & w165 ) | ( w76 & ~w254 ) | ( w165 & ~w254 ) ;
  assign w1406 = w1401 | w1404 ;
  assign w1407 = ( w254 & w339 ) | ( w254 & ~w1404 ) | ( w339 & ~w1404 ) ;
  assign w1408 = w1406 | w1407 ;
  assign w1409 = w1405 | w1408 ;
  assign w1410 = w116 | w899 ;
  assign w1411 = ( ~w116 & w284 ) | ( ~w116 & w1409 ) | ( w284 & w1409 ) ;
  assign w1412 = w1410 | w1411 ;
  assign w1413 = w313 | w470 ;
  assign w1414 = w341 | w593 ;
  assign w1415 = w206 | w1414 ;
  assign w1416 = ( ~w206 & w278 ) | ( ~w206 & w1413 ) | ( w278 & w1413 ) ;
  assign w1417 = w1415 | w1416 ;
  assign w1418 = w359 & ~w817 ;
  assign w1419 = ( w314 & w359 ) | ( w314 & w802 ) | ( w359 & w802 ) ;
  assign w1420 = w1418 & ~w1419 ;
  assign w1421 = w178 | w458 ;
  assign w1422 = w393 | w1128 ;
  assign w1423 = w257 | w1422 ;
  assign w1424 = ( w175 & ~w257 ) | ( w175 & w362 ) | ( ~w257 & w362 ) ;
  assign w1425 = w1423 | w1424 ;
  assign w1426 = w163 | w661 ;
  assign w1427 = ( w87 & ~w661 ) | ( w87 & w1425 ) | ( ~w661 & w1425 ) ;
  assign w1428 = w1426 | w1427 ;
  assign w1429 = ( w315 & w516 ) | ( w315 & ~w626 ) | ( w516 & ~w626 ) ;
  assign w1430 = w1421 | w1428 ;
  assign w1431 = ( w626 & w951 ) | ( w626 & ~w1421 ) | ( w951 & ~w1421 ) ;
  assign w1432 = w1430 | w1431 ;
  assign w1433 = w1429 | w1432 ;
  assign w1434 = ( w530 & ~w1206 ) | ( w530 & w1420 ) | ( ~w1206 & w1420 ) ;
  assign w1435 = w1417 | w1433 ;
  assign w1436 = ( w530 & w1340 ) | ( w530 & ~w1417 ) | ( w1340 & ~w1417 ) ;
  assign w1437 = w1435 | w1436 ;
  assign w1438 = w1434 & ~w1437 ;
  assign w1439 = ( w199 & w209 ) | ( w199 & ~w459 ) | ( w209 & ~w459 ) ;
  assign w1440 = ~w1154 & w1438 ;
  assign w1441 = ( w459 & w628 ) | ( w459 & ~w1154 ) | ( w628 & ~w1154 ) ;
  assign w1442 = w1440 & ~w1441 ;
  assign w1443 = ~w1439 & w1442 ;
  assign w1444 = ( w637 & w674 ) | ( w637 & ~w725 ) | ( w674 & ~w725 ) ;
  assign w1445 = w74 | w467 ;
  assign w1446 = ( ~w467 & w725 ) | ( ~w467 & w980 ) | ( w725 & w980 ) ;
  assign w1447 = w1445 | w1446 ;
  assign w1448 = w1444 | w1447 ;
  assign w1449 = ( w260 & w310 ) | ( w260 & ~w490 ) | ( w310 & ~w490 ) ;
  assign w1450 = w114 | w1448 ;
  assign w1451 = ( ~w114 & w490 ) | ( ~w114 & w764 ) | ( w490 & w764 ) ;
  assign w1452 = w1450 | w1451 ;
  assign w1453 = w1449 | w1452 ;
  assign w1454 = w63 | w680 ;
  assign w1455 = ( ~w63 & w253 ) | ( ~w63 & w1453 ) | ( w253 & w1453 ) ;
  assign w1456 = w1454 | w1455 ;
  assign w1457 = w353 | w681 ;
  assign w1458 = ( w51 & ~w353 ) | ( w51 & w496 ) | ( ~w353 & w496 ) ;
  assign w1459 = w1457 | w1458 ;
  assign w1460 = w56 | w135 ;
  assign w1461 = w258 | w595 ;
  assign w1462 = ( w423 & w625 ) | ( w423 & ~w697 ) | ( w625 & ~w697 ) ;
  assign w1463 = w1245 | w1461 ;
  assign w1464 = ( w697 & w783 ) | ( w697 & ~w1461 ) | ( w783 & ~w1461 ) ;
  assign w1465 = w1463 | w1464 ;
  assign w1466 = w1462 | w1465 ;
  assign w1467 = w495 | w525 ;
  assign w1468 = w1087 | w1467 ;
  assign w1469 = ( w136 & ~w1087 ) | ( w136 & w1466 ) | ( ~w1087 & w1466 ) ;
  assign w1470 = w1468 | w1469 ;
  assign w1471 = ( ~w68 & w208 ) | ( ~w68 & w1470 ) | ( w208 & w1470 ) ;
  assign w1472 = w68 | w1471 ;
  assign w1473 = w271 | w1086 ;
  assign w1474 = w606 | w642 ;
  assign w1475 = w119 | w1474 ;
  assign w1476 = ( ~w119 & w320 ) | ( ~w119 & w1088 ) | ( w320 & w1088 ) ;
  assign w1477 = w1475 | w1476 ;
  assign w1478 = ( w385 & ~w573 ) | ( w385 & w1473 ) | ( ~w573 & w1473 ) ;
  assign w1479 = w609 | w1477 ;
  assign w1480 = ( w573 & ~w609 ) | ( w573 & w837 ) | ( ~w609 & w837 ) ;
  assign w1481 = w1479 | w1480 ;
  assign w1482 = w1478 | w1481 ;
  assign w1483 = ( w838 & w911 ) | ( w838 & ~w1165 ) | ( w911 & ~w1165 ) ;
  assign w1484 = w1472 | w1482 ;
  assign w1485 = ( w1165 & w1265 ) | ( w1165 & ~w1482 ) | ( w1265 & ~w1482 ) ;
  assign w1486 = w1484 | w1485 ;
  assign w1487 = w1483 | w1486 ;
  assign w1488 = ( w144 & w205 ) | ( w144 & ~w409 ) | ( w205 & ~w409 ) ;
  assign w1489 = w59 | w1487 ;
  assign w1490 = ( ~w59 & w409 ) | ( ~w59 & w860 ) | ( w409 & w860 ) ;
  assign w1491 = w1489 | w1490 ;
  assign w1492 = w1488 | w1491 ;
  assign w1493 = ( ~w450 & w641 ) | ( ~w450 & w1492 ) | ( w641 & w1492 ) ;
  assign w1494 = w450 | w1493 ;
  assign w1495 = ( w122 & ~w131 ) | ( w122 & w569 ) | ( ~w131 & w569 ) ;
  assign w1496 = w131 | w1495 ;
  assign w1497 = w1460 | w1496 ;
  assign w1498 = w1456 | w1497 ;
  assign w1499 = ( ~w1456 & w1459 ) | ( ~w1456 & w1494 ) | ( w1459 & w1494 ) ;
  assign w1500 = w1498 | w1499 ;
  assign w1501 = ( w1302 & ~w1400 ) | ( w1302 & w1412 ) | ( ~w1400 & w1412 ) ;
  assign w1502 = w1443 & ~w1500 ;
  assign w1503 = ( w561 & w1400 ) | ( w561 & w1443 ) | ( w1400 & w1443 ) ;
  assign w1504 = w1502 & ~w1503 ;
  assign w1505 = ~w1501 & w1504 ;
  assign w1506 = ( w118 & w392 ) | ( w118 & ~w509 ) | ( w392 & ~w509 ) ;
  assign w1507 = ~w101 & w1505 ;
  assign w1508 = ( ~w101 & w509 ) | ( ~w101 & w787 ) | ( w509 & w787 ) ;
  assign w1509 = w1507 & ~w1508 ;
  assign w1510 = ~w1506 & w1509 ;
  assign w1511 = ( w265 & ~w421 ) | ( w265 & w570 ) | ( ~w421 & w570 ) ;
  assign w1512 = w421 | w1511 ;
  assign w1513 = w496 | w758 ;
  assign w1514 = w226 | w662 ;
  assign w1515 = ( w229 & w266 ) | ( w229 & ~w384 ) | ( w266 & ~w384 ) ;
  assign w1516 = w227 | w1417 ;
  assign w1517 = ( ~w227 & w384 ) | ( ~w227 & w725 ) | ( w384 & w725 ) ;
  assign w1518 = w1516 | w1517 ;
  assign w1519 = w1515 | w1518 ;
  assign w1520 = w467 | w1030 ;
  assign w1521 = w101 | w1520 ;
  assign w1522 = ( ~w101 & w128 ) | ( ~w101 & w1519 ) | ( w128 & w1519 ) ;
  assign w1523 = w1521 | w1522 ;
  assign w1524 = ( w315 & w429 ) | ( w315 & ~w899 ) | ( w429 & ~w899 ) ;
  assign w1525 = w74 | w142 ;
  assign w1526 = ( ~w142 & w899 ) | ( ~w142 & w1031 ) | ( w899 & w1031 ) ;
  assign w1527 = w1525 | w1526 ;
  assign w1528 = w1524 | w1527 ;
  assign w1529 = w95 | w277 ;
  assign w1530 = ( ~w95 & w127 ) | ( ~w95 & w1528 ) | ( w127 & w1528 ) ;
  assign w1531 = w1529 | w1530 ;
  assign w1532 = ( w419 & w512 ) | ( w419 & ~w764 ) | ( w512 & ~w764 ) ;
  assign w1533 = w125 | w1531 ;
  assign w1534 = ( ~w125 & w764 ) | ( ~w125 & w821 ) | ( w764 & w821 ) ;
  assign w1535 = w1533 | w1534 ;
  assign w1536 = w1532 | w1535 ;
  assign w1537 = w1514 | w1536 ;
  assign w1538 = ( w1513 & w1523 ) | ( w1513 & ~w1536 ) | ( w1523 & ~w1536 ) ;
  assign w1539 = w1537 | w1538 ;
  assign w1540 = ( w361 & w385 ) | ( w361 & ~w408 ) | ( w385 & ~w408 ) ;
  assign w1541 = w317 | w1539 ;
  assign w1542 = ( ~w317 & w408 ) | ( ~w317 & w606 ) | ( w408 & w606 ) ;
  assign w1543 = w1541 | w1542 ;
  assign w1544 = w1540 | w1543 ;
  assign w1545 = w571 | w664 ;
  assign w1546 = w144 | w1545 ;
  assign w1547 = ( ~w144 & w252 ) | ( ~w144 & w1544 ) | ( w252 & w1544 ) ;
  assign w1548 = w1546 | w1547 ;
  assign w1549 = ( w230 & w311 ) | ( w230 & ~w351 ) | ( w311 & ~w351 ) ;
  assign w1550 = w76 | w90 ;
  assign w1551 = ( ~w90 & w351 ) | ( ~w90 & w723 ) | ( w351 & w723 ) ;
  assign w1552 = w1550 | w1551 ;
  assign w1553 = w1549 | w1552 ;
  assign w1554 = ( w219 & w254 ) | ( w219 & ~w257 ) | ( w254 & ~w257 ) ;
  assign w1555 = w149 | w1553 ;
  assign w1556 = ( ~w149 & w257 ) | ( ~w149 & w837 ) | ( w257 & w837 ) ;
  assign w1557 = w1555 | w1556 ;
  assign w1558 = w1554 | w1557 ;
  assign w1559 = w783 | w1558 ;
  assign w1560 = w118 | w280 ;
  assign w1561 = w495 | w608 ;
  assign w1562 = w138 | w1561 ;
  assign w1563 = ( w115 & ~w138 ) | ( w115 & w488 ) | ( ~w138 & w488 ) ;
  assign w1564 = w1562 | w1563 ;
  assign w1565 = w340 | w386 ;
  assign w1566 = w275 | w673 ;
  assign w1567 = ( w726 & w1155 ) | ( w726 & ~w1566 ) | ( w1155 & ~w1566 ) ;
  assign w1568 = w1566 | w1567 ;
  assign w1569 = ( w215 & ~w310 ) | ( w215 & w1565 ) | ( ~w310 & w1565 ) ;
  assign w1570 = w1363 | w1568 ;
  assign w1571 = ( w310 & w443 ) | ( w310 & ~w1363 ) | ( w443 & ~w1363 ) ;
  assign w1572 = w1570 | w1571 ;
  assign w1573 = w1569 | w1572 ;
  assign w1574 = ( ~w116 & w1131 ) | ( ~w116 & w1564 ) | ( w1131 & w1564 ) ;
  assign w1575 = w432 | w1573 ;
  assign w1576 = ( w116 & ~w432 ) | ( w116 & w456 ) | ( ~w432 & w456 ) ;
  assign w1577 = w1575 | w1576 ;
  assign w1578 = w1574 | w1577 ;
  assign w1579 = w1461 | w1560 ;
  assign w1580 = w1578 | w1579 ;
  assign w1581 = ( w594 & w1339 ) | ( w594 & ~w1578 ) | ( w1339 & ~w1578 ) ;
  assign w1582 = w1580 | w1581 ;
  assign w1583 = ( ~w199 & w565 ) | ( ~w199 & w1582 ) | ( w565 & w1582 ) ;
  assign w1584 = w199 | w1583 ;
  assign w1585 = ( w287 & w324 ) | ( w287 & ~w505 ) | ( w324 & ~w505 ) ;
  assign w1586 = w285 | w1584 ;
  assign w1587 = ( ~w285 & w505 ) | ( ~w285 & w524 ) | ( w505 & w524 ) ;
  assign w1588 = w1586 | w1587 ;
  assign w1589 = w1585 | w1588 ;
  assign w1590 = w256 | w561 ;
  assign w1591 = ( w259 & ~w449 ) | ( w259 & w1590 ) | ( ~w449 & w1590 ) ;
  assign w1592 = w177 | w264 ;
  assign w1593 = ( ~w264 & w449 ) | ( ~w264 & w1001 ) | ( w449 & w1001 ) ;
  assign w1594 = w1592 | w1593 ;
  assign w1595 = w1591 | w1594 ;
  assign w1596 = ( w98 & w253 ) | ( w98 & ~w352 ) | ( w253 & ~w352 ) ;
  assign w1597 = w1589 | w1595 ;
  assign w1598 = ( w352 & w459 ) | ( w352 & ~w1595 ) | ( w459 & ~w1595 ) ;
  assign w1599 = w1597 | w1598 ;
  assign w1600 = w1596 | w1599 ;
  assign w1601 = ( ~w209 & w636 ) | ( ~w209 & w1559 ) | ( w636 & w1559 ) ;
  assign w1602 = w1548 | w1600 ;
  assign w1603 = ( w209 & w316 ) | ( w209 & ~w1548 ) | ( w316 & ~w1548 ) ;
  assign w1604 = w1602 | w1603 ;
  assign w1605 = w1601 | w1604 ;
  assign w1606 = ( w418 & ~w530 ) | ( w418 & w1512 ) | ( ~w530 & w1512 ) ;
  assign w1607 = w270 | w1605 ;
  assign w1608 = ( ~w270 & w530 ) | ( ~w270 & w1340 ) | ( w530 & w1340 ) ;
  assign w1609 = w1607 | w1608 ;
  assign w1610 = w1606 | w1609 ;
  assign w1611 = w423 | w534 ;
  assign w1612 = w131 | w1611 ;
  assign w1613 = ( ~w131 & w179 ) | ( ~w131 & w1610 ) | ( w179 & w1610 ) ;
  assign w1614 = w1612 | w1613 ;
  assign w1615 = w266 | w531 ;
  assign w1616 = w142 | w312 ;
  assign w1617 = w111 | w724 ;
  assign w1618 = w254 | w1229 ;
  assign w1619 = ( w445 & ~w447 ) | ( w445 & w783 ) | ( ~w447 & w783 ) ;
  assign w1620 = w447 | w1619 ;
  assign w1621 = w122 | w505 ;
  assign w1622 = w1618 | w1621 ;
  assign w1623 = ( w887 & ~w1618 ) | ( w887 & w1620 ) | ( ~w1618 & w1620 ) ;
  assign w1624 = w1622 | w1623 ;
  assign w1625 = w257 | w623 ;
  assign w1626 = w212 | w1625 ;
  assign w1627 = ( w51 & ~w212 ) | ( w51 & w1624 ) | ( ~w212 & w1624 ) ;
  assign w1628 = w1626 | w1627 ;
  assign w1629 = w641 | w664 ;
  assign w1630 = ( w256 & w423 ) | ( w256 & ~w504 ) | ( w423 & ~w504 ) ;
  assign w1631 = w176 | w1461 ;
  assign w1632 = ( ~w176 & w504 ) | ( ~w176 & w697 ) | ( w504 & w697 ) ;
  assign w1633 = w1631 | w1632 ;
  assign w1634 = w1630 | w1633 ;
  assign w1635 = w1514 | w1629 ;
  assign w1636 = w1634 | w1635 ;
  assign w1637 = ( w87 & w1628 ) | ( w87 & ~w1634 ) | ( w1628 & ~w1634 ) ;
  assign w1638 = w1636 | w1637 ;
  assign w1639 = w230 | w1617 ;
  assign w1640 = w126 | w1639 ;
  assign w1641 = ( ~w126 & w742 ) | ( ~w126 & w1638 ) | ( w742 & w1638 ) ;
  assign w1642 = w1640 | w1641 ;
  assign w1643 = w143 | w642 ;
  assign w1644 = ( ~w143 & w269 ) | ( ~w143 & w1642 ) | ( w269 & w1642 ) ;
  assign w1645 = w1643 | w1644 ;
  assign w1646 = w131 | w341 ;
  assign w1647 = w608 | w1031 ;
  assign w1648 = w164 | w1647 ;
  assign w1649 = ( ~w164 & w262 ) | ( ~w164 & w276 ) | ( w262 & w276 ) ;
  assign w1650 = w1648 | w1649 ;
  assign w1651 = w390 | w496 ;
  assign w1652 = w68 | w1651 ;
  assign w1653 = ( ~w68 & w224 ) | ( ~w68 & w1650 ) | ( w224 & w1650 ) ;
  assign w1654 = w1652 | w1653 ;
  assign w1655 = ( w491 & w640 ) | ( w491 & ~w1030 ) | ( w640 & ~w1030 ) ;
  assign w1656 = w311 | w431 ;
  assign w1657 = ( ~w431 & w1030 ) | ( ~w431 & w1274 ) | ( w1030 & w1274 ) ;
  assign w1658 = w1656 | w1657 ;
  assign w1659 = w1655 | w1658 ;
  assign w1660 = w626 | w1001 ;
  assign w1661 = w320 | w1660 ;
  assign w1662 = ( w313 & ~w320 ) | ( w313 & w443 ) | ( ~w320 & w443 ) ;
  assign w1663 = w1661 | w1662 ;
  assign w1664 = ( w76 & ~w605 ) | ( w76 & w1663 ) | ( ~w605 & w1663 ) ;
  assign w1665 = w1654 | w1659 ;
  assign w1666 = ( w605 & w680 ) | ( w605 & ~w1659 ) | ( w680 & ~w1659 ) ;
  assign w1667 = w1665 | w1666 ;
  assign w1668 = w1664 | w1667 ;
  assign w1669 = w458 | w561 ;
  assign w1670 = w1646 | w1669 ;
  assign w1671 = ( w283 & ~w1646 ) | ( w283 & w1668 ) | ( ~w1646 & w1668 ) ;
  assign w1672 = w1670 | w1671 ;
  assign w1673 = ( w354 & w408 ) | ( w354 & ~w465 ) | ( w408 & ~w465 ) ;
  assign w1674 = w56 | w1672 ;
  assign w1675 = ( ~w56 & w465 ) | ( ~w56 & w628 ) | ( w465 & w628 ) ;
  assign w1676 = w1674 | w1675 ;
  assign w1677 = w1673 | w1676 ;
  assign w1678 = ( ~w259 & w488 ) | ( ~w259 & w1677 ) | ( w488 & w1677 ) ;
  assign w1679 = w259 | w1678 ;
  assign w1680 = ( w361 & w418 ) | ( w361 & ~w625 ) | ( w418 & ~w625 ) ;
  assign w1681 = w227 | w260 ;
  assign w1682 = ( ~w260 & w625 ) | ( ~w260 & w1340 ) | ( w625 & w1340 ) ;
  assign w1683 = w1681 | w1682 ;
  assign w1684 = w1680 | w1683 ;
  assign w1685 = w324 | w722 ;
  assign w1686 = ( w255 & ~w324 ) | ( w255 & w421 ) | ( ~w324 & w421 ) ;
  assign w1687 = w1685 | w1686 ;
  assign w1688 = ( ~w199 & w315 ) | ( ~w199 & w1283 ) | ( w315 & w1283 ) ;
  assign w1689 = w199 | w1688 ;
  assign w1690 = w787 | w1687 ;
  assign w1691 = ( w205 & ~w1687 ) | ( w205 & w1689 ) | ( ~w1687 & w1689 ) ;
  assign w1692 = w1690 | w1691 ;
  assign w1693 = ( ~w149 & w1684 ) | ( ~w149 & w1692 ) | ( w1684 & w1692 ) ;
  assign w1694 = w1645 | w1679 ;
  assign w1695 = ( w149 & w214 ) | ( w149 & ~w1645 ) | ( w214 & ~w1645 ) ;
  assign w1696 = w1694 | w1695 ;
  assign w1697 = w1693 | w1696 ;
  assign w1698 = ( w416 & w1276 ) | ( w416 & ~w1615 ) | ( w1276 & ~w1615 ) ;
  assign w1699 = w756 | w1697 ;
  assign w1700 = ( ~w756 & w1615 ) | ( ~w756 & w1616 ) | ( w1615 & w1616 ) ;
  assign w1701 = w1699 | w1700 ;
  assign w1702 = w1698 | w1701 ;
  assign w1703 = ( w310 & w344 ) | ( w310 & ~w345 ) | ( w344 & ~w345 ) ;
  assign w1704 = w120 | w1702 ;
  assign w1705 = ( ~w120 & w345 ) | ( ~w120 & w570 ) | ( w345 & w570 ) ;
  assign w1706 = w1704 | w1705 ;
  assign w1707 = w1703 | w1706 ;
  assign w1708 = w569 | w1130 ;
  assign w1709 = w253 | w1708 ;
  assign w1710 = ( ~w253 & w268 ) | ( ~w253 & w1707 ) | ( w268 & w1707 ) ;
  assign w1711 = w1709 | w1710 ;
  assign w1712 = w101 | w226 ;
  assign w1713 = w56 | w459 ;
  assign w1714 = ( w422 & w492 ) | ( w422 & ~w561 ) | ( w492 & ~w561 ) ;
  assign w1715 = w51 | w199 ;
  assign w1716 = ( ~w199 & w561 ) | ( ~w199 & w860 ) | ( w561 & w860 ) ;
  assign w1717 = w1715 | w1716 ;
  assign w1718 = w1714 | w1717 ;
  assign w1719 = w76 | w1718 ;
  assign w1720 = w1512 | w1719 ;
  assign w1721 = ( w952 & ~w1512 ) | ( w952 & w1713 ) | ( ~w1512 & w1713 ) ;
  assign w1722 = w1720 | w1721 ;
  assign w1723 = ( w419 & w530 ) | ( w419 & ~w593 ) | ( w530 & ~w593 ) ;
  assign w1724 = w208 | w1722 ;
  assign w1725 = ( ~w208 & w593 ) | ( ~w208 & w726 ) | ( w593 & w726 ) ;
  assign w1726 = w1724 | w1725 ;
  assign w1727 = w1723 | w1726 ;
  assign w1728 = ( w637 & ~w724 ) | ( w637 & w1130 ) | ( ~w724 & w1130 ) ;
  assign w1729 = w724 | w1728 ;
  assign w1730 = w284 | w1729 ;
  assign w1731 = ( w283 & w800 ) | ( w283 & ~w1729 ) | ( w800 & ~w1729 ) ;
  assign w1732 = w1730 | w1731 ;
  assign w1733 = w429 | w596 ;
  assign w1734 = w272 | w1733 ;
  assign w1735 = ( ~w272 & w351 ) | ( ~w272 & w1732 ) | ( w351 & w1732 ) ;
  assign w1736 = w1734 | w1735 ;
  assign w1737 = w385 | w605 ;
  assign w1738 = w163 | w1737 ;
  assign w1739 = ( w141 & ~w163 ) | ( w141 & w383 ) | ( ~w163 & w383 ) ;
  assign w1740 = w1738 | w1739 ;
  assign w1741 = w423 | w515 ;
  assign w1742 = w225 | w470 ;
  assign w1743 = ( w104 & ~w225 ) | ( w104 & w281 ) | ( ~w225 & w281 ) ;
  assign w1744 = w1742 | w1743 ;
  assign w1745 = ( w125 & ~w350 ) | ( w125 & w354 ) | ( ~w350 & w354 ) ;
  assign w1746 = w350 | w1745 ;
  assign w1747 = w787 | w1746 ;
  assign w1748 = ( w320 & w1744 ) | ( w320 & ~w1746 ) | ( w1744 & ~w1746 ) ;
  assign w1749 = w1747 | w1748 ;
  assign w1750 = ( w1712 & ~w1740 ) | ( w1712 & w1749 ) | ( ~w1740 & w1749 ) ;
  assign w1751 = w1727 | w1736 ;
  assign w1752 = ( ~w1736 & w1740 ) | ( ~w1736 & w1741 ) | ( w1740 & w1741 ) ;
  assign w1753 = w1751 | w1752 ;
  assign w1754 = w1750 | w1753 ;
  assign w1755 = ~w325 & w359 ;
  assign w1756 = ~w139 & w1755 ;
  assign w1757 = ( ~w139 & w269 ) | ( ~w139 & w1754 ) | ( w269 & w1754 ) ;
  assign w1758 = w1756 & ~w1757 ;
  assign w1759 = w463 | w533 ;
  assign w1760 = w118 | w606 ;
  assign w1761 = w1185 | w1760 ;
  assign w1762 = ( w1185 & w1758 ) | ( w1185 & ~w1759 ) | ( w1758 & ~w1759 ) ;
  assign w1763 = ~w1761 & w1762 ;
  assign w1764 = ( w122 & ~w271 ) | ( w122 & w1763 ) | ( ~w271 & w1763 ) ;
  assign w1765 = ~w122 & w1764 ;
  assign w1766 = ( w128 & w180 ) | ( w128 & ~w223 ) | ( w180 & ~w223 ) ;
  assign w1767 = ~w115 & w1765 ;
  assign w1768 = ( ~w115 & w223 ) | ( ~w115 & w725 ) | ( w223 & w725 ) ;
  assign w1769 = w1767 & ~w1768 ;
  assign w1770 = ~w1766 & w1769 ;
  assign w1771 = ( w362 & w447 ) | ( w362 & ~w516 ) | ( w447 & ~w516 ) ;
  assign w1772 = w175 | w255 ;
  assign w1773 = ( ~w255 & w516 ) | ( ~w255 & w641 ) | ( w516 & w641 ) ;
  assign w1774 = w1772 | w1773 ;
  assign w1775 = w1771 | w1774 ;
  assign w1776 = w90 | w1274 ;
  assign w1777 = ( ~w90 & w342 ) | ( ~w90 & w1775 ) | ( w342 & w1775 ) ;
  assign w1778 = w1776 | w1777 ;
  assign w1779 = ( w256 & w424 ) | ( w256 & ~w488 ) | ( w424 & ~w488 ) ;
  assign w1780 = w59 | w169 ;
  assign w1781 = ( ~w169 & w488 ) | ( ~w169 & w673 ) | ( w488 & w673 ) ;
  assign w1782 = w1780 | w1781 ;
  assign w1783 = w1779 | w1782 ;
  assign w1784 = w443 | w1094 ;
  assign w1785 = w340 | w1784 ;
  assign w1786 = ( w133 & ~w340 ) | ( w133 & w388 ) | ( ~w340 & w388 ) ;
  assign w1787 = w1785 | w1786 ;
  assign w1788 = w227 | w490 ;
  assign w1789 = ( w164 & ~w227 ) | ( w164 & w262 ) | ( ~w227 & w262 ) ;
  assign w1790 = w1788 | w1789 ;
  assign w1791 = w86 | w897 ;
  assign w1792 = ( w74 & ~w86 ) | ( w74 & w495 ) | ( ~w86 & w495 ) ;
  assign w1793 = w1791 | w1792 ;
  assign w1794 = ( ~w221 & w1790 ) | ( ~w221 & w1793 ) | ( w1790 & w1793 ) ;
  assign w1795 = w1404 | w1787 ;
  assign w1796 = ( w221 & w640 ) | ( w221 & ~w1787 ) | ( w640 & ~w1787 ) ;
  assign w1797 = w1795 | w1796 ;
  assign w1798 = w1794 | w1797 ;
  assign w1799 = ( w147 & ~w205 ) | ( w147 & w1783 ) | ( ~w205 & w1783 ) ;
  assign w1800 = w204 | w1798 ;
  assign w1801 = ( ~w204 & w205 ) | ( ~w204 & w314 ) | ( w205 & w314 ) ;
  assign w1802 = w1800 | w1801 ;
  assign w1803 = w1799 | w1802 ;
  assign w1804 = ( w149 & w420 ) | ( w149 & ~w569 ) | ( w420 & ~w569 ) ;
  assign w1805 = w143 | w1803 ;
  assign w1806 = ( ~w143 & w569 ) | ( ~w143 & w1126 ) | ( w569 & w1126 ) ;
  assign w1807 = w1805 | w1806 ;
  assign w1808 = w1804 | w1807 ;
  assign w1809 = ( w662 & w680 ) | ( w662 & ~w764 ) | ( w680 & ~w764 ) ;
  assign w1810 = w113 | w210 ;
  assign w1811 = ( ~w210 & w764 ) | ( ~w210 & w802 ) | ( w764 & w802 ) ;
  assign w1812 = w1810 | w1811 ;
  assign w1813 = w1809 | w1812 ;
  assign w1814 = w418 | w697 ;
  assign w1815 = w260 | w466 ;
  assign w1816 = w201 | w1815 ;
  assign w1817 = ( ~w201 & w209 ) | ( ~w201 & w1814 ) | ( w209 & w1814 ) ;
  assign w1818 = w1816 | w1817 ;
  assign w1819 = w114 | w230 ;
  assign w1820 = w1818 | w1819 ;
  assign w1821 = ( w1808 & w1813 ) | ( w1808 & ~w1818 ) | ( w1813 & ~w1818 ) ;
  assign w1822 = w1820 | w1821 ;
  assign w1823 = w785 | w1207 ;
  assign w1824 = w1822 | w1823 ;
  assign w1825 = ( w1770 & ~w1778 ) | ( w1770 & w1822 ) | ( ~w1778 & w1822 ) ;
  assign w1826 = ~w1824 & w1825 ;
  assign w1827 = ( w103 & w390 ) | ( w103 & ~w504 ) | ( w390 & ~w504 ) ;
  assign w1828 = ~w594 & w1826 ;
  assign w1829 = ( w504 & w567 ) | ( w504 & ~w594 ) | ( w567 & ~w594 ) ;
  assign w1830 = w1828 & ~w1829 ;
  assign w1831 = ~w1827 & w1830 ;
  assign w1832 = w135 | w889 ;
  assign w1833 = ( w135 & ~w309 ) | ( w135 & w1831 ) | ( ~w309 & w1831 ) ;
  assign w1834 = ~w1832 & w1833 ;
  assign w1835 = w662 | w837 ;
  assign w1836 = w163 | w595 ;
  assign w1837 = w124 | w281 ;
  assign w1838 = w1128 | w1229 ;
  assign w1839 = w1837 | w1838 ;
  assign w1840 = ( w133 & w911 ) | ( w133 & ~w1837 ) | ( w911 & ~w1837 ) ;
  assign w1841 = w1839 | w1840 ;
  assign w1842 = w506 | w764 ;
  assign w1843 = w1836 | w1842 ;
  assign w1844 = ( w210 & ~w1836 ) | ( w210 & w1841 ) | ( ~w1836 & w1841 ) ;
  assign w1845 = w1843 | w1844 ;
  assign w1846 = w525 | w697 ;
  assign w1847 = w315 | w1846 ;
  assign w1848 = ( ~w315 & w456 ) | ( ~w315 & w1845 ) | ( w456 & w1845 ) ;
  assign w1849 = w1847 | w1848 ;
  assign w1850 = w512 | w513 ;
  assign w1851 = w339 | w1850 ;
  assign w1852 = ( w199 & ~w339 ) | ( w199 & w350 ) | ( ~w339 & w350 ) ;
  assign w1853 = w1851 | w1852 ;
  assign w1854 = w625 | w725 ;
  assign w1855 = w318 | w1854 ;
  assign w1856 = ( w74 & ~w318 ) | ( w74 & w431 ) | ( ~w318 & w431 ) ;
  assign w1857 = w1855 | w1856 ;
  assign w1858 = w1853 | w1857 ;
  assign w1859 = w493 | w1858 ;
  assign w1860 = ( ~w493 & w514 ) | ( ~w493 & w1040 ) | ( w514 & w1040 ) ;
  assign w1861 = w1859 | w1860 ;
  assign w1862 = ( w104 & w143 ) | ( w104 & ~w278 ) | ( w143 & ~w278 ) ;
  assign w1863 = w168 | w1861 ;
  assign w1864 = ( ~w168 & w278 ) | ( ~w168 & w409 ) | ( w278 & w409 ) ;
  assign w1865 = w1863 | w1864 ;
  assign w1866 = w1862 | w1865 ;
  assign w1867 = w359 & ~w901 ;
  assign w1868 = ~w161 & w1867 ;
  assign w1869 = ( ~w161 & w256 ) | ( ~w161 & w1866 ) | ( w256 & w1866 ) ;
  assign w1870 = w1868 & ~w1869 ;
  assign w1871 = ( w286 & w466 ) | ( w286 & ~w642 ) | ( w466 & ~w642 ) ;
  assign w1872 = w178 | w253 ;
  assign w1873 = ( ~w253 & w642 ) | ( ~w253 & w889 ) | ( w642 & w889 ) ;
  assign w1874 = w1872 | w1873 ;
  assign w1875 = w1871 | w1874 ;
  assign w1876 = ( w257 & w317 ) | ( w257 & ~w567 ) | ( w317 & ~w567 ) ;
  assign w1877 = w59 | w450 ;
  assign w1878 = ( ~w59 & w567 ) | ( ~w59 & w1130 ) | ( w567 & w1130 ) ;
  assign w1879 = w1877 | w1878 ;
  assign w1880 = w1876 | w1879 ;
  assign w1881 = w92 | w128 ;
  assign w1882 = w393 | w606 ;
  assign w1883 = w208 | w504 ;
  assign w1884 = w463 | w787 ;
  assign w1885 = w1126 | w1884 ;
  assign w1886 = ( w203 & w1712 ) | ( w203 & ~w1884 ) | ( w1712 & ~w1884 ) ;
  assign w1887 = w1885 | w1886 ;
  assign w1888 = ( w272 & w490 ) | ( w272 & ~w505 ) | ( w490 & ~w505 ) ;
  assign w1889 = w169 | w1887 ;
  assign w1890 = ( ~w169 & w505 ) | ( ~w169 & w1086 ) | ( w505 & w1086 ) ;
  assign w1891 = w1889 | w1890 ;
  assign w1892 = w1888 | w1891 ;
  assign w1893 = w530 | w571 ;
  assign w1894 = w320 | w1893 ;
  assign w1895 = ( ~w320 & w358 ) | ( ~w320 & w1892 ) | ( w358 & w1892 ) ;
  assign w1896 = w1894 | w1895 ;
  assign w1897 = ( w342 & w388 ) | ( w342 & ~w533 ) | ( w388 & ~w533 ) ;
  assign w1898 = w88 | w119 ;
  assign w1899 = ( ~w119 & w533 ) | ( ~w119 & w980 ) | ( w533 & w980 ) ;
  assign w1900 = w1898 | w1899 ;
  assign w1901 = w1897 | w1900 ;
  assign w1902 = ( ~w411 & w608 ) | ( ~w411 & w1901 ) | ( w608 & w1901 ) ;
  assign w1903 = w411 | w1902 ;
  assign w1904 = w1883 | w1903 ;
  assign w1905 = ( w517 & w1896 ) | ( w517 & ~w1903 ) | ( w1896 & ~w1903 ) ;
  assign w1906 = w1904 | w1905 ;
  assign w1907 = w224 | w413 ;
  assign w1908 = w1617 | w1907 ;
  assign w1909 = ( ~w1617 & w1882 ) | ( ~w1617 & w1906 ) | ( w1882 & w1906 ) ;
  assign w1910 = w1908 | w1909 ;
  assign w1911 = w817 | w860 ;
  assign w1912 = w1881 | w1911 ;
  assign w1913 = ( w313 & ~w1881 ) | ( w313 & w1910 ) | ( ~w1881 & w1910 ) ;
  assign w1914 = w1912 | w1913 ;
  assign w1915 = w175 | w573 ;
  assign w1916 = ( ~w175 & w495 ) | ( ~w175 & w1914 ) | ( w495 & w1914 ) ;
  assign w1917 = w1915 | w1916 ;
  assign w1918 = ( ~w491 & w641 ) | ( ~w491 & w1917 ) | ( w641 & w1917 ) ;
  assign w1919 = w491 | w1918 ;
  assign w1920 = ( w260 & w312 ) | ( w260 & ~w353 ) | ( w312 & ~w353 ) ;
  assign w1921 = w206 | w1919 ;
  assign w1922 = ( ~w206 & w353 ) | ( ~w206 & w470 ) | ( w353 & w470 ) ;
  assign w1923 = w1921 | w1922 ;
  assign w1924 = w1920 | w1923 ;
  assign w1925 = ( ~w1566 & w1849 ) | ( ~w1566 & w1880 ) | ( w1849 & w1880 ) ;
  assign w1926 = w1870 & ~w1924 ;
  assign w1927 = ( w1566 & w1870 ) | ( w1566 & w1875 ) | ( w1870 & w1875 ) ;
  assign w1928 = w1926 & ~w1927 ;
  assign w1929 = ~w1925 & w1928 ;
  assign w1930 = ( ~w311 & w532 ) | ( ~w311 & w1835 ) | ( w532 & w1835 ) ;
  assign w1931 = ~w264 & w1929 ;
  assign w1932 = ( ~w264 & w311 ) | ( ~w264 & w389 ) | ( w311 & w389 ) ;
  assign w1933 = w1931 & ~w1932 ;
  assign w1934 = ~w1930 & w1933 ;
  assign w1935 = ( w122 & w218 ) | ( w122 & ~w227 ) | ( w218 & ~w227 ) ;
  assign w1936 = ~w1064 & w1934 ;
  assign w1937 = ( w227 & w269 ) | ( w227 & ~w1064 ) | ( w269 & ~w1064 ) ;
  assign w1938 = w1936 & ~w1937 ;
  assign w1939 = ~w1935 & w1938 ;
  assign w1940 = w136 | w447 ;
  assign w1941 = ( w63 & ~w389 ) | ( w63 & w1940 ) | ( ~w389 & w1940 ) ;
  assign w1942 = w1275 | w1473 ;
  assign w1943 = ( w389 & w722 ) | ( w389 & ~w1473 ) | ( w722 & ~w1473 ) ;
  assign w1944 = w1942 | w1943 ;
  assign w1945 = w1941 | w1944 ;
  assign w1946 = w260 | w899 ;
  assign w1947 = ( w223 & ~w260 ) | ( w223 & w821 ) | ( ~w260 & w821 ) ;
  assign w1948 = w1946 | w1947 ;
  assign w1949 = w95 | w787 ;
  assign w1950 = ( ~w95 & w265 ) | ( ~w95 & w1948 ) | ( w265 & w1948 ) ;
  assign w1951 = w1949 | w1950 ;
  assign w1952 = w176 | w280 ;
  assign w1953 = ( w104 & ~w176 ) | ( w104 & w269 ) | ( ~w176 & w269 ) ;
  assign w1954 = w1952 | w1953 ;
  assign w1955 = w262 | w674 ;
  assign w1956 = ( w116 & w624 ) | ( w116 & ~w1955 ) | ( w624 & ~w1955 ) ;
  assign w1957 = w1955 | w1956 ;
  assign w1958 = w275 | w511 ;
  assign w1959 = w1746 | w1958 ;
  assign w1960 = ( w128 & ~w1746 ) | ( w128 & w1957 ) | ( ~w1746 & w1957 ) ;
  assign w1961 = w1959 | w1960 ;
  assign w1962 = ( ~w149 & w1237 ) | ( ~w149 & w1961 ) | ( w1237 & w1961 ) ;
  assign w1963 = w1063 | w1379 ;
  assign w1964 = ( w149 & w214 ) | ( w149 & ~w1063 ) | ( w214 & ~w1063 ) ;
  assign w1965 = w1963 | w1964 ;
  assign w1966 = w1962 | w1965 ;
  assign w1967 = ( ~w209 & w1951 ) | ( ~w209 & w1954 ) | ( w1951 & w1954 ) ;
  assign w1968 = w1945 | w1966 ;
  assign w1969 = ( w209 & w316 ) | ( w209 & ~w1945 ) | ( w316 & ~w1945 ) ;
  assign w1970 = w1968 | w1969 ;
  assign w1971 = w1967 | w1970 ;
  assign w1972 = ( w595 & w596 ) | ( w595 & ~w725 ) | ( w596 & ~w725 ) ;
  assign w1973 = w411 | w1971 ;
  assign w1974 = ( ~w411 & w725 ) | ( ~w411 & w1128 ) | ( w725 & w1128 ) ;
  assign w1975 = w1973 | w1974 ;
  assign w1976 = w1972 | w1975 ;
  assign w1977 = w201 | w530 ;
  assign w1978 = w218 | w525 ;
  assign w1979 = w573 | w628 ;
  assign w1980 = ( w723 & w726 ) | ( w723 & ~w821 ) | ( w726 & ~w821 ) ;
  assign w1981 = w284 | w313 ;
  assign w1982 = ( ~w313 & w821 ) | ( ~w313 & w1094 ) | ( w821 & w1094 ) ;
  assign w1983 = w1981 | w1982 ;
  assign w1984 = w1980 | w1983 ;
  assign w1985 = w101 | w285 ;
  assign w1986 = ( ~w101 & w229 ) | ( ~w101 & w1984 ) | ( w229 & w1984 ) ;
  assign w1987 = w1985 | w1986 ;
  assign w1988 = w681 | w1128 ;
  assign w1989 = ( w209 & ~w681 ) | ( w209 & w764 ) | ( ~w681 & w764 ) ;
  assign w1990 = w1988 | w1989 ;
  assign w1991 = w359 & ~w458 ;
  assign w1992 = ( w222 & w359 ) | ( w222 & w420 ) | ( w359 & w420 ) ;
  assign w1993 = w1991 & ~w1992 ;
  assign w1994 = ( w253 & ~w459 ) | ( w253 & w1461 ) | ( ~w459 & w1461 ) ;
  assign w1995 = ~w888 & w1993 ;
  assign w1996 = ( w459 & w642 ) | ( w459 & ~w888 ) | ( w642 & ~w888 ) ;
  assign w1997 = w1995 & ~w1996 ;
  assign w1998 = ~w1994 & w1997 ;
  assign w1999 = ( w259 & w309 ) | ( w259 & ~w324 ) | ( w309 & ~w324 ) ;
  assign w2000 = ~w255 & w1998 ;
  assign w2001 = ( ~w255 & w324 ) | ( ~w255 & w513 ) | ( w324 & w513 ) ;
  assign w2002 = w2000 & ~w2001 ;
  assign w2003 = ~w1999 & w2002 ;
  assign w2004 = ( w283 & ~w361 ) | ( w283 & w899 ) | ( ~w361 & w899 ) ;
  assign w2005 = w361 | w2004 ;
  assign w2006 = w281 | w1130 ;
  assign w2007 = w2005 | w2006 ;
  assign w2008 = ( w98 & w1010 ) | ( w98 & ~w2005 ) | ( w1010 & ~w2005 ) ;
  assign w2009 = w2007 | w2008 ;
  assign w2010 = ( ~w354 & w997 ) | ( ~w354 & w1990 ) | ( w997 & w1990 ) ;
  assign w2011 = w2003 & ~w2009 ;
  assign w2012 = ( w354 & w534 ) | ( w354 & ~w2009 ) | ( w534 & ~w2009 ) ;
  assign w2013 = w2011 & ~w2012 ;
  assign w2014 = ~w2010 & w2013 ;
  assign w2015 = ( w219 & w265 ) | ( w219 & ~w802 ) | ( w265 & ~w802 ) ;
  assign w2016 = ~w84 & w2014 ;
  assign w2017 = ( ~w84 & w802 ) | ( ~w84 & w1229 ) | ( w802 & w1229 ) ;
  assign w2018 = w2016 & ~w2017 ;
  assign w2019 = ~w2015 & w2018 ;
  assign w2020 = w44 | w1030 ;
  assign w2021 = ( w44 & ~w198 ) | ( w44 & w2019 ) | ( ~w198 & w2019 ) ;
  assign w2022 = ~w2020 & w2021 ;
  assign w2023 = w641 | w783 ;
  assign w2024 = w445 | w2023 ;
  assign w2025 = ( w86 & ~w445 ) | ( w86 & w466 ) | ( ~w445 & w466 ) ;
  assign w2026 = w2024 | w2025 ;
  assign w2027 = w511 | w2026 ;
  assign w2028 = ( w225 & w1208 ) | ( w225 & ~w2026 ) | ( w1208 & ~w2026 ) ;
  assign w2029 = w2027 | w2028 ;
  assign w2030 = w385 | w623 ;
  assign w2031 = w911 | w2030 ;
  assign w2032 = ( w353 & ~w911 ) | ( w353 & w2029 ) | ( ~w911 & w2029 ) ;
  assign w2033 = w2031 | w2032 ;
  assign w2034 = ( ~w345 & w524 ) | ( ~w345 & w2033 ) | ( w524 & w2033 ) ;
  assign w2035 = w345 | w2034 ;
  assign w2036 = ( ~w88 & w196 ) | ( ~w88 & w492 ) | ( w196 & w492 ) ;
  assign w2037 = w88 | w2036 ;
  assign w2038 = ( w59 & ~w447 ) | ( w59 & w1276 ) | ( ~w447 & w1276 ) ;
  assign w2039 = w410 | w2037 ;
  assign w2040 = ( ~w410 & w447 ) | ( ~w410 & w664 ) | ( w447 & w664 ) ;
  assign w2041 = w2039 | w2040 ;
  assign w2042 = w2038 | w2041 ;
  assign w2043 = w890 | w1987 ;
  assign w2044 = w2022 & ~w2043 ;
  assign w2045 = ( w2022 & w2035 ) | ( w2022 & w2042 ) | ( w2035 & w2042 ) ;
  assign w2046 = w2044 & ~w2045 ;
  assign w2047 = w1978 | w1979 ;
  assign w2048 = w514 | w2047 ;
  assign w2049 = ( w514 & ~w1977 ) | ( w514 & w2046 ) | ( ~w1977 & w2046 ) ;
  assign w2050 = ~w2048 & w2049 ;
  assign w2051 = w408 | w561 ;
  assign w2052 = w1615 | w2051 ;
  assign w2053 = ( ~w262 & w1615 ) | ( ~w262 & w2050 ) | ( w1615 & w2050 ) ;
  assign w2054 = ~w2052 & w2053 ;
  assign w2055 = ( w275 & w278 ) | ( w275 & ~w418 ) | ( w278 & ~w418 ) ;
  assign w2056 = ~w252 & w2054 ;
  assign w2057 = ( ~w252 & w418 ) | ( ~w252 & w505 ) | ( w418 & w505 ) ;
  assign w2058 = w2056 & ~w2057 ;
  assign w2059 = ~w2055 & w2058 ;
  assign w2060 = w284 | w1128 ;
  assign w2061 = ( w275 & w388 ) | ( w275 & ~w511 ) | ( w388 & ~w511 ) ;
  assign w2062 = w128 | w139 ;
  assign w2063 = ( ~w139 & w511 ) | ( ~w139 & w593 ) | ( w511 & w593 ) ;
  assign w2064 = w2062 | w2063 ;
  assign w2065 = w2061 | w2064 ;
  assign w2066 = ( w131 & ~w223 ) | ( w131 & w2065 ) | ( ~w223 & w2065 ) ;
  assign w2067 = w279 | w2060 ;
  assign w2068 = ( w223 & w1126 ) | ( w223 & ~w2060 ) | ( w1126 & ~w2060 ) ;
  assign w2069 = w2067 | w2068 ;
  assign w2070 = w2066 | w2069 ;
  assign w2071 = ( w179 & w488 ) | ( w179 & ~w889 ) | ( w488 & ~w889 ) ;
  assign w2072 = w165 | w2070 ;
  assign w2073 = ( ~w165 & w889 ) | ( ~w165 & w1153 ) | ( w889 & w1153 ) ;
  assign w2074 = w2072 | w2073 ;
  assign w2075 = w2071 | w2074 ;
  assign w2076 = w534 | w674 ;
  assign w2077 = w456 | w2076 ;
  assign w2078 = ( w98 & ~w456 ) | ( w98 & w491 ) | ( ~w456 & w491 ) ;
  assign w2079 = w2077 | w2078 ;
  assign w2080 = ~w317 & w359 ;
  assign w2081 = ( ~w317 & w318 ) | ( ~w317 & w999 ) | ( w318 & w999 ) ;
  assign w2082 = w2080 & ~w2081 ;
  assign w2083 = ( w219 & w325 ) | ( w219 & ~w449 ) | ( w325 & ~w449 ) ;
  assign w2084 = w136 | w1131 ;
  assign w2085 = ( ~w136 & w449 ) | ( ~w136 & w1031 ) | ( w449 & w1031 ) ;
  assign w2086 = w2084 | w2085 ;
  assign w2087 = w2083 | w2086 ;
  assign w2088 = w342 | w509 ;
  assign w2089 = ( w116 & ~w342 ) | ( w116 & w358 ) | ( ~w342 & w358 ) ;
  assign w2090 = w2088 | w2089 ;
  assign w2091 = w133 | w726 ;
  assign w2092 = w59 | w758 ;
  assign w2093 = w351 | w415 ;
  assign w2094 = ( w180 & ~w351 ) | ( w180 & w352 ) | ( ~w351 & w352 ) ;
  assign w2095 = w2093 | w2094 ;
  assign w2096 = w198 | w431 ;
  assign w2097 = ( ~w118 & w2095 ) | ( ~w118 & w2096 ) | ( w2095 & w2096 ) ;
  assign w2098 = w527 | w1740 ;
  assign w2099 = ( w118 & w606 ) | ( w118 & ~w1740 ) | ( w606 & ~w1740 ) ;
  assign w2100 = w2098 | w2099 ;
  assign w2101 = w2097 | w2100 ;
  assign w2102 = w1363 | w2092 ;
  assign w2103 = ( ~w1363 & w2091 ) | ( ~w1363 & w2101 ) | ( w2091 & w2101 ) ;
  assign w2104 = w2102 | w2103 ;
  assign w2105 = w229 | w625 ;
  assign w2106 = w1713 | w2105 ;
  assign w2107 = ( w119 & ~w1713 ) | ( w119 & w2104 ) | ( ~w1713 & w2104 ) ;
  assign w2108 = w2106 | w2107 ;
  assign w2109 = w465 | w571 ;
  assign w2110 = w167 | w2109 ;
  assign w2111 = ( ~w167 & w430 ) | ( ~w167 & w2108 ) | ( w430 & w2108 ) ;
  assign w2112 = w2110 | w2111 ;
  assign w2113 = ( w1208 & w2082 ) | ( w1208 & ~w2087 ) | ( w2082 & ~w2087 ) ;
  assign w2114 = w1645 | w2112 ;
  assign w2115 = ( w1208 & w2090 ) | ( w1208 & ~w2112 ) | ( w2090 & ~w2112 ) ;
  assign w2116 = w2114 | w2115 ;
  assign w2117 = w2113 & ~w2116 ;
  assign w2118 = ( ~w266 & w731 ) | ( ~w266 & w2079 ) | ( w731 & w2079 ) ;
  assign w2119 = ~w2075 & w2117 ;
  assign w2120 = ( w266 & w561 ) | ( w266 & ~w2075 ) | ( w561 & ~w2075 ) ;
  assign w2121 = w2119 & ~w2120 ;
  assign w2122 = ~w2118 & w2121 ;
  assign w2123 = w178 | w513 ;
  assign w2124 = ( w178 & ~w339 ) | ( w178 & w2122 ) | ( ~w339 & w2122 ) ;
  assign w2125 = ~w2123 & w2124 ;
  assign w2126 = ( w272 & w418 ) | ( w272 & ~w467 ) | ( w418 & ~w467 ) ;
  assign w2127 = ~w68 & w2125 ;
  assign w2128 = ( ~w68 & w467 ) | ( ~w68 & w565 ) | ( w467 & w565 ) ;
  assign w2129 = w2127 & ~w2128 ;
  assign w2130 = ~w2126 & w2129 ;
  assign w2131 = ( w169 & w490 ) | ( w169 & ~w533 ) | ( w490 & ~w533 ) ;
  assign w2132 = w122 | w164 ;
  assign w2133 = ( ~w164 & w533 ) | ( ~w164 & w663 ) | ( w533 & w663 ) ;
  assign w2134 = w2132 | w2133 ;
  assign w2135 = w2131 | w2134 ;
  assign w2136 = ( w209 & w280 ) | ( w209 & ~w496 ) | ( w280 & ~w496 ) ;
  assign w2137 = w113 | w2135 ;
  assign w2138 = ( ~w113 & w496 ) | ( ~w113 & w821 ) | ( w496 & w821 ) ;
  assign w2139 = w2137 | w2138 ;
  assign w2140 = w2136 | w2139 ;
  assign w2141 = ( ~w320 & w637 ) | ( ~w320 & w2140 ) | ( w637 & w2140 ) ;
  assign w2142 = w320 | w2141 ;
  assign w2143 = w271 | w488 ;
  assign w2144 = w1281 | w2143 ;
  assign w2145 = ( w232 & w1276 ) | ( w232 & ~w1281 ) | ( w1276 & ~w1281 ) ;
  assign w2146 = w2144 | w2145 ;
  assign w2147 = w141 | w640 ;
  assign w2148 = w1128 | w1130 ;
  assign w2149 = w2147 | w2148 ;
  assign w2150 = ( w225 & w1837 ) | ( w225 & ~w2147 ) | ( w1837 & ~w2147 ) ;
  assign w2151 = w2149 | w2150 ;
  assign w2152 = ( ~w118 & w409 ) | ( ~w118 & w2151 ) | ( w409 & w2151 ) ;
  assign w2153 = w118 | w2152 ;
  assign w2154 = w256 | w530 ;
  assign w2155 = w181 | w2154 ;
  assign w2156 = ( ~w181 & w1158 ) | ( ~w181 & w2153 ) | ( w1158 & w2153 ) ;
  assign w2157 = w2155 | w2156 ;
  assign w2158 = ( w220 & ~w318 ) | ( w220 & w2146 ) | ( ~w318 & w2146 ) ;
  assign w2159 = w2142 | w2157 ;
  assign w2160 = ( w318 & w783 ) | ( w318 & ~w2142 ) | ( w783 & ~w2142 ) ;
  assign w2161 = w2159 | w2160 ;
  assign w2162 = w2158 | w2161 ;
  assign w2163 = ( w386 & w411 ) | ( w386 & ~w560 ) | ( w411 & ~w560 ) ;
  assign w2164 = w514 | w2162 ;
  assign w2165 = ( ~w514 & w560 ) | ( ~w514 & w605 ) | ( w560 & w605 ) ;
  assign w2166 = w2164 | w2165 ;
  assign w2167 = w2163 | w2166 ;
  assign w2168 = w111 | w642 ;
  assign w2169 = w350 | w561 ;
  assign w2170 = w138 | w506 ;
  assign w2171 = w199 | w2170 ;
  assign w2172 = ( w63 & w2169 ) | ( w63 & ~w2170 ) | ( w2169 & ~w2170 ) ;
  assign w2173 = w2171 | w2172 ;
  assign w2174 = ( w119 & ~w313 ) | ( w119 & w2168 ) | ( ~w313 & w2168 ) ;
  assign w2175 = w1155 | w2173 ;
  assign w2176 = ( w313 & w351 ) | ( w313 & ~w1155 ) | ( w351 & ~w1155 ) ;
  assign w2177 = w2175 | w2176 ;
  assign w2178 = w2174 | w2177 ;
  assign w2179 = ( w359 & ~w383 ) | ( w359 & w524 ) | ( ~w383 & w524 ) ;
  assign w2180 = w135 | w2178 ;
  assign w2181 = ( ~w135 & w524 ) | ( ~w135 & w899 ) | ( w524 & w899 ) ;
  assign w2182 = w2180 | w2181 ;
  assign w2183 = w2179 & ~w2182 ;
  assign w2184 = w606 | w674 ;
  assign w2185 = w206 | w2184 ;
  assign w2186 = ( w81 & ~w206 ) | ( w81 & w420 ) | ( ~w206 & w420 ) ;
  assign w2187 = w2185 | w2186 ;
  assign w2188 = w142 | w317 ;
  assign w2189 = ( ~w142 & w224 ) | ( ~w142 & w2187 ) | ( w224 & w2187 ) ;
  assign w2190 = w2188 | w2189 ;
  assign w2191 = ( w115 & w203 ) | ( w115 & ~w509 ) | ( w203 & ~w509 ) ;
  assign w2192 = w1154 | w1687 ;
  assign w2193 = ( w509 & w1094 ) | ( w509 & ~w1687 ) | ( w1094 & ~w1687 ) ;
  assign w2194 = w2192 | w2193 ;
  assign w2195 = w2191 | w2194 ;
  assign w2196 = w390 | w680 ;
  assign w2197 = w2195 | w2196 ;
  assign w2198 = ( w1940 & w2190 ) | ( w1940 & ~w2195 ) | ( w2190 & ~w2195 ) ;
  assign w2199 = w2197 | w2198 ;
  assign w2200 = w68 | w74 ;
  assign w2201 = w1087 | w2200 ;
  assign w2202 = ( ~w1087 & w2091 ) | ( ~w1087 & w2199 ) | ( w2091 & w2199 ) ;
  assign w2203 = w2201 | w2202 ;
  assign w2204 = ( w269 & w513 ) | ( w269 & ~w596 ) | ( w513 & ~w596 ) ;
  assign w2205 = w178 | w2203 ;
  assign w2206 = ( ~w178 & w596 ) | ( ~w178 & w723 ) | ( w596 & w723 ) ;
  assign w2207 = w2205 | w2206 ;
  assign w2208 = w2204 | w2207 ;
  assign w2209 = ( w388 & w525 ) | ( w388 & ~w569 ) | ( w525 & ~w569 ) ;
  assign w2210 = w223 | w322 ;
  assign w2211 = ( ~w322 & w569 ) | ( ~w322 & w628 ) | ( w569 & w628 ) ;
  assign w2212 = w2210 | w2211 ;
  assign w2213 = w2209 | w2212 ;
  assign w2214 = ( w470 & w512 ) | ( w470 & ~w1031 ) | ( w512 & ~w1031 ) ;
  assign w2215 = w161 | w325 ;
  assign w2216 = ( ~w325 & w1031 ) | ( ~w325 & w1086 ) | ( w1031 & w1086 ) ;
  assign w2217 = w2215 | w2216 ;
  assign w2218 = w2214 | w2217 ;
  assign w2219 = ( w87 & w1280 ) | ( w87 & ~w2213 ) | ( w1280 & ~w2213 ) ;
  assign w2220 = w2183 & ~w2208 ;
  assign w2221 = ( w2183 & w2213 ) | ( w2183 & w2218 ) | ( w2213 & w2218 ) ;
  assign w2222 = w2220 & ~w2221 ;
  assign w2223 = ~w2219 & w2222 ;
  assign w2224 = ( w120 & ~w125 ) | ( w120 & w343 ) | ( ~w125 & w343 ) ;
  assign w2225 = ~w2167 & w2223 ;
  assign w2226 = ( w125 & w515 ) | ( w125 & w2223 ) | ( w515 & w2223 ) ;
  assign w2227 = w2225 & ~w2226 ;
  assign w2228 = ~w2224 & w2227 ;
  assign w2229 = ( w310 & w354 ) | ( w310 & ~w429 ) | ( w354 & ~w429 ) ;
  assign w2230 = ~w98 & w2228 ;
  assign w2231 = ( ~w98 & w429 ) | ( ~w98 & w458 ) | ( w429 & w458 ) ;
  assign w2232 = w2230 & ~w2231 ;
  assign w2233 = ~w2229 & w2232 ;
  assign w2234 = ( w571 & ~w662 ) | ( w571 & w2233 ) | ( ~w662 & w2233 ) ;
  assign w2235 = ~w571 & w2234 ;
  assign w2236 = ( w84 & w530 ) | ( w84 & ~w1094 ) | ( w530 & ~w1094 ) ;
  assign w2237 = w1362 | w1951 ;
  assign w2238 = ( w1094 & w1340 ) | ( w1094 & ~w1362 ) | ( w1340 & ~w1362 ) ;
  assign w2239 = w2237 | w2238 ;
  assign w2240 = w2236 | w2239 ;
  assign w2241 = ( ~w169 & w1154 ) | ( ~w169 & w2147 ) | ( w1154 & w2147 ) ;
  assign w2242 = w326 | w2240 ;
  assign w2243 = ( w169 & ~w326 ) | ( w169 & w1274 ) | ( ~w326 & w1274 ) ;
  assign w2244 = w2242 | w2243 ;
  assign w2245 = w2241 | w2244 ;
  assign w2246 = ( w253 & w344 ) | ( w253 & ~w429 ) | ( w344 & ~w429 ) ;
  assign w2247 = w111 | w2245 ;
  assign w2248 = ( ~w111 & w429 ) | ( ~w111 & w817 ) | ( w429 & w817 ) ;
  assign w2249 = w2247 | w2248 ;
  assign w2250 = w2246 | w2249 ;
  assign w2251 = ( w491 & ~w513 ) | ( w491 & w524 ) | ( ~w513 & w524 ) ;
  assign w2252 = w513 | w2251 ;
  assign w2253 = w383 | w1001 ;
  assign w2254 = ( w343 & w456 ) | ( w343 & ~w2253 ) | ( w456 & ~w2253 ) ;
  assign w2255 = w2253 | w2254 ;
  assign w2256 = ( w126 & w147 ) | ( w126 & ~w1954 ) | ( w147 & ~w1954 ) ;
  assign w2257 = w1954 | w2256 ;
  assign w2258 = ( w759 & ~w784 ) | ( w759 & w1166 ) | ( ~w784 & w1166 ) ;
  assign w2259 = w784 | w2258 ;
  assign w2260 = w2257 | w2259 ;
  assign w2261 = w767 | w2260 ;
  assign w2262 = ( ~w767 & w1494 ) | ( ~w767 & w2255 ) | ( w1494 & w2255 ) ;
  assign w2263 = w2261 | w2262 ;
  assign w2264 = w678 | w2252 ;
  assign w2265 = ( ~w678 & w1713 ) | ( ~w678 & w2263 ) | ( w1713 & w2263 ) ;
  assign w2266 = w2264 | w2265 ;
  assign w2267 = ( ~w257 & w416 ) | ( ~w257 & w1275 ) | ( w416 & w1275 ) ;
  assign w2268 = w2250 | w2266 ;
  assign w2269 = ( w257 & w317 ) | ( w257 & ~w2250 ) | ( w317 & ~w2250 ) ;
  assign w2270 = w2268 | w2269 ;
  assign w2271 = w2267 | w2270 ;
  assign w2272 = ( ~w221 & w723 ) | ( ~w221 & w2271 ) | ( w723 & w2271 ) ;
  assign w2273 = w221 | w2272 ;
  assign w2274 = w127 | w258 ;
  assign w2275 = w1094 | w1126 ;
  assign w2276 = w84 | w2275 ;
  assign w2277 = ( ~w84 & w113 ) | ( ~w84 & w2274 ) | ( w113 & w2274 ) ;
  assign w2278 = w2276 | w2277 ;
  assign w2279 = w1590 | w2147 ;
  assign w2280 = ( ~w1590 & w1882 ) | ( ~w1590 & w2278 ) | ( w1882 & w2278 ) ;
  assign w2281 = w2279 | w2280 ;
  assign w2282 = ( w144 & w164 ) | ( w144 & ~w257 ) | ( w164 & ~w257 ) ;
  assign w2283 = w88 | w2281 ;
  assign w2284 = ( ~w88 & w257 ) | ( ~w88 & w260 ) | ( w257 & w260 ) ;
  assign w2285 = w2283 | w2284 ;
  assign w2286 = w2282 | w2285 ;
  assign w2287 = ~\pi26 & w47 ;
  assign w2288 = \pi23 & w2287 ;
  assign w2289 = ( ~\pi24 & \pi25 ) | ( ~\pi24 & w60 ) | ( \pi25 & w60 ) ;
  assign w2290 = ( \pi23 & w47 ) | ( \pi23 & w2287 ) | ( w47 & w2287 ) ;
  assign w2291 = ( \pi24 & w60 ) | ( \pi24 & ~w112 ) | ( w60 & ~w112 ) ;
  assign w2292 = ( \pi24 & w2290 ) | ( \pi24 & w2291 ) | ( w2290 & w2291 ) ;
  assign w2293 = ( \pi25 & w2290 ) | ( \pi25 & ~w2292 ) | ( w2290 & ~w2292 ) ;
  assign w2294 = ( w2288 & ~w2289 ) | ( w2288 & w2293 ) | ( ~w2289 & w2293 ) ;
  assign w2295 = w116 | w167 ;
  assign w2296 = w724 | w980 ;
  assign w2297 = w420 | w2296 ;
  assign w2298 = ( ~w420 & w565 ) | ( ~w420 & w2295 ) | ( w565 & w2295 ) ;
  assign w2299 = w2297 | w2298 ;
  assign w2300 = ( w263 & w560 ) | ( w263 & ~w573 ) | ( w560 & ~w573 ) ;
  assign w2301 = w205 | w2299 ;
  assign w2302 = ( ~w205 & w573 ) | ( ~w205 & w726 ) | ( w573 & w726 ) ;
  assign w2303 = w2301 | w2302 ;
  assign w2304 = w2300 | w2303 ;
  assign w2305 = ( w169 & ~w625 ) | ( w169 & w837 ) | ( ~w625 & w837 ) ;
  assign w2306 = w625 | w2305 ;
  assign w2307 = ( w199 & w255 ) | ( w199 & ~w506 ) | ( w255 & ~w506 ) ;
  assign w2308 = w63 | w179 ;
  assign w2309 = ( ~w179 & w506 ) | ( ~w179 & w596 ) | ( w506 & w596 ) ;
  assign w2310 = w2308 | w2309 ;
  assign w2311 = w2307 | w2310 ;
  assign w2312 = ( w115 & w341 ) | ( w115 & ~w353 ) | ( w341 & ~w353 ) ;
  assign w2313 = w1093 | w2311 ;
  assign w2314 = ( w353 & w817 ) | ( w353 & ~w2311 ) | ( w817 & ~w2311 ) ;
  assign w2315 = w2313 | w2314 ;
  assign w2316 = w2312 | w2315 ;
  assign w2317 = ( ~w223 & w268 ) | ( ~w223 & w2316 ) | ( w268 & w2316 ) ;
  assign w2318 = w223 | w2317 ;
  assign w2319 = w214 | w456 ;
  assign w2320 = w101 | w764 ;
  assign w2321 = w2319 | w2320 ;
  assign w2322 = ( w98 & w2005 ) | ( w98 & ~w2319 ) | ( w2005 & ~w2319 ) ;
  assign w2323 = w2321 | w2322 ;
  assign w2324 = w409 | w449 ;
  assign w2325 = w163 | w2324 ;
  assign w2326 = ( ~w163 & w384 ) | ( ~w163 & w2323 ) | ( w384 & w2323 ) ;
  assign w2327 = w2325 | w2326 ;
  assign w2328 = w466 | w567 ;
  assign w2329 = w74 | w2328 ;
  assign w2330 = ( ~w74 & w201 ) | ( ~w74 & w1814 ) | ( w201 & w1814 ) ;
  assign w2331 = w2329 | w2330 ;
  assign w2332 = w413 | w505 ;
  assign w2333 = w133 | w2332 ;
  assign w2334 = ( ~w133 & w339 ) | ( ~w133 & w2331 ) | ( w339 & w2331 ) ;
  assign w2335 = w2333 | w2334 ;
  assign w2336 = ( w820 & ~w2060 ) | ( w820 & w2335 ) | ( ~w2060 & w2335 ) ;
  assign w2337 = w2318 | w2327 ;
  assign w2338 = ( w2060 & w2306 ) | ( w2060 & ~w2327 ) | ( w2306 & ~w2327 ) ;
  assign w2339 = w2337 | w2338 ;
  assign w2340 = w2336 | w2339 ;
  assign w2341 = ( w104 & ~w642 ) | ( w104 & w1421 ) | ( ~w642 & w1421 ) ;
  assign w2342 = w82 | w2340 ;
  assign w2343 = ( ~w82 & w642 ) | ( ~w82 & w723 ) | ( w642 & w723 ) ;
  assign w2344 = w2342 | w2343 ;
  assign w2345 = w2341 | w2344 ;
  assign w2346 = ( w272 & w274 ) | ( w272 & ~w386 ) | ( w274 & ~w386 ) ;
  assign w2347 = w225 | w2345 ;
  assign w2348 = ( ~w225 & w386 ) | ( ~w225 & w569 ) | ( w386 & w569 ) ;
  assign w2349 = w2347 | w2348 ;
  assign w2350 = w2346 | w2349 ;
  assign w2351 = w423 | w512 ;
  assign w2352 = w1884 | w2351 ;
  assign w2353 = ( w218 & w624 ) | ( w218 & ~w1884 ) | ( w624 & ~w1884 ) ;
  assign w2354 = w2352 | w2353 ;
  assign w2355 = w470 | w524 ;
  assign w2356 = w254 | w2355 ;
  assign w2357 = ( w215 & ~w254 ) | ( w215 & w358 ) | ( ~w254 & w358 ) ;
  assign w2358 = w2356 | w2357 ;
  assign w2359 = \pi23 ^ \pi25 ;
  assign w2360 = w174 & w2359 ;
  assign w2361 = ~\pi25 & w2360 ;
  assign w2362 = ( \pi24 & ~w2359 ) | ( \pi24 & w2361 ) | ( ~w2359 & w2361 ) ;
  assign w2363 = ( w130 & w2360 ) | ( w130 & ~w2362 ) | ( w2360 & ~w2362 ) ;
  assign w2364 = \pi23 | \pi25 ;
  assign w2365 = \pi24 & w2364 ;
  assign w2366 = ( w174 & ~w2364 ) | ( w174 & w2365 ) | ( ~w2364 & w2365 ) ;
  assign w2367 = ( ~\pi23 & \pi25 ) | ( ~\pi23 & w130 ) | ( \pi25 & w130 ) ;
  assign w2368 = w357 & w2367 ;
  assign w2369 = w2366 | w2368 ;
  assign w2370 = \pi26 ^ w2363 ;
  assign w2371 = ( w2363 & w2369 ) | ( w2363 & w2370 ) | ( w2369 & w2370 ) ;
  assign w2372 = ( w128 & ~w202 ) | ( w128 & w2371 ) | ( ~w202 & w2371 ) ;
  assign w2373 = w202 | w2372 ;
  assign w2374 = w496 | w605 ;
  assign w2375 = ( ~w122 & w344 ) | ( ~w122 & w2374 ) | ( w344 & w2374 ) ;
  assign w2376 = w122 | w2375 ;
  assign w2377 = w351 | w2373 ;
  assign w2378 = ( w350 & ~w2373 ) | ( w350 & w2376 ) | ( ~w2373 & w2376 ) ;
  assign w2379 = w2377 | w2378 ;
  assign w2380 = ( ~w758 & w1301 ) | ( ~w758 & w2354 ) | ( w1301 & w2354 ) ;
  assign w2381 = w2350 | w2379 ;
  assign w2382 = ( w758 & w821 ) | ( w758 & ~w2379 ) | ( w821 & ~w2379 ) ;
  assign w2383 = w2381 | w2382 ;
  assign w2384 = w2380 | w2383 ;
  assign w2385 = w510 | w2294 ;
  assign w2386 = w2286 | w2385 ;
  assign w2387 = ( ~w2286 & w2304 ) | ( ~w2286 & w2384 ) | ( w2304 & w2384 ) ;
  assign w2388 = w2386 | w2387 ;
  assign w2389 = w232 | w626 ;
  assign w2390 = ( ~w232 & w342 ) | ( ~w232 & w2388 ) | ( w342 & w2388 ) ;
  assign w2391 = w2389 | w2390 ;
  assign w2392 = w467 | w534 ;
  assign w2393 = w221 | w2392 ;
  assign w2394 = ( w205 & ~w221 ) | ( w205 & w353 ) | ( ~w221 & w353 ) ;
  assign w2395 = w2393 | w2394 ;
  assign w2396 = ( w119 & w272 ) | ( w119 & ~w456 ) | ( w272 & ~w456 ) ;
  assign w2397 = w115 | w838 ;
  assign w2398 = ( ~w115 & w456 ) | ( ~w115 & w860 ) | ( w456 & w860 ) ;
  assign w2399 = w2397 | w2398 ;
  assign w2400 = w2396 | w2399 ;
  assign w2401 = w209 | w758 ;
  assign w2402 = ( ~w209 & w316 ) | ( ~w209 & w1157 ) | ( w316 & w1157 ) ;
  assign w2403 = w2401 | w2402 ;
  assign w2404 = w255 | w2403 ;
  assign w2405 = ( w124 & w1568 ) | ( w124 & ~w2403 ) | ( w1568 & ~w2403 ) ;
  assign w2406 = w2404 | w2405 ;
  assign w2407 = w626 | w680 ;
  assign w2408 = w181 | w2407 ;
  assign w2409 = ( w141 & ~w181 ) | ( w141 & w2406 ) | ( ~w181 & w2406 ) ;
  assign w2410 = w2408 | w2409 ;
  assign w2411 = ( w1882 & w2169 ) | ( w1882 & ~w2252 ) | ( w2169 & ~w2252 ) ;
  assign w2412 = w2400 | w2410 ;
  assign w2413 = ( w2252 & w2395 ) | ( w2252 & ~w2400 ) | ( w2395 & ~w2400 ) ;
  assign w2414 = w2412 | w2413 ;
  assign w2415 = w2411 | w2414 ;
  assign w2416 = ( w269 & w608 ) | ( w269 & ~w787 ) | ( w608 & ~w787 ) ;
  assign w2417 = w206 | w2415 ;
  assign w2418 = ( ~w206 & w787 ) | ( ~w206 & w1130 ) | ( w787 & w1130 ) ;
  assign w2419 = w2417 | w2418 ;
  assign w2420 = w2416 | w2419 ;
  assign w2421 = ( w262 & w274 ) | ( w262 & ~w341 ) | ( w274 & ~w341 ) ;
  assign w2422 = w143 | w257 ;
  assign w2423 = ( ~w257 & w341 ) | ( ~w257 & w408 ) | ( w341 & w408 ) ;
  assign w2424 = w2422 | w2423 ;
  assign w2425 = w2421 | w2424 ;
  assign w2426 = w135 | w569 ;
  assign w2427 = ( ~w135 & w167 ) | ( ~w135 & w2425 ) | ( w167 & w2425 ) ;
  assign w2428 = w2426 | w2427 ;
  assign w2429 = ( w344 & w429 ) | ( w344 & ~w430 ) | ( w429 & ~w430 ) ;
  assign w2430 = w283 | w324 ;
  assign w2431 = ( ~w324 & w430 ) | ( ~w324 & w664 ) | ( w430 & w664 ) ;
  assign w2432 = w2430 | w2431 ;
  assign w2433 = w2429 | w2432 ;
  assign w2434 = w161 | w2433 ;
  assign w2435 = w420 | w565 ;
  assign w2436 = w229 | w2435 ;
  assign w2437 = ( w138 & ~w229 ) | ( w138 & w315 ) | ( ~w229 & w315 ) ;
  assign w2438 = w2436 | w2437 ;
  assign w2439 = w320 | w674 ;
  assign w2440 = ( ~w320 & w605 ) | ( ~w320 & w2438 ) | ( w605 & w2438 ) ;
  assign w2441 = w2439 | w2440 ;
  assign w2442 = ( ~w68 & w216 ) | ( ~w68 & w2441 ) | ( w216 & w2441 ) ;
  assign w2443 = w2428 | w2434 ;
  assign w2444 = ( w68 & w220 ) | ( w68 & ~w2434 ) | ( w220 & ~w2434 ) ;
  assign w2445 = w2443 | w2444 ;
  assign w2446 = w2442 | w2445 ;
  assign w2447 = ( w125 & w340 ) | ( w125 & ~w413 ) | ( w340 & ~w413 ) ;
  assign w2448 = w911 | w2446 ;
  assign w2449 = ( w413 & ~w911 ) | ( w413 & w1153 ) | ( ~w911 & w1153 ) ;
  assign w2450 = w2448 | w2449 ;
  assign w2451 = w2447 | w2450 ;
  assign w2452 = w567 | w681 ;
  assign w2453 = ( w593 & w897 ) | ( w593 & ~w1274 ) | ( w897 & ~w1274 ) ;
  assign w2454 = w74 | w418 ;
  assign w2455 = ( ~w418 & w1274 ) | ( ~w418 & w1340 ) | ( w1274 & w1340 ) ;
  assign w2456 = w2454 | w2455 ;
  assign w2457 = w2453 | w2456 ;
  assign w2458 = ( w219 & w465 ) | ( w219 & ~w980 ) | ( w465 & ~w980 ) ;
  assign w2459 = w218 | w2457 ;
  assign w2460 = ( ~w218 & w980 ) | ( ~w218 & w1128 ) | ( w980 & w1128 ) ;
  assign w2461 = w2459 | w2460 ;
  assign w2462 = w2458 | w2461 ;
  assign w2463 = w311 | w2452 ;
  assign w2464 = ( w147 & ~w2452 ) | ( w147 & w2462 ) | ( ~w2452 & w2462 ) ;
  assign w2465 = w2463 | w2464 ;
  assign w2466 = w596 | w1229 ;
  assign w2467 = w424 | w2466 ;
  assign w2468 = ( ~w424 & w470 ) | ( ~w424 & w2465 ) | ( w470 & w2465 ) ;
  assign w2469 = w2467 | w2468 ;
  assign w2470 = w284 | w531 ;
  assign w2471 = w263 | w515 ;
  assign w2472 = w56 | w2471 ;
  assign w2473 = ( ~w56 & w111 ) | ( ~w56 & w2470 ) | ( w111 & w2470 ) ;
  assign w2474 = w2472 | w2473 ;
  assign w2475 = ( w345 & w492 ) | ( w345 & ~w802 ) | ( w492 & ~w802 ) ;
  assign w2476 = w116 | w2474 ;
  assign w2477 = ( ~w116 & w802 ) | ( ~w116 & w889 ) | ( w802 & w889 ) ;
  assign w2478 = w2476 | w2477 ;
  assign w2479 = w2475 | w2478 ;
  assign w2480 = w312 | w571 ;
  assign w2481 = ( w88 & w131 ) | ( w88 & ~w223 ) | ( w131 & ~w223 ) ;
  assign w2482 = w289 | w2480 ;
  assign w2483 = ( w223 & w533 ) | ( w223 & ~w2480 ) | ( w533 & ~w2480 ) ;
  assign w2484 = w2482 | w2483 ;
  assign w2485 = w2481 | w2484 ;
  assign w2486 = ( w2469 & w2479 ) | ( w2469 & ~w2485 ) | ( w2479 & ~w2485 ) ;
  assign w2487 = w2420 | w2451 ;
  assign w2488 = ( w1712 & ~w2451 ) | ( w1712 & w2485 ) | ( ~w2451 & w2485 ) ;
  assign w2489 = w2487 | w2488 ;
  assign w2490 = w2486 | w2489 ;
  assign w2491 = ( w164 & ~w201 ) | ( w164 & w1281 ) | ( ~w201 & w1281 ) ;
  assign w2492 = w956 | w2490 ;
  assign w2493 = ( w201 & w459 ) | ( w201 & ~w956 ) | ( w459 & ~w956 ) ;
  assign w2494 = w2492 | w2493 ;
  assign w2495 = w2491 | w2494 ;
  assign w2496 = ( w208 & w309 ) | ( w208 & ~w725 ) | ( w309 & ~w725 ) ;
  assign w2497 = w127 | w2495 ;
  assign w2498 = ( ~w127 & w725 ) | ( ~w127 & w901 ) | ( w725 & w901 ) ;
  assign w2499 = w2497 | w2498 ;
  assign w2500 = w2496 | w2499 ;
  assign w2501 = w144 | w568 ;
  assign w2502 = w1413 | w2501 ;
  assign w2503 = ( w349 & ~w1413 ) | ( w349 & w1940 ) | ( ~w1413 & w1940 ) ;
  assign w2504 = w2502 | w2503 ;
  assign w2505 = ( w90 & w143 ) | ( w90 & ~w511 ) | ( w143 & ~w511 ) ;
  assign w2506 = w1814 | w2504 ;
  assign w2507 = ( w511 & w764 ) | ( w511 & ~w1814 ) | ( w764 & ~w1814 ) ;
  assign w2508 = w2506 | w2507 ;
  assign w2509 = w2505 | w2508 ;
  assign w2510 = ( w272 & w409 ) | ( w272 & ~w534 ) | ( w409 & ~w534 ) ;
  assign w2511 = w84 | w2509 ;
  assign w2512 = ( ~w84 & w534 ) | ( ~w84 & w787 ) | ( w534 & w787 ) ;
  assign w2513 = w2511 | w2512 ;
  assign w2514 = w2510 | w2513 ;
  assign w2515 = w175 | w1153 ;
  assign w2516 = ( ~w175 & w254 ) | ( ~w175 & w2514 ) | ( w254 & w2514 ) ;
  assign w2517 = w2515 | w2516 ;
  assign w2518 = w63 | w445 ;
  assign w2519 = w274 | w897 ;
  assign w2520 = ( w255 & ~w274 ) | ( w255 & w422 ) | ( ~w274 & w422 ) ;
  assign w2521 = w2519 | w2520 ;
  assign w2522 = w116 | w253 ;
  assign w2523 = w641 | w837 ;
  assign w2524 = w515 | w2523 ;
  assign w2525 = ( ~w515 & w570 ) | ( ~w515 & w2522 ) | ( w570 & w2522 ) ;
  assign w2526 = w2524 | w2525 ;
  assign w2527 = w359 & ~w593 ;
  assign w2528 = ~w114 & w2527 ;
  assign w2529 = ( ~w114 & w219 ) | ( ~w114 & w2526 ) | ( w219 & w2526 ) ;
  assign w2530 = w2528 & ~w2529 ;
  assign w2531 = ( w595 & w640 ) | ( w595 & ~w1128 ) | ( w640 & ~w1128 ) ;
  assign w2532 = w179 | w467 ;
  assign w2533 = ( ~w467 & w1128 ) | ( ~w467 & w1229 ) | ( w1128 & w1229 ) ;
  assign w2534 = w2532 | w2533 ;
  assign w2535 = w2531 | w2534 ;
  assign w2536 = w86 | w111 ;
  assign w2537 = w951 | w1086 ;
  assign w2538 = w225 | w2537 ;
  assign w2539 = ( w126 & ~w225 ) | ( w126 & w354 ) | ( ~w225 & w354 ) ;
  assign w2540 = w2538 | w2539 ;
  assign w2541 = w199 | w411 ;
  assign w2542 = w2535 | w2541 ;
  assign w2543 = ( ~w2535 & w2536 ) | ( ~w2535 & w2540 ) | ( w2536 & w2540 ) ;
  assign w2544 = w2542 | w2543 ;
  assign w2545 = w214 | w1275 ;
  assign w2546 = w2544 | w2545 ;
  assign w2547 = ( ~w1157 & w2530 ) | ( ~w1157 & w2544 ) | ( w2530 & w2544 ) ;
  assign w2548 = ~w2546 & w2547 ;
  assign w2549 = w266 | w443 ;
  assign w2550 = w98 | w2549 ;
  assign w2551 = ( w98 & ~w220 ) | ( w98 & w2548 ) | ( ~w220 & w2548 ) ;
  assign w2552 = ~w2550 & w2551 ;
  assign w2553 = ( w270 & ~w423 ) | ( w270 & w2552 ) | ( ~w423 & w2552 ) ;
  assign w2554 = ~w270 & w2553 ;
  assign w2555 = ( w283 & ~w722 ) | ( w283 & w802 ) | ( ~w722 & w802 ) ;
  assign w2556 = w722 | w2555 ;
  assign w2557 = ( ~w419 & w664 ) | ( ~w419 & w2556 ) | ( w664 & w2556 ) ;
  assign w2558 = w419 | w2557 ;
  assign w2559 = w2521 | w2558 ;
  assign w2560 = ( ~w800 & w2554 ) | ( ~w800 & w2558 ) | ( w2554 & w2558 ) ;
  assign w2561 = ~w2559 & w2560 ;
  assign w2562 = w672 | w2112 ;
  assign w2563 = ( ~w609 & w2112 ) | ( ~w609 & w2561 ) | ( w2112 & w2561 ) ;
  assign w2564 = ~w2562 & w2563 ;
  assign w2565 = w311 | w389 ;
  assign w2566 = w1712 | w2565 ;
  assign w2567 = ( w1712 & ~w2518 ) | ( w1712 & w2564 ) | ( ~w2518 & w2564 ) ;
  assign w2568 = ~w2566 & w2567 ;
  assign w2569 = ( w210 & ~w458 ) | ( w210 & w2142 ) | ( ~w458 & w2142 ) ;
  assign w2570 = ~w2517 & w2568 ;
  assign w2571 = ( w458 & w723 ) | ( w458 & ~w2517 ) | ( w723 & ~w2517 ) ;
  assign w2572 = w2570 & ~w2571 ;
  assign w2573 = ~w2569 & w2572 ;
  assign w2574 = ( w322 & w531 ) | ( w322 & ~w628 ) | ( w531 & ~w628 ) ;
  assign w2575 = ~w127 & w2573 ;
  assign w2576 = ( ~w127 & w628 ) | ( ~w127 & w673 ) | ( w628 & w673 ) ;
  assign w2577 = w2575 & ~w2576 ;
  assign w2578 = ~w2574 & w2577 ;
  assign w2579 = w492 | w495 ;
  assign w2580 = w229 | w2579 ;
  assign w2581 = ( w177 & ~w229 ) | ( w177 & w463 ) | ( ~w229 & w463 ) ;
  assign w2582 = w2580 | w2581 ;
  assign w2583 = ( w341 & w352 ) | ( w341 & ~w383 ) | ( w352 & ~w383 ) ;
  assign w2584 = w730 | w2582 ;
  assign w2585 = ( w383 & w697 ) | ( w383 & ~w730 ) | ( w697 & ~w730 ) ;
  assign w2586 = w2584 | w2585 ;
  assign w2587 = w2583 | w2586 ;
  assign w2588 = w465 | w980 ;
  assign w2589 = w286 | w2588 ;
  assign w2590 = ( ~w286 & w445 ) | ( ~w286 & w2587 ) | ( w445 & w2587 ) ;
  assign w2591 = w2589 | w2590 ;
  assign w2592 = ( w232 & w272 ) | ( w232 & ~w386 ) | ( w272 & ~w386 ) ;
  assign w2593 = w168 | w2591 ;
  assign w2594 = ( ~w168 & w386 ) | ( ~w168 & w623 ) | ( w386 & w623 ) ;
  assign w2595 = w2593 | w2594 ;
  assign w2596 = w2592 | w2595 ;
  assign w2597 = w524 | w662 ;
  assign w2598 = w128 | w2597 ;
  assign w2599 = ( ~w128 & w265 ) | ( ~w128 & w2596 ) | ( w265 & w2596 ) ;
  assign w2600 = w2598 | w2599 ;
  assign w2601 = w490 | w608 ;
  assign w2602 = ( w361 & ~w490 ) | ( w361 & w513 ) | ( ~w490 & w513 ) ;
  assign w2603 = w2601 | w2602 ;
  assign w2604 = ( w350 & w351 ) | ( w350 & ~w571 ) | ( w351 & ~w571 ) ;
  assign w2605 = w282 | w2603 ;
  assign w2606 = ( w571 & w1001 ) | ( w571 & ~w2603 ) | ( w1001 & ~w2603 ) ;
  assign w2607 = w2605 | w2606 ;
  assign w2608 = w2604 | w2607 ;
  assign w2609 = w627 | w1977 ;
  assign w2610 = ( ~w627 & w911 ) | ( ~w627 & w2608 ) | ( w911 & w2608 ) ;
  assign w2611 = w2609 | w2610 ;
  assign w2612 = w900 | w1094 ;
  assign w2613 = ( w76 & ~w900 ) | ( w76 & w2611 ) | ( ~w900 & w2611 ) ;
  assign w2614 = w2612 | w2613 ;
  assign w2615 = w821 | w1030 ;
  assign w2616 = w88 | w2615 ;
  assign w2617 = ( ~w88 & w783 ) | ( ~w88 & w2614 ) | ( w783 & w2614 ) ;
  assign w2618 = w2616 | w2617 ;
  assign w2619 = w596 | w664 ;
  assign w2620 = w221 | w2619 ;
  assign w2621 = ( w180 & ~w221 ) | ( w180 & w456 ) | ( ~w221 & w456 ) ;
  assign w2622 = w2620 | w2621 ;
  assign w2623 = ( ~w131 & w680 ) | ( ~w131 & w2622 ) | ( w680 & w2622 ) ;
  assign w2624 = w131 | w2623 ;
  assign w2625 = w133 | w1274 ;
  assign w2626 = w413 | w504 ;
  assign w2627 = ( w429 & w491 ) | ( w429 & ~w516 ) | ( w491 & ~w516 ) ;
  assign w2628 = w274 | w2626 ;
  assign w2629 = ( ~w274 & w516 ) | ( ~w274 & w642 ) | ( w516 & w642 ) ;
  assign w2630 = w2628 | w2629 ;
  assign w2631 = w2627 | w2630 ;
  assign w2632 = ( w208 & ~w209 ) | ( w208 & w264 ) | ( ~w209 & w264 ) ;
  assign w2633 = w338 | w2631 ;
  assign w2634 = ( w209 & w723 ) | ( w209 & ~w2631 ) | ( w723 & ~w2631 ) ;
  assign w2635 = w2633 | w2634 ;
  assign w2636 = w2632 | w2635 ;
  assign w2637 = ( w2552 & ~w2625 ) | ( w2552 & w2636 ) | ( ~w2625 & w2636 ) ;
  assign w2638 = ~w2636 & w2637 ;
  assign w2639 = ( ~w138 & w731 ) | ( ~w138 & w2624 ) | ( w731 & w2624 ) ;
  assign w2640 = ~w2618 & w2638 ;
  assign w2641 = ( w138 & w424 ) | ( w138 & ~w2618 ) | ( w424 & ~w2618 ) ;
  assign w2642 = w2640 & ~w2641 ;
  assign w2643 = ~w2639 & w2642 ;
  assign w2644 = ( w163 & w203 ) | ( w163 & ~w218 ) | ( w203 & ~w218 ) ;
  assign w2645 = ~w2600 & w2643 ;
  assign w2646 = ( w218 & w409 ) | ( w218 & ~w2600 ) | ( w409 & ~w2600 ) ;
  assign w2647 = w2645 & ~w2646 ;
  assign w2648 = ~w2644 & w2647 ;
  assign w2649 = ( w277 & w431 ) | ( w277 & ~w567 ) | ( w431 & ~w567 ) ;
  assign w2650 = ~w275 & w2648 ;
  assign w2651 = ( ~w275 & w567 ) | ( ~w275 & w802 ) | ( w567 & w802 ) ;
  assign w2652 = w2650 & ~w2651 ;
  assign w2653 = ~w2649 & w2652 ;
  assign w2654 = w225 | w311 ;
  assign w2655 = ( w56 & ~w225 ) | ( w56 & w255 ) | ( ~w225 & w255 ) ;
  assign w2656 = w2654 | w2655 ;
  assign w2657 = ( ~w103 & w122 ) | ( ~w103 & w2656 ) | ( w122 & w2656 ) ;
  assign w2658 = w103 | w2657 ;
  assign w2659 = ( w98 & w202 ) | ( w98 & ~w229 ) | ( w202 & ~w229 ) ;
  assign w2660 = w59 | w2658 ;
  assign w2661 = ( ~w59 & w229 ) | ( ~w59 & w980 ) | ( w229 & w980 ) ;
  assign w2662 = w2660 | w2661 ;
  assign w2663 = w2659 | w2662 ;
  assign w2664 = w505 | w951 ;
  assign w2665 = w127 | w2664 ;
  assign w2666 = ( w126 & ~w127 ) | ( w126 & w220 ) | ( ~w127 & w220 ) ;
  assign w2667 = w2665 | w2666 ;
  assign w2668 = w389 | w596 ;
  assign w2669 = w2253 | w2668 ;
  assign w2670 = ( w232 & ~w2253 ) | ( w232 & w2667 ) | ( ~w2253 & w2667 ) ;
  assign w2671 = w2669 | w2670 ;
  assign w2672 = ( w269 & w287 ) | ( w269 & ~w358 ) | ( w287 & ~w358 ) ;
  assign w2673 = w208 | w2671 ;
  assign w2674 = ( ~w208 & w358 ) | ( ~w208 & w625 ) | ( w358 & w625 ) ;
  assign w2675 = w2673 | w2674 ;
  assign w2676 = w2672 | w2675 ;
  assign w2677 = ( w218 & w573 ) | ( w218 & ~w637 ) | ( w573 & ~w637 ) ;
  assign w2678 = w1010 | w1940 ;
  assign w2679 = ( w637 & w640 ) | ( w637 & ~w1940 ) | ( w640 & ~w1940 ) ;
  assign w2680 = w2678 | w2679 ;
  assign w2681 = w2677 | w2680 ;
  assign w2682 = w2663 | w2681 ;
  assign w2683 = w859 | w2682 ;
  assign w2684 = ( w859 & w1228 ) | ( w859 & ~w2676 ) | ( w1228 & ~w2676 ) ;
  assign w2685 = ~w2683 & w2684 ;
  assign w2686 = ( w388 & w530 ) | ( w388 & ~w764 ) | ( w530 & ~w764 ) ;
  assign w2687 = ~w1421 & w2685 ;
  assign w2688 = ( w764 & w1340 ) | ( w764 & ~w1421 ) | ( w1340 & ~w1421 ) ;
  assign w2689 = w2687 & ~w2688 ;
  assign w2690 = ~w2686 & w2689 ;
  assign w2691 = w571 | w726 ;
  assign w2692 = w74 | w2691 ;
  assign w2693 = ( w74 & ~w317 ) | ( w74 & w2690 ) | ( ~w317 & w2690 ) ;
  assign w2694 = ~w2692 & w2693 ;
  assign w2695 = w309 | w897 ;
  assign w2696 = ( w230 & w421 ) | ( w230 & ~w623 ) | ( w421 & ~w623 ) ;
  assign w2697 = w165 | w205 ;
  assign w2698 = ( ~w205 & w623 ) | ( ~w205 & w817 ) | ( w623 & w817 ) ;
  assign w2699 = w2697 | w2698 ;
  assign w2700 = w2696 | w2699 ;
  assign w2701 = w265 | w488 ;
  assign w2702 = ( ~w265 & w352 ) | ( ~w265 & w2700 ) | ( w352 & w2700 ) ;
  assign w2703 = w2701 | w2702 ;
  assign w2704 = w350 | w889 ;
  assign w2705 = w509 | w628 ;
  assign w2706 = w465 | w860 ;
  assign w2707 = w147 | w2706 ;
  assign w2708 = ( ~w147 & w389 ) | ( ~w147 & w2168 ) | ( w389 & w2168 ) ;
  assign w2709 = w2707 | w2708 ;
  assign w2710 = w570 | w1153 ;
  assign w2711 = w199 | w2710 ;
  assign w2712 = ( ~w199 & w325 ) | ( ~w199 & w2709 ) | ( w325 & w2709 ) ;
  assign w2713 = w2711 | w2712 ;
  assign w2714 = ( w59 & w887 ) | ( w59 & ~w1206 ) | ( w887 & ~w1206 ) ;
  assign w2715 = w1206 | w2714 ;
  assign w2716 = ( w223 & w593 ) | ( w223 & ~w1229 ) | ( w593 & ~w1229 ) ;
  assign w2717 = w219 | w2715 ;
  assign w2718 = ( ~w219 & w1229 ) | ( ~w219 & w1274 ) | ( w1229 & w1274 ) ;
  assign w2719 = w2717 | w2718 ;
  assign w2720 = w2716 | w2719 ;
  assign w2721 = w88 | w533 ;
  assign w2722 = w997 | w2721 ;
  assign w2723 = ( w81 & ~w997 ) | ( w81 & w2720 ) | ( ~w997 & w2720 ) ;
  assign w2724 = w2722 | w2723 ;
  assign w2725 = ( w202 & w429 ) | ( w202 & ~w513 ) | ( w429 & ~w513 ) ;
  assign w2726 = w44 | w2724 ;
  assign w2727 = ( ~w44 & w513 ) | ( ~w44 & w531 ) | ( w513 & w531 ) ;
  assign w2728 = w2726 | w2727 ;
  assign w2729 = w2725 | w2728 ;
  assign w2730 = w504 | w625 ;
  assign w2731 = w431 | w2730 ;
  assign w2732 = ( w318 & ~w431 ) | ( w318 & w458 ) | ( ~w431 & w458 ) ;
  assign w2733 = w2731 | w2732 ;
  assign w2734 = w141 | w534 ;
  assign w2735 = ( ~w141 & w524 ) | ( ~w141 & w2733 ) | ( w524 & w2733 ) ;
  assign w2736 = w2734 | w2735 ;
  assign w2737 = ( ~w179 & w800 ) | ( ~w179 & w2736 ) | ( w800 & w2736 ) ;
  assign w2738 = w2713 | w2729 ;
  assign w2739 = ( w179 & w596 ) | ( w179 & ~w2713 ) | ( w596 & ~w2713 ) ;
  assign w2740 = w2738 | w2739 ;
  assign w2741 = w2737 | w2740 ;
  assign w2742 = w351 | w2705 ;
  assign w2743 = w1646 | w2742 ;
  assign w2744 = ( ~w1646 & w2704 ) | ( ~w1646 & w2741 ) | ( w2704 & w2741 ) ;
  assign w2745 = w2743 | w2744 ;
  assign w2746 = ( w139 & w339 ) | ( w139 & ~w418 ) | ( w339 & ~w418 ) ;
  assign w2747 = w84 | w2745 ;
  assign w2748 = ( ~w84 & w418 ) | ( ~w84 & w681 ) | ( w418 & w681 ) ;
  assign w2749 = w2747 | w2748 ;
  assign w2750 = w2746 | w2749 ;
  assign w2751 = ( w169 & w511 ) | ( w169 & ~w561 ) | ( w511 & ~w561 ) ;
  assign w2752 = w98 | w622 ;
  assign w2753 = ( ~w98 & w561 ) | ( ~w98 & w724 ) | ( w561 & w724 ) ;
  assign w2754 = w2752 | w2753 ;
  assign w2755 = w2751 | w2754 ;
  assign w2756 = w344 | w722 ;
  assign w2757 = w2480 | w2756 ;
  assign w2758 = ( w220 & ~w2480 ) | ( w220 & w2755 ) | ( ~w2480 & w2755 ) ;
  assign w2759 = w2757 | w2758 ;
  assign w2760 = w90 | w383 ;
  assign w2761 = ( w149 & ~w176 ) | ( w149 & w229 ) | ( ~w176 & w229 ) ;
  assign w2762 = w176 | w2761 ;
  assign w2763 = ( w180 & w203 ) | ( w180 & ~w345 ) | ( w203 & ~w345 ) ;
  assign w2764 = w1620 | w2762 ;
  assign w2765 = ( w345 & w1126 ) | ( w345 & ~w2762 ) | ( w1126 & ~w2762 ) ;
  assign w2766 = w2764 | w2765 ;
  assign w2767 = w2763 | w2766 ;
  assign w2768 = ( w119 & w221 ) | ( w119 & ~w266 ) | ( w221 & ~w266 ) ;
  assign w2769 = w1456 | w2767 ;
  assign w2770 = ( w266 & w640 ) | ( w266 & ~w2767 ) | ( w640 & ~w2767 ) ;
  assign w2771 = w2769 | w2770 ;
  assign w2772 = w2768 | w2771 ;
  assign w2773 = w138 | w424 ;
  assign w2774 = w952 | w2773 ;
  assign w2775 = ( ~w952 & w2760 ) | ( ~w952 & w2772 ) | ( w2760 & w2772 ) ;
  assign w2776 = w2774 | w2775 ;
  assign w2777 = ( w215 & w388 ) | ( w215 & ~w565 ) | ( w388 & ~w565 ) ;
  assign w2778 = w68 | w2776 ;
  assign w2779 = ( ~w68 & w565 ) | ( ~w68 & w662 ) | ( w565 & w662 ) ;
  assign w2780 = w2778 | w2779 ;
  assign w2781 = w2777 | w2780 ;
  assign w2782 = w56 | w505 ;
  assign w2783 = ( w264 & w525 ) | ( w264 & ~w2782 ) | ( w525 & ~w2782 ) ;
  assign w2784 = w2782 | w2783 ;
  assign w2785 = ( w144 & w413 ) | ( w144 & ~w492 ) | ( w413 & ~w492 ) ;
  assign w2786 = w2781 | w2784 ;
  assign w2787 = ( w492 & w606 ) | ( w492 & ~w2784 ) | ( w606 & ~w2784 ) ;
  assign w2788 = w2786 | w2787 ;
  assign w2789 = w2785 | w2788 ;
  assign w2790 = w2695 | w2703 ;
  assign w2791 = w2789 | w2790 ;
  assign w2792 = ( w2750 & w2759 ) | ( w2750 & ~w2789 ) | ( w2759 & ~w2789 ) ;
  assign w2793 = w2791 | w2792 ;
  assign w2794 = ( ~w466 & w731 ) | ( ~w466 & w999 ) | ( w731 & w999 ) ;
  assign w2795 = w129 | w2793 ;
  assign w2796 = ( ~w129 & w466 ) | ( ~w129 & w1094 ) | ( w466 & w1094 ) ;
  assign w2797 = w2795 | w2796 ;
  assign w2798 = w2794 | w2797 ;
  assign w2799 = ( w358 & w515 ) | ( w358 & ~w568 ) | ( w515 & ~w568 ) ;
  assign w2800 = w259 | w2798 ;
  assign w2801 = ( ~w259 & w568 ) | ( ~w259 & w1001 ) | ( w568 & w1001 ) ;
  assign w2802 = w2800 | w2801 ;
  assign w2803 = w2799 | w2802 ;
  assign w2804 = ( ~w161 & w208 ) | ( ~w161 & w2803 ) | ( w208 & w2803 ) ;
  assign w2805 = w161 | w2804 ;
  assign w2806 = w285 | w504 ;
  assign w2807 = ( w219 & ~w285 ) | ( w219 & w342 ) | ( ~w285 & w342 ) ;
  assign w2808 = w2806 | w2807 ;
  assign w2809 = w608 | w1229 ;
  assign w2810 = w1147 | w2809 ;
  assign w2811 = ( w96 & w530 ) | ( w96 & ~w1147 ) | ( w530 & ~w1147 ) ;
  assign w2812 = w2810 | w2811 ;
  assign w2813 = ( w81 & ~w198 ) | ( w81 & w269 ) | ( ~w198 & w269 ) ;
  assign w2814 = w198 | w2813 ;
  assign w2815 = ( w144 & w512 ) | ( w144 & ~w568 ) | ( w512 & ~w568 ) ;
  assign w2816 = w1420 & ~w2814 ;
  assign w2817 = ( w568 & w1086 ) | ( w568 & ~w2814 ) | ( w1086 & ~w2814 ) ;
  assign w2818 = w2816 & ~w2817 ;
  assign w2819 = ~w2815 & w2818 ;
  assign w2820 = ( ~w999 & w1207 ) | ( ~w999 & w2819 ) | ( w1207 & w2819 ) ;
  assign w2821 = w2428 | w2812 ;
  assign w2822 = ( w1207 & w2705 ) | ( w1207 & ~w2812 ) | ( w2705 & ~w2812 ) ;
  assign w2823 = w2821 | w2822 ;
  assign w2824 = w2820 & ~w2823 ;
  assign w2825 = ( w141 & w386 ) | ( w141 & ~w897 ) | ( w386 & ~w897 ) ;
  assign w2826 = ~w59 & w2824 ;
  assign w2827 = ( ~w59 & w897 ) | ( ~w59 & w1130 ) | ( w897 & w1130 ) ;
  assign w2828 = w2826 & ~w2827 ;
  assign w2829 = ~w2825 & w2828 ;
  assign w2830 = \pi25 & w71 ;
  assign w2831 = \pi24 & w2830 ;
  assign w2832 = \pi23 ^ \pi24 ;
  assign w2833 = ( \pi24 & \pi25 ) | ( \pi24 & \pi26 ) | ( \pi25 & \pi26 ) ;
  assign w2834 = ( ~\pi26 & w2832 ) | ( ~\pi26 & w2833 ) | ( w2832 & w2833 ) ;
  assign w2835 = w145 & ~w2833 ;
  assign w2836 = ( w2831 & ~w2834 ) | ( w2831 & w2835 ) | ( ~w2834 & w2835 ) ;
  assign w2837 = ( w418 & w605 ) | ( w418 & ~w889 ) | ( w605 & ~w889 ) ;
  assign w2838 = w147 | w277 ;
  assign w2839 = ( ~w277 & w889 ) | ( ~w277 & w1340 ) | ( w889 & w1340 ) ;
  assign w2840 = w2838 | w2839 ;
  assign w2841 = w2837 | w2840 ;
  assign w2842 = w495 | w1031 ;
  assign w2843 = w2841 | w2842 ;
  assign w2844 = ( w84 & w2625 ) | ( w84 & ~w2841 ) | ( w2625 & ~w2841 ) ;
  assign w2845 = w2843 | w2844 ;
  assign w2846 = ( w384 & w390 ) | ( w384 & ~w787 ) | ( w390 & ~w787 ) ;
  assign w2847 = w252 | w2845 ;
  assign w2848 = ( ~w252 & w787 ) | ( ~w252 & w901 ) | ( w787 & w901 ) ;
  assign w2849 = w2847 | w2848 ;
  assign w2850 = w2846 | w2849 ;
  assign w2851 = w232 | w567 ;
  assign w2852 = w2319 | w2851 ;
  assign w2853 = ( w51 & ~w2319 ) | ( w51 & w2403 ) | ( ~w2319 & w2403 ) ;
  assign w2854 = w2852 | w2853 ;
  assign w2855 = w287 | w449 ;
  assign w2856 = w1836 | w2855 ;
  assign w2857 = ( w226 & ~w1836 ) | ( w226 & w2854 ) | ( ~w1836 & w2854 ) ;
  assign w2858 = w2856 | w2857 ;
  assign w2859 = w2836 | w2858 ;
  assign w2860 = ( w2781 & w2850 ) | ( w2781 & ~w2858 ) | ( w2850 & ~w2858 ) ;
  assign w2861 = w2859 | w2860 ;
  assign w2862 = ( ~w415 & w1208 ) | ( ~w415 & w2808 ) | ( w1208 & w2808 ) ;
  assign w2863 = w2829 & ~w2861 ;
  assign w2864 = ( w415 & w524 ) | ( w415 & w2829 ) | ( w524 & w2829 ) ;
  assign w2865 = w2863 & ~w2864 ;
  assign w2866 = ~w2862 & w2865 ;
  assign w2867 = ( w175 & w625 ) | ( w175 & ~w641 ) | ( w625 & ~w641 ) ;
  assign w2868 = ~w956 & w2866 ;
  assign w2869 = ( w641 & ~w956 ) | ( w641 & w1030 ) | ( ~w956 & w1030 ) ;
  assign w2870 = w2868 & ~w2869 ;
  assign w2871 = ~w2867 & w2870 ;
  assign w2872 = w206 | w1274 ;
  assign w2873 = w120 | w143 ;
  assign w2874 = w342 | w889 ;
  assign w2875 = ( w310 & ~w342 ) | ( w310 & w511 ) | ( ~w342 & w511 ) ;
  assign w2876 = w2874 | w2875 ;
  assign w2877 = w2873 | w2876 ;
  assign w2878 = ( w103 & w317 ) | ( w103 & ~w663 ) | ( w317 & ~w663 ) ;
  assign w2879 = w1154 | w2877 ;
  assign w2880 = ( w663 & w821 ) | ( w663 & ~w1154 ) | ( w821 & ~w1154 ) ;
  assign w2881 = w2879 | w2880 ;
  assign w2882 = w2878 | w2881 ;
  assign w2883 = w431 | w725 ;
  assign w2884 = w199 | w2883 ;
  assign w2885 = ( ~w199 & w229 ) | ( ~w199 & w2882 ) | ( w229 & w2882 ) ;
  assign w2886 = w2884 | w2885 ;
  assign w2887 = w390 | w569 ;
  assign w2888 = ( ~w390 & w430 ) | ( ~w390 & w517 ) | ( w430 & w517 ) ;
  assign w2889 = w2887 | w2888 ;
  assign w2890 = w386 | w623 ;
  assign w2891 = w122 | w2890 ;
  assign w2892 = ( w84 & ~w122 ) | ( w84 & w384 ) | ( ~w122 & w384 ) ;
  assign w2893 = w2891 | w2892 ;
  assign w2894 = ( ~w389 & w493 ) | ( ~w389 & w2893 ) | ( w493 & w2893 ) ;
  assign w2895 = w2558 | w2889 ;
  assign w2896 = ( w389 & w596 ) | ( w389 & ~w2889 ) | ( w596 & ~w2889 ) ;
  assign w2897 = w2895 | w2896 ;
  assign w2898 = w2894 | w2897 ;
  assign w2899 = w2872 | w2898 ;
  assign w2900 = ( w1282 & w2886 ) | ( w1282 & ~w2898 ) | ( w2886 & ~w2898 ) ;
  assign w2901 = w2899 | w2900 ;
  assign w2902 = w230 | w312 ;
  assign w2903 = w507 | w2902 ;
  assign w2904 = ( ~w507 & w2782 ) | ( ~w507 & w2901 ) | ( w2782 & w2901 ) ;
  assign w2905 = w2903 | w2904 ;
  assign w2906 = w530 | w570 ;
  assign w2907 = w221 | w2906 ;
  assign w2908 = ( ~w221 & w281 ) | ( ~w221 & w2905 ) | ( w281 & w2905 ) ;
  assign w2909 = w2907 | w2908 ;
  assign w2910 = w837 | w1031 ;
  assign w2911 = w392 | w2910 ;
  assign w2912 = ( w286 & ~w392 ) | ( w286 & w758 ) | ( ~w392 & w758 ) ;
  assign w2913 = w2911 | w2912 ;
  assign w2914 = ( ~w358 & w680 ) | ( ~w358 & w2913 ) | ( w680 & w2913 ) ;
  assign w2915 = w358 | w2914 ;
  assign w2916 = ( w565 & w567 ) | ( w565 & ~w568 ) | ( w567 & ~w568 ) ;
  assign w2917 = w59 | w420 ;
  assign w2918 = ( ~w420 & w568 ) | ( ~w420 & w673 ) | ( w568 & w673 ) ;
  assign w2919 = w2917 | w2918 ;
  assign w2920 = w2916 | w2919 ;
  assign w2921 = ( ~w114 & w353 ) | ( ~w114 & w2920 ) | ( w353 & w2920 ) ;
  assign w2922 = w114 | w2921 ;
  assign w2923 = w223 | w491 ;
  assign w2924 = w68 | w2923 ;
  assign w2925 = ( ~w68 & w220 ) | ( ~w68 & w410 ) | ( w220 & w410 ) ;
  assign w2926 = w2924 | w2925 ;
  assign w2927 = w177 | w178 ;
  assign w2928 = w2922 | w2927 ;
  assign w2929 = ( w2915 & ~w2922 ) | ( w2915 & w2926 ) | ( ~w2922 & w2926 ) ;
  assign w2930 = w2928 | w2929 ;
  assign w2931 = w514 | w2060 ;
  assign w2932 = ( ~w514 & w1265 ) | ( ~w514 & w2930 ) | ( w1265 & w2930 ) ;
  assign w2933 = w2931 | w2932 ;
  assign w2934 = ( w383 & w408 ) | ( w383 & ~w488 ) | ( w408 & ~w488 ) ;
  assign w2935 = w638 | w2933 ;
  assign w2936 = ( w488 & ~w638 ) | ( w488 & w724 ) | ( ~w638 & w724 ) ;
  assign w2937 = w2935 | w2936 ;
  assign w2938 = w2934 | w2937 ;
  assign w2939 = w255 | w1646 ;
  assign w2940 = ( w124 & w1461 ) | ( w124 & ~w1646 ) | ( w1461 & ~w1646 ) ;
  assign w2941 = w2939 | w2940 ;
  assign w2942 = w509 | w1094 ;
  assign w2943 = w661 | w2942 ;
  assign w2944 = ( w116 & ~w661 ) | ( w116 & w2941 ) | ( ~w661 & w2941 ) ;
  assign w2945 = w2943 | w2944 ;
  assign w2946 = w95 | w2597 ;
  assign w2947 = ( ~w95 & w98 ) | ( ~w95 & w2945 ) | ( w98 & w2945 ) ;
  assign w2948 = w2946 | w2947 ;
  assign w2949 = ~w275 & w359 ;
  assign w2950 = w259 | w1126 ;
  assign w2951 = w135 | w2950 ;
  assign w2952 = ( ~w135 & w203 ) | ( ~w135 & w2147 ) | ( w203 & w2147 ) ;
  assign w2953 = w2951 | w2952 ;
  assign w2954 = ~w901 & w2949 ;
  assign w2955 = ( w169 & w2949 ) | ( w169 & w2953 ) | ( w2949 & w2953 ) ;
  assign w2956 = w2954 & ~w2955 ;
  assign w2957 = w101 | w309 ;
  assign w2958 = w2956 & ~w2957 ;
  assign w2959 = ( w1759 & w2948 ) | ( w1759 & w2956 ) | ( w2948 & w2956 ) ;
  assign w2960 = w2958 & ~w2959 ;
  assign w2961 = w467 | w674 ;
  assign w2962 = w2938 | w2961 ;
  assign w2963 = ( ~w2909 & w2938 ) | ( ~w2909 & w2960 ) | ( w2938 & w2960 ) ;
  assign w2964 = ~w2962 & w2963 ;
  assign w2965 = w532 | w1979 ;
  assign w2966 = ( w532 & ~w1618 ) | ( w532 & w2964 ) | ( ~w1618 & w2964 ) ;
  assign w2967 = ~w2965 & w2966 ;
  assign w2968 = w266 | w414 ;
  assign w2969 = ( w414 & ~w2374 ) | ( w414 & w2967 ) | ( ~w2374 & w2967 ) ;
  assign w2970 = ~w2968 & w2969 ;
  assign w2971 = w115 | w315 ;
  assign w2972 = ( w115 & ~w256 ) | ( w115 & w2970 ) | ( ~w256 & w2970 ) ;
  assign w2973 = ~w2971 & w2972 ;
  assign w2974 = w2871 & w2973 ;
  assign w2975 = ( w2694 & w2973 ) | ( w2694 & ~w2974 ) | ( w2973 & ~w2974 ) ;
  assign w2976 = ( w2653 & w2871 ) | ( w2653 & w2975 ) | ( w2871 & w2975 ) ;
  assign w2977 = ( w2694 & ~w2805 ) | ( w2694 & w2976 ) | ( ~w2805 & w2976 ) ;
  assign w2978 = ( w2578 & w2653 ) | ( w2578 & w2977 ) | ( w2653 & w2977 ) ;
  assign w2979 = ( ~w2500 & w2578 ) | ( ~w2500 & w2978 ) | ( w2578 & w2978 ) ;
  assign w2980 = ( w2391 & w2500 ) | ( w2391 & ~w2979 ) | ( w2500 & ~w2979 ) ;
  assign w2981 = ( w2273 & w2391 ) | ( w2273 & w2980 ) | ( w2391 & w2980 ) ;
  assign w2982 = ( ~w2235 & w2273 ) | ( ~w2235 & w2981 ) | ( w2273 & w2981 ) ;
  assign w2983 = ( w2130 & w2235 ) | ( w2130 & ~w2982 ) | ( w2235 & ~w2982 ) ;
  assign w2984 = ( w2059 & w2130 ) | ( w2059 & w2983 ) | ( w2130 & w2983 ) ;
  assign w2985 = ( ~w1976 & w2059 ) | ( ~w1976 & w2984 ) | ( w2059 & w2984 ) ;
  assign w2986 = ( w1939 & ~w1976 ) | ( w1939 & w2985 ) | ( ~w1976 & w2985 ) ;
  assign w2987 = ( w1834 & w1939 ) | ( w1834 & w2986 ) | ( w1939 & w2986 ) ;
  assign w2988 = ( ~w1711 & w1834 ) | ( ~w1711 & w2987 ) | ( w1834 & w2987 ) ;
  assign w2989 = ( w1614 & w1711 ) | ( w1614 & ~w2988 ) | ( w1711 & ~w2988 ) ;
  assign w2990 = ( ~w1510 & w1614 ) | ( ~w1510 & w2989 ) | ( w1614 & w2989 ) ;
  assign w2991 = ( w1399 & ~w1510 ) | ( w1399 & w2990 ) | ( ~w1510 & w2990 ) ;
  assign w2992 = ( ~w1264 & w1399 ) | ( ~w1264 & w2991 ) | ( w1399 & w2991 ) ;
  assign w2993 = ( w1205 & ~w1264 ) | ( w1205 & w2992 ) | ( ~w1264 & w2992 ) ;
  assign w2994 = ( w1085 & w1205 ) | ( w1085 & w2993 ) | ( w1205 & w2993 ) ;
  assign w2995 = ( w979 & w1085 ) | ( w979 & w2994 ) | ( w1085 & w2994 ) ;
  assign w2996 = ( ~w883 & w979 ) | ( ~w883 & w2995 ) | ( w979 & w2995 ) ;
  assign w2997 = ( w721 & ~w883 ) | ( w721 & w2996 ) | ( ~w883 & w2996 ) ;
  assign w2998 = ( w592 & w721 ) | ( w592 & w2997 ) | ( w721 & w2997 ) ;
  assign w2999 = ( ~w381 & w592 ) | ( ~w381 & w2998 ) | ( w592 & w2998 ) ;
  assign w3000 = w311 | w662 ;
  assign w3001 = ( w180 & ~w311 ) | ( w180 & w465 ) | ( ~w311 & w465 ) ;
  assign w3002 = w3000 | w3001 ;
  assign w3003 = w560 | w1094 ;
  assign w3004 = w3002 | w3003 ;
  assign w3005 = ( w420 & w2168 ) | ( w420 & ~w3002 ) | ( w2168 & ~w3002 ) ;
  assign w3006 = w3004 | w3005 ;
  assign w3007 = ( w320 & w640 ) | ( w320 & ~w680 ) | ( w640 & ~w680 ) ;
  assign w3008 = w287 | w3006 ;
  assign w3009 = ( ~w287 & w680 ) | ( ~w287 & w783 ) | ( w680 & w783 ) ;
  assign w3010 = w3008 | w3009 ;
  assign w3011 = w3007 | w3010 ;
  assign w3012 = w352 | w570 ;
  assign w3013 = w98 | w3012 ;
  assign w3014 = ( w63 & ~w98 ) | ( w63 & w118 ) | ( ~w98 & w118 ) ;
  assign w3015 = w3013 | w3014 ;
  assign w3016 = ( w74 & w463 ) | ( w74 & ~w492 ) | ( w463 & ~w492 ) ;
  assign w3017 = w3011 | w3015 ;
  assign w3018 = ( w492 & w725 ) | ( w492 & ~w3015 ) | ( w725 & ~w3015 ) ;
  assign w3019 = w3017 | w3018 ;
  assign w3020 = w3016 | w3019 ;
  assign w3021 = ( w258 & ~w283 ) | ( w258 & w2306 ) | ( ~w283 & w2306 ) ;
  assign w3022 = w1206 | w3020 ;
  assign w3023 = ( w283 & w342 ) | ( w283 & ~w1206 ) | ( w342 & ~w1206 ) ;
  assign w3024 = w3022 | w3023 ;
  assign w3025 = w3021 | w3024 ;
  assign w3026 = ( w256 & w318 ) | ( w256 & ~w641 ) | ( w318 & ~w641 ) ;
  assign w3027 = w219 | w3025 ;
  assign w3028 = ( ~w219 & w641 ) | ( ~w219 & w724 ) | ( w641 & w724 ) ;
  assign w3029 = w3027 | w3028 ;
  assign w3030 = w3026 | w3029 ;
  assign w3031 = ( ~w259 & w309 ) | ( ~w259 & w3030 ) | ( w309 & w3030 ) ;
  assign w3032 = w259 | w3031 ;
  assign w3033 = ( w569 & w758 ) | ( w569 & ~w821 ) | ( w758 & ~w821 ) ;
  assign w3034 = w430 | w459 ;
  assign w3035 = ( ~w459 & w821 ) | ( ~w459 & w1001 ) | ( w821 & w1001 ) ;
  assign w3036 = w3034 | w3035 ;
  assign w3037 = w3033 | w3036 ;
  assign w3038 = w504 | w515 ;
  assign w3039 = w2319 | w3038 ;
  assign w3040 = ( w252 & w1460 ) | ( w252 & ~w2319 ) | ( w1460 & ~w2319 ) ;
  assign w3041 = w3039 | w3040 ;
  assign w3042 = w263 | w723 ;
  assign w3043 = w209 | w3042 ;
  assign w3044 = ( ~w209 & w260 ) | ( ~w209 & w3041 ) | ( w260 & w3041 ) ;
  assign w3045 = w3043 | w3044 ;
  assign w3046 = w2091 | w3037 ;
  assign w3047 = w270 | w3046 ;
  assign w3048 = ( ~w270 & w1978 ) | ( ~w270 & w3045 ) | ( w1978 & w3045 ) ;
  assign w3049 = w3047 | w3048 ;
  assign w3050 = ( w232 & ~w596 ) | ( w232 & w1882 ) | ( ~w596 & w1882 ) ;
  assign w3051 = w532 | w3049 ;
  assign w3052 = ( ~w532 & w596 ) | ( ~w532 & w623 ) | ( w596 & w623 ) ;
  assign w3053 = w3051 | w3052 ;
  assign w3054 = w3050 | w3053 ;
  assign w3055 = ( w467 & w488 ) | ( w467 & ~w595 ) | ( w488 & ~w595 ) ;
  assign w3056 = w226 | w3054 ;
  assign w3057 = ( ~w226 & w595 ) | ( ~w226 & w673 ) | ( w595 & w673 ) ;
  assign w3058 = w3056 | w3057 ;
  assign w3059 = w3055 | w3058 ;
  assign w3060 = ( w143 & w265 ) | ( w143 & ~w286 ) | ( w265 & ~w286 ) ;
  assign w3061 = w68 | w2521 ;
  assign w3062 = ( ~w68 & w286 ) | ( ~w68 & w315 ) | ( w286 & w315 ) ;
  assign w3063 = w3061 | w3062 ;
  assign w3064 = w3060 | w3063 ;
  assign w3065 = w359 & ~w1030 ;
  assign w3066 = ( w359 & w516 ) | ( w359 & w3064 ) | ( w516 & w3064 ) ;
  assign w3067 = w3065 & ~w3066 ;
  assign w3068 = w271 | w530 ;
  assign w3069 = w119 | w3068 ;
  assign w3070 = ( ~w119 & w229 ) | ( ~w119 & w638 ) | ( w229 & w638 ) ;
  assign w3071 = w3069 | w3070 ;
  assign w3072 = w88 | w389 ;
  assign w3073 = ( w81 & ~w88 ) | ( w81 & w149 ) | ( ~w88 & w149 ) ;
  assign w3074 = w3072 | w3073 ;
  assign w3075 = ( w203 & w322 ) | ( w203 & ~w339 ) | ( w322 & ~w339 ) ;
  assign w3076 = w414 | w3074 ;
  assign w3077 = ( w339 & w509 ) | ( w339 & ~w3074 ) | ( w509 & ~w3074 ) ;
  assign w3078 = w3076 | w3077 ;
  assign w3079 = w3075 | w3078 ;
  assign w3080 = ( w1880 & w3071 ) | ( w1880 & ~w3079 ) | ( w3071 & ~w3079 ) ;
  assign w3081 = ~w3059 & w3067 ;
  assign w3082 = ( w222 & w3067 ) | ( w222 & w3079 ) | ( w3067 & w3079 ) ;
  assign w3083 = w3081 & ~w3082 ;
  assign w3084 = ~w3080 & w3083 ;
  assign w3085 = ( ~w104 & w594 ) | ( ~w104 & w1421 ) | ( w594 & w1421 ) ;
  assign w3086 = ~w3032 & w3084 ;
  assign w3087 = ( w104 & w506 ) | ( w104 & w3084 ) | ( w506 & w3084 ) ;
  assign w3088 = w3086 & ~w3087 ;
  assign w3089 = ~w3085 & w3088 ;
  assign w3090 = ( w310 & w344 ) | ( w310 & ~w358 ) | ( w344 & ~w358 ) ;
  assign w3091 = ~w175 & w3089 ;
  assign w3092 = ( ~w175 & w358 ) | ( ~w175 & w1229 ) | ( w358 & w1229 ) ;
  assign w3093 = w3091 & ~w3092 ;
  assign w3094 = ~w3090 & w3093 ;
  assign w3095 = w381 ^ w2999 ;
  assign w3096 = w3094 ^ w3095 ;
  assign w3097 = ( \pi29 & ~\pi30 ) | ( \pi29 & \pi31 ) | ( ~\pi30 & \pi31 ) ;
  assign w3098 = \pi30 & w3097 ;
  assign w3099 = ( \pi30 & \pi31 ) | ( \pi30 & ~w381 ) | ( \pi31 & ~w381 ) ;
  assign w3100 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w3099 ) | ( \pi30 & w3099 ) ;
  assign w3101 = ( \pi29 & ~\pi30 ) | ( \pi29 & w3099 ) | ( ~\pi30 & w3099 ) ;
  assign w3102 = ( ~\pi30 & w592 ) | ( ~\pi30 & w3101 ) | ( w592 & w3101 ) ;
  assign w3103 = ( w3094 & ~w3101 ) | ( w3094 & w3102 ) | ( ~w3101 & w3102 ) ;
  assign w3104 = \pi31 | w3103 ;
  assign w3105 = ( w3100 & w3102 ) | ( w3100 & ~w3104 ) | ( w3102 & ~w3104 ) ;
  assign w3106 = ( w37 & w3096 ) | ( w37 & w3105 ) | ( w3096 & w3105 ) ;
  assign w3107 = w3105 | w3106 ;
  assign w3108 = ( w256 & w257 ) | ( w256 & ~w274 ) | ( w257 & ~w274 ) ;
  assign w3109 = w223 | w2893 ;
  assign w3110 = ( ~w223 & w274 ) | ( ~w223 & w344 ) | ( w274 & w344 ) ;
  assign w3111 = w3109 | w3110 ;
  assign w3112 = w3108 | w3111 ;
  assign w3113 = ( ~w488 & w628 ) | ( ~w488 & w3112 ) | ( w628 & w3112 ) ;
  assign w3114 = w488 | w3113 ;
  assign w3115 = w309 | w1153 ;
  assign w3116 = w525 | w723 ;
  assign w3117 = w165 | w3116 ;
  assign w3118 = ( w164 & ~w165 ) | ( w164 & w390 ) | ( ~w165 & w390 ) ;
  assign w3119 = w3117 | w3118 ;
  assign w3120 = w663 | w3119 ;
  assign w3121 = ( w161 & w3115 ) | ( w161 & ~w3119 ) | ( w3115 & ~w3119 ) ;
  assign w3122 = w3120 | w3121 ;
  assign w3123 = ( w267 & ~w268 ) | ( w267 & w1835 ) | ( ~w268 & w1835 ) ;
  assign w3124 = w3114 | w3122 ;
  assign w3125 = ( w268 & w449 ) | ( w268 & ~w3122 ) | ( w449 & ~w3122 ) ;
  assign w3126 = w3124 | w3125 ;
  assign w3127 = w3123 | w3126 ;
  assign w3128 = ( w509 & ~w567 ) | ( w509 & w1166 ) | ( ~w567 & w1166 ) ;
  assign w3129 = w532 | w3127 ;
  assign w3130 = ( ~w532 & w567 ) | ( ~w532 & w674 ) | ( w567 & w674 ) ;
  assign w3131 = w3129 | w3130 ;
  assign w3132 = w3128 | w3131 ;
  assign w3133 = ( w490 & w640 ) | ( w490 & ~w642 ) | ( w640 & ~w642 ) ;
  assign w3134 = w258 | w388 ;
  assign w3135 = ( ~w388 & w642 ) | ( ~w388 & w764 ) | ( w642 & w764 ) ;
  assign w3136 = w3134 | w3135 ;
  assign w3137 = w3133 | w3136 ;
  assign w3138 = w131 | w1030 ;
  assign w3139 = ( ~w131 & w175 ) | ( ~w131 & w3137 ) | ( w175 & w3137 ) ;
  assign w3140 = w3138 | w3139 ;
  assign w3141 = w103 | w1274 ;
  assign w3142 = ( ~w103 & w565 ) | ( ~w103 & w2760 ) | ( w565 & w2760 ) ;
  assign w3143 = w3141 | w3142 ;
  assign w3144 = ( w360 & w575 ) | ( w360 & w1473 ) | ( w575 & w1473 ) ;
  assign w3145 = w360 & ~w3144 ;
  assign w3146 = ( w493 & ~w3143 ) | ( w493 & w3145 ) | ( ~w3143 & w3145 ) ;
  assign w3147 = w950 | w2420 ;
  assign w3148 = ( w493 & ~w950 ) | ( w493 & w2782 ) | ( ~w950 & w2782 ) ;
  assign w3149 = w3147 | w3148 ;
  assign w3150 = w3146 & ~w3149 ;
  assign w3151 = ( w310 & ~w421 ) | ( w310 & w3140 ) | ( ~w421 & w3140 ) ;
  assign w3152 = ~w3132 & w3150 ;
  assign w3153 = ( w421 & w511 ) | ( w421 & ~w3132 ) | ( w511 & ~w3132 ) ;
  assign w3154 = w3152 & ~w3153 ;
  assign w3155 = ~w3151 & w3154 ;
  assign w3156 = w340 | w1128 ;
  assign w3157 = w178 | w3156 ;
  assign w3158 = ( w178 & ~w219 ) | ( w178 & w3155 ) | ( ~w219 & w3155 ) ;
  assign w3159 = ~w3157 & w3158 ;
  assign w3160 = w531 | w802 ;
  assign w3161 = w178 | w3160 ;
  assign w3162 = ( w116 & ~w178 ) | ( w116 & w456 ) | ( ~w178 & w456 ) ;
  assign w3163 = w3161 | w3162 ;
  assign w3164 = ( w120 & w311 ) | ( w120 & ~w312 ) | ( w311 & ~w312 ) ;
  assign w3165 = w103 | w3163 ;
  assign w3166 = ( ~w103 & w312 ) | ( ~w103 & w1274 ) | ( w312 & w1274 ) ;
  assign w3167 = w3165 | w3166 ;
  assign w3168 = w3164 | w3167 ;
  assign w3169 = w345 | w980 ;
  assign w3170 = w111 | w3169 ;
  assign w3171 = ( ~w111 & w272 ) | ( ~w111 & w3168 ) | ( w272 & w3168 ) ;
  assign w3172 = w3170 | w3171 ;
  assign w3173 = ( w496 & w640 ) | ( w496 & ~w642 ) | ( w640 & ~w642 ) ;
  assign w3174 = w495 | w3172 ;
  assign w3175 = ( ~w495 & w642 ) | ( ~w495 & w764 ) | ( w642 & w764 ) ;
  assign w3176 = w3174 | w3175 ;
  assign w3177 = w3173 | w3176 ;
  assign w3178 = w415 | w524 ;
  assign w3179 = w1884 | w3178 ;
  assign w3180 = ( ~w1884 & w2695 ) | ( ~w1884 & w3177 ) | ( w2695 & w3177 ) ;
  assign w3181 = w3179 | w3180 ;
  assign w3182 = ( w84 & w104 ) | ( w84 & ~w149 ) | ( w104 & ~w149 ) ;
  assign w3183 = w1945 | w3181 ;
  assign w3184 = ( w149 & w205 ) | ( w149 & ~w1945 ) | ( w205 & ~w1945 ) ;
  assign w3185 = w3183 | w3184 ;
  assign w3186 = w3182 | w3185 ;
  assign w3187 = w505 | w673 ;
  assign w3188 = w142 | w3187 ;
  assign w3189 = ( ~w142 & w269 ) | ( ~w142 & w3186 ) | ( w269 & w3186 ) ;
  assign w3190 = w3188 | w3189 ;
  assign w3191 = ( w263 & w459 ) | ( w263 & ~w723 ) | ( w459 & ~w723 ) ;
  assign w3192 = w144 | w2274 ;
  assign w3193 = ( ~w144 & w723 ) | ( ~w144 & w1229 ) | ( w723 & w1229 ) ;
  assign w3194 = w3192 | w3193 ;
  assign w3195 = w3191 | w3194 ;
  assign w3196 = w139 | w988 ;
  assign w3197 = w131 | w281 ;
  assign w3198 = ( ~w131 & w175 ) | ( ~w131 & w3196 ) | ( w175 & w3196 ) ;
  assign w3199 = w3197 | w3198 ;
  assign w3200 = w257 | w2452 ;
  assign w3201 = ( w147 & ~w2452 ) | ( w147 & w3199 ) | ( ~w2452 & w3199 ) ;
  assign w3202 = w3200 | w3201 ;
  assign w3203 = w1979 | w2808 ;
  assign w3204 = w3195 | w3203 ;
  assign w3205 = ( w1158 & ~w3195 ) | ( w1158 & w3202 ) | ( ~w3195 & w3202 ) ;
  assign w3206 = w3204 | w3205 ;
  assign w3207 = w1276 | w1835 ;
  assign w3208 = ( ~w1276 & w1400 ) | ( ~w1276 & w3206 ) | ( w1400 & w3206 ) ;
  assign w3209 = w3207 | w3208 ;
  assign w3210 = w95 | w220 ;
  assign w3211 = ( ~w95 & w165 ) | ( ~w95 & w3209 ) | ( w165 & w3209 ) ;
  assign w3212 = w3210 | w3211 ;
  assign w3213 = w421 | w860 ;
  assign w3214 = w624 | w3213 ;
  assign w3215 = ( w322 & w432 ) | ( w322 & ~w624 ) | ( w432 & ~w624 ) ;
  assign w3216 = w3214 | w3215 ;
  assign w3217 = w697 | w2169 ;
  assign w3218 = ( w164 & ~w2169 ) | ( w164 & w3216 ) | ( ~w2169 & w3216 ) ;
  assign w3219 = w3217 | w3218 ;
  assign w3220 = ( ~w225 & w1152 ) | ( ~w225 & w3219 ) | ( w1152 & w3219 ) ;
  assign w3221 = w1523 | w3212 ;
  assign w3222 = ( w225 & w511 ) | ( w225 & ~w1523 ) | ( w511 & ~w1523 ) ;
  assign w3223 = w3221 | w3222 ;
  assign w3224 = w3220 | w3223 ;
  assign w3225 = ( w326 & w1265 ) | ( w326 & ~w2060 ) | ( w1265 & ~w2060 ) ;
  assign w3226 = w3190 | w3224 ;
  assign w3227 = ( w1340 & w2060 ) | ( w1340 & ~w3190 ) | ( w2060 & ~w3190 ) ;
  assign w3228 = w3226 | w3227 ;
  assign w3229 = w3225 | w3228 ;
  assign w3230 = ( w253 & w393 ) | ( w253 & ~w458 ) | ( w393 & ~w458 ) ;
  assign w3231 = w133 | w3229 ;
  assign w3232 = ( ~w133 & w458 ) | ( ~w133 & w491 ) | ( w458 & w491 ) ;
  assign w3233 = w3231 | w3232 ;
  assign w3234 = w3230 | w3233 ;
  assign w3235 = ( w317 & w445 ) | ( w317 & ~w459 ) | ( w445 & ~w459 ) ;
  assign w3236 = w96 | w286 ;
  assign w3237 = ( ~w286 & w459 ) | ( ~w286 & w530 ) | ( w459 & w530 ) ;
  assign w3238 = w3236 | w3237 ;
  assign w3239 = w3235 | w3238 ;
  assign w3240 = ( w350 & w463 ) | ( w350 & ~w505 ) | ( w463 & ~w505 ) ;
  assign w3241 = w227 | w3239 ;
  assign w3242 = ( ~w227 & w505 ) | ( ~w227 & w516 ) | ( w505 & w516 ) ;
  assign w3243 = w3241 | w3242 ;
  assign w3244 = w3240 | w3243 ;
  assign w3245 = w512 | w901 ;
  assign w3246 = w283 | w3245 ;
  assign w3247 = ( w169 & ~w283 ) | ( w169 & w392 ) | ( ~w283 & w392 ) ;
  assign w3248 = w3246 | w3247 ;
  assign w3249 = ( ~w280 & w456 ) | ( ~w280 & w3248 ) | ( w456 & w3248 ) ;
  assign w3250 = w280 | w3249 ;
  assign w3251 = w139 | w419 ;
  assign w3252 = w593 | w1274 ;
  assign w3253 = w198 | w3252 ;
  assign w3254 = ( ~w198 & w470 ) | ( ~w198 & w3251 ) | ( w470 & w3251 ) ;
  assign w3255 = w3253 | w3254 ;
  assign w3256 = ( w309 & w722 ) | ( w309 & ~w817 ) | ( w722 & ~w817 ) ;
  assign w3257 = w759 | w3255 ;
  assign w3258 = ( ~w759 & w817 ) | ( ~w759 & w1030 ) | ( w817 & w1030 ) ;
  assign w3259 = w3257 | w3258 ;
  assign w3260 = w3256 | w3259 ;
  assign w3261 = w1165 | w2760 ;
  assign w3262 = w672 | w3261 ;
  assign w3263 = ( ~w672 & w1087 ) | ( ~w672 & w3260 ) | ( w1087 & w3260 ) ;
  assign w3264 = w3262 | w3263 ;
  assign w3265 = ( ~w310 & w326 ) | ( ~w310 & w822 ) | ( w326 & w822 ) ;
  assign w3266 = w3250 | w3264 ;
  assign w3267 = ( w310 & w511 ) | ( w310 & ~w3250 ) | ( w511 & ~w3250 ) ;
  assign w3268 = w3266 | w3267 ;
  assign w3269 = w3265 | w3268 ;
  assign w3270 = w409 | w663 ;
  assign w3271 = w104 | w3270 ;
  assign w3272 = ( ~w104 & w232 ) | ( ~w104 & w3269 ) | ( w232 & w3269 ) ;
  assign w3273 = w3271 | w3272 ;
  assign w3274 = w318 | w390 ;
  assign w3275 = w510 | w3274 ;
  assign w3276 = ( w76 & w168 ) | ( w76 & ~w510 ) | ( w168 & ~w510 ) ;
  assign w3277 = w3275 | w3276 ;
  assign w3278 = ( w178 & w215 ) | ( w178 & ~w255 ) | ( w215 & ~w255 ) ;
  assign w3279 = w133 | w3277 ;
  assign w3280 = ( ~w133 & w255 ) | ( ~w133 & w354 ) | ( w255 & w354 ) ;
  assign w3281 = w3279 | w3280 ;
  assign w3282 = w3278 | w3281 ;
  assign w3283 = w202 | w277 ;
  assign w3284 = ( ~w202 & w252 ) | ( ~w202 & w3282 ) | ( w252 & w3282 ) ;
  assign w3285 = w3283 | w3284 ;
  assign w3286 = w314 | w1031 ;
  assign w3287 = w122 | w3286 ;
  assign w3288 = ( ~w122 & w258 ) | ( ~w122 & w507 ) | ( w258 & w507 ) ;
  assign w3289 = w3287 | w3288 ;
  assign w3290 = ( w742 & ~w1460 ) | ( w742 & w3289 ) | ( ~w1460 & w3289 ) ;
  assign w3291 = w1595 | w3285 ;
  assign w3292 = ( w1460 & ~w1595 ) | ( w1460 & w1882 ) | ( ~w1595 & w1882 ) ;
  assign w3293 = w3291 | w3292 ;
  assign w3294 = w3290 | w3293 ;
  assign w3295 = ( w63 & w111 ) | ( w63 & ~w311 ) | ( w111 & ~w311 ) ;
  assign w3296 = w1281 | w3294 ;
  assign w3297 = ( w311 & w513 ) | ( w311 & ~w1281 ) | ( w513 & ~w1281 ) ;
  assign w3298 = w3296 | w3297 ;
  assign w3299 = w3295 | w3298 ;
  assign w3300 = ( w313 & w413 ) | ( w313 & ~w623 ) | ( w413 & ~w623 ) ;
  assign w3301 = w201 | w214 ;
  assign w3302 = ( ~w214 & w623 ) | ( ~w214 & w764 ) | ( w623 & w764 ) ;
  assign w3303 = w3301 | w3302 ;
  assign w3304 = w3300 | w3303 ;
  assign w3305 = ( w138 & w225 ) | ( w138 & ~w837 ) | ( w225 & ~w837 ) ;
  assign w3306 = w68 | w3304 ;
  assign w3307 = ( ~w68 & w837 ) | ( ~w68 & w1126 ) | ( w837 & w1126 ) ;
  assign w3308 = w3306 | w3307 ;
  assign w3309 = w3305 | w3308 ;
  assign w3310 = w595 | w802 ;
  assign w3311 = w161 | w3310 ;
  assign w3312 = ( ~w161 & w322 ) | ( ~w161 & w3309 ) | ( w322 & w3309 ) ;
  assign w3313 = w3311 | w3312 ;
  assign w3314 = ( w465 & w680 ) | ( w465 & ~w681 ) | ( w680 & ~w681 ) ;
  assign w3315 = w98 | w1566 ;
  assign w3316 = ( ~w98 & w681 ) | ( ~w98 & w1153 ) | ( w681 & w1153 ) ;
  assign w3317 = w3315 | w3316 ;
  assign w3318 = w3314 | w3317 ;
  assign w3319 = ( ~w59 & w423 ) | ( ~w59 & w3318 ) | ( w423 & w3318 ) ;
  assign w3320 = w59 | w3319 ;
  assign w3321 = ( w320 & w385 ) | ( w320 & ~w605 ) | ( w385 & ~w605 ) ;
  assign w3322 = w210 | w3320 ;
  assign w3323 = ( ~w210 & w605 ) | ( ~w210 & w674 ) | ( w605 & w674 ) ;
  assign w3324 = w3322 | w3323 ;
  assign w3325 = w3321 | w3324 ;
  assign w3326 = ( w3244 & ~w3313 ) | ( w3244 & w3325 ) | ( ~w3313 & w3325 ) ;
  assign w3327 = w3273 | w3299 ;
  assign w3328 = ( w87 & ~w3299 ) | ( w87 & w3313 ) | ( ~w3299 & w3313 ) ;
  assign w3329 = w3327 | w3328 ;
  assign w3330 = w3326 | w3329 ;
  assign w3331 = w627 | w723 ;
  assign w3332 = ( ~w627 & w1615 ) | ( ~w627 & w3330 ) | ( w1615 & w3330 ) ;
  assign w3333 = w3331 | w3332 ;
  assign w3334 = w128 | w345 ;
  assign w3335 = ( ~w128 & w226 ) | ( ~w128 & w3333 ) | ( w226 & w3333 ) ;
  assign w3336 = w3334 | w3335 ;
  assign w3337 = ( ~\pi20 & w3234 ) | ( ~\pi20 & w3336 ) | ( w3234 & w3336 ) ;
  assign w3338 = w3107 ^ w3337 ;
  assign w3339 = w3159 ^ w3338 ;
  assign w3340 = ( w263 & w277 ) | ( w263 & ~w389 ) | ( w277 & ~w389 ) ;
  assign w3341 = w124 | w147 ;
  assign w3342 = ( ~w147 & w389 ) | ( ~w147 & w663 ) | ( w389 & w663 ) ;
  assign w3343 = w3341 | w3342 ;
  assign w3344 = w3340 | w3343 ;
  assign w3345 = w167 | w802 ;
  assign w3346 = ( ~w167 & w640 ) | ( ~w167 & w3344 ) | ( w640 & w3344 ) ;
  assign w3347 = w3345 | w3346 ;
  assign w3348 = w232 | w1422 ;
  assign w3349 = ( w175 & ~w232 ) | ( w175 & w255 ) | ( ~w232 & w255 ) ;
  assign w3350 = w3348 | w3349 ;
  assign w3351 = w201 | w673 ;
  assign w3352 = ( ~w201 & w341 ) | ( ~w201 & w536 ) | ( w341 & w536 ) ;
  assign w3353 = w3351 | w3352 ;
  assign w3354 = ( w202 & ~w253 ) | ( w202 & w1154 ) | ( ~w253 & w1154 ) ;
  assign w3355 = w468 | w1087 ;
  assign w3356 = ( w253 & w350 ) | ( w253 & ~w1087 ) | ( w350 & ~w1087 ) ;
  assign w3357 = w3355 | w3356 ;
  assign w3358 = w3354 | w3357 ;
  assign w3359 = ( w3002 & w3353 ) | ( w3002 & ~w3358 ) | ( w3353 & ~w3358 ) ;
  assign w3360 = w3358 | w3359 ;
  assign w3361 = w2196 | w3347 ;
  assign w3362 = ( ~w3347 & w3350 ) | ( ~w3347 & w3360 ) | ( w3350 & w3360 ) ;
  assign w3363 = w3361 | w3362 ;
  assign w3364 = w273 | w340 ;
  assign w3365 = ( ~w273 & w784 ) | ( ~w273 & w3363 ) | ( w784 & w3363 ) ;
  assign w3366 = w3364 | w3365 ;
  assign w3367 = ( w339 & w567 ) | ( w339 & ~w637 ) | ( w567 & ~w637 ) ;
  assign w3368 = w161 | w3366 ;
  assign w3369 = ( ~w161 & w637 ) | ( ~w161 & w642 ) | ( w637 & w642 ) ;
  assign w3370 = w3368 | w3369 ;
  assign w3371 = w3367 | w3370 ;
  assign w3372 = ( w525 & w560 ) | ( w525 & ~w817 ) | ( w560 & ~w817 ) ;
  assign w3373 = w281 | w317 ;
  assign w3374 = ( ~w317 & w817 ) | ( ~w317 & w1274 ) | ( w817 & w1274 ) ;
  assign w3375 = w3373 | w3374 ;
  assign w3376 = w3372 | w3375 ;
  assign w3377 = w252 | w641 ;
  assign w3378 = ( ~w252 & w524 ) | ( ~w252 & w3376 ) | ( w524 & w3376 ) ;
  assign w3379 = w3377 | w3378 ;
  assign w3380 = ( w262 & w725 ) | ( w262 & ~w951 ) | ( w725 & ~w951 ) ;
  assign w3381 = w111 | w731 ;
  assign w3382 = ( ~w111 & w951 ) | ( ~w111 & w980 ) | ( w951 & w980 ) ;
  assign w3383 = w3381 | w3382 ;
  assign w3384 = w3380 | w3383 ;
  assign w3385 = w530 | w3384 ;
  assign w3386 = ( ~w179 & w198 ) | ( ~w179 & w2782 ) | ( w198 & w2782 ) ;
  assign w3387 = w179 | w3386 ;
  assign w3388 = w447 | w488 ;
  assign w3389 = w3387 | w3388 ;
  assign w3390 = ( w385 & w3385 ) | ( w385 & ~w3387 ) | ( w3385 & ~w3387 ) ;
  assign w3391 = w3389 | w3390 ;
  assign w3392 = ( w96 & w416 ) | ( w96 & ~w1513 ) | ( w416 & ~w1513 ) ;
  assign w3393 = w3379 | w3391 ;
  assign w3394 = ( w1513 & w1560 ) | ( w1513 & ~w3379 ) | ( w1560 & ~w3379 ) ;
  assign w3395 = w3393 | w3394 ;
  assign w3396 = w3392 | w3395 ;
  assign w3397 = ( w208 & ~w383 ) | ( w208 & w742 ) | ( ~w383 & w742 ) ;
  assign w3398 = w507 | w3396 ;
  assign w3399 = ( w383 & w445 ) | ( w383 & ~w507 ) | ( w445 & ~w507 ) ;
  assign w3400 = w3398 | w3399 ;
  assign w3401 = w3397 | w3400 ;
  assign w3402 = ( w215 & w388 ) | ( w215 & ~w429 ) | ( w388 & ~w429 ) ;
  assign w3403 = ~w136 & w1993 ;
  assign w3404 = ( ~w136 & w429 ) | ( ~w136 & w431 ) | ( w429 & w431 ) ;
  assign w3405 = w3403 & ~w3404 ;
  assign w3406 = ~w3402 & w3405 ;
  assign w3407 = ( w523 & w2327 ) | ( w523 & w3406 ) | ( w2327 & w3406 ) ;
  assign w3408 = w3371 | w3401 ;
  assign w3409 = ( ~w886 & w3401 ) | ( ~w886 & w3406 ) | ( w3401 & w3406 ) ;
  assign w3410 = ~w3408 & w3409 ;
  assign w3411 = ~w3407 & w3410 ;
  assign w3412 = ( w144 & w203 ) | ( w144 & ~w310 ) | ( w203 & ~w310 ) ;
  assign w3413 = ~w572 & w3411 ;
  assign w3414 = ( w310 & w511 ) | ( w310 & ~w572 ) | ( w511 & ~w572 ) ;
  assign w3415 = w3413 & ~w3414 ;
  assign w3416 = ~w3412 & w3415 ;
  assign w3417 = w128 | w596 ;
  assign w3418 = ( w128 & ~w210 ) | ( w128 & w3416 ) | ( ~w210 & w3416 ) ;
  assign w3419 = ~w3417 & w3418 ;
  assign w3420 = w592 ^ w2997 ;
  assign w3421 = w721 ^ w3420 ;
  assign w3422 = ( \pi29 & \pi31 ) | ( \pi29 & w721 ) | ( \pi31 & w721 ) ;
  assign w3423 = ( \pi29 & ~\pi30 ) | ( \pi29 & w3422 ) | ( ~\pi30 & w3422 ) ;
  assign w3424 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w3422 ) | ( \pi30 & w3422 ) ;
  assign w3425 = ( \pi29 & w883 ) | ( \pi29 & ~w3424 ) | ( w883 & ~w3424 ) ;
  assign w3426 = ( w592 & w3424 ) | ( w592 & w3425 ) | ( w3424 & w3425 ) ;
  assign w3427 = ~\pi31 & w3426 ;
  assign w3428 = ( w3423 & ~w3425 ) | ( w3423 & w3427 ) | ( ~w3425 & w3427 ) ;
  assign w3429 = ( w37 & w3421 ) | ( w37 & w3428 ) | ( w3421 & w3428 ) ;
  assign w3430 = w3428 | w3429 ;
  assign w3431 = ( w3234 & w3419 ) | ( w3234 & ~w3430 ) | ( w3419 & ~w3430 ) ;
  assign w3432 = w3234 ^ w3336 ;
  assign w3433 = \pi20 ^ w3432 ;
  assign w3434 = w381 ^ w2998 ;
  assign w3435 = w592 ^ w3434 ;
  assign w3436 = ( \pi29 & \pi31 ) | ( \pi29 & w592 ) | ( \pi31 & w592 ) ;
  assign w3437 = ( \pi29 & ~\pi30 ) | ( \pi29 & w3436 ) | ( ~\pi30 & w3436 ) ;
  assign w3438 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w3436 ) | ( \pi30 & w3436 ) ;
  assign w3439 = ( ~\pi29 & w721 ) | ( ~\pi29 & w3438 ) | ( w721 & w3438 ) ;
  assign w3440 = ( w381 & ~w3438 ) | ( w381 & w3439 ) | ( ~w3438 & w3439 ) ;
  assign w3441 = \pi31 | w3440 ;
  assign w3442 = ( w3437 & w3439 ) | ( w3437 & ~w3441 ) | ( w3439 & ~w3441 ) ;
  assign w3443 = ( w37 & ~w3435 ) | ( w37 & w3442 ) | ( ~w3435 & w3442 ) ;
  assign w3444 = w3442 | w3443 ;
  assign w3445 = ( w3431 & w3433 ) | ( w3431 & ~w3444 ) | ( w3433 & ~w3444 ) ;
  assign w3446 = \pi28 ^ \pi29 ;
  assign w3447 = \pi26 ^ \pi27 ;
  assign w3448 = w3446 & w3447 ;
  assign w3449 = ( w466 & w663 ) | ( w466 & ~w1030 ) | ( w663 & ~w1030 ) ;
  assign w3450 = w225 | w354 ;
  assign w3451 = ( ~w354 & w1030 ) | ( ~w354 & w1086 ) | ( w1030 & w1086 ) ;
  assign w3452 = w3450 | w3451 ;
  assign w3453 = w3449 | w3452 ;
  assign w3454 = w324 | w758 ;
  assign w3455 = w3453 | w3454 ;
  assign w3456 = ( w169 & w2470 ) | ( w169 & ~w3453 ) | ( w2470 & ~w3453 ) ;
  assign w3457 = w3455 | w3456 ;
  assign w3458 = w114 | w569 ;
  assign w3459 = ( ~w114 & w383 ) | ( ~w114 & w3457 ) | ( w383 & w3457 ) ;
  assign w3460 = w3458 | w3459 ;
  assign w3461 = ( w422 & w458 ) | ( w422 & ~w511 ) | ( w458 & ~w511 ) ;
  assign w3462 = w115 | w283 ;
  assign w3463 = ( ~w283 & w511 ) | ( ~w283 & w533 ) | ( w511 & w533 ) ;
  assign w3464 = w3462 | w3463 ;
  assign w3465 = w3461 | w3464 ;
  assign w3466 = w175 | w697 ;
  assign w3467 = ( ~w175 & w567 ) | ( ~w175 & w3465 ) | ( w567 & w3465 ) ;
  assign w3468 = w3466 | w3467 ;
  assign w3469 = w124 | w1340 ;
  assign w3470 = ( ~w124 & w409 ) | ( ~w124 & w2626 ) | ( w409 & w2626 ) ;
  assign w3471 = w3469 | w3470 ;
  assign w3472 = w122 | w642 ;
  assign w3473 = ( ~w122 & w505 ) | ( ~w122 & w956 ) | ( w505 & w956 ) ;
  assign w3474 = w3472 | w3473 ;
  assign w3475 = w362 | w897 ;
  assign w3476 = w74 | w3475 ;
  assign w3477 = ( ~w74 & w257 ) | ( ~w74 & w3474 ) | ( w257 & w3474 ) ;
  assign w3478 = w3476 | w3477 ;
  assign w3479 = w316 | w421 ;
  assign w3480 = ( w316 & w359 ) | ( w316 & ~w3478 ) | ( w359 & ~w3478 ) ;
  assign w3481 = ~w3479 & w3480 ;
  assign w3482 = w273 | w623 ;
  assign w3483 = w3468 | w3482 ;
  assign w3484 = ( w3468 & ~w3471 ) | ( w3468 & w3481 ) | ( ~w3471 & w3481 ) ;
  assign w3485 = ~w3483 & w3484 ;
  assign w3486 = ( w320 & w445 ) | ( w320 & ~w456 ) | ( w445 & ~w456 ) ;
  assign w3487 = ~w103 & w3485 ;
  assign w3488 = ( ~w103 & w456 ) | ( ~w103 & w889 ) | ( w456 & w889 ) ;
  assign w3489 = w3487 & ~w3488 ;
  assign w3490 = ~w3486 & w3489 ;
  assign w3491 = w84 | w764 ;
  assign w3492 = ( ~w84 & w674 ) | ( ~w84 & w2147 ) | ( w674 & w2147 ) ;
  assign w3493 = w3491 | w3492 ;
  assign w3494 = w230 | w318 ;
  assign w3495 = w980 | w3494 ;
  assign w3496 = ( w282 & w388 ) | ( w282 & ~w3494 ) | ( w388 & ~w3494 ) ;
  assign w3497 = w3495 | w3496 ;
  assign w3498 = w722 | w1094 ;
  assign w3499 = w165 | w3498 ;
  assign w3500 = ( ~w165 & w512 ) | ( ~w165 & w3497 ) | ( w512 & w3497 ) ;
  assign w3501 = w3499 | w3500 ;
  assign w3502 = w104 | w264 ;
  assign w3503 = ( w82 & ~w264 ) | ( w82 & w514 ) | ( ~w264 & w514 ) ;
  assign w3504 = w3502 | w3503 ;
  assign w3505 = w350 | w468 ;
  assign w3506 = ( w253 & ~w468 ) | ( w253 & w3504 ) | ( ~w468 & w3504 ) ;
  assign w3507 = w3505 | w3506 ;
  assign w3508 = w315 | w951 ;
  assign w3509 = w3507 | w3508 ;
  assign w3510 = ( w1158 & w3501 ) | ( w1158 & ~w3507 ) | ( w3501 & ~w3507 ) ;
  assign w3511 = w3509 | w3510 ;
  assign w3512 = w1565 | w3493 ;
  assign w3513 = ( w887 & ~w3493 ) | ( w887 & w3511 ) | ( ~w3493 & w3511 ) ;
  assign w3514 = w3512 | w3513 ;
  assign w3515 = w88 | w286 ;
  assign w3516 = w731 | w3515 ;
  assign w3517 = ( ~w731 & w1207 ) | ( ~w731 & w3514 ) | ( w1207 & w3514 ) ;
  assign w3518 = w3516 | w3517 ;
  assign w3519 = w393 | w491 ;
  assign w3520 = w180 | w3519 ;
  assign w3521 = ( ~w180 & w203 ) | ( ~w180 & w3518 ) | ( w203 & w3518 ) ;
  assign w3522 = w3520 | w3521 ;
  assign w3523 = w339 | w608 ;
  assign w3524 = ( ~w339 & w534 ) | ( ~w339 & w1166 ) | ( w534 & w1166 ) ;
  assign w3525 = w3523 | w3524 ;
  assign w3526 = ( w111 & w219 ) | ( w111 & ~w570 ) | ( w219 & ~w570 ) ;
  assign w3527 = w51 | w3525 ;
  assign w3528 = ( ~w51 & w570 ) | ( ~w51 & w726 ) | ( w570 & w726 ) ;
  assign w3529 = w3527 | w3528 ;
  assign w3530 = w3526 | w3529 ;
  assign w3531 = w2873 | w3530 ;
  assign w3532 = w3490 & ~w3531 ;
  assign w3533 = ( w3320 & w3490 ) | ( w3320 & w3522 ) | ( w3490 & w3522 ) ;
  assign w3534 = w3532 & ~w3533 ;
  assign w3535 = w223 | w224 ;
  assign w3536 = w3460 | w3535 ;
  assign w3537 = ( ~w1979 & w3460 ) | ( ~w1979 & w3534 ) | ( w3460 & w3534 ) ;
  assign w3538 = ~w3536 & w3537 ;
  assign w3539 = w490 | w998 ;
  assign w3540 = ( ~w488 & w998 ) | ( ~w488 & w3538 ) | ( w998 & w3538 ) ;
  assign w3541 = ~w3539 & w3540 ;
  assign w3542 = w459 | w787 ;
  assign w3543 = w822 | w3542 ;
  assign w3544 = ( ~w202 & w822 ) | ( ~w202 & w3541 ) | ( w822 & w3541 ) ;
  assign w3545 = ~w3543 & w3544 ;
  assign w3546 = w277 | w516 ;
  assign w3547 = ( w277 & ~w285 ) | ( w277 & w3545 ) | ( ~w285 & w3545 ) ;
  assign w3548 = ~w3546 & w3547 ;
  assign w3549 = ~w3446 & w3447 ;
  assign w3550 = ( w253 & w496 ) | ( w253 & ~w533 ) | ( w496 & ~w533 ) ;
  assign w3551 = w86 | w230 ;
  assign w3552 = ( ~w230 & w533 ) | ( ~w230 & w722 ) | ( w533 & w722 ) ;
  assign w3553 = w3551 | w3552 ;
  assign w3554 = w3550 | w3553 ;
  assign w3555 = w1030 | w3554 ;
  assign w3556 = w802 | w1126 ;
  assign w3557 = w139 | w3556 ;
  assign w3558 = ( ~w139 & w278 ) | ( ~w139 & w2169 ) | ( w278 & w2169 ) ;
  assign w3559 = w3557 | w3558 ;
  assign w3560 = w524 | w1001 ;
  assign w3561 = ( ~w524 & w628 ) | ( ~w524 & w3559 ) | ( w628 & w3559 ) ;
  assign w3562 = w3560 | w3561 ;
  assign w3563 = w449 | w723 ;
  assign w3564 = ( w315 & ~w449 ) | ( w315 & w513 ) | ( ~w449 & w513 ) ;
  assign w3565 = w3563 | w3564 ;
  assign w3566 = w567 | w764 ;
  assign w3567 = w210 | w3566 ;
  assign w3568 = ( w124 & ~w210 ) | ( w124 & w385 ) | ( ~w210 & w385 ) ;
  assign w3569 = w3567 | w3568 ;
  assign w3570 = ( w218 & w466 ) | ( w218 & ~w470 ) | ( w466 & ~w470 ) ;
  assign w3571 = w410 | w3569 ;
  assign w3572 = ( w470 & w637 ) | ( w470 & ~w3569 ) | ( w637 & ~w3569 ) ;
  assign w3573 = w3571 | w3572 ;
  assign w3574 = w3570 | w3573 ;
  assign w3575 = w430 | w595 ;
  assign w3576 = w205 | w3575 ;
  assign w3577 = ( ~w205 & w429 ) | ( ~w205 & w3574 ) | ( w429 & w3574 ) ;
  assign w3578 = w3576 | w3577 ;
  assign w3579 = ( w120 & w149 ) | ( w120 & ~w214 ) | ( w149 & ~w214 ) ;
  assign w3580 = w3565 | w3578 ;
  assign w3581 = ( w214 & w311 ) | ( w214 & ~w3565 ) | ( w311 & ~w3565 ) ;
  assign w3582 = w3580 | w3581 ;
  assign w3583 = w3579 | w3582 ;
  assign w3584 = w1069 | w1617 ;
  assign w3585 = w3562 | w3584 ;
  assign w3586 = ( w572 & ~w3562 ) | ( w572 & w3583 ) | ( ~w3562 & w3583 ) ;
  assign w3587 = w3585 | w3586 ;
  assign w3588 = w135 | w314 ;
  assign w3589 = ( ~w135 & w284 ) | ( ~w135 & w3587 ) | ( w284 & w3587 ) ;
  assign w3590 = w3588 | w3589 ;
  assign w3591 = ( w318 & w342 ) | ( w318 & ~w390 ) | ( w342 & ~w390 ) ;
  assign w3592 = w203 | w1566 ;
  assign w3593 = ( ~w203 & w390 ) | ( ~w203 & w509 ) | ( w390 & w509 ) ;
  assign w3594 = w3592 | w3593 ;
  assign w3595 = w3591 | w3594 ;
  assign w3596 = w266 | w787 ;
  assign w3597 = w180 | w3596 ;
  assign w3598 = ( ~w180 & w215 ) | ( ~w180 & w3595 ) | ( w215 & w3595 ) ;
  assign w3599 = w3597 | w3598 ;
  assign w3600 = ( w226 & w255 ) | ( w226 & ~w277 ) | ( w255 & ~w277 ) ;
  assign w3601 = w63 | w116 ;
  assign w3602 = ( ~w116 & w277 ) | ( ~w116 & w506 ) | ( w277 & w506 ) ;
  assign w3603 = w3601 | w3602 ;
  assign w3604 = w3600 | w3603 ;
  assign w3605 = ( ~w491 & w2091 ) | ( ~w491 & w3604 ) | ( w2091 & w3604 ) ;
  assign w3606 = w620 | w3599 ;
  assign w3607 = ( w491 & w534 ) | ( w491 & ~w3599 ) | ( w534 & ~w3599 ) ;
  assign w3608 = w3606 | w3607 ;
  assign w3609 = w3605 | w3608 ;
  assign w3610 = ( ~w273 & w1302 ) | ( ~w273 & w3609 ) | ( w1302 & w3609 ) ;
  assign w3611 = w3482 | w3610 ;
  assign w3612 = ( w201 & w352 ) | ( w201 & ~w411 ) | ( w352 & ~w411 ) ;
  assign w3613 = w127 | w3611 ;
  assign w3614 = ( ~w127 & w411 ) | ( ~w127 & w573 ) | ( w411 & w573 ) ;
  assign w3615 = w3613 | w3614 ;
  assign w3616 = w3612 | w3615 ;
  assign w3617 = ( w225 & ~w420 ) | ( w225 & w725 ) | ( ~w420 & w725 ) ;
  assign w3618 = w420 | w3617 ;
  assign w3619 = ( w142 & w143 ) | ( w142 & ~w419 ) | ( w143 & ~w419 ) ;
  assign w3620 = w988 | w3618 ;
  assign w3621 = ( w419 & w1086 ) | ( w419 & ~w3618 ) | ( w1086 & ~w3618 ) ;
  assign w3622 = w3620 | w3621 ;
  assign w3623 = w3619 | w3622 ;
  assign w3624 = ( w223 & ~w860 ) | ( w223 & w2092 ) | ( ~w860 & w2092 ) ;
  assign w3625 = w3616 | w3623 ;
  assign w3626 = ( w860 & w980 ) | ( w860 & ~w3623 ) | ( w980 & ~w3623 ) ;
  assign w3627 = w3625 | w3626 ;
  assign w3628 = w3624 | w3627 ;
  assign w3629 = ( w88 & ~w114 ) | ( w88 & w322 ) | ( ~w114 & w322 ) ;
  assign w3630 = w114 | w3629 ;
  assign w3631 = w316 | w3630 ;
  assign w3632 = ( w268 & w3387 ) | ( w268 & ~w3630 ) | ( w3387 & ~w3630 ) ;
  assign w3633 = w3631 | w3632 ;
  assign w3634 = w528 | w1629 ;
  assign w3635 = w3633 | w3634 ;
  assign w3636 = ( w462 & w3628 ) | ( w462 & ~w3633 ) | ( w3628 & ~w3633 ) ;
  assign w3637 = w3635 | w3636 ;
  assign w3638 = ( w1051 & ~w1283 ) | ( w1051 & w3555 ) | ( ~w1283 & w3555 ) ;
  assign w3639 = w3590 | w3637 ;
  assign w3640 = ( w1283 & w1565 ) | ( w1283 & ~w3590 ) | ( w1565 & ~w3590 ) ;
  assign w3641 = w3639 | w3640 ;
  assign w3642 = w3638 | w3641 ;
  assign w3643 = ( w169 & w317 ) | ( w169 & ~w358 ) | ( w317 & ~w358 ) ;
  assign w3644 = w167 | w3642 ;
  assign w3645 = ( ~w167 & w358 ) | ( ~w167 & w490 ) | ( w358 & w490 ) ;
  assign w3646 = w3644 | w3645 ;
  assign w3647 = w3643 | w3646 ;
  assign w3648 = ( \pi26 & \pi27 ) | ( \pi26 & w42 ) | ( \pi27 & w42 ) ;
  assign w3649 = w42 ^ w3648 ;
  assign w3650 = w723 | w802 ;
  assign w3651 = w362 | w3650 ;
  assign w3652 = ( w316 & ~w362 ) | ( w316 & w571 ) | ( ~w362 & w571 ) ;
  assign w3653 = w3651 | w3652 ;
  assign w3654 = ( w203 & w466 ) | ( w203 & ~w641 ) | ( w466 & ~w641 ) ;
  assign w3655 = w86 | w3653 ;
  assign w3656 = ( ~w86 & w641 ) | ( ~w86 & w1153 ) | ( w641 & w1153 ) ;
  assign w3657 = w3655 | w3656 ;
  assign w3658 = w3654 | w3657 ;
  assign w3659 = w210 | w899 ;
  assign w3660 = w1513 | w3659 ;
  assign w3661 = ( ~w1513 & w2079 ) | ( ~w1513 & w3658 ) | ( w2079 & w3658 ) ;
  assign w3662 = w3660 | w3661 ;
  assign w3663 = ( w317 & ~w341 ) | ( w317 & w1615 ) | ( ~w341 & w1615 ) ;
  assign w3664 = w414 | w3662 ;
  assign w3665 = ( w341 & ~w414 ) | ( w341 & w628 ) | ( ~w414 & w628 ) ;
  assign w3666 = w3664 | w3665 ;
  assign w3667 = w3663 | w3666 ;
  assign w3668 = w570 | w1340 ;
  assign w3669 = w310 | w3668 ;
  assign w3670 = ( w82 & ~w310 ) | ( w82 & w506 ) | ( ~w310 & w506 ) ;
  assign w3671 = w3669 | w3670 ;
  assign w3672 = ( ~w415 & w424 ) | ( ~w415 & w3671 ) | ( w424 & w3671 ) ;
  assign w3673 = w415 | w3672 ;
  assign w3674 = w625 | w787 ;
  assign w3675 = w490 | w3674 ;
  assign w3676 = ( w344 & ~w490 ) | ( w344 & w495 ) | ( ~w490 & w495 ) ;
  assign w3677 = w3675 | w3676 ;
  assign w3678 = w422 | w1031 ;
  assign w3679 = w2704 | w3678 ;
  assign w3680 = ( w325 & w2358 ) | ( w325 & ~w2704 ) | ( w2358 & ~w2704 ) ;
  assign w3681 = w3679 | w3680 ;
  assign w3682 = ( w459 & w465 ) | ( w459 & ~w567 ) | ( w465 & ~w567 ) ;
  assign w3683 = w3677 | w3681 ;
  assign w3684 = ( w567 & w980 ) | ( w567 & ~w3677 ) | ( w980 & ~w3677 ) ;
  assign w3685 = w3683 | w3684 ;
  assign w3686 = w3682 | w3685 ;
  assign w3687 = w322 | w533 ;
  assign w3688 = w101 | w3687 ;
  assign w3689 = ( ~w101 & w320 ) | ( ~w101 & w3686 ) | ( w320 & w3686 ) ;
  assign w3690 = w3688 | w3689 ;
  assign w3691 = w386 | w467 ;
  assign w3692 = ( w342 & ~w386 ) | ( w342 & w420 ) | ( ~w386 & w420 ) ;
  assign w3693 = w3691 | w3692 ;
  assign w3694 = w345 | w389 ;
  assign w3695 = w1883 | w3694 ;
  assign w3696 = ( w59 & w1363 ) | ( w59 & ~w1883 ) | ( w1363 & ~w1883 ) ;
  assign w3697 = w3695 | w3696 ;
  assign w3698 = ( ~w1990 & w3673 ) | ( ~w1990 & w3697 ) | ( w3673 & w3697 ) ;
  assign w3699 = w196 | w3690 ;
  assign w3700 = ( w1990 & ~w3690 ) | ( w1990 & w3693 ) | ( ~w3690 & w3693 ) ;
  assign w3701 = w3699 | w3700 ;
  assign w3702 = w3698 | w3701 ;
  assign w3703 = ( w103 & ~w214 ) | ( w103 & w1736 ) | ( ~w214 & w1736 ) ;
  assign w3704 = w3667 | w3702 ;
  assign w3705 = ( w214 & w262 ) | ( w214 & ~w3667 ) | ( w262 & ~w3667 ) ;
  assign w3706 = w3704 | w3705 ;
  assign w3707 = w3703 | w3706 ;
  assign w3708 = ( w286 & w513 ) | ( w286 & ~w697 ) | ( w513 & ~w697 ) ;
  assign w3709 = w285 | w3707 ;
  assign w3710 = ( ~w285 & w697 ) | ( ~w285 & w1126 ) | ( w697 & w1126 ) ;
  assign w3711 = w3709 | w3710 ;
  assign w3712 = w3708 | w3711 ;
  assign w3713 = w51 | w783 ;
  assign w3714 = ( ~w51 & w488 ) | ( ~w51 & w3712 ) | ( w488 & w3712 ) ;
  assign w3715 = w3713 | w3714 ;
  assign w3716 = ( \pi26 & \pi27 ) | ( \pi26 & \pi28 ) | ( \pi27 & \pi28 ) ;
  assign w3717 = \pi28 ^ w3716 ;
  assign w3718 = w3647 & ~w3649 ;
  assign w3719 = w3715 & w3717 ;
  assign w3720 = ( w3647 & ~w3718 ) | ( w3647 & w3719 ) | ( ~w3718 & w3719 ) ;
  assign w3721 = ( w381 & ~w2999 ) | ( w381 & w3094 ) | ( ~w2999 & w3094 ) ;
  assign w3722 = ( w3094 & ~w3647 ) | ( w3094 & w3721 ) | ( ~w3647 & w3721 ) ;
  assign w3723 = ( w3647 & w3715 ) | ( w3647 & ~w3722 ) | ( w3715 & ~w3722 ) ;
  assign w3724 = w3548 ^ w3723 ;
  assign w3725 = w3715 ^ w3724 ;
  assign w3726 = w3548 | w3549 ;
  assign w3727 = ~w3720 & w3725 ;
  assign w3728 = ( w3448 & w3720 ) | ( w3448 & ~w3727 ) | ( w3720 & ~w3727 ) ;
  assign w3729 = ( ~w3548 & w3726 ) | ( ~w3548 & w3728 ) | ( w3726 & w3728 ) ;
  assign w3730 = \pi29 ^ w3729 ;
  assign w3731 = ( w3339 & ~w3445 ) | ( w3339 & w3730 ) | ( ~w3445 & w3730 ) ;
  assign w3732 = ( w3107 & w3159 ) | ( w3107 & w3337 ) | ( w3159 & w3337 ) ;
  assign w3733 = ( w509 & w511 ) | ( w509 & ~w663 ) | ( w511 & ~w663 ) ;
  assign w3734 = w210 | w385 ;
  assign w3735 = ( ~w385 & w663 ) | ( ~w385 & w1086 ) | ( w663 & w1086 ) ;
  assign w3736 = w3734 | w3735 ;
  assign w3737 = w3733 | w3736 ;
  assign w3738 = w223 | w353 ;
  assign w3739 = w44 | w3738 ;
  assign w3740 = ( ~w44 & w118 ) | ( ~w44 & w3737 ) | ( w118 & w3737 ) ;
  assign w3741 = w3739 | w3740 ;
  assign w3742 = ( w133 & w147 ) | ( w133 & ~w340 ) | ( w147 & ~w340 ) ;
  assign w3743 = w101 | w177 ;
  assign w3744 = ( ~w101 & w340 ) | ( ~w101 & w560 ) | ( w340 & w560 ) ;
  assign w3745 = w3743 | w3744 ;
  assign w3746 = w3742 | w3745 ;
  assign w3747 = ( ~w221 & w571 ) | ( ~w221 & w3746 ) | ( w571 & w3746 ) ;
  assign w3748 = w221 | w3747 ;
  assign w3749 = w725 | w3565 ;
  assign w3750 = ( w74 & w1496 ) | ( w74 & ~w3565 ) | ( w1496 & ~w3565 ) ;
  assign w3751 = w3749 | w3750 ;
  assign w3752 = w209 | w389 ;
  assign w3753 = w144 | w3752 ;
  assign w3754 = ( ~w144 & w203 ) | ( ~w144 & w3751 ) | ( w203 & w3751 ) ;
  assign w3755 = w3753 | w3754 ;
  assign w3756 = ( w281 & w344 ) | ( w281 & ~w354 ) | ( w344 & ~w354 ) ;
  assign w3757 = w143 | w3755 ;
  assign w3758 = ( ~w143 & w354 ) | ( ~w143 & w361 ) | ( w354 & w361 ) ;
  assign w3759 = w3757 | w3758 ;
  assign w3760 = w3756 | w3759 ;
  assign w3761 = ( ~w59 & w637 ) | ( ~w59 & w3760 ) | ( w637 & w3760 ) ;
  assign w3762 = w59 | w3761 ;
  assign w3763 = ( ~w218 & w2703 ) | ( ~w218 & w3741 ) | ( w2703 & w3741 ) ;
  assign w3764 = w3748 | w3762 ;
  assign w3765 = ( w218 & w219 ) | ( w218 & ~w3748 ) | ( w219 & ~w3748 ) ;
  assign w3766 = w3764 | w3765 ;
  assign w3767 = w3763 | w3766 ;
  assign w3768 = ( w104 & w256 ) | ( w104 & ~w419 ) | ( w256 & ~w419 ) ;
  assign w3769 = w1566 | w3767 ;
  assign w3770 = ( w419 & w625 ) | ( w419 & ~w1566 ) | ( w625 & ~w1566 ) ;
  assign w3771 = w3769 | w3770 ;
  assign w3772 = w3768 | w3771 ;
  assign w3773 = w463 | w662 ;
  assign w3774 = w322 | w3773 ;
  assign w3775 = ( ~w322 & w415 ) | ( ~w322 & w3772 ) | ( w415 & w3772 ) ;
  assign w3776 = w3774 | w3775 ;
  assign w3777 = w206 | w1094 ;
  assign w3778 = ( w257 & w408 ) | ( w257 & ~w458 ) | ( w408 & ~w458 ) ;
  assign w3779 = w229 | w3777 ;
  assign w3780 = ( ~w229 & w458 ) | ( ~w229 & w1229 ) | ( w458 & w1229 ) ;
  assign w3781 = w3779 | w3780 ;
  assign w3782 = w3778 | w3781 ;
  assign w3783 = w504 | w642 ;
  assign w3784 = w254 | w3783 ;
  assign w3785 = ( w198 & ~w254 ) | ( w198 & w287 ) | ( ~w254 & w287 ) ;
  assign w3786 = w3784 | w3785 ;
  assign w3787 = w951 | w1030 ;
  assign w3788 = w1413 | w3787 ;
  assign w3789 = ( w126 & w492 ) | ( w126 & ~w1413 ) | ( w492 & ~w1413 ) ;
  assign w3790 = w3788 | w3789 ;
  assign w3791 = ( ~w116 & w3786 ) | ( ~w116 & w3790 ) | ( w3786 & w3790 ) ;
  assign w3792 = w1357 | w3782 ;
  assign w3793 = ( w116 & w456 ) | ( w116 & ~w3782 ) | ( w456 & ~w3782 ) ;
  assign w3794 = w3792 | w3793 ;
  assign w3795 = w3791 | w3794 ;
  assign w3796 = ( w1069 & w1400 ) | ( w1069 & ~w1977 ) | ( w1400 & ~w1977 ) ;
  assign w3797 = w3776 | w3795 ;
  assign w3798 = ( w141 & w1977 ) | ( w141 & ~w3795 ) | ( w1977 & ~w3795 ) ;
  assign w3799 = w3797 | w3798 ;
  assign w3800 = w3796 | w3799 ;
  assign w3801 = ( w120 & w180 ) | ( w120 & ~w447 ) | ( w180 & ~w447 ) ;
  assign w3802 = w84 | w3800 ;
  assign w3803 = ( ~w84 & w447 ) | ( ~w84 & w860 ) | ( w447 & w860 ) ;
  assign w3804 = w3802 | w3803 ;
  assign w3805 = w3801 | w3804 ;
  assign w3806 = ( w3159 & ~w3732 ) | ( w3159 & w3805 ) | ( ~w3732 & w3805 ) ;
  assign w3807 = w3732 ^ w3805 ;
  assign w3808 = w3159 ^ w3807 ;
  assign w3809 = w3647 ^ w3721 ;
  assign w3810 = w3094 ^ w3809 ;
  assign w3811 = ~w37 & w3810 ;
  assign w3812 = ~w381 & w3098 ;
  assign w3813 = ( w3810 & ~w3811 ) | ( w3810 & w3812 ) | ( ~w3811 & w3812 ) ;
  assign w3814 = ( \pi29 & \pi30 ) | ( \pi29 & w3647 ) | ( \pi30 & w3647 ) ;
  assign w3815 = \pi31 | w3814 ;
  assign w3816 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w3094 ) | ( \pi30 & w3094 ) ;
  assign w3817 = ( \pi29 & \pi31 ) | ( \pi29 & w3816 ) | ( \pi31 & w3816 ) ;
  assign w3818 = ( w3813 & w3815 ) | ( w3813 & ~w3817 ) | ( w3815 & ~w3817 ) ;
  assign w3819 = w3731 ^ w3808 ;
  assign w3820 = w3818 ^ w3819 ;
  assign w3821 = w141 | w262 ;
  assign w3822 = ( w81 & ~w141 ) | ( w81 & w163 ) | ( ~w141 & w163 ) ;
  assign w3823 = w3821 | w3822 ;
  assign w3824 = w118 | w569 ;
  assign w3825 = ( ~w118 & w490 ) | ( ~w118 & w3823 ) | ( w490 & w3823 ) ;
  assign w3826 = w3824 | w3825 ;
  assign w3827 = ( w560 & w561 ) | ( w560 & ~w674 ) | ( w561 & ~w674 ) ;
  assign w3828 = ( ~w533 & w674 ) | ( ~w533 & w764 ) | ( w674 & w764 ) ;
  assign w3829 = w2721 | w3828 ;
  assign w3830 = w3827 | w3829 ;
  assign w3831 = ( ~w199 & w628 ) | ( ~w199 & w3830 ) | ( w628 & w3830 ) ;
  assign w3832 = w199 | w3831 ;
  assign w3833 = ( w119 & w208 ) | ( w119 & ~w505 ) | ( w208 & ~w505 ) ;
  assign w3834 = w90 | w910 ;
  assign w3835 = ( ~w90 & w505 ) | ( ~w90 & w641 ) | ( w505 & w641 ) ;
  assign w3836 = w3834 | w3835 ;
  assign w3837 = w3833 | w3836 ;
  assign w3838 = ( w218 & w318 ) | ( w218 & ~w390 ) | ( w318 & ~w390 ) ;
  assign w3839 = w3832 | w3837 ;
  assign w3840 = ( w390 & w637 ) | ( w390 & ~w3832 ) | ( w637 & ~w3832 ) ;
  assign w3841 = w3839 | w3840 ;
  assign w3842 = w3838 | w3841 ;
  assign w3843 = w2704 | w3826 ;
  assign w3844 = ( w731 & ~w3826 ) | ( w731 & w3842 ) | ( ~w3826 & w3842 ) ;
  assign w3845 = w3843 | w3844 ;
  assign w3846 = w817 | w1401 ;
  assign w3847 = w514 | w3846 ;
  assign w3848 = ( ~w514 & w1166 ) | ( ~w514 & w3845 ) | ( w1166 & w3845 ) ;
  assign w3849 = w3847 | w3848 ;
  assign w3850 = w419 | w511 ;
  assign w3851 = w116 | w3850 ;
  assign w3852 = ( ~w116 & w149 ) | ( ~w116 & w3849 ) | ( w149 & w3849 ) ;
  assign w3853 = w3851 | w3852 ;
  assign w3854 = w353 | w626 ;
  assign w3855 = w179 | w3854 ;
  assign w3856 = ( w131 & ~w179 ) | ( w131 & w221 ) | ( ~w179 & w221 ) ;
  assign w3857 = w3855 | w3856 ;
  assign w3858 = w470 | w568 ;
  assign w3859 = w325 | w3858 ;
  assign w3860 = ( ~w325 & w430 ) | ( ~w325 & w3857 ) | ( w430 & w3857 ) ;
  assign w3861 = w3859 | w3860 ;
  assign w3862 = ( w84 & w257 ) | ( w84 & ~w362 ) | ( w257 & ~w362 ) ;
  assign w3863 = w594 | w3196 ;
  assign w3864 = ( w362 & w525 ) | ( w362 & ~w594 ) | ( w525 & ~w594 ) ;
  assign w3865 = w3863 | w3864 ;
  assign w3866 = w3862 | w3865 ;
  assign w3867 = w415 | w1030 ;
  assign w3868 = ( ~w415 & w571 ) | ( ~w415 & w759 ) | ( w571 & w759 ) ;
  assign w3869 = w3867 | w3868 ;
  assign w3870 = ( w1128 & ~w1837 ) | ( w1128 & w3869 ) | ( ~w1837 & w3869 ) ;
  assign w3871 = w1837 | w3870 ;
  assign w3872 = ( ~w258 & w886 ) | ( ~w258 & w2631 ) | ( w886 & w2631 ) ;
  assign w3873 = w3866 | w3871 ;
  assign w3874 = ( w258 & w606 ) | ( w258 & ~w3871 ) | ( w606 & ~w3871 ) ;
  assign w3875 = w3873 | w3874 ;
  assign w3876 = w3872 | w3875 ;
  assign w3877 = ( w309 & w384 ) | ( w309 & ~w422 ) | ( w384 & ~w422 ) ;
  assign w3878 = w253 | w3876 ;
  assign w3879 = ( ~w253 & w422 ) | ( ~w253 & w899 ) | ( w422 & w899 ) ;
  assign w3880 = w3878 | w3879 ;
  assign w3881 = w3877 | w3880 ;
  assign w3882 = w567 | w951 ;
  assign w3883 = w101 | w3882 ;
  assign w3884 = ( ~w101 & w315 ) | ( ~w101 & w1618 ) | ( w315 & w1618 ) ;
  assign w3885 = w3883 | w3884 ;
  assign w3886 = ( w202 & w530 ) | ( w202 & ~w664 ) | ( w530 & ~w664 ) ;
  assign w3887 = w51 | w3885 ;
  assign w3888 = ( ~w51 & w664 ) | ( ~w51 & w1130 ) | ( w664 & w1130 ) ;
  assign w3889 = w3887 | w3888 ;
  assign w3890 = w3886 | w3889 ;
  assign w3891 = ( w113 & ~w165 ) | ( w113 & w463 ) | ( ~w165 & w463 ) ;
  assign w3892 = w165 | w3891 ;
  assign w3893 = w449 | w3892 ;
  assign w3894 = ( w268 & w3890 ) | ( w268 & ~w3892 ) | ( w3890 & ~w3892 ) ;
  assign w3895 = w3893 | w3894 ;
  assign w3896 = w956 | w2873 ;
  assign w3897 = w3895 | w3896 ;
  assign w3898 = ( w3861 & w3881 ) | ( w3861 & ~w3895 ) | ( w3881 & ~w3895 ) ;
  assign w3899 = w3897 | w3898 ;
  assign w3900 = ( w354 & ~w459 ) | ( w354 & w1814 ) | ( ~w459 & w1814 ) ;
  assign w3901 = w3853 | w3899 ;
  assign w3902 = ( w459 & w534 ) | ( w459 & ~w3899 ) | ( w534 & ~w3899 ) ;
  assign w3903 = w3901 | w3902 ;
  assign w3904 = w3900 | w3903 ;
  assign w3905 = w259 | w392 ;
  assign w3906 = ( ~w259 & w275 ) | ( ~w259 & w3904 ) | ( w275 & w3904 ) ;
  assign w3907 = w3905 | w3906 ;
  assign w3908 = w3548 | w3717 ;
  assign w3909 = w3649 & w3715 ;
  assign w3910 = ( ~w3548 & w3908 ) | ( ~w3548 & w3909 ) | ( w3908 & w3909 ) ;
  assign w3911 = ( ~w3548 & w3715 ) | ( ~w3548 & w3723 ) | ( w3715 & w3723 ) ;
  assign w3912 = w3548 ^ w3911 ;
  assign w3913 = w3907 ^ w3912 ;
  assign w3914 = ~w3549 & w3907 ;
  assign w3915 = ~w3910 & w3913 ;
  assign w3916 = ( w3448 & w3910 ) | ( w3448 & ~w3915 ) | ( w3910 & ~w3915 ) ;
  assign w3917 = ( w3907 & ~w3914 ) | ( w3907 & w3916 ) | ( ~w3914 & w3916 ) ;
  assign w3918 = \pi29 ^ w3917 ;
  assign w3919 = ~\pi25 & w137 ;
  assign w3920 = \pi26 ^ w3919 ;
  assign w3921 = \pi24 ^ \pi25 ;
  assign w3922 = ( \pi26 & w62 ) | ( \pi26 & ~w3921 ) | ( w62 & ~w3921 ) ;
  assign w3923 = ( w3919 & w3920 ) | ( w3919 & ~w3922 ) | ( w3920 & ~w3922 ) ;
  assign w3924 = \pi26 & w62 ;
  assign w3925 = ( w62 & ~w137 ) | ( w62 & w3924 ) | ( ~w137 & w3924 ) ;
  assign w3926 = ( w62 & w801 ) | ( w62 & w3925 ) | ( w801 & w3925 ) ;
  assign w3927 = ( \pi25 & w3925 ) | ( \pi25 & w3926 ) | ( w3925 & w3926 ) ;
  assign w3928 = w445 | w783 ;
  assign w3929 = w838 | w3928 ;
  assign w3930 = ( w468 & ~w838 ) | ( w468 & w1131 ) | ( ~w838 & w1131 ) ;
  assign w3931 = w3929 | w3930 ;
  assign w3932 = w229 | w664 ;
  assign w3933 = ( ~w229 & w595 ) | ( ~w229 & w3931 ) | ( w595 & w3931 ) ;
  assign w3934 = w3932 | w3933 ;
  assign w3935 = w259 | w1153 ;
  assign w3936 = ( ~w259 & w316 ) | ( ~w259 & w3934 ) | ( w316 & w3934 ) ;
  assign w3937 = w3935 | w3936 ;
  assign w3938 = w488 | w2294 ;
  assign w3939 = w2695 | w3938 ;
  assign w3940 = ( w86 & w96 ) | ( w86 & ~w2695 ) | ( w96 & ~w2695 ) ;
  assign w3941 = w3939 | w3940 ;
  assign w3942 = w51 | w571 ;
  assign w3943 = w3941 | w3942 ;
  assign w3944 = ( w2373 & w3937 ) | ( w2373 & ~w3941 ) | ( w3937 & ~w3941 ) ;
  assign w3945 = w3943 | w3944 ;
  assign w3946 = \pi26 | w102 ;
  assign w3947 = ( w99 & w102 ) | ( w99 & w3946 ) | ( w102 & w3946 ) ;
  assign w3948 = ( ~\pi25 & w43 ) | ( ~\pi25 & w3947 ) | ( w43 & w3947 ) ;
  assign w3949 = ( \pi25 & w102 ) | ( \pi25 & w3948 ) | ( w102 & w3948 ) ;
  assign w3950 = ( w43 & w102 ) | ( w43 & w3946 ) | ( w102 & w3946 ) ;
  assign w3951 = ( \pi24 & w102 ) | ( \pi24 & w3950 ) | ( w102 & w3950 ) ;
  assign w3952 = ( \pi25 & w3950 ) | ( \pi25 & w3951 ) | ( w3950 & w3951 ) ;
  assign w3953 = ( \pi23 & w3950 ) | ( \pi23 & w3952 ) | ( w3950 & w3952 ) ;
  assign w3954 = ( \pi24 & ~\pi25 ) | ( \pi24 & w43 ) | ( ~\pi25 & w43 ) ;
  assign w3955 = ( \pi23 & ~\pi26 ) | ( \pi23 & w3954 ) | ( ~\pi26 & w3954 ) ;
  assign w3956 = ( \pi23 & ~\pi24 ) | ( \pi23 & w3955 ) | ( ~\pi24 & w3955 ) ;
  assign w3957 = ~\pi23 & w3956 ;
  assign w3958 = ( w43 & w102 ) | ( w43 & ~w3957 ) | ( w102 & ~w3957 ) ;
  assign w3959 = w3945 | w3958 ;
  assign w3960 = ~w278 & w3927 ;
  assign w3961 = ( ~w278 & w312 ) | ( ~w278 & w3959 ) | ( w312 & w3959 ) ;
  assign w3962 = w3960 & ~w3961 ;
  assign w3963 = \pi25 ^ \pi26 ;
  assign w3964 = w2832 & ~w3963 ;
  assign w3965 = w95 | w259 ;
  assign w3966 = ( ~w144 & w2760 ) | ( ~w144 & w3115 ) | ( w2760 & w3115 ) ;
  assign w3967 = w1513 | w1881 ;
  assign w3968 = ( w144 & w568 ) | ( w144 & ~w1881 ) | ( w568 & ~w1881 ) ;
  assign w3969 = w3967 | w3968 ;
  assign w3970 = w3966 | w3969 ;
  assign w3971 = w787 | w860 ;
  assign w3972 = w3965 | w3971 ;
  assign w3973 = ( w164 & ~w3965 ) | ( w164 & w3970 ) | ( ~w3965 & w3970 ) ;
  assign w3974 = w3972 | w3973 ;
  assign w3975 = ( w142 & w325 ) | ( w142 & ~w491 ) | ( w325 & ~w491 ) ;
  assign w3976 = w133 | w3974 ;
  assign w3977 = ( ~w133 & w491 ) | ( ~w133 & w680 ) | ( w491 & w680 ) ;
  assign w3978 = w3976 | w3977 ;
  assign w3979 = w3975 | w3978 ;
  assign w3980 = ( ~w345 & w430 ) | ( ~w345 & w3979 ) | ( w430 & w3979 ) ;
  assign w3981 = w345 | w3980 ;
  assign w3982 = w505 | w897 ;
  assign w3983 = w362 | w3982 ;
  assign w3984 = ( w76 & ~w362 ) | ( w76 & w384 ) | ( ~w362 & w384 ) ;
  assign w3985 = w3983 | w3984 ;
  assign w3986 = ( \pi24 & \pi26 ) | ( \pi24 & w123 ) | ( \pi26 & w123 ) ;
  assign w3987 = w123 & ~w3986 ;
  assign w3988 = ( \pi25 & w2832 ) | ( \pi25 & w3987 ) | ( w2832 & w3987 ) ;
  assign w3989 = \pi26 ^ w2832 ;
  assign w3990 = ( \pi26 & w3988 ) | ( \pi26 & w3989 ) | ( w3988 & w3989 ) ;
  assign w3991 = w75 & w3990 ;
  assign w3992 = ( \pi25 & ~w2832 ) | ( \pi25 & w3987 ) | ( ~w2832 & w3987 ) ;
  assign w3993 = ( w3987 & w3991 ) | ( w3987 & ~w3992 ) | ( w3991 & ~w3992 ) ;
  assign w3994 = w421 | w3993 ;
  assign w3995 = ( w351 & ~w421 ) | ( w351 & w1094 ) | ( ~w421 & w1094 ) ;
  assign w3996 = w3994 | w3995 ;
  assign w3997 = ( ~w131 & w998 ) | ( ~w131 & w3996 ) | ( w998 & w3996 ) ;
  assign w3998 = w514 | w759 ;
  assign w3999 = ( w131 & w316 ) | ( w131 & ~w759 ) | ( w316 & ~w759 ) ;
  assign w4000 = w3998 | w3999 ;
  assign w4001 = w3997 | w4000 ;
  assign w4002 = ( ~w358 & w1783 ) | ( ~w358 & w3985 ) | ( w1783 & w3985 ) ;
  assign w4003 = w3981 | w4001 ;
  assign w4004 = ( w358 & w470 ) | ( w358 & ~w4001 ) | ( w470 & ~w4001 ) ;
  assign w4005 = w4003 | w4004 ;
  assign w4006 = w4002 | w4005 ;
  assign w4007 = ( w419 & w465 ) | ( w419 & ~w490 ) | ( w465 & ~w490 ) ;
  assign w4008 = w255 | w4006 ;
  assign w4009 = ( ~w255 & w490 ) | ( ~w255 & w623 ) | ( w490 & w623 ) ;
  assign w4010 = w4008 | w4009 ;
  assign w4011 = w4007 | w4010 ;
  assign w4012 = w571 | w901 ;
  assign w4013 = w277 | w4012 ;
  assign w4014 = ( ~w277 & w531 ) | ( ~w277 & w4011 ) | ( w531 & w4011 ) ;
  assign w4015 = w4013 | w4014 ;
  assign w4016 = ( w314 & w415 ) | ( w314 & ~w504 ) | ( w415 & ~w504 ) ;
  assign w4017 = w220 | w2872 ;
  assign w4018 = ( ~w220 & w504 ) | ( ~w220 & w524 ) | ( w504 & w524 ) ;
  assign w4019 = w4017 | w4018 ;
  assign w4020 = w4016 | w4019 ;
  assign w4021 = w569 | w802 ;
  assign w4022 = w111 | w4021 ;
  assign w4023 = ( ~w111 & w223 ) | ( ~w111 & w4020 ) | ( w223 & w4020 ) ;
  assign w4024 = w4022 | w4023 ;
  assign w4025 = ( ~w253 & w783 ) | ( ~w253 & w4024 ) | ( w783 & w4024 ) ;
  assign w4026 = w253 | w4025 ;
  assign w4027 = \pi25 | \pi26 ;
  assign w4028 = \pi24 | w4027 ;
  assign w4029 = w75 ^ w4028 ;
  assign w4030 = \pi23 & w80 ;
  assign w4031 = ( w80 & w4027 ) | ( w80 & w4030 ) | ( w4027 & w4030 ) ;
  assign w4032 = ( w75 & w4029 ) | ( w75 & w4031 ) | ( w4029 & w4031 ) ;
  assign w4033 = w443 | w1514 ;
  assign w4034 = ( w359 & ~w1181 ) | ( w359 & w1514 ) | ( ~w1181 & w1514 ) ;
  assign w4035 = ~w4033 & w4034 ;
  assign w4036 = ( ~w1069 & w2873 ) | ( ~w1069 & w4035 ) | ( w2873 & w4035 ) ;
  assign w4037 = w4015 | w4026 ;
  assign w4038 = ( w2873 & ~w4026 ) | ( w2873 & w4032 ) | ( ~w4026 & w4032 ) ;
  assign w4039 = w4037 | w4038 ;
  assign w4040 = w4036 & ~w4039 ;
  assign w4041 = w1031 | w2705 ;
  assign w4042 = w517 | w4041 ;
  assign w4043 = ( w517 & ~w731 ) | ( w517 & w4040 ) | ( ~w731 & w4040 ) ;
  assign w4044 = ~w4042 & w4043 ;
  assign w4045 = ( w322 & w447 ) | ( w322 & ~w533 ) | ( w447 & ~w533 ) ;
  assign w4046 = ~w265 & w4044 ;
  assign w4047 = ( ~w265 & w533 ) | ( ~w265 & w1001 ) | ( w533 & w1001 ) ;
  assign w4048 = w4046 & ~w4047 ;
  assign w4049 = ~w4045 & w4048 ;
  assign w4050 = ( \pi24 & ~\pi25 ) | ( \pi24 & \pi26 ) | ( ~\pi25 & \pi26 ) ;
  assign w4051 = ( \pi23 & \pi24 ) | ( \pi23 & w4050 ) | ( \pi24 & w4050 ) ;
  assign w4052 = w4050 ^ w4051 ;
  assign w4053 = \pi23 | \pi26 ;
  assign w4054 = ( \pi23 & \pi24 ) | ( \pi23 & ~w4053 ) | ( \pi24 & ~w4053 ) ;
  assign w4055 = ( \pi25 & \pi26 ) | ( \pi25 & ~w4054 ) | ( \pi26 & ~w4054 ) ;
  assign w4056 = \pi25 ^ w4055 ;
  assign w4057 = w137 & w4056 ;
  assign w4058 = ( w280 & w495 ) | ( w280 & ~w625 ) | ( w495 & ~w625 ) ;
  assign w4059 = w177 | w229 ;
  assign w4060 = ( ~w229 & w625 ) | ( ~w229 & w980 ) | ( w625 & w980 ) ;
  assign w4061 = w4059 | w4060 ;
  assign w4062 = w4058 | w4061 ;
  assign w4063 = w595 | w722 ;
  assign w4064 = w215 | w4063 ;
  assign w4065 = ( ~w215 & w445 ) | ( ~w215 & w4062 ) | ( w445 & w4062 ) ;
  assign w4066 = w4064 | w4065 ;
  assign w4067 = \pi23 & \pi26 ;
  assign w4068 = \pi25 & w4067 ;
  assign w4069 = ( \pi25 & w145 ) | ( \pi25 & ~w4067 ) | ( w145 & ~w4067 ) ;
  assign w4070 = w4067 ^ w4069 ;
  assign w4071 = ( w55 & w4069 ) | ( w55 & ~w4070 ) | ( w4069 & ~w4070 ) ;
  assign w4072 = ( ~\pi23 & w2833 ) | ( ~\pi23 & w4068 ) | ( w2833 & w4068 ) ;
  assign w4073 = ( w4068 & w4071 ) | ( w4068 & ~w4072 ) | ( w4071 & ~w4072 ) ;
  assign w4074 = w272 | w899 ;
  assign w4075 = ( w116 & ~w272 ) | ( w116 & w393 ) | ( ~w272 & w393 ) ;
  assign w4076 = w4074 | w4075 ;
  assign w4077 = w386 | w390 ;
  assign w4078 = w125 | w4077 ;
  assign w4079 = ( ~w125 & w353 ) | ( ~w125 & w4076 ) | ( w353 & w4076 ) ;
  assign w4080 = w4078 | w4079 ;
  assign w4081 = w83 & w93 ;
  assign w4082 = \pi26 & w4081 ;
  assign w4083 = ( ~\pi23 & \pi24 ) | ( ~\pi23 & \pi26 ) | ( \pi24 & \pi26 ) ;
  assign w4084 = ( \pi26 & w71 ) | ( \pi26 & ~w4083 ) | ( w71 & ~w4083 ) ;
  assign w4085 = \pi24 ^ w4083 ;
  assign w4086 = ( \pi23 & \pi26 ) | ( \pi23 & ~w4081 ) | ( \pi26 & ~w4081 ) ;
  assign w4087 = ( ~\pi23 & w4085 ) | ( ~\pi23 & w4086 ) | ( w4085 & w4086 ) ;
  assign w4088 = ( \pi23 & \pi26 ) | ( \pi23 & w93 ) | ( \pi26 & w93 ) ;
  assign w4089 = \pi25 ^ w4081 ;
  assign w4090 = w4088 ^ w4089 ;
  assign w4091 = ( w4084 & w4087 ) | ( w4084 & ~w4090 ) | ( w4087 & ~w4090 ) ;
  assign w4092 = ( w71 & w4082 ) | ( w71 & ~w4091 ) | ( w4082 & ~w4091 ) ;
  assign w4093 = ( w354 & w429 ) | ( w354 & ~w534 ) | ( w429 & ~w534 ) ;
  assign w4094 = w274 | w4080 ;
  assign w4095 = ( ~w274 & w534 ) | ( ~w274 & w4092 ) | ( w534 & w4092 ) ;
  assign w4096 = w4094 | w4095 ;
  assign w4097 = w4093 | w4096 ;
  assign w4098 = ( w265 & w359 ) | ( w265 & ~w4097 ) | ( w359 & ~w4097 ) ;
  assign w4099 = ~w265 & w4098 ;
  assign w4100 = w48 ^ w145 ;
  assign w4101 = ( w71 & w145 ) | ( w71 & w4100 ) | ( w145 & w4100 ) ;
  assign w4102 = w149 | w409 ;
  assign w4103 = ( w88 & ~w149 ) | ( w88 & w257 ) | ( ~w149 & w257 ) ;
  assign w4104 = w4102 | w4103 ;
  assign w4105 = w3493 | w4104 ;
  assign w4106 = ( w414 & ~w449 ) | ( w414 & w1837 ) | ( ~w449 & w1837 ) ;
  assign w4107 = w4099 & ~w4105 ;
  assign w4108 = ( w449 & w4101 ) | ( w449 & ~w4105 ) | ( w4101 & ~w4105 ) ;
  assign w4109 = w4107 & ~w4108 ;
  assign w4110 = ~w4106 & w4109 ;
  assign w4111 = w314 | w3996 ;
  assign w4112 = ( w220 & w2872 ) | ( w220 & ~w3996 ) | ( w2872 & ~w3996 ) ;
  assign w4113 = w4111 | w4112 ;
  assign w4114 = ( w90 & w169 ) | ( w90 & ~w860 ) | ( w169 & ~w860 ) ;
  assign w4115 = w624 | w4113 ;
  assign w4116 = ( ~w624 & w860 ) | ( ~w624 & w4032 ) | ( w860 & w4032 ) ;
  assign w4117 = w4115 | w4116 ;
  assign w4118 = w4114 | w4117 ;
  assign w4119 = ( w459 & w509 ) | ( w459 & ~w758 ) | ( w509 & ~w758 ) ;
  assign w4120 = w76 | w4118 ;
  assign w4121 = ( ~w76 & w758 ) | ( ~w76 & w1031 ) | ( w758 & w1031 ) ;
  assign w4122 = w4120 | w4121 ;
  assign w4123 = w4119 | w4122 ;
  assign w4124 = w120 | w515 ;
  assign w4125 = ( ~w120 & w164 ) | ( ~w120 & w4123 ) | ( w164 & w4123 ) ;
  assign w4126 = w4124 | w4125 ;
  assign w4127 = w837 | w4073 ;
  assign w4128 = w4126 | w4127 ;
  assign w4129 = ( ~w63 & w4110 ) | ( ~w63 & w4126 ) | ( w4110 & w4126 ) ;
  assign w4130 = ~w4128 & w4129 ;
  assign w4131 = w571 | w1001 ;
  assign w4132 = w3941 | w4131 ;
  assign w4133 = ( w609 & w3890 ) | ( w609 & ~w3941 ) | ( w3890 & ~w3941 ) ;
  assign w4134 = w4132 | w4133 ;
  assign w4135 = w98 | w129 ;
  assign w4136 = ( ~w129 & w1069 ) | ( ~w129 & w4134 ) | ( w1069 & w4134 ) ;
  assign w4137 = w4135 | w4136 ;
  assign w4138 = ( w468 & ~w593 ) | ( w468 & w4066 ) | ( ~w593 & w4066 ) ;
  assign w4139 = w4130 & ~w4137 ;
  assign w4140 = ( w593 & w4057 ) | ( w593 & ~w4137 ) | ( w4057 & ~w4137 ) ;
  assign w4141 = w4139 & ~w4140 ;
  assign w4142 = ~w4138 & w4141 ;
  assign w4143 = \pi25 ^ w57 ;
  assign w4144 = w4049 | w4052 ;
  assign w4145 = ~w4142 & w4143 ;
  assign w4146 = ( ~w4049 & w4144 ) | ( ~w4049 & w4145 ) | ( w4144 & w4145 ) ;
  assign w4147 = w2832 & w3963 ;
  assign w4148 = ( ~w3548 & w3907 ) | ( ~w3548 & w3911 ) | ( w3907 & w3911 ) ;
  assign w4149 = ( w3907 & ~w4049 ) | ( w3907 & w4148 ) | ( ~w4049 & w4148 ) ;
  assign w4150 = ( w4049 & w4142 ) | ( w4049 & ~w4149 ) | ( w4142 & ~w4149 ) ;
  assign w4151 = w3962 ^ w4150 ;
  assign w4152 = w4142 ^ w4151 ;
  assign w4153 = w4147 | w4152 ;
  assign w4154 = w3962 & ~w4146 ;
  assign w4155 = ( w3964 & w4146 ) | ( w3964 & ~w4154 ) | ( w4146 & ~w4154 ) ;
  assign w4156 = ( ~w4152 & w4153 ) | ( ~w4152 & w4155 ) | ( w4153 & w4155 ) ;
  assign w4157 = \pi26 ^ w4156 ;
  assign w4158 = w3820 ^ w4157 ;
  assign w4159 = w3918 ^ w4158 ;
  assign w4160 = w3647 & ~w3717 ;
  assign w4161 = ~w3094 & w3649 ;
  assign w4162 = ( w3647 & ~w4160 ) | ( w3647 & w4161 ) | ( ~w4160 & w4161 ) ;
  assign w4163 = w3647 ^ w3722 ;
  assign w4164 = w3715 ^ w4163 ;
  assign w4165 = ~w3549 & w3715 ;
  assign w4166 = ~w4162 & w4164 ;
  assign w4167 = ( w3448 & w4162 ) | ( w3448 & ~w4166 ) | ( w4162 & ~w4166 ) ;
  assign w4168 = ( w3715 & ~w4165 ) | ( w3715 & w4167 ) | ( ~w4165 & w4167 ) ;
  assign w4169 = \pi29 ^ w4168 ;
  assign w4170 = w3431 ^ w3444 ;
  assign w4171 = w3433 ^ w4170 ;
  assign w4172 = w3234 ^ w3430 ;
  assign w4173 = w3419 ^ w4172 ;
  assign w4174 = w385 | w596 ;
  assign w4175 = w341 | w1031 ;
  assign w4176 = ( w149 & ~w341 ) | ( w149 & w353 ) | ( ~w341 & w353 ) ;
  assign w4177 = w4175 | w4176 ;
  assign w4178 = ( w225 & w226 ) | ( w225 & ~w260 ) | ( w226 & ~w260 ) ;
  assign w4179 = w139 | w209 ;
  assign w4180 = ( ~w209 & w260 ) | ( ~w209 & w802 ) | ( w260 & w802 ) ;
  assign w4181 = w4179 | w4180 ;
  assign w4182 = w4178 | w4181 ;
  assign w4183 = w113 | w1126 ;
  assign w4184 = w4177 | w4183 ;
  assign w4185 = ( w3015 & ~w4177 ) | ( w3015 & w4182 ) | ( ~w4177 & w4182 ) ;
  assign w4186 = w4184 | w4185 ;
  assign w4187 = w890 | w4186 ;
  assign w4188 = w3981 | w4187 ;
  assign w4189 = ( ~w2304 & w3490 ) | ( ~w2304 & w3981 ) | ( w3490 & w3981 ) ;
  assign w4190 = ~w4188 & w4189 ;
  assign w4191 = w1208 | w4174 ;
  assign w4192 = w2618 | w4191 ;
  assign w4193 = ( ~w507 & w2618 ) | ( ~w507 & w4190 ) | ( w2618 & w4190 ) ;
  assign w4194 = ~w4192 & w4193 ;
  assign w4195 = w311 | w1130 ;
  assign w4196 = w268 | w4195 ;
  assign w4197 = ( w268 & ~w274 ) | ( w268 & w4194 ) | ( ~w274 & w4194 ) ;
  assign w4198 = ~w4196 & w4197 ;
  assign w4199 = w951 | w1001 ;
  assign w4200 = w136 | w4199 ;
  assign w4201 = ( ~w136 & w385 ) | ( ~w136 & w1095 ) | ( w385 & w1095 ) ;
  assign w4202 = w4200 | w4201 ;
  assign w4203 = ( ~w51 & w362 ) | ( ~w51 & w4202 ) | ( w362 & w4202 ) ;
  assign w4204 = w51 | w4203 ;
  assign w4205 = w565 | w1835 ;
  assign w4206 = ( w220 & w1165 ) | ( w220 & ~w1835 ) | ( w1165 & ~w1835 ) ;
  assign w4207 = w4205 | w4206 ;
  assign w4208 = w392 | w505 ;
  assign w4209 = ( w122 & ~w392 ) | ( w122 & w408 ) | ( ~w392 & w408 ) ;
  assign w4210 = w4208 | w4209 ;
  assign w4211 = ( w104 & ~w118 ) | ( w104 & w4210 ) | ( ~w118 & w4210 ) ;
  assign w4212 = w264 | w1741 ;
  assign w4213 = ( w118 & w409 ) | ( w118 & ~w1741 ) | ( w409 & ~w1741 ) ;
  assign w4214 = w4212 | w4213 ;
  assign w4215 = w4211 | w4214 ;
  assign w4216 = ( ~w488 & w1280 ) | ( ~w488 & w4215 ) | ( w1280 & w4215 ) ;
  assign w4217 = w4204 | w4207 ;
  assign w4218 = ( w488 & w490 ) | ( w488 & ~w4207 ) | ( w490 & ~w4207 ) ;
  assign w4219 = w4217 | w4218 ;
  assign w4220 = w4216 | w4219 ;
  assign w4221 = w317 | w1126 ;
  assign w4222 = w1166 | w4221 ;
  assign w4223 = ( w90 & ~w1166 ) | ( w90 & w4220 ) | ( ~w1166 & w4220 ) ;
  assign w4224 = w4222 | w4223 ;
  assign w4225 = ( w525 & w596 ) | ( w525 & ~w697 ) | ( w596 & ~w697 ) ;
  assign w4226 = w175 | w4224 ;
  assign w4227 = ( ~w175 & w697 ) | ( ~w175 & w1130 ) | ( w697 & w1130 ) ;
  assign w4228 = w4226 | w4227 ;
  assign w4229 = w4225 | w4228 ;
  assign w4230 = w161 | w1229 ;
  assign w4231 = ( w139 & ~w161 ) | ( w139 & w901 ) | ( ~w161 & w901 ) ;
  assign w4232 = w4230 | w4231 ;
  assign w4233 = w260 | w593 ;
  assign w4234 = ( w259 & ~w260 ) | ( w259 & w384 ) | ( ~w260 & w384 ) ;
  assign w4235 = w4233 | w4234 ;
  assign w4236 = ( w2480 & w3493 ) | ( w2480 & ~w4232 ) | ( w3493 & ~w4232 ) ;
  assign w4237 = w3628 | w4229 ;
  assign w4238 = ( ~w4229 & w4232 ) | ( ~w4229 & w4235 ) | ( w4232 & w4235 ) ;
  assign w4239 = w4237 | w4238 ;
  assign w4240 = w4236 | w4239 ;
  assign w4241 = w784 | w1064 ;
  assign w4242 = w212 | w4241 ;
  assign w4243 = ( ~w212 & w450 ) | ( ~w212 & w4240 ) | ( w450 & w4240 ) ;
  assign w4244 = w4242 | w4243 ;
  assign w4245 = ( w341 & w388 ) | ( w341 & ~w393 ) | ( w388 & ~w393 ) ;
  assign w4246 = w311 | w4244 ;
  assign w4247 = ( ~w311 & w393 ) | ( ~w311 & w1128 ) | ( w393 & w1128 ) ;
  assign w4248 = w4246 | w4247 ;
  assign w4249 = w4245 | w4248 ;
  assign w4250 = ( w176 & w310 ) | ( w176 & ~w431 ) | ( w310 & ~w431 ) ;
  assign w4251 = w115 | w4249 ;
  assign w4252 = ( ~w115 & w431 ) | ( ~w115 & w495 ) | ( w431 & w495 ) ;
  assign w4253 = w4251 | w4252 ;
  assign w4254 = w4250 | w4253 ;
  assign w4255 = ( \pi17 & w4198 ) | ( \pi17 & ~w4254 ) | ( w4198 & ~w4254 ) ;
  assign w4256 = w883 ^ w2996 ;
  assign w4257 = w721 ^ w4256 ;
  assign w4258 = ( \pi30 & \pi31 ) | ( \pi30 & ~w883 ) | ( \pi31 & ~w883 ) ;
  assign w4259 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w4258 ) | ( \pi30 & w4258 ) ;
  assign w4260 = ( \pi29 & ~\pi30 ) | ( \pi29 & w4258 ) | ( ~\pi30 & w4258 ) ;
  assign w4261 = ( ~\pi30 & w979 ) | ( ~\pi30 & w4260 ) | ( w979 & w4260 ) ;
  assign w4262 = ( w721 & w4260 ) | ( w721 & ~w4261 ) | ( w4260 & ~w4261 ) ;
  assign w4263 = ~\pi31 & w4262 ;
  assign w4264 = ( w4259 & w4261 ) | ( w4259 & w4263 ) | ( w4261 & w4263 ) ;
  assign w4265 = ( w37 & ~w4257 ) | ( w37 & w4264 ) | ( ~w4257 & w4264 ) ;
  assign w4266 = w4264 | w4265 ;
  assign w4267 = ( w3234 & w4255 ) | ( w3234 & ~w4266 ) | ( w4255 & ~w4266 ) ;
  assign w4268 = w4255 ^ w4266 ;
  assign w4269 = w3234 ^ w4268 ;
  assign w4270 = w4198 ^ w4254 ;
  assign w4271 = \pi17 ^ w4270 ;
  assign w4272 = w883 ^ w2995 ;
  assign w4273 = w979 ^ w4272 ;
  assign w4274 = w37 | w4273 ;
  assign w4275 = w1085 & w3098 ;
  assign w4276 = ( ~w4273 & w4274 ) | ( ~w4273 & w4275 ) | ( w4274 & w4275 ) ;
  assign w4277 = ( \pi29 & \pi30 ) | ( \pi29 & ~w883 ) | ( \pi30 & ~w883 ) ;
  assign w4278 = \pi31 | w4277 ;
  assign w4279 = ( \pi29 & ~\pi30 ) | ( \pi29 & w979 ) | ( ~\pi30 & w979 ) ;
  assign w4280 = ( \pi29 & \pi31 ) | ( \pi29 & ~w4279 ) | ( \pi31 & ~w4279 ) ;
  assign w4281 = ( w4276 & w4278 ) | ( w4276 & ~w4280 ) | ( w4278 & ~w4280 ) ;
  assign w4282 = ( w209 & w465 ) | ( w209 & ~w723 ) | ( w465 & ~w723 ) ;
  assign w4283 = w208 | w264 ;
  assign w4284 = ( ~w208 & w723 ) | ( ~w208 & w980 ) | ( w723 & w980 ) ;
  assign w4285 = w4283 | w4284 ;
  assign w4286 = w4282 | w4285 ;
  assign w4287 = ( w59 & ~w350 ) | ( w59 & w2168 ) | ( ~w350 & w2168 ) ;
  assign w4288 = w997 | w4286 ;
  assign w4289 = ( w350 & w443 ) | ( w350 & ~w997 ) | ( w443 & ~w997 ) ;
  assign w4290 = w4288 | w4289 ;
  assign w4291 = w4287 | w4290 ;
  assign w4292 = ( w214 & ~w889 ) | ( w214 & w1153 ) | ( ~w889 & w1153 ) ;
  assign w4293 = w889 | w4292 ;
  assign w4294 = ( w386 & w424 ) | ( w386 & ~w531 ) | ( w424 & ~w531 ) ;
  assign w4295 = w178 | w4293 ;
  assign w4296 = ( ~w178 & w531 ) | ( ~w178 & w802 ) | ( w531 & w802 ) ;
  assign w4297 = w4295 | w4296 ;
  assign w4298 = w4294 | w4297 ;
  assign w4299 = ( ~w495 & w2213 ) | ( ~w495 & w4298 ) | ( w2213 & w4298 ) ;
  assign w4300 = w2286 | w2400 ;
  assign w4301 = ( w495 & w513 ) | ( w495 & ~w2400 ) | ( w513 & ~w2400 ) ;
  assign w4302 = w4300 | w4301 ;
  assign w4303 = w4299 | w4302 ;
  assign w4304 = w204 | w2565 ;
  assign w4305 = ( ~w204 & w900 ) | ( ~w204 & w4303 ) | ( w900 & w4303 ) ;
  assign w4306 = w4304 | w4305 ;
  assign w4307 = ( w163 & w674 ) | ( w163 & ~w722 ) | ( w674 & ~w722 ) ;
  assign w4308 = w104 | w4306 ;
  assign w4309 = ( ~w104 & w722 ) | ( ~w104 & w1128 ) | ( w722 & w1128 ) ;
  assign w4310 = w4308 | w4309 ;
  assign w4311 = w4307 | w4310 ;
  assign w4312 = w496 | w897 ;
  assign w4313 = ( w352 & ~w496 ) | ( w352 & w697 ) | ( ~w496 & w697 ) ;
  assign w4314 = w4312 | w4313 ;
  assign w4315 = ( ~w268 & w431 ) | ( ~w268 & w4314 ) | ( w431 & w4314 ) ;
  assign w4316 = w268 | w4315 ;
  assign w4317 = ( w126 & ~w320 ) | ( w126 & w2873 ) | ( ~w320 & w2873 ) ;
  assign w4318 = w2087 | w4316 ;
  assign w4319 = ( w320 & w787 ) | ( w320 & ~w4316 ) | ( w787 & ~w4316 ) ;
  assign w4320 = w4318 | w4319 ;
  assign w4321 = w4317 | w4320 ;
  assign w4322 = w210 | w340 ;
  assign w4323 = w81 | w4322 ;
  assign w4324 = ( ~w81 & w90 ) | ( ~w81 & w4321 ) | ( w90 & w4321 ) ;
  assign w4325 = w4323 | w4324 ;
  assign w4326 = w419 | w641 ;
  assign w4327 = w63 | w4326 ;
  assign w4328 = ( ~w63 & w287 ) | ( ~w63 & w4325 ) | ( w287 & w4325 ) ;
  assign w4329 = w4327 | w4328 ;
  assign w4330 = ( w74 & w280 ) | ( w74 & ~w345 ) | ( w280 & ~w345 ) ;
  assign w4331 = w536 | w2434 ;
  assign w4332 = ( w345 & ~w536 ) | ( w345 & w567 ) | ( ~w536 & w567 ) ;
  assign w4333 = w4331 | w4332 ;
  assign w4334 = w4330 | w4333 ;
  assign w4335 = ( ~w2625 & w4291 ) | ( ~w2625 & w4334 ) | ( w4291 & w4334 ) ;
  assign w4336 = w4311 | w4329 ;
  assign w4337 = ( w2625 & w2762 ) | ( w2625 & ~w4329 ) | ( w2762 & ~w4329 ) ;
  assign w4338 = w4336 | w4337 ;
  assign w4339 = w4335 | w4338 ;
  assign w4340 = w421 | w458 ;
  assign w4341 = w2812 | w4340 ;
  assign w4342 = ( w1835 & ~w2812 ) | ( w1835 & w4339 ) | ( ~w2812 & w4339 ) ;
  assign w4343 = w4341 | w4342 ;
  assign w4344 = ( w285 & w310 ) | ( w285 & ~w385 ) | ( w310 & ~w385 ) ;
  assign w4345 = w205 | w4343 ;
  assign w4346 = ( ~w205 & w385 ) | ( ~w205 & w724 ) | ( w385 & w724 ) ;
  assign w4347 = w4345 | w4346 ;
  assign w4348 = w4344 | w4347 ;
  assign w4349 = w673 | w901 ;
  assign w4350 = ( ~w673 & w783 ) | ( ~w673 & w4348 ) | ( w783 & w4348 ) ;
  assign w4351 = w4349 | w4350 ;
  assign w4352 = w119 | w125 ;
  assign w4353 = w392 | w764 ;
  assign w4354 = w225 | w4353 ;
  assign w4355 = ( ~w225 & w226 ) | ( ~w225 & w4352 ) | ( w226 & w4352 ) ;
  assign w4356 = w4354 | w4355 ;
  assign w4357 = ( ~w422 & w424 ) | ( ~w422 & w4356 ) | ( w424 & w4356 ) ;
  assign w4358 = w422 | w4357 ;
  assign w4359 = ( w393 & w411 ) | ( w393 & ~w418 ) | ( w411 & ~w418 ) ;
  assign w4360 = w142 | w258 ;
  assign w4361 = ( ~w258 & w418 ) | ( ~w258 & w897 ) | ( w418 & w897 ) ;
  assign w4362 = w4360 | w4361 ;
  assign w4363 = w4359 | w4362 ;
  assign w4364 = w98 | w1130 ;
  assign w4365 = ( ~w98 & w281 ) | ( ~w98 & w2814 ) | ( w281 & w2814 ) ;
  assign w4366 = w4364 | w4365 ;
  assign w4367 = ( w784 & ~w1979 ) | ( w784 & w4366 ) | ( ~w1979 & w4366 ) ;
  assign w4368 = w4291 | w4358 ;
  assign w4369 = ( w1979 & ~w4358 ) | ( w1979 & w4363 ) | ( ~w4358 & w4363 ) ;
  assign w4370 = w4368 | w4369 ;
  assign w4371 = w4367 | w4370 ;
  assign w4372 = ( w68 & w115 ) | ( w68 & ~w260 ) | ( w115 & ~w260 ) ;
  assign w4373 = w1265 | w4371 ;
  assign w4374 = ( w260 & w286 ) | ( w260 & ~w1265 ) | ( w286 & ~w1265 ) ;
  assign w4375 = w4373 | w4374 ;
  assign w4376 = w4372 | w4375 ;
  assign w4377 = w175 | w951 ;
  assign w4378 = ( ~w175 & w358 ) | ( ~w175 & w4376 ) | ( w358 & w4376 ) ;
  assign w4379 = w4377 | w4378 ;
  assign w4380 = ( w322 & ~w324 ) | ( w322 & w361 ) | ( ~w324 & w361 ) ;
  assign w4381 = w324 | w4380 ;
  assign w4382 = w127 | w467 ;
  assign w4383 = ( w63 & ~w127 ) | ( w63 & w314 ) | ( ~w127 & w314 ) ;
  assign w4384 = w4382 | w4383 ;
  assign w4385 = ( w133 & ~w180 ) | ( w133 & w4293 ) | ( ~w180 & w4293 ) ;
  assign w4386 = w1069 | w2762 ;
  assign w4387 = ( w180 & w345 ) | ( w180 & ~w2762 ) | ( w345 & ~w2762 ) ;
  assign w4388 = w4386 | w4387 ;
  assign w4389 = w4385 | w4388 ;
  assign w4390 = ( w3555 & w4384 ) | ( w3555 & ~w4389 ) | ( w4384 & ~w4389 ) ;
  assign w4391 = w4389 | w4390 ;
  assign w4392 = w90 | w561 ;
  assign w4393 = w2872 | w4392 ;
  assign w4394 = ( ~w2872 & w4381 ) | ( ~w2872 & w4391 ) | ( w4381 & w4391 ) ;
  assign w4395 = w4393 | w4394 ;
  assign w4396 = ( w255 & w504 ) | ( w255 & ~w525 ) | ( w504 & ~w525 ) ;
  assign w4397 = w118 | w4395 ;
  assign w4398 = ( ~w118 & w525 ) | ( ~w118 & w568 ) | ( w525 & w568 ) ;
  assign w4399 = w4397 | w4398 ;
  assign w4400 = w4396 | w4399 ;
  assign w4401 = ( w116 & w265 ) | ( w116 & ~w277 ) | ( w265 & ~w277 ) ;
  assign w4402 = w103 | w1646 ;
  assign w4403 = ( ~w103 & w277 ) | ( ~w103 & w447 ) | ( w277 & w447 ) ;
  assign w4404 = w4402 | w4403 ;
  assign w4405 = w4401 | w4404 ;
  assign w4406 = ( w124 & w386 ) | ( w124 & ~w596 ) | ( w386 & ~w596 ) ;
  assign w4407 = w88 | w4405 ;
  assign w4408 = ( ~w88 & w596 ) | ( ~w88 & w625 ) | ( w596 & w625 ) ;
  assign w4409 = w4407 | w4408 ;
  assign w4410 = w4406 | w4409 ;
  assign w4411 = ( w310 & w419 ) | ( w310 & ~w787 ) | ( w419 & ~w787 ) ;
  assign w4412 = w280 | w4410 ;
  assign w4413 = ( ~w280 & w787 ) | ( ~w280 & w802 ) | ( w787 & w802 ) ;
  assign w4414 = w4412 | w4413 ;
  assign w4415 = w4411 | w4414 ;
  assign w4416 = w256 | w637 ;
  assign w4417 = ( ~w256 & w420 ) | ( ~w256 & w2480 ) | ( w420 & w2480 ) ;
  assign w4418 = w4416 | w4417 ;
  assign w4419 = w663 | w664 ;
  assign w4420 = w2147 | w4419 ;
  assign w4421 = ( w511 & ~w2147 ) | ( w511 & w4418 ) | ( ~w2147 & w4418 ) ;
  assign w4422 = w4420 | w4421 ;
  assign w4423 = w257 | w725 ;
  assign w4424 = w147 | w4423 ;
  assign w4425 = ( ~w147 & w210 ) | ( ~w147 & w2452 ) | ( w210 & w2452 ) ;
  assign w4426 = w4424 | w4425 ;
  assign w4427 = ( w167 & ~w325 ) | ( w167 & w2873 ) | ( ~w325 & w2873 ) ;
  assign w4428 = w4422 | w4426 ;
  assign w4429 = ( w325 & w509 ) | ( w325 & ~w4426 ) | ( w509 & ~w4426 ) ;
  assign w4430 = w4428 | w4429 ;
  assign w4431 = w4427 | w4430 ;
  assign w4432 = w2252 | w4415 ;
  assign w4433 = ( w4400 & ~w4415 ) | ( w4400 & w4431 ) | ( ~w4415 & w4431 ) ;
  assign w4434 = w4432 | w4433 ;
  assign w4435 = ( w84 & ~w488 ) | ( w84 & w1207 ) | ( ~w488 & w1207 ) ;
  assign w4436 = w4379 | w4434 ;
  assign w4437 = ( w488 & w490 ) | ( w488 & ~w4434 ) | ( w490 & ~w4434 ) ;
  assign w4438 = w4436 | w4437 ;
  assign w4439 = w4435 | w4438 ;
  assign w4440 = ( w161 & w259 ) | ( w161 & ~w680 ) | ( w259 & ~w680 ) ;
  assign w4441 = w51 | w4439 ;
  assign w4442 = ( ~w51 & w680 ) | ( ~w51 & w697 ) | ( w680 & w697 ) ;
  assign w4443 = w4441 | w4442 ;
  assign w4444 = w4440 | w4443 ;
  assign w4445 = ( w422 & w458 ) | ( w422 & ~w492 ) | ( w458 & ~w492 ) ;
  assign w4446 = w51 | w271 ;
  assign w4447 = ( ~w271 & w492 ) | ( ~w271 & w1274 ) | ( w492 & w1274 ) ;
  assign w4448 = w4446 | w4447 ;
  assign w4449 = w4445 | w4448 ;
  assign w4450 = ( ~w350 & w565 ) | ( ~w350 & w4449 ) | ( w565 & w4449 ) ;
  assign w4451 = w350 | w4450 ;
  assign w4452 = ( w229 & w315 ) | ( w229 & ~w681 ) | ( w315 & ~w681 ) ;
  assign w4453 = w138 | w1161 ;
  assign w4454 = ( ~w138 & w681 ) | ( ~w138 & w1340 ) | ( w681 & w1340 ) ;
  assign w4455 = w4453 | w4454 ;
  assign w4456 = w4452 | w4455 ;
  assign w4457 = w209 | w232 ;
  assign w4458 = w1064 | w4457 ;
  assign w4459 = ( w178 & ~w1064 ) | ( w178 & w4456 ) | ( ~w1064 & w4456 ) ;
  assign w4460 = w4458 | w4459 ;
  assign w4461 = w218 | w821 ;
  assign w4462 = ( w218 & w359 ) | ( w218 & ~w4460 ) | ( w359 & ~w4460 ) ;
  assign w4463 = ~w4461 & w4462 ;
  assign w4464 = w68 | w275 ;
  assign w4465 = w512 | w4235 ;
  assign w4466 = ( w283 & w2295 ) | ( w283 & ~w4235 ) | ( w2295 & ~w4235 ) ;
  assign w4467 = w4465 | w4466 ;
  assign w4468 = w325 | w1031 ;
  assign w4469 = w101 | w4468 ;
  assign w4470 = ( ~w101 & w309 ) | ( ~w101 & w4467 ) | ( w309 & w4467 ) ;
  assign w4471 = w4469 | w4470 ;
  assign w4472 = w164 | w429 ;
  assign w4473 = w4464 | w4472 ;
  assign w4474 = ( w141 & ~w4464 ) | ( w141 & w4471 ) | ( ~w4464 & w4471 ) ;
  assign w4475 = w4473 | w4474 ;
  assign w4476 = w124 | w513 ;
  assign w4477 = w432 | w4476 ;
  assign w4478 = ( ~w432 & w4314 ) | ( ~w432 & w4475 ) | ( w4314 & w4475 ) ;
  assign w4479 = w4477 | w4478 ;
  assign w4480 = ( w115 & ~w413 ) | ( w115 & w1590 ) | ( ~w413 & w1590 ) ;
  assign w4481 = w3460 | w4479 ;
  assign w4482 = ( w413 & w421 ) | ( w413 & ~w3460 ) | ( w421 & ~w3460 ) ;
  assign w4483 = w4481 | w4482 ;
  assign w4484 = w4480 | w4483 ;
  assign w4485 = ( w226 & w253 ) | ( w226 & ~w278 ) | ( w253 & ~w278 ) ;
  assign w4486 = w176 | w4484 ;
  assign w4487 = ( ~w176 & w278 ) | ( ~w176 & w1001 ) | ( w278 & w1001 ) ;
  assign w4488 = w4486 | w4487 ;
  assign w4489 = w4485 | w4488 ;
  assign w4490 = ( w120 & w131 ) | ( w120 & ~w223 ) | ( w131 & ~w223 ) ;
  assign w4491 = w2395 | w3385 ;
  assign w4492 = ( w223 & w311 ) | ( w223 & ~w2395 ) | ( w311 & ~w2395 ) ;
  assign w4493 = w4491 | w4492 ;
  assign w4494 = w4490 | w4493 ;
  assign w4495 = w998 | w1363 ;
  assign w4496 = w594 | w4495 ;
  assign w4497 = ( ~w594 & w838 ) | ( ~w594 & w4494 ) | ( w838 & w4494 ) ;
  assign w4498 = w4496 | w4497 ;
  assign w4499 = ( w342 & w511 ) | ( w342 & ~w596 ) | ( w511 & ~w596 ) ;
  assign w4500 = w122 | w4498 ;
  assign w4501 = ( ~w122 & w596 ) | ( ~w122 & w674 ) | ( w596 & w674 ) ;
  assign w4502 = w4500 | w4501 ;
  assign w4503 = w4499 | w4502 ;
  assign w4504 = ( w322 & w605 ) | ( w322 & ~w608 ) | ( w605 & ~w608 ) ;
  assign w4505 = w74 | w4503 ;
  assign w4506 = ( ~w74 & w608 ) | ( ~w74 & w640 ) | ( w608 & w640 ) ;
  assign w4507 = w4505 | w4506 ;
  assign w4508 = w4504 | w4507 ;
  assign w4509 = ( w84 & w136 ) | ( w84 & ~w219 ) | ( w136 & ~w219 ) ;
  assign w4510 = w82 | w514 ;
  assign w4511 = ( w219 & w341 ) | ( w219 & ~w514 ) | ( w341 & ~w514 ) ;
  assign w4512 = w4510 | w4511 ;
  assign w4513 = w4509 | w4512 ;
  assign w4514 = ( w133 & w623 ) | ( w133 & ~w837 ) | ( w623 & ~w837 ) ;
  assign w4515 = w118 | w4513 ;
  assign w4516 = ( ~w118 & w837 ) | ( ~w118 & w1229 ) | ( w837 & w1229 ) ;
  assign w4517 = w4515 | w4516 ;
  assign w4518 = w4514 | w4517 ;
  assign w4519 = w4451 | w4518 ;
  assign w4520 = w4508 | w4519 ;
  assign w4521 = ( w4463 & ~w4489 ) | ( w4463 & w4508 ) | ( ~w4489 & w4508 ) ;
  assign w4522 = ~w4520 & w4521 ;
  assign w4523 = w267 | w3178 ;
  assign w4524 = ( w267 & ~w785 ) | ( w267 & w4522 ) | ( ~w785 & w4522 ) ;
  assign w4525 = ~w4523 & w4524 ;
  assign w4526 = ( w318 & w388 ) | ( w318 & ~w488 ) | ( w388 & ~w488 ) ;
  assign w4527 = ~w214 & w4525 ;
  assign w4528 = ( ~w214 & w488 ) | ( ~w214 & w567 ) | ( w488 & w567 ) ;
  assign w4529 = w4527 & ~w4528 ;
  assign w4530 = ~w4526 & w4529 ;
  assign w4531 = ( \pi14 & ~w4444 ) | ( \pi14 & w4530 ) | ( ~w4444 & w4530 ) ;
  assign w4532 = w1085 ^ w2993 ;
  assign w4533 = w1205 ^ w4532 ;
  assign w4534 = ( \pi29 & \pi31 ) | ( \pi29 & w1205 ) | ( \pi31 & w1205 ) ;
  assign w4535 = ( \pi29 & ~\pi30 ) | ( \pi29 & w4534 ) | ( ~\pi30 & w4534 ) ;
  assign w4536 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w4534 ) | ( \pi30 & w4534 ) ;
  assign w4537 = ( \pi29 & w1264 ) | ( \pi29 & ~w4536 ) | ( w1264 & ~w4536 ) ;
  assign w4538 = ( w1085 & w4536 ) | ( w1085 & w4537 ) | ( w4536 & w4537 ) ;
  assign w4539 = ~\pi31 & w4538 ;
  assign w4540 = ( w4535 & ~w4537 ) | ( w4535 & w4539 ) | ( ~w4537 & w4539 ) ;
  assign w4541 = ( w37 & w4533 ) | ( w37 & w4540 ) | ( w4533 & w4540 ) ;
  assign w4542 = w4540 | w4541 ;
  assign w4543 = ( w4351 & w4531 ) | ( w4351 & ~w4542 ) | ( w4531 & ~w4542 ) ;
  assign w4544 = ( w4198 & w4351 ) | ( w4198 & ~w4543 ) | ( w4351 & ~w4543 ) ;
  assign w4545 = ( w4271 & w4281 ) | ( w4271 & w4544 ) | ( w4281 & w4544 ) ;
  assign w4546 = w381 | w3717 ;
  assign w4547 = w592 & w3649 ;
  assign w4548 = ( ~w381 & w4546 ) | ( ~w381 & w4547 ) | ( w4546 & w4547 ) ;
  assign w4549 = w3094 | w3549 ;
  assign w4550 = w3096 | w4548 ;
  assign w4551 = ( w3448 & w4548 ) | ( w3448 & w4550 ) | ( w4548 & w4550 ) ;
  assign w4552 = ( ~w3094 & w4549 ) | ( ~w3094 & w4551 ) | ( w4549 & w4551 ) ;
  assign w4553 = \pi29 ^ w4552 ;
  assign w4554 = ( w4269 & w4545 ) | ( w4269 & w4553 ) | ( w4545 & w4553 ) ;
  assign w4555 = ( w4173 & ~w4267 ) | ( w4173 & w4554 ) | ( ~w4267 & w4554 ) ;
  assign w4556 = ( w4169 & w4171 ) | ( w4169 & w4555 ) | ( w4171 & w4555 ) ;
  assign w4557 = w3339 ^ w3730 ;
  assign w4558 = w3445 ^ w4557 ;
  assign w4559 = w4049 | w4143 ;
  assign w4560 = w3907 & w4052 ;
  assign w4561 = ( ~w4049 & w4559 ) | ( ~w4049 & w4560 ) | ( w4559 & w4560 ) ;
  assign w4562 = w4049 ^ w4149 ;
  assign w4563 = w4142 ^ w4562 ;
  assign w4564 = ~w4147 & w4563 ;
  assign w4565 = w4142 & ~w4561 ;
  assign w4566 = ( w3964 & w4561 ) | ( w3964 & ~w4565 ) | ( w4561 & ~w4565 ) ;
  assign w4567 = ( w4563 & ~w4564 ) | ( w4563 & w4566 ) | ( ~w4564 & w4566 ) ;
  assign w4568 = \pi26 ^ w4567 ;
  assign w4569 = ( w4556 & ~w4558 ) | ( w4556 & w4568 ) | ( ~w4558 & w4568 ) ;
  assign w4570 = ( \pi23 & \pi25 ) | ( \pi23 & w2832 ) | ( \pi25 & w2832 ) ;
  assign w4571 = \pi26 ^ w4570 ;
  assign w4572 = w112 & w4571 ;
  assign w4573 = ( \pi26 & w65 ) | ( \pi26 & w4572 ) | ( w65 & w4572 ) ;
  assign w4574 = ~\pi23 & w97 ;
  assign w4575 = \pi26 | w4574 ;
  assign w4576 = ( \pi24 & ~\pi25 ) | ( \pi24 & w97 ) | ( ~\pi25 & w97 ) ;
  assign w4577 = ( \pi23 & w137 ) | ( \pi23 & w4576 ) | ( w137 & w4576 ) ;
  assign w4578 = w4576 | w4577 ;
  assign w4579 = ( \pi25 & ~\pi26 ) | ( \pi25 & w4578 ) | ( ~\pi26 & w4578 ) ;
  assign w4580 = w4575 & w4579 ;
  assign w4581 = w384 | w4580 ;
  assign w4582 = w144 | w4581 ;
  assign w4583 = ( w113 & ~w144 ) | ( w113 & w287 ) | ( ~w144 & w287 ) ;
  assign w4584 = w4582 | w4583 ;
  assign w4585 = ( ~w127 & w362 ) | ( ~w127 & w4584 ) | ( w362 & w4584 ) ;
  assign w4586 = w127 | w4585 ;
  assign w4587 = ( w98 & ~w101 ) | ( w98 & w2452 ) | ( ~w101 & w2452 ) ;
  assign w4588 = w1069 | w4586 ;
  assign w4589 = ( w101 & ~w1069 ) | ( w101 & w4573 ) | ( ~w1069 & w4573 ) ;
  assign w4590 = w4588 | w4589 ;
  assign w4591 = w4587 | w4590 ;
  assign w4592 = ( w256 & ~w465 ) | ( w256 & w1814 ) | ( ~w465 & w1814 ) ;
  assign w4593 = w1401 | w4591 ;
  assign w4594 = ( w465 & w593 ) | ( w465 & ~w1401 ) | ( w593 & ~w1401 ) ;
  assign w4595 = w4593 | w4594 ;
  assign w4596 = w4592 | w4595 ;
  assign w4597 = w278 | w4057 ;
  assign w4598 = ( ~w278 & w605 ) | ( ~w278 & w4596 ) | ( w605 & w4596 ) ;
  assign w4599 = w4597 | w4598 ;
  assign w4600 = w3927 & ~w4599 ;
  assign w4601 = ( w3962 & w4142 ) | ( w3962 & w4150 ) | ( w4142 & w4150 ) ;
  assign w4602 = ( w3962 & w4600 ) | ( w3962 & w4601 ) | ( w4600 & w4601 ) ;
  assign w4603 = w4600 | w4602 ;
  assign w4604 = ( \pi21 & ~\pi22 ) | ( \pi21 & \pi23 ) | ( ~\pi22 & \pi23 ) ;
  assign w4605 = ( \pi20 & \pi21 ) | ( \pi20 & w4604 ) | ( \pi21 & w4604 ) ;
  assign w4606 = w4604 ^ w4605 ;
  assign w4607 = \pi22 ^ \pi23 ;
  assign w4608 = \pi20 ^ \pi21 ;
  assign w4609 = w4607 & w4608 ;
  assign w4610 = ~w4600 & w4606 ;
  assign w4611 = w4609 | w4610 ;
  assign w4612 = ( ~w4603 & w4610 ) | ( ~w4603 & w4611 ) | ( w4610 & w4611 ) ;
  assign w4613 = \pi23 ^ w4612 ;
  assign w4614 = w4159 ^ w4613 ;
  assign w4615 = w4569 ^ w4614 ;
  assign w4616 = w4169 ^ w4555 ;
  assign w4617 = w4171 ^ w4616 ;
  assign w4618 = w3548 | w4052 ;
  assign w4619 = w3907 & w4143 ;
  assign w4620 = ( ~w3548 & w4618 ) | ( ~w3548 & w4619 ) | ( w4618 & w4619 ) ;
  assign w4621 = w4049 ^ w4148 ;
  assign w4622 = w3907 ^ w4621 ;
  assign w4623 = w4147 | w4622 ;
  assign w4624 = w4049 & ~w4620 ;
  assign w4625 = ( w3964 & w4620 ) | ( w3964 & ~w4624 ) | ( w4620 & ~w4624 ) ;
  assign w4626 = ( ~w4622 & w4623 ) | ( ~w4622 & w4625 ) | ( w4623 & w4625 ) ;
  assign w4627 = \pi26 ^ w4626 ;
  assign w4628 = w3548 | w4143 ;
  assign w4629 = w3715 & w4052 ;
  assign w4630 = ( ~w3548 & w4628 ) | ( ~w3548 & w4629 ) | ( w4628 & w4629 ) ;
  assign w4631 = w3913 | w4147 ;
  assign w4632 = w3907 | w4630 ;
  assign w4633 = ( w3964 & w4630 ) | ( w3964 & w4632 ) | ( w4630 & w4632 ) ;
  assign w4634 = ( ~w3913 & w4631 ) | ( ~w3913 & w4633 ) | ( w4631 & w4633 ) ;
  assign w4635 = \pi26 ^ w4634 ;
  assign w4636 = w4173 ^ w4554 ;
  assign w4637 = w4267 ^ w4636 ;
  assign w4638 = w381 | w3649 ;
  assign w4639 = ~w3094 & w3717 ;
  assign w4640 = ( ~w381 & w4638 ) | ( ~w381 & w4639 ) | ( w4638 & w4639 ) ;
  assign w4641 = ~w3549 & w3647 ;
  assign w4642 = w3810 | w4640 ;
  assign w4643 = ( w3448 & w4640 ) | ( w3448 & w4642 ) | ( w4640 & w4642 ) ;
  assign w4644 = ( w3647 & ~w4641 ) | ( w3647 & w4643 ) | ( ~w4641 & w4643 ) ;
  assign w4645 = \pi29 ^ w4644 ;
  assign w4646 = ( w4635 & ~w4637 ) | ( w4635 & w4645 ) | ( ~w4637 & w4645 ) ;
  assign w4647 = ( w4617 & w4627 ) | ( w4617 & w4646 ) | ( w4627 & w4646 ) ;
  assign w4648 = w4558 ^ w4568 ;
  assign w4649 = w4556 ^ w4648 ;
  assign w4650 = ( \pi20 & \pi21 ) | ( \pi20 & \pi22 ) | ( \pi21 & \pi22 ) ;
  assign w4651 = \pi22 ^ w4650 ;
  assign w4652 = ~w4600 & w4651 ;
  assign w4653 = ( ~w3962 & w4606 ) | ( ~w3962 & w4652 ) | ( w4606 & w4652 ) ;
  assign w4654 = ( ~w3962 & w4601 ) | ( ~w3962 & w4653 ) | ( w4601 & w4653 ) ;
  assign w4655 = ( w4600 & w4601 ) | ( w4600 & w4609 ) | ( w4601 & w4609 ) ;
  assign w4656 = ( w4652 & ~w4654 ) | ( w4652 & w4655 ) | ( ~w4654 & w4655 ) ;
  assign w4657 = w3962 & w4600 ;
  assign w4658 = ( w4653 & w4656 ) | ( w4653 & ~w4657 ) | ( w4656 & ~w4657 ) ;
  assign w4659 = \pi23 ^ w4658 ;
  assign w4660 = ( w4647 & ~w4649 ) | ( w4647 & w4659 ) | ( ~w4649 & w4659 ) ;
  assign w4661 = w4635 ^ w4637 ;
  assign w4662 = w4645 ^ w4661 ;
  assign w4663 = w4351 ^ w4543 ;
  assign w4664 = w4198 ^ w4663 ;
  assign w4665 = w979 ^ w2994 ;
  assign w4666 = w1085 ^ w4665 ;
  assign w4667 = ~w37 & w4666 ;
  assign w4668 = w1205 & w3098 ;
  assign w4669 = ( w4666 & ~w4667 ) | ( w4666 & w4668 ) | ( ~w4667 & w4668 ) ;
  assign w4670 = ( \pi29 & \pi30 ) | ( \pi29 & w979 ) | ( \pi30 & w979 ) ;
  assign w4671 = \pi31 | w4670 ;
  assign w4672 = ( \pi29 & ~\pi30 ) | ( \pi29 & w1085 ) | ( ~\pi30 & w1085 ) ;
  assign w4673 = ( \pi29 & \pi31 ) | ( \pi29 & ~w4672 ) | ( \pi31 & ~w4672 ) ;
  assign w4674 = ( w4669 & w4671 ) | ( w4669 & ~w4673 ) | ( w4671 & ~w4673 ) ;
  assign w4675 = w883 | w3649 ;
  assign w4676 = w721 & w3717 ;
  assign w4677 = ( ~w883 & w4675 ) | ( ~w883 & w4676 ) | ( w4675 & w4676 ) ;
  assign w4678 = w592 & ~w3549 ;
  assign w4679 = w3421 | w4677 ;
  assign w4680 = ( w3448 & w4677 ) | ( w3448 & w4679 ) | ( w4677 & w4679 ) ;
  assign w4681 = ( w592 & ~w4678 ) | ( w592 & w4680 ) | ( ~w4678 & w4680 ) ;
  assign w4682 = \pi29 ^ w4681 ;
  assign w4683 = ( ~w4664 & w4674 ) | ( ~w4664 & w4682 ) | ( w4674 & w4682 ) ;
  assign w4684 = w4281 ^ w4544 ;
  assign w4685 = w4271 ^ w4684 ;
  assign w4686 = w592 & ~w3717 ;
  assign w4687 = w721 & w3649 ;
  assign w4688 = ( w592 & ~w4686 ) | ( w592 & w4687 ) | ( ~w4686 & w4687 ) ;
  assign w4689 = w381 | w3549 ;
  assign w4690 = w3435 & ~w4688 ;
  assign w4691 = ( w3448 & w4688 ) | ( w3448 & ~w4690 ) | ( w4688 & ~w4690 ) ;
  assign w4692 = ( ~w381 & w4689 ) | ( ~w381 & w4691 ) | ( w4689 & w4691 ) ;
  assign w4693 = \pi29 ^ w4692 ;
  assign w4694 = ( w4683 & w4685 ) | ( w4683 & w4693 ) | ( w4685 & w4693 ) ;
  assign w4695 = w4269 ^ w4553 ;
  assign w4696 = w4545 ^ w4695 ;
  assign w4697 = w3647 & ~w4052 ;
  assign w4698 = w3715 & w4143 ;
  assign w4699 = ( w3647 & ~w4697 ) | ( w3647 & w4698 ) | ( ~w4697 & w4698 ) ;
  assign w4700 = w3725 | w4147 ;
  assign w4701 = w3548 & ~w4699 ;
  assign w4702 = ( w3964 & w4699 ) | ( w3964 & ~w4701 ) | ( w4699 & ~w4701 ) ;
  assign w4703 = ( ~w3725 & w4700 ) | ( ~w3725 & w4702 ) | ( w4700 & w4702 ) ;
  assign w4704 = \pi26 ^ w4703 ;
  assign w4705 = ( w4694 & w4696 ) | ( w4694 & w4704 ) | ( w4696 & w4704 ) ;
  assign w4706 = ~w4607 & w4608 ;
  assign w4707 = w4049 | w4606 ;
  assign w4708 = ~w4142 & w4651 ;
  assign w4709 = ( ~w4049 & w4707 ) | ( ~w4049 & w4708 ) | ( w4707 & w4708 ) ;
  assign w4710 = w3962 | w4706 ;
  assign w4711 = w4152 & ~w4709 ;
  assign w4712 = ( w4609 & w4709 ) | ( w4609 & ~w4711 ) | ( w4709 & ~w4711 ) ;
  assign w4713 = ( ~w3962 & w4710 ) | ( ~w3962 & w4712 ) | ( w4710 & w4712 ) ;
  assign w4714 = \pi23 ^ w4713 ;
  assign w4715 = ( ~w4662 & w4705 ) | ( ~w4662 & w4714 ) | ( w4705 & w4714 ) ;
  assign w4716 = ~w4142 & w4606 ;
  assign w4717 = ( ~w4600 & w4706 ) | ( ~w4600 & w4716 ) | ( w4706 & w4716 ) ;
  assign w4718 = w4651 | w4717 ;
  assign w4719 = ( ~w3962 & w4717 ) | ( ~w3962 & w4718 ) | ( w4717 & w4718 ) ;
  assign w4720 = w4716 | w4719 ;
  assign w4721 = w3962 ^ w4601 ;
  assign w4722 = w4600 ^ w4721 ;
  assign w4723 = w4627 ^ w4646 ;
  assign w4724 = w4617 ^ w4723 ;
  assign w4725 = ~w4720 & w4722 ;
  assign w4726 = ( w4609 & w4720 ) | ( w4609 & ~w4725 ) | ( w4720 & ~w4725 ) ;
  assign w4727 = \pi23 ^ w4726 ;
  assign w4728 = ( w4715 & w4724 ) | ( w4715 & w4727 ) | ( w4724 & w4727 ) ;
  assign w4729 = \pi23 ^ w4647 ;
  assign w4730 = w4649 ^ w4729 ;
  assign w4731 = w4658 ^ w4730 ;
  assign w4732 = w4609 & w4722 ;
  assign w4733 = ( w4609 & w4720 ) | ( w4609 & ~w4732 ) | ( w4720 & ~w4732 ) ;
  assign w4734 = w4715 ^ w4733 ;
  assign w4735 = \pi23 ^ w4724 ;
  assign w4736 = w4734 ^ w4735 ;
  assign w4737 = w4696 ^ w4704 ;
  assign w4738 = w4694 ^ w4737 ;
  assign w4739 = w4683 ^ w4693 ;
  assign w4740 = w4685 ^ w4739 ;
  assign w4741 = w3647 & ~w4143 ;
  assign w4742 = ~w3094 & w4052 ;
  assign w4743 = ( w3647 & ~w4741 ) | ( w3647 & w4742 ) | ( ~w4741 & w4742 ) ;
  assign w4744 = w4147 | w4164 ;
  assign w4745 = w3715 | w4743 ;
  assign w4746 = ( w3964 & w4743 ) | ( w3964 & w4745 ) | ( w4743 & w4745 ) ;
  assign w4747 = ( ~w4164 & w4744 ) | ( ~w4164 & w4746 ) | ( w4744 & w4746 ) ;
  assign w4748 = \pi26 ^ w4747 ;
  assign w4749 = w4664 ^ w4682 ;
  assign w4750 = w4674 ^ w4749 ;
  assign w4751 = w4351 ^ w4542 ;
  assign w4752 = w4531 ^ w4751 ;
  assign w4753 = w4444 ^ w4530 ;
  assign w4754 = \pi14 ^ w4753 ;
  assign w4755 = ( w312 & w525 ) | ( w312 & ~w623 ) | ( w525 & ~w623 ) ;
  assign w4756 = w124 | w164 ;
  assign w4757 = ( ~w164 & w623 ) | ( ~w164 & w642 ) | ( w623 & w642 ) ;
  assign w4758 = w4756 | w4757 ;
  assign w4759 = w4755 | w4758 ;
  assign w4760 = ( ~w384 & w673 ) | ( ~w384 & w4759 ) | ( w673 & w4759 ) ;
  assign w4761 = w384 | w4760 ;
  assign w4762 = w315 | w443 ;
  assign w4763 = ( ~w315 & w316 ) | ( ~w315 & w1421 ) | ( w316 & w1421 ) ;
  assign w4764 = w4762 | w4763 ;
  assign w4765 = ( w127 & w568 ) | ( w127 & ~w573 ) | ( w568 & ~w573 ) ;
  assign w4766 = w2470 | w4764 ;
  assign w4767 = ( w573 & w901 ) | ( w573 & ~w2470 ) | ( w901 & ~w2470 ) ;
  assign w4768 = w4766 | w4767 ;
  assign w4769 = w4765 | w4768 ;
  assign w4770 = ( ~w122 & w888 ) | ( ~w122 & w988 ) | ( w888 & w988 ) ;
  assign w4771 = w110 | w4769 ;
  assign w4772 = ( w122 & w505 ) | ( w122 & ~w4769 ) | ( w505 & ~w4769 ) ;
  assign w4773 = w4771 | w4772 ;
  assign w4774 = w4770 | w4773 ;
  assign w4775 = w144 | w203 ;
  assign w4776 = w1884 | w4775 ;
  assign w4777 = ( ~w1884 & w2705 ) | ( ~w1884 & w4774 ) | ( w2705 & w4774 ) ;
  assign w4778 = w4776 | w4777 ;
  assign w4779 = ( w141 & w229 ) | ( w141 & ~w268 ) | ( w229 & ~w268 ) ;
  assign w4780 = w4174 | w4778 ;
  assign w4781 = ( w268 & w593 ) | ( w268 & ~w4174 ) | ( w593 & ~w4174 ) ;
  assign w4782 = w4780 | w4781 ;
  assign w4783 = w4779 | w4782 ;
  assign w4784 = w318 | w353 ;
  assign w4785 = ( w362 & w511 ) | ( w362 & ~w1094 ) | ( w511 & ~w1094 ) ;
  assign w4786 = w84 | w285 ;
  assign w4787 = ( ~w285 & w1094 ) | ( ~w285 & w1340 ) | ( w1094 & w1340 ) ;
  assign w4788 = w4786 | w4787 ;
  assign w4789 = w4785 | w4788 ;
  assign w4790 = w210 | w388 ;
  assign w4791 = w131 | w4790 ;
  assign w4792 = ( ~w131 & w163 ) | ( ~w131 & w4789 ) | ( w163 & w4789 ) ;
  assign w4793 = w4791 | w4792 ;
  assign w4794 = w226 | w980 ;
  assign w4795 = ( w179 & ~w226 ) | ( w179 & w257 ) | ( ~w226 & w257 ) ;
  assign w4796 = w4794 | w4795 ;
  assign w4797 = w725 | w4464 ;
  assign w4798 = ( w1814 & ~w4464 ) | ( w1814 & w4796 ) | ( ~w4464 & w4796 ) ;
  assign w4799 = w4797 | w4798 ;
  assign w4800 = w432 | w4799 ;
  assign w4801 = ( w279 & w4793 ) | ( w279 & ~w4799 ) | ( w4793 & ~w4799 ) ;
  assign w4802 = w4800 | w4801 ;
  assign w4803 = w952 | w4784 ;
  assign w4804 = ( ~w952 & w2306 ) | ( ~w952 & w4802 ) | ( w2306 & w4802 ) ;
  assign w4805 = w4803 | w4804 ;
  assign w4806 = w466 | w560 ;
  assign w4807 = w326 | w4806 ;
  assign w4808 = ( w258 & ~w326 ) | ( w258 & w4805 ) | ( ~w326 & w4805 ) ;
  assign w4809 = w4807 | w4808 ;
  assign w4810 = ( w165 & w408 ) | ( w165 & ~w606 ) | ( w408 & ~w606 ) ;
  assign w4811 = w119 | w4809 ;
  assign w4812 = ( ~w119 & w606 ) | ( ~w119 & w802 ) | ( w606 & w802 ) ;
  assign w4813 = w4811 | w4812 ;
  assign w4814 = w4810 | w4813 ;
  assign w4815 = w561 | w680 ;
  assign w4816 = w175 | w4815 ;
  assign w4817 = ( w135 & ~w175 ) | ( w135 & w534 ) | ( ~w175 & w534 ) ;
  assign w4818 = w4816 | w4817 ;
  assign w4819 = ( w232 & w389 ) | ( w232 & ~w465 ) | ( w389 & ~w465 ) ;
  assign w4820 = w51 | w4818 ;
  assign w4821 = ( ~w51 & w465 ) | ( ~w51 & w567 ) | ( w465 & w567 ) ;
  assign w4822 = w4820 | w4821 ;
  assign w4823 = w4819 | w4822 ;
  assign w4824 = ( w147 & w205 ) | ( w147 & ~w272 ) | ( w205 & ~w272 ) ;
  assign w4825 = w572 | w4823 ;
  assign w4826 = ( w272 & ~w572 ) | ( w272 & w1031 ) | ( ~w572 & w1031 ) ;
  assign w4827 = w4825 | w4826 ;
  assign w4828 = w4824 | w4827 ;
  assign w4829 = ( ~w224 & w383 ) | ( ~w224 & w4828 ) | ( w383 & w4828 ) ;
  assign w4830 = w224 | w4829 ;
  assign w4831 = ( w59 & ~w496 ) | ( w59 & w1276 ) | ( ~w496 & w1276 ) ;
  assign w4832 = w410 | w4830 ;
  assign w4833 = ( ~w410 & w496 ) | ( ~w410 & w899 ) | ( w496 & w899 ) ;
  assign w4834 = w4832 | w4833 ;
  assign w4835 = w4831 | w4834 ;
  assign w4836 = ( ~w1617 & w4761 ) | ( ~w1617 & w4835 ) | ( w4761 & w4835 ) ;
  assign w4837 = w4783 | w4814 ;
  assign w4838 = ( w1617 & w1990 ) | ( w1617 & ~w4814 ) | ( w1990 & ~w4814 ) ;
  assign w4839 = w4837 | w4838 ;
  assign w4840 = w4836 | w4839 ;
  assign w4841 = ( w56 & w286 ) | ( w56 & ~w445 ) | ( w286 & ~w445 ) ;
  assign w4842 = w416 | w4840 ;
  assign w4843 = ( ~w416 & w445 ) | ( ~w416 & w674 ) | ( w445 & w674 ) ;
  assign w4844 = w4842 | w4843 ;
  assign w4845 = w4841 | w4844 ;
  assign w4846 = ( w221 & w253 ) | ( w221 & ~w265 ) | ( w253 & ~w265 ) ;
  assign w4847 = w215 | w4845 ;
  assign w4848 = ( ~w215 & w265 ) | ( ~w215 & w533 ) | ( w265 & w533 ) ;
  assign w4849 = w4847 | w4848 ;
  assign w4850 = w4846 | w4849 ;
  assign w4851 = w1264 ^ w2991 ;
  assign w4852 = w1399 ^ w4851 ;
  assign w4853 = ( \pi29 & \pi31 ) | ( \pi29 & w1399 ) | ( \pi31 & w1399 ) ;
  assign w4854 = ( \pi29 & ~\pi30 ) | ( \pi29 & w4853 ) | ( ~\pi30 & w4853 ) ;
  assign w4855 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w4853 ) | ( \pi30 & w4853 ) ;
  assign w4856 = ( \pi29 & w1510 ) | ( \pi29 & ~w4855 ) | ( w1510 & ~w4855 ) ;
  assign w4857 = ( ~w1264 & w4855 ) | ( ~w1264 & w4856 ) | ( w4855 & w4856 ) ;
  assign w4858 = ~\pi31 & w4857 ;
  assign w4859 = ( w4854 & ~w4856 ) | ( w4854 & w4858 ) | ( ~w4856 & w4858 ) ;
  assign w4860 = ( w37 & ~w4852 ) | ( w37 & w4859 ) | ( ~w4852 & w4859 ) ;
  assign w4861 = w4859 | w4860 ;
  assign w4862 = ( ~w4444 & w4850 ) | ( ~w4444 & w4861 ) | ( w4850 & w4861 ) ;
  assign w4863 = w1264 ^ w2992 ;
  assign w4864 = w1205 ^ w4863 ;
  assign w4865 = ( \pi30 & \pi31 ) | ( \pi30 & ~w1264 ) | ( \pi31 & ~w1264 ) ;
  assign w4866 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w4865 ) | ( \pi30 & w4865 ) ;
  assign w4867 = ( \pi29 & ~\pi30 ) | ( \pi29 & w4865 ) | ( ~\pi30 & w4865 ) ;
  assign w4868 = ( ~\pi30 & w1399 ) | ( ~\pi30 & w4867 ) | ( w1399 & w4867 ) ;
  assign w4869 = ( w1205 & w4867 ) | ( w1205 & ~w4868 ) | ( w4867 & ~w4868 ) ;
  assign w4870 = ~\pi31 & w4869 ;
  assign w4871 = ( w4866 & w4868 ) | ( w4866 & w4870 ) | ( w4868 & w4870 ) ;
  assign w4872 = ( w37 & ~w4864 ) | ( w37 & w4871 ) | ( ~w4864 & w4871 ) ;
  assign w4873 = w4871 | w4872 ;
  assign w4874 = ( w4754 & w4862 ) | ( w4754 & w4873 ) | ( w4862 & w4873 ) ;
  assign w4875 = w883 | w3717 ;
  assign w4876 = w979 & w3649 ;
  assign w4877 = ( ~w883 & w4875 ) | ( ~w883 & w4876 ) | ( w4875 & w4876 ) ;
  assign w4878 = w721 & ~w3549 ;
  assign w4879 = w4257 & ~w4877 ;
  assign w4880 = ( w3448 & w4877 ) | ( w3448 & ~w4879 ) | ( w4877 & ~w4879 ) ;
  assign w4881 = ( w721 & ~w4878 ) | ( w721 & w4880 ) | ( ~w4878 & w4880 ) ;
  assign w4882 = \pi29 ^ w4881 ;
  assign w4883 = ( w4752 & w4874 ) | ( w4752 & w4882 ) | ( w4874 & w4882 ) ;
  assign w4884 = w381 | w4052 ;
  assign w4885 = ~w3094 & w4143 ;
  assign w4886 = ( ~w381 & w4884 ) | ( ~w381 & w4885 ) | ( w4884 & w4885 ) ;
  assign w4887 = w3810 & ~w4147 ;
  assign w4888 = w3647 | w4886 ;
  assign w4889 = ( w3964 & w4886 ) | ( w3964 & w4888 ) | ( w4886 & w4888 ) ;
  assign w4890 = ( w3810 & ~w4887 ) | ( w3810 & w4889 ) | ( ~w4887 & w4889 ) ;
  assign w4891 = \pi26 ^ w4890 ;
  assign w4892 = ( ~w4750 & w4883 ) | ( ~w4750 & w4891 ) | ( w4883 & w4891 ) ;
  assign w4893 = ( w4740 & w4748 ) | ( w4740 & w4892 ) | ( w4748 & w4892 ) ;
  assign w4894 = w4049 | w4651 ;
  assign w4895 = w3907 & w4606 ;
  assign w4896 = ( ~w4049 & w4894 ) | ( ~w4049 & w4895 ) | ( w4894 & w4895 ) ;
  assign w4897 = w4142 | w4706 ;
  assign w4898 = w4563 | w4896 ;
  assign w4899 = ( w4609 & w4896 ) | ( w4609 & w4898 ) | ( w4896 & w4898 ) ;
  assign w4900 = ( ~w4142 & w4897 ) | ( ~w4142 & w4899 ) | ( w4897 & w4899 ) ;
  assign w4901 = \pi23 ^ w4900 ;
  assign w4902 = ( w4738 & w4893 ) | ( w4738 & w4901 ) | ( w4893 & w4901 ) ;
  assign w4903 = ( \pi18 & ~\pi19 ) | ( \pi18 & \pi20 ) | ( ~\pi19 & \pi20 ) ;
  assign w4904 = ( \pi17 & \pi18 ) | ( \pi17 & w4903 ) | ( \pi18 & w4903 ) ;
  assign w4905 = w4903 ^ w4904 ;
  assign w4906 = \pi19 ^ \pi20 ;
  assign w4907 = \pi17 ^ \pi18 ;
  assign w4908 = w4906 & w4907 ;
  assign w4909 = ~w4600 & w4905 ;
  assign w4910 = w4908 | w4909 ;
  assign w4911 = ( ~w4603 & w4909 ) | ( ~w4603 & w4910 ) | ( w4909 & w4910 ) ;
  assign w4912 = \pi20 ^ w4911 ;
  assign w4913 = w4662 ^ w4714 ;
  assign w4914 = w4705 ^ w4913 ;
  assign w4915 = ( w4902 & w4912 ) | ( w4902 & ~w4914 ) | ( w4912 & ~w4914 ) ;
  assign w4916 = w4912 ^ w4914 ;
  assign w4917 = w4902 ^ w4916 ;
  assign w4918 = w4738 ^ w4901 ;
  assign w4919 = w4893 ^ w4918 ;
  assign w4920 = w3548 | w4606 ;
  assign w4921 = w3907 & w4651 ;
  assign w4922 = ( ~w3548 & w4920 ) | ( ~w3548 & w4921 ) | ( w4920 & w4921 ) ;
  assign w4923 = w4049 | w4706 ;
  assign w4924 = w4622 & ~w4922 ;
  assign w4925 = ( w4609 & w4922 ) | ( w4609 & ~w4924 ) | ( w4922 & ~w4924 ) ;
  assign w4926 = ( ~w4049 & w4923 ) | ( ~w4049 & w4925 ) | ( w4923 & w4925 ) ;
  assign w4927 = \pi23 ^ w4926 ;
  assign w4928 = w4748 ^ w4892 ;
  assign w4929 = w4740 ^ w4928 ;
  assign w4930 = w4750 ^ w4891 ;
  assign w4931 = w4883 ^ w4930 ;
  assign w4932 = w979 & ~w3717 ;
  assign w4933 = w1085 & w3649 ;
  assign w4934 = ( w979 & ~w4932 ) | ( w979 & w4933 ) | ( ~w4932 & w4933 ) ;
  assign w4935 = w883 | w3549 ;
  assign w4936 = w4273 & ~w4934 ;
  assign w4937 = ( w3448 & w4934 ) | ( w3448 & ~w4936 ) | ( w4934 & ~w4936 ) ;
  assign w4938 = ( ~w883 & w4935 ) | ( ~w883 & w4937 ) | ( w4935 & w4937 ) ;
  assign w4939 = \pi29 ^ w4938 ;
  assign w4940 = w4862 ^ w4873 ;
  assign w4941 = w4754 ^ w4940 ;
  assign w4942 = w4850 ^ w4861 ;
  assign w4943 = w4444 ^ w4942 ;
  assign w4944 = w505 | w1086 ;
  assign w4945 = w220 | w4944 ;
  assign w4946 = ( w127 & ~w220 ) | ( w127 & w384 ) | ( ~w220 & w384 ) ;
  assign w4947 = w4945 | w4946 ;
  assign w4948 = ( w51 & w219 ) | ( w51 & ~w681 ) | ( w219 & ~w681 ) ;
  assign w4949 = w3965 | w4947 ;
  assign w4950 = ( w681 & w1340 ) | ( w681 & ~w4947 ) | ( w1340 & ~w4947 ) ;
  assign w4951 = w4949 | w4950 ;
  assign w4952 = w4948 | w4951 ;
  assign w4953 = w284 | w286 ;
  assign w4954 = w414 | w4953 ;
  assign w4955 = ( ~w414 & w1265 ) | ( ~w414 & w4952 ) | ( w1265 & w4952 ) ;
  assign w4956 = w4954 | w4955 ;
  assign w4957 = w465 | w897 ;
  assign w4958 = ( ~w465 & w593 ) | ( ~w465 & w4956 ) | ( w593 & w4956 ) ;
  assign w4959 = w4957 | w4958 ;
  assign w4960 = w88 | w2093 ;
  assign w4961 = ( ~w88 & w98 ) | ( ~w88 & w1759 ) | ( w98 & w1759 ) ;
  assign w4962 = w4960 | w4961 ;
  assign w4963 = ( ~w128 & w309 ) | ( ~w128 & w4962 ) | ( w309 & w4962 ) ;
  assign w4964 = w128 | w4963 ;
  assign w4965 = w353 | w470 ;
  assign w4966 = w206 | w4965 ;
  assign w4967 = ( ~w206 & w215 ) | ( ~w206 & w1363 ) | ( w215 & w1363 ) ;
  assign w4968 = w4966 | w4967 ;
  assign w4969 = w142 | w837 ;
  assign w4970 = ( ~w142 & w516 ) | ( ~w142 & w4968 ) | ( w516 & w4968 ) ;
  assign w4971 = w4969 | w4970 ;
  assign w4972 = ( w119 & ~w124 ) | ( w119 & w3251 ) | ( ~w124 & w3251 ) ;
  assign w4973 = w4964 | w4971 ;
  assign w4974 = ( w124 & w266 ) | ( w124 & ~w4971 ) | ( w266 & ~w4971 ) ;
  assign w4975 = w4973 | w4974 ;
  assign w4976 = w4972 | w4975 ;
  assign w4977 = ( w272 & w361 ) | ( w272 & ~w392 ) | ( w361 & ~w392 ) ;
  assign w4978 = w103 | w4976 ;
  assign w4979 = ( ~w103 & w392 ) | ( ~w103 & w1128 ) | ( w392 & w1128 ) ;
  assign w4980 = w4978 | w4979 ;
  assign w4981 = w4977 | w4980 ;
  assign w4982 = ( ~w208 & w697 ) | ( ~w208 & w4981 ) | ( w697 & w4981 ) ;
  assign w4983 = w208 | w4982 ;
  assign w4984 = ( w265 & ~w324 ) | ( w265 & w389 ) | ( ~w324 & w389 ) ;
  assign w4985 = w324 | w4984 ;
  assign w4986 = ( w118 & ~w409 ) | ( w118 & w4985 ) | ( ~w409 & w4985 ) ;
  assign w4987 = w999 | w2518 ;
  assign w4988 = ( w409 & w1094 ) | ( w409 & ~w2518 ) | ( w1094 & ~w2518 ) ;
  assign w4989 = w4987 | w4988 ;
  assign w4990 = w4986 | w4989 ;
  assign w4991 = ( w285 & w386 ) | ( w285 & ~w424 ) | ( w386 & ~w424 ) ;
  assign w4992 = w227 | w4990 ;
  assign w4993 = ( ~w227 & w424 ) | ( ~w227 & w512 ) | ( w424 & w512 ) ;
  assign w4994 = w4992 | w4993 ;
  assign w4995 = w4991 | w4994 ;
  assign w4996 = ( w1654 & ~w4422 ) | ( w1654 & w4959 ) | ( ~w4422 & w4959 ) ;
  assign w4997 = w3059 | w4983 ;
  assign w4998 = ( w4422 & ~w4983 ) | ( w4422 & w4995 ) | ( ~w4983 & w4995 ) ;
  assign w4999 = w4997 | w4998 ;
  assign w5000 = w4996 | w4999 ;
  assign w5001 = w764 | w1126 ;
  assign w5002 = w176 | w5001 ;
  assign w5003 = ( ~w176 & w565 ) | ( ~w176 & w5000 ) | ( w565 & w5000 ) ;
  assign w5004 = w5002 | w5003 ;
  assign w5005 = w511 | w758 ;
  assign w5006 = ( w265 & ~w511 ) | ( w265 & w565 ) | ( ~w511 & w565 ) ;
  assign w5007 = w5005 | w5006 ;
  assign w5008 = ( w164 & w458 ) | ( w164 & ~w504 ) | ( w458 & ~w504 ) ;
  assign w5009 = w627 | w5007 ;
  assign w5010 = ( w504 & w525 ) | ( w504 & ~w5007 ) | ( w525 & ~w5007 ) ;
  assign w5011 = w5009 | w5010 ;
  assign w5012 = w5008 | w5011 ;
  assign w5013 = w393 | w408 ;
  assign w5014 = w911 | w5013 ;
  assign w5015 = ( w113 & ~w911 ) | ( w113 & w5012 ) | ( ~w911 & w5012 ) ;
  assign w5016 = w5014 | w5015 ;
  assign w5017 = w726 | w860 ;
  assign w5018 = w262 | w5017 ;
  assign w5019 = ( w202 & ~w262 ) | ( w202 & w392 ) | ( ~w262 & w392 ) ;
  assign w5020 = w5018 | w5019 ;
  assign w5021 = w167 | w227 ;
  assign w5022 = w671 | w5021 ;
  assign w5023 = ( ~w671 & w5016 ) | ( ~w671 & w5020 ) | ( w5016 & w5020 ) ;
  assign w5024 = w5022 | w5023 ;
  assign w5025 = ( ~w1712 & w1713 ) | ( ~w1712 & w5024 ) | ( w1713 & w5024 ) ;
  assign w5026 = w1712 | w5025 ;
  assign w5027 = ( w141 & ~w313 ) | ( w141 & w1064 ) | ( ~w313 & w1064 ) ;
  assign w5028 = w343 | w5026 ;
  assign w5029 = ( w313 & ~w343 ) | ( w313 & w623 ) | ( ~w343 & w623 ) ;
  assign w5030 = w5028 | w5029 ;
  assign w5031 = w5027 | w5030 ;
  assign w5032 = ( w318 & w362 ) | ( w318 & ~w817 ) | ( w362 & ~w817 ) ;
  assign w5033 = w128 | w5031 ;
  assign w5034 = ( ~w128 & w817 ) | ( ~w128 & w1229 ) | ( w817 & w1229 ) ;
  assign w5035 = w5033 | w5034 ;
  assign w5036 = w5032 | w5035 ;
  assign w5037 = w280 | w837 ;
  assign w5038 = ( w98 & ~w280 ) | ( w98 & w492 ) | ( ~w280 & w492 ) ;
  assign w5039 = w5037 | w5038 ;
  assign w5040 = w680 | w783 ;
  assign w5041 = w390 | w5040 ;
  assign w5042 = ( ~w390 & w608 ) | ( ~w390 & w1131 ) | ( w608 & w1131 ) ;
  assign w5043 = w5041 | w5042 ;
  assign w5044 = ( w119 & w266 ) | ( w119 & ~w467 ) | ( w266 & ~w467 ) ;
  assign w5045 = w3762 | w5043 ;
  assign w5046 = ( w467 & w674 ) | ( w467 & ~w5043 ) | ( w674 & ~w5043 ) ;
  assign w5047 = w5045 | w5046 ;
  assign w5048 = w5044 | w5047 ;
  assign w5049 = w2253 | w5039 ;
  assign w5050 = w5048 | w5049 ;
  assign w5051 = ( w3172 & w5036 ) | ( w3172 & ~w5048 ) | ( w5036 & ~w5048 ) ;
  assign w5052 = w5050 | w5051 ;
  assign w5053 = ( w82 & ~w257 ) | ( w82 & w410 ) | ( ~w257 & w410 ) ;
  assign w5054 = w4959 | w5052 ;
  assign w5055 = ( w257 & w317 ) | ( w257 & ~w4959 ) | ( w317 & ~w4959 ) ;
  assign w5056 = w5054 | w5055 ;
  assign w5057 = w5053 | w5056 ;
  assign w5058 = ( w268 & w418 ) | ( w268 & ~w506 ) | ( w418 & ~w506 ) ;
  assign w5059 = w260 | w5057 ;
  assign w5060 = ( ~w260 & w506 ) | ( ~w260 & w596 ) | ( w506 & w596 ) ;
  assign w5061 = w5059 | w5060 ;
  assign w5062 = w5058 | w5061 ;
  assign w5063 = w423 | w951 ;
  assign w5064 = w320 | w5063 ;
  assign w5065 = ( ~w320 & w325 ) | ( ~w320 & w5062 ) | ( w325 & w5062 ) ;
  assign w5066 = w5064 | w5065 ;
  assign w5067 = ( ~\pi11 & w5004 ) | ( ~\pi11 & w5066 ) | ( w5004 & w5066 ) ;
  assign w5068 = w1399 ^ w2990 ;
  assign w5069 = w1510 ^ w5068 ;
  assign w5070 = ( \pi29 & \pi31 ) | ( \pi29 & ~w1510 ) | ( \pi31 & ~w1510 ) ;
  assign w5071 = ( \pi29 & ~\pi30 ) | ( \pi29 & w5070 ) | ( ~\pi30 & w5070 ) ;
  assign w5072 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w5070 ) | ( \pi30 & w5070 ) ;
  assign w5073 = ( ~\pi29 & w1614 ) | ( ~\pi29 & w5072 ) | ( w1614 & w5072 ) ;
  assign w5074 = ( w1399 & w5072 ) | ( w1399 & ~w5073 ) | ( w5072 & ~w5073 ) ;
  assign w5075 = ~\pi31 & w5074 ;
  assign w5076 = ( w5071 & w5073 ) | ( w5071 & w5075 ) | ( w5073 & w5075 ) ;
  assign w5077 = ( w37 & ~w5069 ) | ( w37 & w5076 ) | ( ~w5069 & w5076 ) ;
  assign w5078 = w5076 | w5077 ;
  assign w5079 = ( ~w4444 & w5067 ) | ( ~w4444 & w5078 ) | ( w5067 & w5078 ) ;
  assign w5080 = w5067 ^ w5078 ;
  assign w5081 = w4444 ^ w5080 ;
  assign w5082 = w5004 ^ w5066 ;
  assign w5083 = \pi11 ^ w5082 ;
  assign w5084 = w1614 ^ w2989 ;
  assign w5085 = w1510 ^ w5084 ;
  assign w5086 = w37 | w5085 ;
  assign w5087 = w1711 & w3098 ;
  assign w5088 = ( ~w5085 & w5086 ) | ( ~w5085 & w5087 ) | ( w5086 & w5087 ) ;
  assign w5089 = ( \pi29 & \pi30 ) | ( \pi29 & ~w1510 ) | ( \pi30 & ~w1510 ) ;
  assign w5090 = \pi31 | w5089 ;
  assign w5091 = ( \pi29 & ~\pi30 ) | ( \pi29 & w1614 ) | ( ~\pi30 & w1614 ) ;
  assign w5092 = ( \pi29 & \pi31 ) | ( \pi29 & ~w5091 ) | ( \pi31 & ~w5091 ) ;
  assign w5093 = ( w5088 & w5090 ) | ( w5088 & ~w5092 ) | ( w5090 & ~w5092 ) ;
  assign w5094 = w179 | w568 ;
  assign w5095 = w74 | w5094 ;
  assign w5096 = ( ~w74 & w81 ) | ( ~w74 & w1208 ) | ( w81 & w1208 ) ;
  assign w5097 = w5095 | w5096 ;
  assign w5098 = ( ~w252 & w422 ) | ( ~w252 & w1560 ) | ( w422 & w1560 ) ;
  assign w5099 = w252 | w5098 ;
  assign w5100 = w139 | w229 ;
  assign w5101 = w936 | w5100 ;
  assign w5102 = ( ~w936 & w1363 ) | ( ~w936 & w5099 ) | ( w1363 & w5099 ) ;
  assign w5103 = w5101 | w5102 ;
  assign w5104 = ( w3748 & ~w5097 ) | ( w3748 & w5103 ) | ( ~w5097 & w5103 ) ;
  assign w5105 = w1628 | w1679 ;
  assign w5106 = ( ~w1628 & w1977 ) | ( ~w1628 & w5097 ) | ( w1977 & w5097 ) ;
  assign w5107 = w5105 | w5106 ;
  assign w5108 = w5104 | w5107 ;
  assign w5109 = ( w138 & w424 ) | ( w138 & ~w513 ) | ( w424 & ~w513 ) ;
  assign w5110 = w782 | w5108 ;
  assign w5111 = ( w513 & ~w782 ) | ( w513 & w1094 ) | ( ~w782 & w1094 ) ;
  assign w5112 = w5110 | w5111 ;
  assign w5113 = w5109 | w5112 ;
  assign w5114 = ( w309 & w534 ) | ( w309 & ~w681 ) | ( w534 & ~w681 ) ;
  assign w5115 = w272 | w5113 ;
  assign w5116 = ( ~w272 & w681 ) | ( ~w272 & w837 ) | ( w681 & w837 ) ;
  assign w5117 = w5115 | w5116 ;
  assign w5118 = w5114 | w5117 ;
  assign w5119 = ( w269 & w312 ) | ( w269 & ~w322 ) | ( w312 & ~w322 ) ;
  assign w5120 = w1154 | w2376 ;
  assign w5121 = ( w322 & w421 ) | ( w322 & ~w1154 ) | ( w421 & ~w1154 ) ;
  assign w5122 = w5120 | w5121 ;
  assign w5123 = w5119 | w5122 ;
  assign w5124 = ( ~w225 & w343 ) | ( ~w225 & w661 ) | ( w343 & w661 ) ;
  assign w5125 = w4451 | w5123 ;
  assign w5126 = ( w225 & w511 ) | ( w225 & ~w4451 ) | ( w511 & ~w4451 ) ;
  assign w5127 = w5125 | w5126 ;
  assign w5128 = w5124 | w5127 ;
  assign w5129 = w386 | w573 ;
  assign w5130 = w3251 | w5129 ;
  assign w5131 = ( w203 & ~w3251 ) | ( w203 & w5128 ) | ( ~w3251 & w5128 ) ;
  assign w5132 = w5130 | w5131 ;
  assign w5133 = ( w254 & w277 ) | ( w254 & ~w641 ) | ( w277 & ~w641 ) ;
  assign w5134 = w175 | w5132 ;
  assign w5135 = ( ~w175 & w641 ) | ( ~w175 & w1001 ) | ( w641 & w1001 ) ;
  assign w5136 = w5134 | w5135 ;
  assign w5137 = w5133 | w5136 ;
  assign w5138 = ( w268 & w311 ) | ( w268 & ~w459 ) | ( w311 & ~w459 ) ;
  assign w5139 = w141 | w2536 ;
  assign w5140 = ( ~w141 & w459 ) | ( ~w141 & w1031 ) | ( w459 & w1031 ) ;
  assign w5141 = w5139 | w5140 ;
  assign w5142 = w5138 | w5141 ;
  assign w5143 = ( w339 & w413 ) | ( w339 & ~w505 ) | ( w413 & ~w505 ) ;
  assign w5144 = w133 | w310 ;
  assign w5145 = ( ~w310 & w505 ) | ( ~w310 & w681 ) | ( w505 & w681 ) ;
  assign w5146 = w5144 | w5145 ;
  assign w5147 = w5143 | w5146 ;
  assign w5148 = w901 | w980 ;
  assign w5149 = w352 | w5148 ;
  assign w5150 = ( ~w352 & w608 ) | ( ~w352 & w5147 ) | ( w608 & w5147 ) ;
  assign w5151 = w5149 | w5150 ;
  assign w5152 = ( w214 & w443 ) | ( w214 & ~w449 ) | ( w443 & ~w449 ) ;
  assign w5153 = w147 | w206 ;
  assign w5154 = ( ~w206 & w449 ) | ( ~w206 & w758 ) | ( w449 & w758 ) ;
  assign w5155 = w5153 | w5154 ;
  assign w5156 = w5152 | w5155 ;
  assign w5157 = ( ~w221 & w359 ) | ( ~w221 & w431 ) | ( w359 & w431 ) ;
  assign w5158 = w119 | w5156 ;
  assign w5159 = ( ~w119 & w431 ) | ( ~w119 & w662 ) | ( w431 & w662 ) ;
  assign w5160 = w5158 | w5159 ;
  assign w5161 = w5157 & ~w5160 ;
  assign w5162 = w447 | w456 ;
  assign w5163 = w115 | w5162 ;
  assign w5164 = ( w103 & ~w115 ) | ( w103 & w265 ) | ( ~w115 & w265 ) ;
  assign w5165 = w5163 | w5164 ;
  assign w5166 = ( ~w205 & w1157 ) | ( ~w205 & w5165 ) | ( w1157 & w5165 ) ;
  assign w5167 = ~w1044 & w5161 ;
  assign w5168 = ( w205 & w595 ) | ( w205 & ~w1044 ) | ( w595 & ~w1044 ) ;
  assign w5169 = w5167 & ~w5168 ;
  assign w5170 = ~w5166 & w5169 ;
  assign w5171 = ( w76 & w138 ) | ( w76 & ~w409 ) | ( w138 & ~w409 ) ;
  assign w5172 = ~w5151 & w5170 ;
  assign w5173 = ( w409 & w626 ) | ( w409 & ~w5151 ) | ( w626 & ~w5151 ) ;
  assign w5174 = w5172 & ~w5173 ;
  assign w5175 = ~w5171 & w5174 ;
  assign w5176 = ( w470 & w571 ) | ( w470 & ~w628 ) | ( w571 & ~w628 ) ;
  assign w5177 = ~w144 & w5175 ;
  assign w5178 = ( ~w144 & w628 ) | ( ~w144 & w1130 ) | ( w628 & w1130 ) ;
  assign w5179 = w5177 & ~w5178 ;
  assign w5180 = ~w5176 & w5179 ;
  assign w5181 = w530 | w569 ;
  assign w5182 = w256 | w5181 ;
  assign w5183 = ( ~w256 & w430 ) | ( ~w256 & w1181 ) | ( w430 & w1181 ) ;
  assign w5184 = w5182 | w5183 ;
  assign w5185 = w280 | w314 ;
  assign w5186 = w1401 | w5185 ;
  assign w5187 = ( w98 & ~w1401 ) | ( w98 & w5184 ) | ( ~w1401 & w5184 ) ;
  assign w5188 = w5186 | w5187 ;
  assign w5189 = w44 | w722 ;
  assign w5190 = ( ~w44 & w531 ) | ( ~w44 & w5188 ) | ( w531 & w5188 ) ;
  assign w5191 = w5189 | w5190 ;
  assign w5192 = ( w340 & w512 ) | ( w340 & ~w1086 ) | ( w512 & ~w1086 ) ;
  assign w5193 = ( ~w232 & w1086 ) | ( ~w232 & w1094 ) | ( w1086 & w1094 ) ;
  assign w5194 = w4457 | w5193 ;
  assign w5195 = w5192 | w5194 ;
  assign w5196 = w128 | w525 ;
  assign w5197 = ( ~w128 & w281 ) | ( ~w128 & w5195 ) | ( w281 & w5195 ) ;
  assign w5198 = w5196 | w5197 ;
  assign w5199 = ( w262 & w390 ) | ( w262 & ~w392 ) | ( w390 & ~w392 ) ;
  assign w5200 = w124 | w638 ;
  assign w5201 = ( ~w124 & w392 ) | ( ~w124 & w860 ) | ( w392 & w860 ) ;
  assign w5202 = w5200 | w5201 ;
  assign w5203 = w5199 | w5202 ;
  assign w5204 = ( w5142 & w5198 ) | ( w5142 & ~w5203 ) | ( w5198 & ~w5203 ) ;
  assign w5205 = w5180 & ~w5191 ;
  assign w5206 = ( w1875 & ~w5191 ) | ( w1875 & w5203 ) | ( ~w5191 & w5203 ) ;
  assign w5207 = w5205 & ~w5206 ;
  assign w5208 = ~w5204 & w5207 ;
  assign w5209 = ( w324 & w606 ) | ( w324 & ~w723 ) | ( w606 & ~w723 ) ;
  assign w5210 = ~w5137 & w5208 ;
  assign w5211 = ( w723 & w1126 ) | ( w723 & w5208 ) | ( w1126 & w5208 ) ;
  assign w5212 = w5210 & ~w5211 ;
  assign w5213 = ~w5209 & w5212 ;
  assign w5214 = ( w176 & w320 ) | ( w176 & ~w423 ) | ( w320 & ~w423 ) ;
  assign w5215 = ~w114 & w5213 ;
  assign w5216 = ( ~w114 & w423 ) | ( ~w114 & w673 ) | ( w423 & w673 ) ;
  assign w5217 = w5215 & ~w5216 ;
  assign w5218 = ~w5214 & w5217 ;
  assign w5219 = w411 | w449 ;
  assign w5220 = w199 | w5219 ;
  assign w5221 = ( ~w199 & w268 ) | ( ~w199 & w2091 ) | ( w268 & w2091 ) ;
  assign w5222 = w5220 | w5221 ;
  assign w5223 = ( w122 & w342 ) | ( w122 & ~w351 ) | ( w342 & ~w351 ) ;
  assign w5224 = w81 | w5222 ;
  assign w5225 = ( ~w81 & w351 ) | ( ~w81 & w899 ) | ( w351 & w899 ) ;
  assign w5226 = w5224 | w5225 ;
  assign w5227 = w5223 | w5226 ;
  assign w5228 = w165 | w1130 ;
  assign w5229 = ( ~w165 & w443 ) | ( ~w165 & w5227 ) | ( w443 & w5227 ) ;
  assign w5230 = w5228 | w5229 ;
  assign w5231 = ( w161 & w219 ) | ( w161 & ~w226 ) | ( w219 & ~w226 ) ;
  assign w5232 = w638 | w956 ;
  assign w5233 = ( w226 & w257 ) | ( w226 & ~w956 ) | ( w257 & ~w956 ) ;
  assign w5234 = w5232 | w5233 ;
  assign w5235 = w5231 | w5234 ;
  assign w5236 = ( w202 & ~w422 ) | ( w202 & w1154 ) | ( ~w422 & w1154 ) ;
  assign w5237 = w177 | w1087 ;
  assign w5238 = ( w422 & w512 ) | ( w422 & ~w1087 ) | ( w512 & ~w1087 ) ;
  assign w5239 = w5237 | w5238 ;
  assign w5240 = w5236 | w5239 ;
  assign w5241 = ( ~w205 & w887 ) | ( ~w205 & w5240 ) | ( w887 & w5240 ) ;
  assign w5242 = w5230 | w5235 ;
  assign w5243 = ( w205 & w595 ) | ( w205 & ~w5235 ) | ( w595 & ~w5235 ) ;
  assign w5244 = w5242 | w5243 ;
  assign w5245 = w5241 | w5244 ;
  assign w5246 = ( w886 & w1616 ) | ( w886 & ~w2452 ) | ( w1616 & ~w2452 ) ;
  assign w5247 = w627 | w5245 ;
  assign w5248 = ( ~w627 & w1340 ) | ( ~w627 & w2452 ) | ( w1340 & w2452 ) ;
  assign w5249 = w5247 | w5248 ;
  assign w5250 = w5246 | w5249 ;
  assign w5251 = ( w266 & w287 ) | ( w266 & ~w419 ) | ( w287 & ~w419 ) ;
  assign w5252 = w127 | w5250 ;
  assign w5253 = ( ~w127 & w419 ) | ( ~w127 & w516 ) | ( w419 & w516 ) ;
  assign w5254 = w5252 | w5253 ;
  assign w5255 = w5251 | w5254 ;
  assign w5256 = w1031 | w2626 ;
  assign w5257 = ( w608 & w1129 ) | ( w608 & ~w2626 ) | ( w1129 & ~w2626 ) ;
  assign w5258 = w5256 | w5257 ;
  assign w5259 = w90 | w286 ;
  assign w5260 = w672 | w5259 ;
  assign w5261 = ( w74 & ~w672 ) | ( w74 & w5258 ) | ( ~w672 & w5258 ) ;
  assign w5262 = w5260 | w5261 ;
  assign w5263 = w362 | w490 ;
  assign w5264 = w259 | w5263 ;
  assign w5265 = ( ~w259 & w269 ) | ( ~w259 & w5262 ) | ( w269 & w5262 ) ;
  assign w5266 = w5264 | w5265 ;
  assign w5267 = w593 | w674 ;
  assign w5268 = w124 | w5267 ;
  assign w5269 = ( ~w124 & w260 ) | ( ~w124 & w1276 ) | ( w260 & w1276 ) ;
  assign w5270 = w5268 | w5269 ;
  assign w5271 = w568 | w722 ;
  assign w5272 = w322 | w5271 ;
  assign w5273 = ( ~w322 & w345 ) | ( ~w322 & w5270 ) | ( w345 & w5270 ) ;
  assign w5274 = w5272 | w5273 ;
  assign w5275 = ( w169 & ~w561 ) | ( w169 & w3353 ) | ( ~w561 & w3353 ) ;
  assign w5276 = w3401 | w5274 ;
  assign w5277 = ( w561 & w724 ) | ( w561 & ~w5274 ) | ( w724 & ~w5274 ) ;
  assign w5278 = w5276 | w5277 ;
  assign w5279 = w5275 | w5278 ;
  assign w5280 = w3535 | w5266 ;
  assign w5281 = ( w1618 & ~w5266 ) | ( w1618 & w5279 ) | ( ~w5266 & w5279 ) ;
  assign w5282 = w5280 | w5281 ;
  assign w5283 = w120 | w311 ;
  assign w5284 = w5255 | w5283 ;
  assign w5285 = ( w1283 & ~w5255 ) | ( w1283 & w5282 ) | ( ~w5255 & w5282 ) ;
  assign w5286 = w5284 | w5285 ;
  assign w5287 = w392 | w837 ;
  assign w5288 = w64 | w5287 ;
  assign w5289 = ( ~w64 & w318 ) | ( ~w64 & w5286 ) | ( w318 & w5286 ) ;
  assign w5290 = w5288 | w5289 ;
  assign w5291 = w167 | w423 ;
  assign w5292 = ( ~w167 & w278 ) | ( ~w167 & w5290 ) | ( w278 & w5290 ) ;
  assign w5293 = w5291 | w5292 ;
  assign w5294 = ( \pi08 & w5218 ) | ( \pi08 & ~w5293 ) | ( w5218 & ~w5293 ) ;
  assign w5295 = w1711 ^ w2987 ;
  assign w5296 = w1834 ^ w5295 ;
  assign w5297 = ( \pi29 & \pi31 ) | ( \pi29 & ~w1834 ) | ( \pi31 & ~w1834 ) ;
  assign w5298 = ( \pi29 & ~\pi30 ) | ( \pi29 & w5297 ) | ( ~\pi30 & w5297 ) ;
  assign w5299 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w5297 ) | ( \pi30 & w5297 ) ;
  assign w5300 = ( \pi29 & w1939 ) | ( \pi29 & ~w5299 ) | ( w1939 & ~w5299 ) ;
  assign w5301 = ( w1711 & w5299 ) | ( w1711 & w5300 ) | ( w5299 & w5300 ) ;
  assign w5302 = ~\pi31 & w5301 ;
  assign w5303 = ( w5298 & ~w5300 ) | ( w5298 & w5302 ) | ( ~w5300 & w5302 ) ;
  assign w5304 = ( w37 & w5296 ) | ( w37 & w5303 ) | ( w5296 & w5303 ) ;
  assign w5305 = w5303 | w5304 ;
  assign w5306 = ( w5004 & w5294 ) | ( w5004 & ~w5305 ) | ( w5294 & ~w5305 ) ;
  assign w5307 = ( w5004 & ~w5118 ) | ( w5004 & w5306 ) | ( ~w5118 & w5306 ) ;
  assign w5308 = ( w5083 & ~w5093 ) | ( w5083 & w5307 ) | ( ~w5093 & w5307 ) ;
  assign w5309 = w1264 | w3649 ;
  assign w5310 = w1205 & w3717 ;
  assign w5311 = ( ~w1264 & w5309 ) | ( ~w1264 & w5310 ) | ( w5309 & w5310 ) ;
  assign w5312 = w1085 & ~w3549 ;
  assign w5313 = w4533 | w5311 ;
  assign w5314 = ( w3448 & w5311 ) | ( w3448 & w5313 ) | ( w5311 & w5313 ) ;
  assign w5315 = ( w1085 & ~w5312 ) | ( w1085 & w5314 ) | ( ~w5312 & w5314 ) ;
  assign w5316 = \pi29 ^ w5315 ;
  assign w5317 = ( w5081 & w5308 ) | ( w5081 & ~w5316 ) | ( w5308 & ~w5316 ) ;
  assign w5318 = ( w4943 & ~w5079 ) | ( w4943 & w5317 ) | ( ~w5079 & w5317 ) ;
  assign w5319 = ( w4939 & w4941 ) | ( w4939 & ~w5318 ) | ( w4941 & ~w5318 ) ;
  assign w5320 = w4752 ^ w4882 ;
  assign w5321 = w4874 ^ w5320 ;
  assign w5322 = w381 | w4143 ;
  assign w5323 = w592 & w4052 ;
  assign w5324 = ( ~w381 & w5322 ) | ( ~w381 & w5323 ) | ( w5322 & w5323 ) ;
  assign w5325 = w3096 & ~w4147 ;
  assign w5326 = w3094 & ~w5324 ;
  assign w5327 = ( w3964 & w5324 ) | ( w3964 & ~w5326 ) | ( w5324 & ~w5326 ) ;
  assign w5328 = ( w3096 & ~w5325 ) | ( w3096 & w5327 ) | ( ~w5325 & w5327 ) ;
  assign w5329 = \pi26 ^ w5328 ;
  assign w5330 = ( w5319 & w5321 ) | ( w5319 & w5329 ) | ( w5321 & w5329 ) ;
  assign w5331 = w3548 | w4651 ;
  assign w5332 = w3715 & w4606 ;
  assign w5333 = ( ~w3548 & w5331 ) | ( ~w3548 & w5332 ) | ( w5331 & w5332 ) ;
  assign w5334 = w3907 & ~w4706 ;
  assign w5335 = w3913 & ~w5333 ;
  assign w5336 = ( w4609 & w5333 ) | ( w4609 & ~w5335 ) | ( w5333 & ~w5335 ) ;
  assign w5337 = ( w3907 & ~w5334 ) | ( w3907 & w5336 ) | ( ~w5334 & w5336 ) ;
  assign w5338 = \pi23 ^ w5337 ;
  assign w5339 = ( ~w4931 & w5330 ) | ( ~w4931 & w5338 ) | ( w5330 & w5338 ) ;
  assign w5340 = ( w4927 & w4929 ) | ( w4927 & w5339 ) | ( w4929 & w5339 ) ;
  assign w5341 = w4919 ^ w5340 ;
  assign w5342 = ( \pi17 & \pi18 ) | ( \pi17 & \pi19 ) | ( \pi18 & \pi19 ) ;
  assign w5343 = \pi19 ^ w5342 ;
  assign w5344 = ~w4600 & w5343 ;
  assign w5345 = ( ~w3962 & w4905 ) | ( ~w3962 & w5344 ) | ( w4905 & w5344 ) ;
  assign w5346 = ( ~w3962 & w4601 ) | ( ~w3962 & w5345 ) | ( w4601 & w5345 ) ;
  assign w5347 = ( w4600 & w4601 ) | ( w4600 & w4908 ) | ( w4601 & w4908 ) ;
  assign w5348 = ( w5344 & ~w5346 ) | ( w5344 & w5347 ) | ( ~w5346 & w5347 ) ;
  assign w5349 = ( ~w4657 & w5345 ) | ( ~w4657 & w5348 ) | ( w5345 & w5348 ) ;
  assign w5350 = \pi20 ^ w5349 ;
  assign w5351 = ( w4919 & w5340 ) | ( w4919 & w5350 ) | ( w5340 & w5350 ) ;
  assign w5352 = w4931 ^ w5338 ;
  assign w5353 = w5330 ^ w5352 ;
  assign w5354 = w5321 ^ w5329 ;
  assign w5355 = w5319 ^ w5354 ;
  assign w5356 = w4939 ^ w5318 ;
  assign w5357 = w4941 ^ w5356 ;
  assign w5358 = w592 & ~w4143 ;
  assign w5359 = w721 & w4052 ;
  assign w5360 = ( w592 & ~w5358 ) | ( w592 & w5359 ) | ( ~w5358 & w5359 ) ;
  assign w5361 = w3435 | w4147 ;
  assign w5362 = w381 & ~w5360 ;
  assign w5363 = ( w3964 & w5360 ) | ( w3964 & ~w5362 ) | ( w5360 & ~w5362 ) ;
  assign w5364 = ( ~w3435 & w5361 ) | ( ~w3435 & w5363 ) | ( w5361 & w5363 ) ;
  assign w5365 = \pi26 ^ w5364 ;
  assign w5366 = w883 | w4052 ;
  assign w5367 = w721 & w4143 ;
  assign w5368 = ( ~w883 & w5366 ) | ( ~w883 & w5367 ) | ( w5366 & w5367 ) ;
  assign w5369 = w3421 & ~w4147 ;
  assign w5370 = w592 | w5368 ;
  assign w5371 = ( w3964 & w5368 ) | ( w3964 & w5370 ) | ( w5368 & w5370 ) ;
  assign w5372 = ( w3421 & ~w5369 ) | ( w3421 & w5371 ) | ( ~w5369 & w5371 ) ;
  assign w5373 = \pi26 ^ w5372 ;
  assign w5374 = w4943 ^ w5317 ;
  assign w5375 = w5079 ^ w5374 ;
  assign w5376 = w1085 & ~w3717 ;
  assign w5377 = w1205 & w3649 ;
  assign w5378 = ( w1085 & ~w5376 ) | ( w1085 & w5377 ) | ( ~w5376 & w5377 ) ;
  assign w5379 = w979 & ~w3549 ;
  assign w5380 = w4666 | w5378 ;
  assign w5381 = ( w3448 & w5378 ) | ( w3448 & w5380 ) | ( w5378 & w5380 ) ;
  assign w5382 = ( w979 & ~w5379 ) | ( w979 & w5381 ) | ( ~w5379 & w5381 ) ;
  assign w5383 = \pi29 ^ w5382 ;
  assign w5384 = ( w5373 & w5375 ) | ( w5373 & w5383 ) | ( w5375 & w5383 ) ;
  assign w5385 = ( ~w5357 & w5365 ) | ( ~w5357 & w5384 ) | ( w5365 & w5384 ) ;
  assign w5386 = w3647 & ~w4606 ;
  assign w5387 = w3715 & w4651 ;
  assign w5388 = ( w3647 & ~w5386 ) | ( w3647 & w5387 ) | ( ~w5386 & w5387 ) ;
  assign w5389 = w3548 | w4706 ;
  assign w5390 = w3725 & ~w5388 ;
  assign w5391 = ( w4609 & w5388 ) | ( w4609 & ~w5390 ) | ( w5388 & ~w5390 ) ;
  assign w5392 = ( ~w3548 & w5389 ) | ( ~w3548 & w5391 ) | ( w5389 & w5391 ) ;
  assign w5393 = \pi23 ^ w5392 ;
  assign w5394 = ( w5355 & w5385 ) | ( w5355 & w5393 ) | ( w5385 & w5393 ) ;
  assign w5395 = ~w4906 & w4907 ;
  assign w5396 = w4049 | w4905 ;
  assign w5397 = ~w4142 & w5343 ;
  assign w5398 = ( ~w4049 & w5396 ) | ( ~w4049 & w5397 ) | ( w5396 & w5397 ) ;
  assign w5399 = w3962 | w5395 ;
  assign w5400 = w4152 & ~w5398 ;
  assign w5401 = ( w4908 & w5398 ) | ( w4908 & ~w5400 ) | ( w5398 & ~w5400 ) ;
  assign w5402 = ( ~w3962 & w5399 ) | ( ~w3962 & w5401 ) | ( w5399 & w5401 ) ;
  assign w5403 = \pi20 ^ w5402 ;
  assign w5404 = ( ~w5353 & w5394 ) | ( ~w5353 & w5403 ) | ( w5394 & w5403 ) ;
  assign w5405 = ~w4142 & w4905 ;
  assign w5406 = ( ~w4600 & w5395 ) | ( ~w4600 & w5405 ) | ( w5395 & w5405 ) ;
  assign w5407 = w5343 | w5406 ;
  assign w5408 = ( ~w3962 & w5406 ) | ( ~w3962 & w5407 ) | ( w5406 & w5407 ) ;
  assign w5409 = w5405 | w5408 ;
  assign w5410 = w4927 ^ w5339 ;
  assign w5411 = w4929 ^ w5410 ;
  assign w5412 = w4722 & ~w5409 ;
  assign w5413 = ( w4908 & w5409 ) | ( w4908 & ~w5412 ) | ( w5409 & ~w5412 ) ;
  assign w5414 = \pi20 ^ w5413 ;
  assign w5415 = ( w5404 & w5411 ) | ( w5404 & w5414 ) | ( w5411 & w5414 ) ;
  assign w5416 = w5355 ^ w5393 ;
  assign w5417 = w5385 ^ w5416 ;
  assign w5418 = w3647 & ~w4651 ;
  assign w5419 = ~w3094 & w4606 ;
  assign w5420 = ( w3647 & ~w5418 ) | ( w3647 & w5419 ) | ( ~w5418 & w5419 ) ;
  assign w5421 = w3715 & ~w4706 ;
  assign w5422 = w4164 & ~w5420 ;
  assign w5423 = ( w4609 & w5420 ) | ( w4609 & ~w5422 ) | ( w5420 & ~w5422 ) ;
  assign w5424 = ( w3715 & ~w5421 ) | ( w3715 & w5423 ) | ( ~w5421 & w5423 ) ;
  assign w5425 = \pi23 ^ w5424 ;
  assign w5426 = w5365 ^ w5384 ;
  assign w5427 = w5357 ^ w5426 ;
  assign w5428 = w5373 ^ w5375 ;
  assign w5429 = w5383 ^ w5428 ;
  assign w5430 = w5118 ^ w5306 ;
  assign w5431 = w5004 ^ w5430 ;
  assign w5432 = w1614 ^ w2988 ;
  assign w5433 = w1711 ^ w5432 ;
  assign w5434 = w37 | w5433 ;
  assign w5435 = ~w1834 & w3098 ;
  assign w5436 = ( ~w5433 & w5434 ) | ( ~w5433 & w5435 ) | ( w5434 & w5435 ) ;
  assign w5437 = ( \pi29 & \pi30 ) | ( \pi29 & w1614 ) | ( \pi30 & w1614 ) ;
  assign w5438 = \pi31 | w5437 ;
  assign w5439 = ( \pi29 & ~\pi30 ) | ( \pi29 & w1711 ) | ( ~\pi30 & w1711 ) ;
  assign w5440 = ( \pi29 & \pi31 ) | ( \pi29 & ~w5439 ) | ( \pi31 & ~w5439 ) ;
  assign w5441 = ( w5436 & w5438 ) | ( w5436 & ~w5440 ) | ( w5438 & ~w5440 ) ;
  assign w5442 = w1399 & ~w3717 ;
  assign w5443 = ~w1510 & w3649 ;
  assign w5444 = ( w1399 & ~w5442 ) | ( w1399 & w5443 ) | ( ~w5442 & w5443 ) ;
  assign w5445 = w1264 | w3549 ;
  assign w5446 = w4852 & ~w5444 ;
  assign w5447 = ( w3448 & w5444 ) | ( w3448 & ~w5446 ) | ( w5444 & ~w5446 ) ;
  assign w5448 = ( ~w1264 & w5445 ) | ( ~w1264 & w5447 ) | ( w5445 & w5447 ) ;
  assign w5449 = \pi29 ^ w5448 ;
  assign w5450 = ( w5431 & w5441 ) | ( w5431 & w5449 ) | ( w5441 & w5449 ) ;
  assign w5451 = w5093 ^ w5307 ;
  assign w5452 = w5083 ^ w5451 ;
  assign w5453 = w1264 | w3717 ;
  assign w5454 = w1399 & w3649 ;
  assign w5455 = ( ~w1264 & w5453 ) | ( ~w1264 & w5454 ) | ( w5453 & w5454 ) ;
  assign w5456 = w1205 & ~w3549 ;
  assign w5457 = w4864 & ~w5455 ;
  assign w5458 = ( w3448 & w5455 ) | ( w3448 & ~w5457 ) | ( w5455 & ~w5457 ) ;
  assign w5459 = ( w1205 & ~w5456 ) | ( w1205 & w5458 ) | ( ~w5456 & w5458 ) ;
  assign w5460 = \pi29 ^ w5459 ;
  assign w5461 = ( w5450 & w5452 ) | ( w5450 & w5460 ) | ( w5452 & w5460 ) ;
  assign w5462 = w5081 ^ w5316 ;
  assign w5463 = w5308 ^ w5462 ;
  assign w5464 = w883 | w4143 ;
  assign w5465 = w979 & w4052 ;
  assign w5466 = ( ~w883 & w5464 ) | ( ~w883 & w5465 ) | ( w5464 & w5465 ) ;
  assign w5467 = w4147 | w4257 ;
  assign w5468 = w721 | w5466 ;
  assign w5469 = ( w3964 & w5466 ) | ( w3964 & w5468 ) | ( w5466 & w5468 ) ;
  assign w5470 = ( ~w4257 & w5467 ) | ( ~w4257 & w5469 ) | ( w5467 & w5469 ) ;
  assign w5471 = \pi26 ^ w5470 ;
  assign w5472 = ( w5461 & w5463 ) | ( w5461 & w5471 ) | ( w5463 & w5471 ) ;
  assign w5473 = w381 | w4606 ;
  assign w5474 = ~w3094 & w4651 ;
  assign w5475 = ( ~w381 & w5473 ) | ( ~w381 & w5474 ) | ( w5473 & w5474 ) ;
  assign w5476 = w3647 & ~w4706 ;
  assign w5477 = w3810 | w5475 ;
  assign w5478 = ( w4609 & w5475 ) | ( w4609 & w5477 ) | ( w5475 & w5477 ) ;
  assign w5479 = ( w3647 & ~w5476 ) | ( w3647 & w5478 ) | ( ~w5476 & w5478 ) ;
  assign w5480 = \pi23 ^ w5479 ;
  assign w5481 = ( w5429 & w5472 ) | ( w5429 & w5480 ) | ( w5472 & w5480 ) ;
  assign w5482 = ( w5425 & ~w5427 ) | ( w5425 & w5481 ) | ( ~w5427 & w5481 ) ;
  assign w5483 = w4049 | w5343 ;
  assign w5484 = w3907 & w4905 ;
  assign w5485 = ( ~w4049 & w5483 ) | ( ~w4049 & w5484 ) | ( w5483 & w5484 ) ;
  assign w5486 = w4142 | w5395 ;
  assign w5487 = w4563 | w5485 ;
  assign w5488 = ( w4908 & w5485 ) | ( w4908 & w5487 ) | ( w5485 & w5487 ) ;
  assign w5489 = ( ~w4142 & w5486 ) | ( ~w4142 & w5488 ) | ( w5486 & w5488 ) ;
  assign w5490 = \pi20 ^ w5489 ;
  assign w5491 = ( w5417 & w5482 ) | ( w5417 & w5490 ) | ( w5482 & w5490 ) ;
  assign w5492 = ( \pi15 & ~\pi16 ) | ( \pi15 & \pi17 ) | ( ~\pi16 & \pi17 ) ;
  assign w5493 = ( \pi14 & \pi15 ) | ( \pi14 & w5492 ) | ( \pi15 & w5492 ) ;
  assign w5494 = w5492 ^ w5493 ;
  assign w5495 = \pi16 ^ \pi17 ;
  assign w5496 = \pi14 ^ \pi15 ;
  assign w5497 = w5495 & w5496 ;
  assign w5498 = ~w4600 & w5494 ;
  assign w5499 = w5497 | w5498 ;
  assign w5500 = ( ~w4603 & w5498 ) | ( ~w4603 & w5499 ) | ( w5498 & w5499 ) ;
  assign w5501 = \pi17 ^ w5500 ;
  assign w5502 = w5353 ^ w5403 ;
  assign w5503 = w5394 ^ w5502 ;
  assign w5504 = ( w5491 & w5501 ) | ( w5491 & ~w5503 ) | ( w5501 & ~w5503 ) ;
  assign w5505 = w4722 & w4908 ;
  assign w5506 = ( w4908 & w5409 ) | ( w4908 & ~w5505 ) | ( w5409 & ~w5505 ) ;
  assign w5507 = w5404 ^ w5506 ;
  assign w5508 = \pi20 ^ w5411 ;
  assign w5509 = w5507 ^ w5508 ;
  assign w5510 = w5501 ^ w5503 ;
  assign w5511 = w5491 ^ w5510 ;
  assign w5512 = w5417 ^ w5490 ;
  assign w5513 = w5482 ^ w5512 ;
  assign w5514 = w5425 ^ w5481 ;
  assign w5515 = w5427 ^ w5514 ;
  assign w5516 = w3548 | w4905 ;
  assign w5517 = w3907 & w5343 ;
  assign w5518 = ( ~w3548 & w5516 ) | ( ~w3548 & w5517 ) | ( w5516 & w5517 ) ;
  assign w5519 = w4049 | w5395 ;
  assign w5520 = w4622 & ~w5518 ;
  assign w5521 = ( w4908 & w5518 ) | ( w4908 & ~w5520 ) | ( w5518 & ~w5520 ) ;
  assign w5522 = ( ~w4049 & w5519 ) | ( ~w4049 & w5521 ) | ( w5519 & w5521 ) ;
  assign w5523 = \pi20 ^ w5522 ;
  assign w5524 = w5429 ^ w5480 ;
  assign w5525 = w5472 ^ w5524 ;
  assign w5526 = w5463 ^ w5471 ;
  assign w5527 = w5461 ^ w5526 ;
  assign w5528 = w5450 ^ w5460 ;
  assign w5529 = w5452 ^ w5528 ;
  assign w5530 = w979 & ~w4143 ;
  assign w5531 = w1085 & w4052 ;
  assign w5532 = ( w979 & ~w5530 ) | ( w979 & w5531 ) | ( ~w5530 & w5531 ) ;
  assign w5533 = w4147 | w4273 ;
  assign w5534 = w883 & ~w5532 ;
  assign w5535 = ( w3964 & w5532 ) | ( w3964 & ~w5534 ) | ( w5532 & ~w5534 ) ;
  assign w5536 = ( ~w4273 & w5533 ) | ( ~w4273 & w5535 ) | ( w5533 & w5535 ) ;
  assign w5537 = \pi26 ^ w5536 ;
  assign w5538 = w5431 ^ w5449 ;
  assign w5539 = w5441 ^ w5538 ;
  assign w5540 = w5294 ^ w5305 ;
  assign w5541 = w5004 ^ w5540 ;
  assign w5542 = w5218 ^ w5293 ;
  assign w5543 = \pi08 ^ w5542 ;
  assign w5544 = w169 | w490 ;
  assign w5545 = ( ~w169 & w278 ) | ( ~w169 & w532 ) | ( w278 & w532 ) ;
  assign w5546 = w5544 | w5545 ;
  assign w5547 = w492 | w1030 ;
  assign w5548 = w1413 | w5547 ;
  assign w5549 = ( ~w1413 & w3693 ) | ( ~w1413 & w5546 ) | ( w3693 & w5546 ) ;
  assign w5550 = w5548 | w5549 ;
  assign w5551 = w495 | w817 ;
  assign w5552 = w136 | w5551 ;
  assign w5553 = ( ~w136 & w309 ) | ( ~w136 & w5550 ) | ( w309 & w5550 ) ;
  assign w5554 = w5552 | w5553 ;
  assign w5555 = w466 | w997 ;
  assign w5556 = ( ~w997 & w1616 ) | ( ~w997 & w5554 ) | ( w1616 & w5554 ) ;
  assign w5557 = w5555 | w5556 ;
  assign w5558 = ( w534 & w662 ) | ( w534 & ~w899 ) | ( w662 & ~w899 ) ;
  assign w5559 = w443 | w5557 ;
  assign w5560 = ( ~w443 & w899 ) | ( ~w443 & w1229 ) | ( w899 & w1229 ) ;
  assign w5561 = w5559 | w5560 ;
  assign w5562 = w5558 | w5561 ;
  assign w5563 = ( w271 & w351 ) | ( w271 & ~w447 ) | ( w351 & ~w447 ) ;
  assign w5564 = w269 | w5235 ;
  assign w5565 = ( ~w269 & w447 ) | ( ~w269 & w664 ) | ( w447 & w664 ) ;
  assign w5566 = w5564 | w5565 ;
  assign w5567 = w5563 | w5566 ;
  assign w5568 = w5198 | w5567 ;
  assign w5569 = w5562 | w5568 ;
  assign w5570 = ( w836 & w3299 ) | ( w836 & ~w5562 ) | ( w3299 & ~w5562 ) ;
  assign w5571 = w5569 | w5570 ;
  assign w5572 = w572 | w2200 ;
  assign w5573 = ( ~w572 & w2760 ) | ( ~w572 & w5571 ) | ( w2760 & w5571 ) ;
  assign w5574 = w5572 | w5573 ;
  assign w5575 = ( w149 & w341 ) | ( w149 & ~w344 ) | ( w341 & ~w344 ) ;
  assign w5576 = w81 | w5574 ;
  assign w5577 = ( ~w81 & w344 ) | ( ~w81 & w567 ) | ( w344 & w567 ) ;
  assign w5578 = w5576 | w5577 ;
  assign w5579 = w5575 | w5578 ;
  assign w5580 = w144 | w605 ;
  assign w5581 = ( ~w144 & w265 ) | ( ~w144 & w5579 ) | ( w265 & w5579 ) ;
  assign w5582 = w5580 | w5581 ;
  assign w5583 = ( w268 & w316 ) | ( w268 & ~w504 ) | ( w316 & ~w504 ) ;
  assign w5584 = w125 | w214 ;
  assign w5585 = ( ~w214 & w504 ) | ( ~w214 & w821 ) | ( w504 & w821 ) ;
  assign w5586 = w5584 | w5585 ;
  assign w5587 = w5583 | w5586 ;
  assign w5588 = w179 | w673 ;
  assign w5589 = ( ~w179 & w534 ) | ( ~w179 & w5587 ) | ( w534 & w5587 ) ;
  assign w5590 = w5588 | w5589 ;
  assign w5591 = ( w178 & ~w263 ) | ( w178 & w312 ) | ( ~w263 & w312 ) ;
  assign w5592 = w263 | w5591 ;
  assign w5593 = ( w139 & w220 ) | ( w139 & ~w351 ) | ( w220 & ~w351 ) ;
  assign w5594 = w95 | w5592 ;
  assign w5595 = ( ~w95 & w351 ) | ( ~w95 & w424 ) | ( w351 & w424 ) ;
  assign w5596 = w5594 | w5595 ;
  assign w5597 = w5593 | w5596 ;
  assign w5598 = ( w128 & w269 ) | ( w128 & ~w899 ) | ( w269 & ~w899 ) ;
  assign w5599 = w51 | w5597 ;
  assign w5600 = ( ~w51 & w899 ) | ( ~w51 & w980 ) | ( w899 & w980 ) ;
  assign w5601 = w5599 | w5600 ;
  assign w5602 = w5598 | w5601 ;
  assign w5603 = ( w350 & w445 ) | ( w350 & ~w511 ) | ( w445 & ~w511 ) ;
  assign w5604 = w104 | w257 ;
  assign w5605 = ( ~w257 & w511 ) | ( ~w257 & w951 ) | ( w511 & w951 ) ;
  assign w5606 = w5604 | w5605 ;
  assign w5607 = w5603 | w5606 ;
  assign w5608 = w205 | w5607 ;
  assign w5609 = w120 | w606 ;
  assign w5610 = ( ~w120 & w163 ) | ( ~w120 & w5608 ) | ( w163 & w5608 ) ;
  assign w5611 = w5609 | w5610 ;
  assign w5612 = w204 | w1265 ;
  assign w5613 = w5611 | w5612 ;
  assign w5614 = ( w64 & w5602 ) | ( w64 & ~w5611 ) | ( w5602 & ~w5611 ) ;
  assign w5615 = w5613 | w5614 ;
  assign w5616 = ( w122 & w506 ) | ( w122 & ~w623 ) | ( w506 & ~w623 ) ;
  assign w5617 = w88 | w5615 ;
  assign w5618 = ( ~w88 & w623 ) | ( ~w88 & w626 ) | ( w623 & w626 ) ;
  assign w5619 = w5617 | w5618 ;
  assign w5620 = w5616 | w5619 ;
  assign w5621 = w525 | w1153 ;
  assign w5622 = w113 | w5621 ;
  assign w5623 = ( ~w113 & w492 ) | ( ~w113 & w5620 ) | ( w492 & w5620 ) ;
  assign w5624 = w5622 | w5623 ;
  assign w5625 = ( w198 & ~w314 ) | ( w198 & w443 ) | ( ~w314 & w443 ) ;
  assign w5626 = w314 | w5625 ;
  assign w5627 = w622 | w5626 ;
  assign w5628 = w5624 | w5627 ;
  assign w5629 = ( w3071 & w4489 ) | ( w3071 & ~w5624 ) | ( w4489 & ~w5624 ) ;
  assign w5630 = w5628 | w5629 ;
  assign w5631 = ( w517 & ~w2782 ) | ( w517 & w5590 ) | ( ~w2782 & w5590 ) ;
  assign w5632 = w3011 | w5630 ;
  assign w5633 = ( w860 & w2782 ) | ( w860 & ~w3011 ) | ( w2782 & ~w3011 ) ;
  assign w5634 = w5632 | w5633 ;
  assign w5635 = w5631 | w5634 ;
  assign w5636 = ( w224 & w315 ) | ( w224 & ~w456 ) | ( w315 & ~w456 ) ;
  assign w5637 = w143 | w5635 ;
  assign w5638 = ( ~w143 & w456 ) | ( ~w143 & w723 ) | ( w456 & w723 ) ;
  assign w5639 = w5637 | w5638 ;
  assign w5640 = w5636 | w5639 ;
  assign w5641 = w44 | w628 ;
  assign w5642 = ( ~w44 & w208 ) | ( ~w44 & w5640 ) | ( w208 & w5640 ) ;
  assign w5643 = w5641 | w5642 ;
  assign w5644 = ( \pi02 & \pi05 ) | ( \pi02 & ~w5643 ) | ( \pi05 & ~w5643 ) ;
  assign w5645 = w2059 ^ w2984 ;
  assign w5646 = w1976 ^ w5645 ;
  assign w5647 = ( \pi30 & \pi31 ) | ( \pi30 & ~w2059 ) | ( \pi31 & ~w2059 ) ;
  assign w5648 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w5647 ) | ( \pi30 & w5647 ) ;
  assign w5649 = ( \pi29 & ~\pi30 ) | ( \pi29 & w5647 ) | ( ~\pi30 & w5647 ) ;
  assign w5650 = ( \pi30 & w2130 ) | ( \pi30 & ~w5649 ) | ( w2130 & ~w5649 ) ;
  assign w5651 = ( w1976 & w5649 ) | ( w1976 & w5650 ) | ( w5649 & w5650 ) ;
  assign w5652 = ~\pi31 & w5651 ;
  assign w5653 = ( w5648 & ~w5650 ) | ( w5648 & w5652 ) | ( ~w5650 & w5652 ) ;
  assign w5654 = ( w37 & w5646 ) | ( w37 & w5653 ) | ( w5646 & w5653 ) ;
  assign w5655 = w5653 | w5654 ;
  assign w5656 = ( w5218 & ~w5644 ) | ( w5218 & w5655 ) | ( ~w5644 & w5655 ) ;
  assign w5657 = ( w5218 & w5582 ) | ( w5218 & w5656 ) | ( w5582 & w5656 ) ;
  assign w5658 = w1939 ^ w2986 ;
  assign w5659 = w1834 ^ w5658 ;
  assign w5660 = ( \pi30 & \pi31 ) | ( \pi30 & ~w1939 ) | ( \pi31 & ~w1939 ) ;
  assign w5661 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w5660 ) | ( \pi30 & w5660 ) ;
  assign w5662 = ( \pi29 & ~\pi30 ) | ( \pi29 & w5660 ) | ( ~\pi30 & w5660 ) ;
  assign w5663 = ( ~\pi30 & w1976 ) | ( ~\pi30 & w5662 ) | ( w1976 & w5662 ) ;
  assign w5664 = ( w1834 & ~w5662 ) | ( w1834 & w5663 ) | ( ~w5662 & w5663 ) ;
  assign w5665 = \pi31 | w5664 ;
  assign w5666 = ( w5661 & w5663 ) | ( w5661 & ~w5665 ) | ( w5663 & ~w5665 ) ;
  assign w5667 = ( w37 & ~w5659 ) | ( w37 & w5666 ) | ( ~w5659 & w5666 ) ;
  assign w5668 = w5666 | w5667 ;
  assign w5669 = ( w5543 & w5657 ) | ( w5543 & w5668 ) | ( w5657 & w5668 ) ;
  assign w5670 = w1614 & ~w3649 ;
  assign w5671 = ~w1510 & w3717 ;
  assign w5672 = ( w1614 & ~w5670 ) | ( w1614 & w5671 ) | ( ~w5670 & w5671 ) ;
  assign w5673 = w1399 & ~w3549 ;
  assign w5674 = w5069 & ~w5672 ;
  assign w5675 = ( w3448 & w5672 ) | ( w3448 & ~w5674 ) | ( w5672 & ~w5674 ) ;
  assign w5676 = ( w1399 & ~w5673 ) | ( w1399 & w5675 ) | ( ~w5673 & w5675 ) ;
  assign w5677 = \pi29 ^ w5676 ;
  assign w5678 = ( w5541 & w5669 ) | ( w5541 & w5677 ) | ( w5669 & w5677 ) ;
  assign w5679 = w1085 & ~w4143 ;
  assign w5680 = w1205 & w4052 ;
  assign w5681 = ( w1085 & ~w5679 ) | ( w1085 & w5680 ) | ( ~w5679 & w5680 ) ;
  assign w5682 = ~w4147 & w4666 ;
  assign w5683 = w979 | w5681 ;
  assign w5684 = ( w3964 & w5681 ) | ( w3964 & w5683 ) | ( w5681 & w5683 ) ;
  assign w5685 = ( w4666 & ~w5682 ) | ( w4666 & w5684 ) | ( ~w5682 & w5684 ) ;
  assign w5686 = \pi26 ^ w5685 ;
  assign w5687 = ( w5539 & w5678 ) | ( w5539 & w5686 ) | ( w5678 & w5686 ) ;
  assign w5688 = ( w5529 & w5537 ) | ( w5529 & w5687 ) | ( w5537 & w5687 ) ;
  assign w5689 = w381 | w4651 ;
  assign w5690 = w592 & w4606 ;
  assign w5691 = ( ~w381 & w5689 ) | ( ~w381 & w5690 ) | ( w5689 & w5690 ) ;
  assign w5692 = w3094 | w4706 ;
  assign w5693 = w3096 | w5691 ;
  assign w5694 = ( w4609 & w5691 ) | ( w4609 & w5693 ) | ( w5691 & w5693 ) ;
  assign w5695 = ( ~w3094 & w5692 ) | ( ~w3094 & w5694 ) | ( w5692 & w5694 ) ;
  assign w5696 = \pi23 ^ w5695 ;
  assign w5697 = ( w5527 & w5688 ) | ( w5527 & w5696 ) | ( w5688 & w5696 ) ;
  assign w5698 = w3548 | w5343 ;
  assign w5699 = w3715 & w4905 ;
  assign w5700 = ( ~w3548 & w5698 ) | ( ~w3548 & w5699 ) | ( w5698 & w5699 ) ;
  assign w5701 = w3907 & ~w5395 ;
  assign w5702 = w3913 & ~w5700 ;
  assign w5703 = ( w4908 & w5700 ) | ( w4908 & ~w5702 ) | ( w5700 & ~w5702 ) ;
  assign w5704 = ( w3907 & ~w5701 ) | ( w3907 & w5703 ) | ( ~w5701 & w5703 ) ;
  assign w5705 = \pi20 ^ w5704 ;
  assign w5706 = ( w5525 & w5697 ) | ( w5525 & w5705 ) | ( w5697 & w5705 ) ;
  assign w5707 = ( ~w5515 & w5523 ) | ( ~w5515 & w5706 ) | ( w5523 & w5706 ) ;
  assign w5708 = w5513 ^ w5707 ;
  assign w5709 = ( \pi14 & \pi15 ) | ( \pi14 & \pi16 ) | ( \pi15 & \pi16 ) ;
  assign w5710 = \pi16 ^ w5709 ;
  assign w5711 = ~w4600 & w5710 ;
  assign w5712 = ( ~w3962 & w5494 ) | ( ~w3962 & w5711 ) | ( w5494 & w5711 ) ;
  assign w5713 = ( ~w3962 & w4601 ) | ( ~w3962 & w5712 ) | ( w4601 & w5712 ) ;
  assign w5714 = ( w4600 & w4601 ) | ( w4600 & w5497 ) | ( w4601 & w5497 ) ;
  assign w5715 = ( w5711 & ~w5713 ) | ( w5711 & w5714 ) | ( ~w5713 & w5714 ) ;
  assign w5716 = ( ~w4657 & w5712 ) | ( ~w4657 & w5715 ) | ( w5712 & w5715 ) ;
  assign w5717 = \pi17 ^ w5716 ;
  assign w5718 = ( w5513 & w5707 ) | ( w5513 & w5717 ) | ( w5707 & w5717 ) ;
  assign w5719 = w5525 ^ w5705 ;
  assign w5720 = w5697 ^ w5719 ;
  assign w5721 = w5527 ^ w5696 ;
  assign w5722 = w5688 ^ w5721 ;
  assign w5723 = w592 & ~w4651 ;
  assign w5724 = w721 & w4606 ;
  assign w5725 = ( w592 & ~w5723 ) | ( w592 & w5724 ) | ( ~w5723 & w5724 ) ;
  assign w5726 = w381 | w4706 ;
  assign w5727 = w3435 & ~w5725 ;
  assign w5728 = ( w4609 & w5725 ) | ( w4609 & ~w5727 ) | ( w5725 & ~w5727 ) ;
  assign w5729 = ( ~w381 & w5726 ) | ( ~w381 & w5728 ) | ( w5726 & w5728 ) ;
  assign w5730 = \pi23 ^ w5729 ;
  assign w5731 = w5537 ^ w5687 ;
  assign w5732 = w5529 ^ w5731 ;
  assign w5733 = w5539 ^ w5686 ;
  assign w5734 = w5678 ^ w5733 ;
  assign w5735 = w1614 & ~w3717 ;
  assign w5736 = w1711 & w3649 ;
  assign w5737 = ( w1614 & ~w5735 ) | ( w1614 & w5736 ) | ( ~w5735 & w5736 ) ;
  assign w5738 = w1510 | w3549 ;
  assign w5739 = w5085 & ~w5737 ;
  assign w5740 = ( w3448 & w5737 ) | ( w3448 & ~w5739 ) | ( w5737 & ~w5739 ) ;
  assign w5741 = ( ~w1510 & w5738 ) | ( ~w1510 & w5740 ) | ( w5738 & w5740 ) ;
  assign w5742 = \pi29 ^ w5741 ;
  assign w5743 = w5657 ^ w5668 ;
  assign w5744 = w5543 ^ w5743 ;
  assign w5745 = w5582 ^ w5656 ;
  assign w5746 = w5218 ^ w5745 ;
  assign w5747 = w1939 ^ w2985 ;
  assign w5748 = w1976 ^ w5747 ;
  assign w5749 = ~w37 & w5748 ;
  assign w5750 = ~w2059 & w3098 ;
  assign w5751 = ( w5748 & ~w5749 ) | ( w5748 & w5750 ) | ( ~w5749 & w5750 ) ;
  assign w5752 = ( \pi29 & \pi30 ) | ( \pi29 & ~w1939 ) | ( \pi30 & ~w1939 ) ;
  assign w5753 = \pi31 | w5752 ;
  assign w5754 = ( \pi29 & ~\pi30 ) | ( \pi29 & w1976 ) | ( ~\pi30 & w1976 ) ;
  assign w5755 = ( \pi29 & \pi31 ) | ( \pi29 & ~w5754 ) | ( \pi31 & ~w5754 ) ;
  assign w5756 = ( w5751 & w5753 ) | ( w5751 & ~w5755 ) | ( w5753 & ~w5755 ) ;
  assign w5757 = w5644 ^ w5655 ;
  assign w5758 = w5218 ^ w5757 ;
  assign w5759 = w164 | w626 ;
  assign w5760 = ( w122 & ~w164 ) | ( w122 & w271 ) | ( ~w164 & w271 ) ;
  assign w5761 = w5759 | w5760 ;
  assign w5762 = ( ~w339 & w384 ) | ( ~w339 & w5761 ) | ( w384 & w5761 ) ;
  assign w5763 = w3523 | w5762 ;
  assign w5764 = ( w218 & w277 ) | ( w218 & ~w637 ) | ( w277 & ~w637 ) ;
  assign w5765 = w59 | w147 ;
  assign w5766 = ( ~w147 & w637 ) | ( ~w147 & w673 ) | ( w637 & w673 ) ;
  assign w5767 = w5765 | w5766 ;
  assign w5768 = w5764 | w5767 ;
  assign w5769 = ( w314 & w463 ) | ( w314 & ~w724 ) | ( w463 & ~w724 ) ;
  assign w5770 = w252 | w5768 ;
  assign w5771 = ( ~w252 & w724 ) | ( ~w252 & w1130 ) | ( w724 & w1130 ) ;
  assign w5772 = w5770 | w5771 ;
  assign w5773 = w5769 | w5772 ;
  assign w5774 = ( w139 & w210 ) | ( w139 & ~w229 ) | ( w210 & ~w229 ) ;
  assign w5775 = w1363 | w5007 ;
  assign w5776 = ( w229 & w725 ) | ( w229 & ~w5007 ) | ( w725 & ~w5007 ) ;
  assign w5777 = w5775 | w5776 ;
  assign w5778 = w5774 | w5777 ;
  assign w5779 = ( w3690 & w5773 ) | ( w3690 & ~w5778 ) | ( w5773 & ~w5778 ) ;
  assign w5780 = ~w2208 & w2552 ;
  assign w5781 = ( w1108 & w2552 ) | ( w1108 & w5778 ) | ( w2552 & w5778 ) ;
  assign w5782 = w5780 & ~w5781 ;
  assign w5783 = ~w5779 & w5782 ;
  assign w5784 = w1051 | w4784 ;
  assign w5785 = w5763 | w5784 ;
  assign w5786 = ( ~w624 & w5763 ) | ( ~w624 & w5783 ) | ( w5763 & w5783 ) ;
  assign w5787 = ~w5785 & w5786 ;
  assign w5788 = w221 | w516 ;
  assign w5789 = w44 | w5788 ;
  assign w5790 = ( w44 & ~w95 ) | ( w44 & w5787 ) | ( ~w95 & w5787 ) ;
  assign w5791 = ~w5789 & w5790 ;
  assign w5792 = ( w463 & w491 ) | ( w463 & ~w1030 ) | ( w491 & ~w1030 ) ;
  assign w5793 = w210 | w413 ;
  assign w5794 = ( ~w413 & w1030 ) | ( ~w413 & w1086 ) | ( w1030 & w1086 ) ;
  assign w5795 = w5793 | w5794 ;
  assign w5796 = w5792 | w5795 ;
  assign w5797 = ( w390 & w408 ) | ( w390 & ~w409 ) | ( w408 & ~w409 ) ;
  assign w5798 = w167 | w5796 ;
  assign w5799 = ( ~w167 & w409 ) | ( ~w167 & w567 ) | ( w409 & w567 ) ;
  assign w5800 = w5798 | w5799 ;
  assign w5801 = w5797 | w5800 ;
  assign w5802 = w221 | w724 ;
  assign w5803 = ( ~w221 & w419 ) | ( ~w221 & w5801 ) | ( w419 & w5801 ) ;
  assign w5804 = w5802 | w5803 ;
  assign w5805 = w203 | w697 ;
  assign w5806 = w144 | w5805 ;
  assign w5807 = ( ~w144 & w164 ) | ( ~w144 & w624 ) | ( w164 & w624 ) ;
  assign w5808 = w5806 | w5807 ;
  assign w5809 = ( w177 & w178 ) | ( w177 & ~w496 ) | ( w178 & ~w496 ) ;
  assign w5810 = w307 | w5808 ;
  assign w5811 = ( w496 & w899 ) | ( w496 & ~w5808 ) | ( w899 & ~w5808 ) ;
  assign w5812 = w5810 | w5811 ;
  assign w5813 = w5809 | w5812 ;
  assign w5814 = w3037 | w5804 ;
  assign w5815 = w5813 | w5814 ;
  assign w5816 = ( w2750 & w4358 ) | ( w2750 & ~w5813 ) | ( w4358 & ~w5813 ) ;
  assign w5817 = w5815 | w5816 ;
  assign w5818 = w416 | w609 ;
  assign w5819 = ( ~w416 & w450 ) | ( ~w416 & w5817 ) | ( w450 & w5817 ) ;
  assign w5820 = w5818 | w5819 ;
  assign w5821 = ( w118 & w224 ) | ( w118 & ~w530 ) | ( w224 & ~w530 ) ;
  assign w5822 = w742 | w5820 ;
  assign w5823 = ( w530 & ~w742 ) | ( w530 & w1340 ) | ( ~w742 & w1340 ) ;
  assign w5824 = w5822 | w5823 ;
  assign w5825 = w5821 | w5824 ;
  assign w5826 = w802 | w901 ;
  assign w5827 = w443 | w5826 ;
  assign w5828 = ( ~w443 & w595 ) | ( ~w443 & w5825 ) | ( w595 & w5825 ) ;
  assign w5829 = w5827 | w5828 ;
  assign w5830 = w218 | w787 ;
  assign w5831 = w164 | w5830 ;
  assign w5832 = ( ~w164 & w205 ) | ( ~w164 & w1461 ) | ( w205 & w1461 ) ;
  assign w5833 = w5831 | w5832 ;
  assign w5834 = w640 | w1030 ;
  assign w5835 = w98 | w5834 ;
  assign w5836 = ( ~w98 & w286 ) | ( ~w98 & w5833 ) | ( w286 & w5833 ) ;
  assign w5837 = w5835 | w5836 ;
  assign w5838 = w219 | w1229 ;
  assign w5839 = ( ~w219 & w223 ) | ( ~w219 & w5099 ) | ( w223 & w5099 ) ;
  assign w5840 = w5838 | w5839 ;
  assign w5841 = w277 | w385 ;
  assign w5842 = w5142 | w5841 ;
  assign w5843 = ( w1473 & ~w5142 ) | ( w1473 & w5840 ) | ( ~w5142 & w5840 ) ;
  assign w5844 = w5842 | w5843 ;
  assign w5845 = ( ~w149 & w999 ) | ( ~w149 & w1051 ) | ( w999 & w1051 ) ;
  assign w5846 = w450 | w5844 ;
  assign w5847 = ( w149 & w214 ) | ( w149 & ~w450 ) | ( w214 & ~w450 ) ;
  assign w5848 = w5846 | w5847 ;
  assign w5849 = w5845 | w5848 ;
  assign w5850 = ( w203 & w257 ) | ( w203 & ~w445 ) | ( w257 & ~w445 ) ;
  assign w5851 = w201 | w5849 ;
  assign w5852 = ( ~w201 & w445 ) | ( ~w201 & w764 ) | ( w445 & w764 ) ;
  assign w5853 = w5851 | w5852 ;
  assign w5854 = w5850 | w5853 ;
  assign w5855 = ( w470 & w697 ) | ( w470 & ~w724 ) | ( w697 & ~w724 ) ;
  assign w5856 = w180 | w594 ;
  assign w5857 = ( ~w180 & w724 ) | ( ~w180 & w1094 ) | ( w724 & w1094 ) ;
  assign w5858 = w5856 | w5857 ;
  assign w5859 = w5855 | w5858 ;
  assign w5860 = w608 | w4464 ;
  assign w5861 = ( w76 & w4352 ) | ( w76 & ~w4464 ) | ( w4352 & ~w4464 ) ;
  assign w5862 = w5860 | w5861 ;
  assign w5863 = ( w74 & w101 ) | ( w74 & ~w309 ) | ( w101 & ~w309 ) ;
  assign w5864 = w5859 | w5862 ;
  assign w5865 = ( w309 & w567 ) | ( w309 & ~w5862 ) | ( w567 & ~w5862 ) ;
  assign w5866 = w5864 | w5865 ;
  assign w5867 = w5863 | w5866 ;
  assign w5868 = ( ~w315 & w5837 ) | ( ~w315 & w5867 ) | ( w5837 & w5867 ) ;
  assign w5869 = w2886 | w5854 ;
  assign w5870 = ( w315 & w316 ) | ( w315 & ~w2886 ) | ( w316 & ~w2886 ) ;
  assign w5871 = w5869 | w5870 ;
  assign w5872 = w5868 | w5871 ;
  assign w5873 = w176 | w1324 ;
  assign w5874 = ( ~w1324 & w4784 ) | ( ~w1324 & w5872 ) | ( w4784 & w5872 ) ;
  assign w5875 = w5873 | w5874 ;
  assign w5876 = w488 | w901 ;
  assign w5877 = ( ~w488 & w568 ) | ( ~w488 & w5875 ) | ( w568 & w5875 ) ;
  assign w5878 = w5876 | w5877 ;
  assign w5879 = w2273 ^ w2980 ;
  assign w5880 = w2391 ^ w5879 ;
  assign w5881 = ( \pi29 & \pi31 ) | ( \pi29 & w2391 ) | ( \pi31 & w2391 ) ;
  assign w5882 = ( \pi29 & ~\pi30 ) | ( \pi29 & w5881 ) | ( ~\pi30 & w5881 ) ;
  assign w5883 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w5881 ) | ( \pi30 & w5881 ) ;
  assign w5884 = ( ~\pi29 & w2500 ) | ( ~\pi29 & w5883 ) | ( w2500 & w5883 ) ;
  assign w5885 = ( w2273 & w5883 ) | ( w2273 & ~w5884 ) | ( w5883 & ~w5884 ) ;
  assign w5886 = ~\pi31 & w5885 ;
  assign w5887 = ( w5882 & w5884 ) | ( w5882 & w5886 ) | ( w5884 & w5886 ) ;
  assign w5888 = ( w37 & w5880 ) | ( w37 & w5887 ) | ( w5880 & w5887 ) ;
  assign w5889 = w5887 | w5888 ;
  assign w5890 = ( \pi02 & w5878 ) | ( \pi02 & w5889 ) | ( w5878 & w5889 ) ;
  assign w5891 = ( \pi02 & w5829 ) | ( \pi02 & w5890 ) | ( w5829 & w5890 ) ;
  assign w5892 = ( \pi02 & ~w5791 ) | ( \pi02 & w5891 ) | ( ~w5791 & w5891 ) ;
  assign w5893 = \pi02 ^ w5643 ;
  assign w5894 = \pi05 ^ w5893 ;
  assign w5895 = w2059 ^ w2983 ;
  assign w5896 = w2130 ^ w5895 ;
  assign w5897 = ( \pi29 & \pi31 ) | ( \pi29 & ~w2130 ) | ( \pi31 & ~w2130 ) ;
  assign w5898 = ( \pi29 & ~\pi30 ) | ( \pi29 & w5897 ) | ( ~\pi30 & w5897 ) ;
  assign w5899 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w5897 ) | ( \pi30 & w5897 ) ;
  assign w5900 = ( \pi29 & w2235 ) | ( \pi29 & ~w5899 ) | ( w2235 & ~w5899 ) ;
  assign w5901 = ( ~w2059 & w5899 ) | ( ~w2059 & w5900 ) | ( w5899 & w5900 ) ;
  assign w5902 = ~\pi31 & w5901 ;
  assign w5903 = ( w5898 & ~w5900 ) | ( w5898 & w5902 ) | ( ~w5900 & w5902 ) ;
  assign w5904 = ( w37 & ~w5896 ) | ( w37 & w5903 ) | ( ~w5896 & w5903 ) ;
  assign w5905 = w5903 | w5904 ;
  assign w5906 = ( w5892 & w5894 ) | ( w5892 & w5905 ) | ( w5894 & w5905 ) ;
  assign w5907 = w1939 | w3649 ;
  assign w5908 = ~w1834 & w3717 ;
  assign w5909 = ( ~w1939 & w5907 ) | ( ~w1939 & w5908 ) | ( w5907 & w5908 ) ;
  assign w5910 = w1711 & ~w3549 ;
  assign w5911 = w5296 | w5909 ;
  assign w5912 = ( w3448 & w5909 ) | ( w3448 & w5911 ) | ( w5909 & w5911 ) ;
  assign w5913 = ( w1711 & ~w5910 ) | ( w1711 & w5912 ) | ( ~w5910 & w5912 ) ;
  assign w5914 = \pi29 ^ w5913 ;
  assign w5915 = ( ~w5758 & w5906 ) | ( ~w5758 & w5914 ) | ( w5906 & w5914 ) ;
  assign w5916 = ( w5746 & w5756 ) | ( w5746 & w5915 ) | ( w5756 & w5915 ) ;
  assign w5917 = ( w5742 & w5744 ) | ( w5742 & w5916 ) | ( w5744 & w5916 ) ;
  assign w5918 = w5541 ^ w5677 ;
  assign w5919 = w5669 ^ w5918 ;
  assign w5920 = w1264 | w4052 ;
  assign w5921 = w1205 & w4143 ;
  assign w5922 = ( ~w1264 & w5920 ) | ( ~w1264 & w5921 ) | ( w5920 & w5921 ) ;
  assign w5923 = ~w4147 & w4533 ;
  assign w5924 = w1085 | w5922 ;
  assign w5925 = ( w3964 & w5922 ) | ( w3964 & w5924 ) | ( w5922 & w5924 ) ;
  assign w5926 = ( w4533 & ~w5923 ) | ( w4533 & w5925 ) | ( ~w5923 & w5925 ) ;
  assign w5927 = \pi26 ^ w5926 ;
  assign w5928 = ( w5917 & w5919 ) | ( w5917 & w5927 ) | ( w5919 & w5927 ) ;
  assign w5929 = w883 | w4606 ;
  assign w5930 = w721 & w4651 ;
  assign w5931 = ( ~w883 & w5929 ) | ( ~w883 & w5930 ) | ( w5929 & w5930 ) ;
  assign w5932 = w592 & ~w4706 ;
  assign w5933 = w3421 | w5931 ;
  assign w5934 = ( w4609 & w5931 ) | ( w4609 & w5933 ) | ( w5931 & w5933 ) ;
  assign w5935 = ( w592 & ~w5932 ) | ( w592 & w5934 ) | ( ~w5932 & w5934 ) ;
  assign w5936 = \pi23 ^ w5935 ;
  assign w5937 = ( w5734 & w5928 ) | ( w5734 & w5936 ) | ( w5928 & w5936 ) ;
  assign w5938 = ( w5730 & w5732 ) | ( w5730 & w5937 ) | ( w5732 & w5937 ) ;
  assign w5939 = w3647 & ~w4905 ;
  assign w5940 = w3715 & w5343 ;
  assign w5941 = ( w3647 & ~w5939 ) | ( w3647 & w5940 ) | ( ~w5939 & w5940 ) ;
  assign w5942 = w3548 | w5395 ;
  assign w5943 = w3725 & ~w5941 ;
  assign w5944 = ( w4908 & w5941 ) | ( w4908 & ~w5943 ) | ( w5941 & ~w5943 ) ;
  assign w5945 = ( ~w3548 & w5942 ) | ( ~w3548 & w5944 ) | ( w5942 & w5944 ) ;
  assign w5946 = \pi20 ^ w5945 ;
  assign w5947 = ( w5722 & w5938 ) | ( w5722 & w5946 ) | ( w5938 & w5946 ) ;
  assign w5948 = ~w5495 & w5496 ;
  assign w5949 = w4049 | w5494 ;
  assign w5950 = ~w4142 & w5710 ;
  assign w5951 = ( ~w4049 & w5949 ) | ( ~w4049 & w5950 ) | ( w5949 & w5950 ) ;
  assign w5952 = w3962 | w5948 ;
  assign w5953 = w4152 & ~w5951 ;
  assign w5954 = ( w5497 & w5951 ) | ( w5497 & ~w5953 ) | ( w5951 & ~w5953 ) ;
  assign w5955 = ( ~w3962 & w5952 ) | ( ~w3962 & w5954 ) | ( w5952 & w5954 ) ;
  assign w5956 = \pi17 ^ w5955 ;
  assign w5957 = ( w5720 & w5947 ) | ( w5720 & w5956 ) | ( w5947 & w5956 ) ;
  assign w5958 = ~w4142 & w5494 ;
  assign w5959 = ( ~w4600 & w5948 ) | ( ~w4600 & w5958 ) | ( w5948 & w5958 ) ;
  assign w5960 = w5710 | w5959 ;
  assign w5961 = ( ~w3962 & w5959 ) | ( ~w3962 & w5960 ) | ( w5959 & w5960 ) ;
  assign w5962 = w5958 | w5961 ;
  assign w5963 = w5523 ^ w5706 ;
  assign w5964 = w5515 ^ w5963 ;
  assign w5965 = w4722 & ~w5962 ;
  assign w5966 = ( w5497 & w5962 ) | ( w5497 & ~w5965 ) | ( w5962 & ~w5965 ) ;
  assign w5967 = \pi17 ^ w5966 ;
  assign w5968 = ( w5957 & ~w5964 ) | ( w5957 & w5967 ) | ( ~w5964 & w5967 ) ;
  assign w5969 = w5722 ^ w5946 ;
  assign w5970 = w5938 ^ w5969 ;
  assign w5971 = w5730 ^ w5937 ;
  assign w5972 = w5732 ^ w5971 ;
  assign w5973 = w3647 & ~w5343 ;
  assign w5974 = ~w3094 & w4905 ;
  assign w5975 = ( w3647 & ~w5973 ) | ( w3647 & w5974 ) | ( ~w5973 & w5974 ) ;
  assign w5976 = w3715 & ~w5395 ;
  assign w5977 = w4164 & ~w5975 ;
  assign w5978 = ( w4908 & w5975 ) | ( w4908 & ~w5977 ) | ( w5975 & ~w5977 ) ;
  assign w5979 = ( w3715 & ~w5976 ) | ( w3715 & w5978 ) | ( ~w5976 & w5978 ) ;
  assign w5980 = \pi20 ^ w5979 ;
  assign w5981 = w5734 ^ w5936 ;
  assign w5982 = w5928 ^ w5981 ;
  assign w5983 = w5919 ^ w5927 ;
  assign w5984 = w5917 ^ w5983 ;
  assign w5985 = w5742 ^ w5916 ;
  assign w5986 = w5744 ^ w5985 ;
  assign w5987 = w1264 | w4143 ;
  assign w5988 = w1399 & w4052 ;
  assign w5989 = ( ~w1264 & w5987 ) | ( ~w1264 & w5988 ) | ( w5987 & w5988 ) ;
  assign w5990 = w4147 | w4864 ;
  assign w5991 = w1205 | w5989 ;
  assign w5992 = ( w3964 & w5989 ) | ( w3964 & w5991 ) | ( w5989 & w5991 ) ;
  assign w5993 = ( ~w4864 & w5990 ) | ( ~w4864 & w5992 ) | ( w5990 & w5992 ) ;
  assign w5994 = \pi26 ^ w5993 ;
  assign w5995 = w5746 ^ w5915 ;
  assign w5996 = w5756 ^ w5995 ;
  assign w5997 = w1711 & ~w3717 ;
  assign w5998 = ~w1834 & w3649 ;
  assign w5999 = ( w1711 & ~w5997 ) | ( w1711 & w5998 ) | ( ~w5997 & w5998 ) ;
  assign w6000 = w1614 & ~w3549 ;
  assign w6001 = w5433 & ~w5999 ;
  assign w6002 = ( w3448 & w5999 ) | ( w3448 & ~w6001 ) | ( w5999 & ~w6001 ) ;
  assign w6003 = ( w1614 & ~w6000 ) | ( w1614 & w6002 ) | ( ~w6000 & w6002 ) ;
  assign w6004 = \pi29 ^ w6003 ;
  assign w6005 = w1399 & ~w4143 ;
  assign w6006 = ~w1510 & w4052 ;
  assign w6007 = ( w1399 & ~w6005 ) | ( w1399 & w6006 ) | ( ~w6005 & w6006 ) ;
  assign w6008 = w4147 | w4852 ;
  assign w6009 = w1264 & ~w6007 ;
  assign w6010 = ( w3964 & w6007 ) | ( w3964 & ~w6009 ) | ( w6007 & ~w6009 ) ;
  assign w6011 = ( ~w4852 & w6008 ) | ( ~w4852 & w6010 ) | ( w6008 & w6010 ) ;
  assign w6012 = \pi26 ^ w6011 ;
  assign w6013 = ( w5996 & w6004 ) | ( w5996 & w6012 ) | ( w6004 & w6012 ) ;
  assign w6014 = ( w5986 & w5994 ) | ( w5986 & w6013 ) | ( w5994 & w6013 ) ;
  assign w6015 = w883 | w4651 ;
  assign w6016 = w979 & w4606 ;
  assign w6017 = ( ~w883 & w6015 ) | ( ~w883 & w6016 ) | ( w6015 & w6016 ) ;
  assign w6018 = w721 & ~w4706 ;
  assign w6019 = w4257 & ~w6017 ;
  assign w6020 = ( w4609 & w6017 ) | ( w4609 & ~w6019 ) | ( w6017 & ~w6019 ) ;
  assign w6021 = ( w721 & ~w6018 ) | ( w721 & w6020 ) | ( ~w6018 & w6020 ) ;
  assign w6022 = \pi23 ^ w6021 ;
  assign w6023 = ( w5984 & w6014 ) | ( w5984 & w6022 ) | ( w6014 & w6022 ) ;
  assign w6024 = w381 | w4905 ;
  assign w6025 = ~w3094 & w5343 ;
  assign w6026 = ( ~w381 & w6024 ) | ( ~w381 & w6025 ) | ( w6024 & w6025 ) ;
  assign w6027 = w3647 & ~w5395 ;
  assign w6028 = w3810 | w6026 ;
  assign w6029 = ( w4908 & w6026 ) | ( w4908 & w6028 ) | ( w6026 & w6028 ) ;
  assign w6030 = ( w3647 & ~w6027 ) | ( w3647 & w6029 ) | ( ~w6027 & w6029 ) ;
  assign w6031 = \pi20 ^ w6030 ;
  assign w6032 = ( w5982 & w6023 ) | ( w5982 & w6031 ) | ( w6023 & w6031 ) ;
  assign w6033 = ( w5972 & w5980 ) | ( w5972 & w6032 ) | ( w5980 & w6032 ) ;
  assign w6034 = w4049 | w5710 ;
  assign w6035 = w3907 & w5494 ;
  assign w6036 = ( ~w4049 & w6034 ) | ( ~w4049 & w6035 ) | ( w6034 & w6035 ) ;
  assign w6037 = w4142 | w5948 ;
  assign w6038 = w4563 | w6036 ;
  assign w6039 = ( w5497 & w6036 ) | ( w5497 & w6038 ) | ( w6036 & w6038 ) ;
  assign w6040 = ( ~w4142 & w6037 ) | ( ~w4142 & w6039 ) | ( w6037 & w6039 ) ;
  assign w6041 = \pi17 ^ w6040 ;
  assign w6042 = ( w5970 & w6033 ) | ( w5970 & w6041 ) | ( w6033 & w6041 ) ;
  assign w6043 = \pi13 ^ \pi14 ;
  assign w6044 = \pi11 ^ \pi12 ;
  assign w6045 = w6043 & w6044 ;
  assign w6046 = ( \pi12 & ~\pi13 ) | ( \pi12 & \pi14 ) | ( ~\pi13 & \pi14 ) ;
  assign w6047 = ( \pi11 & \pi12 ) | ( \pi11 & w6046 ) | ( \pi12 & w6046 ) ;
  assign w6048 = w6046 ^ w6047 ;
  assign w6049 = ~w4600 & w6048 ;
  assign w6050 = w6045 | w6049 ;
  assign w6051 = ( ~w4603 & w6049 ) | ( ~w4603 & w6050 ) | ( w6049 & w6050 ) ;
  assign w6052 = \pi14 ^ w6051 ;
  assign w6053 = w5720 ^ w5956 ;
  assign w6054 = w5947 ^ w6053 ;
  assign w6055 = ( w6042 & w6052 ) | ( w6042 & w6054 ) | ( w6052 & w6054 ) ;
  assign w6056 = w4722 & w5497 ;
  assign w6057 = ( w5497 & w5962 ) | ( w5497 & ~w6056 ) | ( w5962 & ~w6056 ) ;
  assign w6058 = w5957 ^ w6057 ;
  assign w6059 = \pi17 ^ w5964 ;
  assign w6060 = w6058 ^ w6059 ;
  assign w6061 = w6052 ^ w6054 ;
  assign w6062 = w6042 ^ w6061 ;
  assign w6063 = w3548 | w5494 ;
  assign w6064 = w3907 & w5710 ;
  assign w6065 = ( ~w3548 & w6063 ) | ( ~w3548 & w6064 ) | ( w6063 & w6064 ) ;
  assign w6066 = w4049 | w5948 ;
  assign w6067 = w4622 & ~w6065 ;
  assign w6068 = ( w5497 & w6065 ) | ( w5497 & ~w6067 ) | ( w6065 & ~w6067 ) ;
  assign w6069 = ( ~w4049 & w6066 ) | ( ~w4049 & w6068 ) | ( w6066 & w6068 ) ;
  assign w6070 = \pi17 ^ w6069 ;
  assign w6071 = w5980 ^ w6032 ;
  assign w6072 = w5972 ^ w6071 ;
  assign w6073 = w5982 ^ w6031 ;
  assign w6074 = w6023 ^ w6073 ;
  assign w6075 = w5984 ^ w6022 ;
  assign w6076 = w6014 ^ w6075 ;
  assign w6077 = w979 & ~w4651 ;
  assign w6078 = w1085 & w4606 ;
  assign w6079 = ( w979 & ~w6077 ) | ( w979 & w6078 ) | ( ~w6077 & w6078 ) ;
  assign w6080 = w883 | w4706 ;
  assign w6081 = w4273 & ~w6079 ;
  assign w6082 = ( w4609 & w6079 ) | ( w4609 & ~w6081 ) | ( w6079 & ~w6081 ) ;
  assign w6083 = ( ~w883 & w6080 ) | ( ~w883 & w6082 ) | ( w6080 & w6082 ) ;
  assign w6084 = \pi23 ^ w6083 ;
  assign w6085 = w5994 ^ w6013 ;
  assign w6086 = w5986 ^ w6085 ;
  assign w6087 = w5996 ^ w6012 ;
  assign w6088 = w6004 ^ w6087 ;
  assign w6089 = w5892 ^ w5905 ;
  assign w6090 = w5894 ^ w6089 ;
  assign w6091 = w5791 ^ w5891 ;
  assign w6092 = \pi02 ^ w6091 ;
  assign w6093 = w2130 ^ w2982 ;
  assign w6094 = w2235 ^ w6093 ;
  assign w6095 = ~w37 & w6094 ;
  assign w6096 = w2273 & w3098 ;
  assign w6097 = ( w6094 & ~w6095 ) | ( w6094 & w6096 ) | ( ~w6095 & w6096 ) ;
  assign w6098 = ( \pi29 & \pi30 ) | ( \pi29 & ~w2130 ) | ( \pi30 & ~w2130 ) ;
  assign w6099 = \pi31 | w6098 ;
  assign w6100 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w2235 ) | ( \pi30 & w2235 ) ;
  assign w6101 = ( \pi29 & \pi31 ) | ( \pi29 & w6100 ) | ( \pi31 & w6100 ) ;
  assign w6102 = ( w6097 & w6099 ) | ( w6097 & ~w6101 ) | ( w6099 & ~w6101 ) ;
  assign w6103 = w5829 ^ w5890 ;
  assign w6104 = \pi02 ^ w6103 ;
  assign w6105 = w2273 ^ w2981 ;
  assign w6106 = w2235 ^ w6105 ;
  assign w6107 = w37 | w6106 ;
  assign w6108 = w2391 & w3098 ;
  assign w6109 = ( ~w6106 & w6107 ) | ( ~w6106 & w6108 ) | ( w6107 & w6108 ) ;
  assign w6110 = ( \pi29 & \pi30 ) | ( \pi29 & ~w2235 ) | ( \pi30 & ~w2235 ) ;
  assign w6111 = \pi31 | w6110 ;
  assign w6112 = ( \pi29 & ~\pi30 ) | ( \pi29 & w2273 ) | ( ~\pi30 & w2273 ) ;
  assign w6113 = ( \pi29 & \pi31 ) | ( \pi29 & ~w6112 ) | ( \pi31 & ~w6112 ) ;
  assign w6114 = ( w6109 & w6111 ) | ( w6109 & ~w6113 ) | ( w6111 & ~w6113 ) ;
  assign w6115 = w5878 ^ w5889 ;
  assign w6116 = \pi02 ^ w6115 ;
  assign w6117 = ( w504 & w681 ) | ( w504 & ~w899 ) | ( w681 & ~w899 ) ;
  assign w6118 = w458 | w496 ;
  assign w6119 = ( ~w496 & w899 ) | ( ~w496 & w1340 ) | ( w899 & w1340 ) ;
  assign w6120 = w6118 | w6119 ;
  assign w6121 = w6117 | w6120 ;
  assign w6122 = ( ~w561 & w4363 ) | ( ~w561 & w6121 ) | ( w4363 & w6121 ) ;
  assign w6123 = w888 | w1849 ;
  assign w6124 = ( w561 & w817 ) | ( w561 & ~w888 ) | ( w817 & ~w888 ) ;
  assign w6125 = w6123 | w6124 ;
  assign w6126 = w6122 | w6125 ;
  assign w6127 = ( w88 & ~w149 ) | ( w88 & w1165 ) | ( ~w149 & w1165 ) ;
  assign w6128 = w82 | w6126 ;
  assign w6129 = ( ~w82 & w149 ) | ( ~w82 & w623 ) | ( w149 & w623 ) ;
  assign w6130 = w6128 | w6129 ;
  assign w6131 = w6127 | w6130 ;
  assign w6132 = w802 | w821 ;
  assign w6133 = w230 | w6132 ;
  assign w6134 = ( ~w230 & w354 ) | ( ~w230 & w6131 ) | ( w354 & w6131 ) ;
  assign w6135 = w6133 | w6134 ;
  assign w6136 = w723 | w1126 ;
  assign w6137 = w180 | w6136 ;
  assign w6138 = ( w147 & ~w180 ) | ( w147 & w662 ) | ( ~w180 & w662 ) ;
  assign w6139 = w6137 | w6138 ;
  assign w6140 = w127 | w515 ;
  assign w6141 = ( w90 & ~w127 ) | ( w90 & w252 ) | ( ~w127 & w252 ) ;
  assign w6142 = w6140 | w6141 ;
  assign w6143 = ( w268 & w316 ) | ( w268 & ~w351 ) | ( w316 & ~w351 ) ;
  assign w6144 = w95 | w698 ;
  assign w6145 = w5595 | w6144 ;
  assign w6146 = w6143 | w6145 ;
  assign w6147 = w6142 | w6146 ;
  assign w6148 = ( ~w1759 & w4475 ) | ( ~w1759 & w6147 ) | ( w4475 & w6147 ) ;
  assign w6149 = w4508 | w6135 ;
  assign w6150 = ( w1759 & ~w6135 ) | ( w1759 & w6139 ) | ( ~w6135 & w6139 ) ;
  assign w6151 = w6149 | w6150 ;
  assign w6152 = w6148 | w6151 ;
  assign w6153 = ( w361 & ~w385 ) | ( w361 & w742 ) | ( ~w385 & w742 ) ;
  assign w6154 = w450 | w6152 ;
  assign w6155 = ( w385 & w408 ) | ( w385 & ~w450 ) | ( w408 & ~w450 ) ;
  assign w6156 = w6154 | w6155 ;
  assign w6157 = w6153 | w6156 ;
  assign w6158 = ( w225 & w255 ) | ( w225 & ~w280 ) | ( w255 & ~w280 ) ;
  assign w6159 = w104 | w6157 ;
  assign w6160 = ( ~w104 & w280 ) | ( ~w104 & w430 ) | ( w280 & w430 ) ;
  assign w6161 = w6159 | w6160 ;
  assign w6162 = w6158 | w6161 ;
  assign w6163 = w2391 ^ w2979 ;
  assign w6164 = w2500 ^ w6163 ;
  assign w6165 = w37 | w6164 ;
  assign w6166 = ~w2578 & w3098 ;
  assign w6167 = ( ~w6164 & w6165 ) | ( ~w6164 & w6166 ) | ( w6165 & w6166 ) ;
  assign w6168 = ( \pi29 & \pi30 ) | ( \pi29 & w2391 ) | ( \pi30 & w2391 ) ;
  assign w6169 = \pi31 | w6168 ;
  assign w6170 = ( \pi29 & ~\pi30 ) | ( \pi29 & w2500 ) | ( ~\pi30 & w2500 ) ;
  assign w6171 = ( \pi29 & \pi31 ) | ( \pi29 & ~w6170 ) | ( \pi31 & ~w6170 ) ;
  assign w6172 = ( w6167 & w6169 ) | ( w6167 & ~w6171 ) | ( w6169 & ~w6171 ) ;
  assign w6173 = ( w260 & ~w386 ) | ( w260 & w531 ) | ( ~w386 & w531 ) ;
  assign w6174 = w386 | w6173 ;
  assign w6175 = ( w142 & w516 ) | ( w142 & ~w837 ) | ( w516 & ~w837 ) ;
  assign w6176 = w133 | w6174 ;
  assign w6177 = ( ~w133 & w837 ) | ( ~w133 & w1229 ) | ( w837 & w1229 ) ;
  assign w6178 = w6176 | w6177 ;
  assign w6179 = w6175 | w6178 ;
  assign w6180 = w1629 | w2705 ;
  assign w6181 = w6179 | w6180 ;
  assign w6182 = ( w64 & w4204 ) | ( w64 & ~w6179 ) | ( w4204 & ~w6179 ) ;
  assign w6183 = w6181 | w6182 ;
  assign w6184 = ( w163 & w642 ) | ( w163 & ~w674 ) | ( w642 & ~w674 ) ;
  assign w6185 = w74 | w6183 ;
  assign w6186 = ( ~w74 & w674 ) | ( ~w74 & w787 ) | ( w674 & w787 ) ;
  assign w6187 = w6185 | w6186 ;
  assign w6188 = w6184 | w6187 ;
  assign w6189 = ( ~w44 & w568 ) | ( ~w44 & w6188 ) | ( w568 & w6188 ) ;
  assign w6190 = w44 | w6189 ;
  assign w6191 = w899 | w1086 ;
  assign w6192 = w280 | w6191 ;
  assign w6193 = ( ~w280 & w416 ) | ( ~w280 & w524 ) | ( w416 & w524 ) ;
  assign w6194 = w6192 | w6193 ;
  assign w6195 = ( w86 & w255 ) | ( w86 & ~w495 ) | ( w255 & ~w495 ) ;
  assign w6196 = ( w495 & w506 ) | ( w495 & ~w514 ) | ( w506 & ~w514 ) ;
  assign w6197 = w4510 | w6196 ;
  assign w6198 = w6195 | w6197 ;
  assign w6199 = w456 | w1154 ;
  assign w6200 = ( w266 & ~w1154 ) | ( w266 & w6198 ) | ( ~w1154 & w6198 ) ;
  assign w6201 = w6199 | w6200 ;
  assign w6202 = ( w890 & ~w1741 ) | ( w890 & w6194 ) | ( ~w1741 & w6194 ) ;
  assign w6203 = w250 | w6201 ;
  assign w6204 = ( w1741 & w1759 ) | ( w1741 & ~w6201 ) | ( w1759 & ~w6201 ) ;
  assign w6205 = w6203 | w6204 ;
  assign w6206 = w6202 | w6205 ;
  assign w6207 = ( w444 & ~w1814 ) | ( w444 & w5016 ) | ( ~w1814 & w5016 ) ;
  assign w6208 = w6190 | w6206 ;
  assign w6209 = ( w1814 & w4464 ) | ( w1814 & ~w6206 ) | ( w4464 & ~w6206 ) ;
  assign w6210 = w6208 | w6209 ;
  assign w6211 = w6207 | w6210 ;
  assign w6212 = w169 | w257 ;
  assign w6213 = w120 | w6212 ;
  assign w6214 = ( ~w120 & w144 ) | ( ~w120 & w6211 ) | ( w144 & w6211 ) ;
  assign w6215 = w6213 | w6214 ;
  assign w6216 = ( ~w175 & w492 ) | ( ~w175 & w6215 ) | ( w492 & w6215 ) ;
  assign w6217 = w175 | w6216 ;
  assign w6218 = w2578 ^ w2978 ;
  assign w6219 = w2500 ^ w6218 ;
  assign w6220 = ~w37 & w6219 ;
  assign w6221 = ~w2653 & w3098 ;
  assign w6222 = ( w6219 & ~w6220 ) | ( w6219 & w6221 ) | ( ~w6220 & w6221 ) ;
  assign w6223 = ( \pi29 & \pi30 ) | ( \pi29 & w2500 ) | ( \pi30 & w2500 ) ;
  assign w6224 = \pi31 | w6223 ;
  assign w6225 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w2578 ) | ( \pi30 & w2578 ) ;
  assign w6226 = ( \pi29 & \pi31 ) | ( \pi29 & w6225 ) | ( \pi31 & w6225 ) ;
  assign w6227 = ( w6222 & w6224 ) | ( w6222 & ~w6226 ) | ( w6224 & ~w6226 ) ;
  assign w6228 = w220 | w783 ;
  assign w6229 = ( ~w220 & w318 ) | ( ~w220 & w2274 ) | ( w318 & w2274 ) ;
  assign w6230 = w6228 | w6229 ;
  assign w6231 = w260 | w271 ;
  assign w6232 = w64 | w6231 ;
  assign w6233 = ( ~w64 & w259 ) | ( ~w64 & w6230 ) | ( w259 & w6230 ) ;
  assign w6234 = w6232 | w6233 ;
  assign w6235 = w680 | w817 ;
  assign w6236 = w224 | w6235 ;
  assign w6237 = ( ~w224 & w463 ) | ( ~w224 & w6234 ) | ( w463 & w6234 ) ;
  assign w6238 = w6236 | w6237 ;
  assign w6239 = w312 | w465 ;
  assign w6240 = ( ~w312 & w386 ) | ( ~w312 & w514 ) | ( w386 & w514 ) ;
  assign w6241 = w6239 | w6240 ;
  assign w6242 = w488 | w764 ;
  assign w6243 = ( ~w488 & w726 ) | ( ~w488 & w1881 ) | ( w726 & w1881 ) ;
  assign w6244 = w6242 | w6243 ;
  assign w6245 = ( w176 & w256 ) | ( w176 & ~w495 ) | ( w256 & ~w495 ) ;
  assign w6246 = w136 | w6244 ;
  assign w6247 = ( ~w136 & w495 ) | ( ~w136 & w504 ) | ( w495 & w504 ) ;
  assign w6248 = w6246 | w6247 ;
  assign w6249 = w6245 | w6248 ;
  assign w6250 = ( w638 & ~w731 ) | ( w638 & w6241 ) | ( ~w731 & w6241 ) ;
  assign w6251 = w5097 | w6249 ;
  assign w6252 = ( w389 & w731 ) | ( w389 & ~w5097 ) | ( w731 & ~w5097 ) ;
  assign w6253 = w6251 | w6252 ;
  assign w6254 = w6250 | w6253 ;
  assign w6255 = ( w341 & w354 ) | ( w341 & ~w408 ) | ( w354 & ~w408 ) ;
  assign w6256 = w122 | w6254 ;
  assign w6257 = ( ~w122 & w408 ) | ( ~w122 & w787 ) | ( w408 & w787 ) ;
  assign w6258 = w6256 | w6257 ;
  assign w6259 = w6255 | w6258 ;
  assign w6260 = w254 | w951 ;
  assign w6261 = ( ~w254 & w722 ) | ( ~w254 & w6259 ) | ( w722 & w6259 ) ;
  assign w6262 = w6260 | w6261 ;
  assign w6263 = w311 | w561 ;
  assign w6264 = ( ~w311 & w324 ) | ( ~w311 & w2252 ) | ( w324 & w2252 ) ;
  assign w6265 = w6263 | w6264 ;
  assign w6266 = ( w125 & w142 ) | ( w125 & ~w143 ) | ( w142 & ~w143 ) ;
  assign w6267 = w2479 | w6265 ;
  assign w6268 = ( w143 & w821 ) | ( w143 & ~w6265 ) | ( w821 & ~w6265 ) ;
  assign w6269 = w6267 | w6268 ;
  assign w6270 = w6266 | w6269 ;
  assign w6271 = ( ~w3866 & w6238 ) | ( ~w3866 & w6270 ) | ( w6238 & w6270 ) ;
  assign w6272 = w5180 & ~w6262 ;
  assign w6273 = ( w340 & w3866 ) | ( w340 & w5180 ) | ( w3866 & w5180 ) ;
  assign w6274 = w6272 & ~w6273 ;
  assign w6275 = ~w6271 & w6274 ;
  assign w6276 = ( w202 & w353 ) | ( w202 & ~w430 ) | ( w353 & ~w430 ) ;
  assign w6277 = ~w165 & w6275 ;
  assign w6278 = ( ~w165 & w430 ) | ( ~w165 & w837 ) | ( w430 & w837 ) ;
  assign w6279 = w6277 & ~w6278 ;
  assign w6280 = ~w6276 & w6279 ;
  assign w6281 = w2578 ^ w2977 ;
  assign w6282 = w2653 ^ w6281 ;
  assign w6283 = w37 | w6282 ;
  assign w6284 = ~w2694 & w3098 ;
  assign w6285 = ( ~w6282 & w6283 ) | ( ~w6282 & w6284 ) | ( w6283 & w6284 ) ;
  assign w6286 = ( \pi29 & \pi30 ) | ( \pi29 & ~w2578 ) | ( \pi30 & ~w2578 ) ;
  assign w6287 = \pi31 | w6286 ;
  assign w6288 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w2653 ) | ( \pi30 & w2653 ) ;
  assign w6289 = ( \pi29 & \pi31 ) | ( \pi29 & w6288 ) | ( \pi31 & w6288 ) ;
  assign w6290 = ( w6285 & w6287 ) | ( w6285 & ~w6289 ) | ( w6287 & ~w6289 ) ;
  assign w6291 = ( w388 & w429 ) | ( w388 & ~w431 ) | ( w429 & ~w431 ) ;
  assign w6292 = w203 | w3494 ;
  assign w6293 = ( ~w203 & w431 ) | ( ~w203 & w1153 ) | ( w431 & w1153 ) ;
  assign w6294 = w6292 | w6293 ;
  assign w6295 = w6291 | w6294 ;
  assign w6296 = w90 | w421 ;
  assign w6297 = w1131 | w6296 ;
  assign w6298 = ( ~w1131 & w1560 ) | ( ~w1131 & w6295 ) | ( w1560 & w6295 ) ;
  assign w6299 = w6297 | w6298 ;
  assign w6300 = ( w313 & w325 ) | ( w313 & ~w392 ) | ( w325 & ~w392 ) ;
  assign w6301 = w312 | w6299 ;
  assign w6302 = ( ~w312 & w392 ) | ( ~w312 & w424 ) | ( w392 & w424 ) ;
  assign w6303 = w6301 | w6302 ;
  assign w6304 = w6300 | w6303 ;
  assign w6305 = ( w287 & w345 ) | ( w287 & ~w422 ) | ( w345 & ~w422 ) ;
  assign w6306 = w128 | w838 ;
  assign w6307 = ( ~w128 & w422 ) | ( ~w128 & w515 ) | ( w422 & w515 ) ;
  assign w6308 = w6306 | w6307 ;
  assign w6309 = w6305 | w6308 ;
  assign w6310 = w198 | w530 ;
  assign w6311 = ( w131 & ~w198 ) | ( w131 & w285 ) | ( ~w198 & w285 ) ;
  assign w6312 = w6310 | w6311 ;
  assign w6313 = w262 | w316 ;
  assign w6314 = w1620 | w6313 ;
  assign w6315 = ( w609 & ~w1620 ) | ( w609 & w4352 ) | ( ~w1620 & w4352 ) ;
  assign w6316 = w6314 | w6315 ;
  assign w6317 = ( w6309 & w6312 ) | ( w6309 & ~w6316 ) | ( w6312 & ~w6316 ) ;
  assign w6318 = w6316 | w6317 ;
  assign w6319 = ( ~w495 & w2695 ) | ( ~w495 & w6318 ) | ( w2695 & w6318 ) ;
  assign w6320 = w2350 | w6304 ;
  assign w6321 = ( w495 & w513 ) | ( w495 & ~w6304 ) | ( w513 & ~w6304 ) ;
  assign w6322 = w6320 | w6321 ;
  assign w6323 = w6319 | w6322 ;
  assign w6324 = ( w1166 & w1185 ) | ( w1166 & ~w1566 ) | ( w1185 & ~w1566 ) ;
  assign w6325 = w998 | w6323 ;
  assign w6326 = ( w340 & ~w998 ) | ( w340 & w1566 ) | ( ~w998 & w1566 ) ;
  assign w6327 = w6325 | w6326 ;
  assign w6328 = w6324 | w6327 ;
  assign w6329 = ( w281 & w490 ) | ( w281 & ~w570 ) | ( w490 & ~w570 ) ;
  assign w6330 = w135 | w6328 ;
  assign w6331 = ( ~w135 & w570 ) | ( ~w135 & w628 ) | ( w570 & w628 ) ;
  assign w6332 = w6330 | w6331 ;
  assign w6333 = w6329 | w6332 ;
  assign w6334 = ( ~w2694 & w2805 ) | ( ~w2694 & w2871 ) | ( w2805 & w2871 ) ;
  assign w6335 = ~w2694 & w2973 ;
  assign w6336 = w6334 | w6335 ;
  assign w6337 = w2653 ^ w2805 ;
  assign w6338 = w6336 ^ w6337 ;
  assign w6339 = w37 | w6338 ;
  assign w6340 = w2805 & w3098 ;
  assign w6341 = ( ~w6338 & w6339 ) | ( ~w6338 & w6340 ) | ( w6339 & w6340 ) ;
  assign w6342 = ( \pi29 & \pi30 ) | ( \pi29 & ~w2653 ) | ( \pi30 & ~w2653 ) ;
  assign w6343 = \pi31 | w6342 ;
  assign w6344 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w2694 ) | ( \pi30 & w2694 ) ;
  assign w6345 = ( \pi29 & \pi31 ) | ( \pi29 & w6344 ) | ( \pi31 & w6344 ) ;
  assign w6346 = ( w6341 & w6343 ) | ( w6341 & ~w6345 ) | ( w6343 & ~w6345 ) ;
  assign w6347 = ( w269 & w283 ) | ( w269 & ~w310 ) | ( w283 & ~w310 ) ;
  assign w6348 = w178 | w282 ;
  assign w6349 = ( ~w178 & w310 ) | ( ~w178 & w1128 ) | ( w310 & w1128 ) ;
  assign w6350 = w6348 | w6349 ;
  assign w6351 = w6347 | w6350 ;
  assign w6352 = ( w114 & ~w135 ) | ( w114 & w533 ) | ( ~w135 & w533 ) ;
  assign w6353 = w135 | w6352 ;
  assign w6354 = w605 | w680 ;
  assign w6355 = w2760 | w6354 ;
  assign w6356 = ( w76 & w1565 ) | ( w76 & ~w2760 ) | ( w1565 & ~w2760 ) ;
  assign w6357 = w6355 | w6356 ;
  assign w6358 = ( ~w352 & w359 ) | ( ~w352 & w637 ) | ( w359 & w637 ) ;
  assign w6359 = w3965 | w6357 ;
  assign w6360 = ( w637 & w725 ) | ( w637 & ~w3965 ) | ( w725 & ~w3965 ) ;
  assign w6361 = w6359 | w6360 ;
  assign w6362 = w6358 & ~w6361 ;
  assign w6363 = w176 | w420 ;
  assign w6364 = ( w101 & ~w176 ) | ( w101 & w342 ) | ( ~w176 & w342 ) ;
  assign w6365 = w6363 | w6364 ;
  assign w6366 = w351 | w560 ;
  assign w6367 = w2536 | w6366 ;
  assign w6368 = ( w1155 & ~w2536 ) | ( w1155 & w6365 ) | ( ~w2536 & w6365 ) ;
  assign w6369 = w6367 | w6368 ;
  assign w6370 = ( w209 & w316 ) | ( w209 & ~w322 ) | ( w316 & ~w322 ) ;
  assign w6371 = w672 | w6369 ;
  assign w6372 = ( w322 & w421 ) | ( w322 & ~w672 ) | ( w421 & ~w672 ) ;
  assign w6373 = w6371 | w6372 ;
  assign w6374 = w6370 | w6373 ;
  assign w6375 = ( w204 & ~w224 ) | ( w204 & w1566 ) | ( ~w224 & w1566 ) ;
  assign w6376 = w6362 & ~w6374 ;
  assign w6377 = ( w224 & w413 ) | ( w224 & ~w6374 ) | ( w413 & ~w6374 ) ;
  assign w6378 = w6376 & ~w6377 ;
  assign w6379 = ~w6375 & w6378 ;
  assign w6380 = w951 | w1126 ;
  assign w6381 = w167 | w6380 ;
  assign w6382 = ( w167 & ~w515 ) | ( w167 & w6379 ) | ( ~w515 & w6379 ) ;
  assign w6383 = ~w6381 & w6382 ;
  assign w6384 = ( w470 & ~w531 ) | ( w470 & w6383 ) | ( ~w531 & w6383 ) ;
  assign w6385 = ~w470 & w6384 ;
  assign w6386 = ( ~w113 & w210 ) | ( ~w113 & w900 ) | ( w210 & w900 ) ;
  assign w6387 = w113 | w6386 ;
  assign w6388 = w1659 | w6387 ;
  assign w6389 = ( w1247 & w2759 ) | ( w1247 & ~w6387 ) | ( w2759 & ~w6387 ) ;
  assign w6390 = w6388 | w6389 ;
  assign w6391 = w2091 | w6353 ;
  assign w6392 = w6385 & ~w6391 ;
  assign w6393 = ( w1492 & w6385 ) | ( w1492 & w6390 ) | ( w6385 & w6390 ) ;
  assign w6394 = w6392 & ~w6393 ;
  assign w6395 = ( w254 & w315 ) | ( w254 & ~w445 ) | ( w315 & ~w445 ) ;
  assign w6396 = ~w6351 & w6394 ;
  assign w6397 = ( w445 & w1130 ) | ( w445 & ~w6351 ) | ( w1130 & ~w6351 ) ;
  assign w6398 = w6396 & ~w6397 ;
  assign w6399 = ~w6395 & w6398 ;
  assign w6400 = ( w565 & ~w662 ) | ( w565 & w6399 ) | ( ~w662 & w6399 ) ;
  assign w6401 = ~w565 & w6400 ;
  assign w6402 = w889 | w1340 ;
  assign w6403 = w76 | w6402 ;
  assign w6404 = ( ~w76 & w282 ) | ( ~w76 & w605 ) | ( w282 & w605 ) ;
  assign w6405 = w6403 | w6404 ;
  assign w6406 = w361 | w567 ;
  assign w6407 = w315 | w6406 ;
  assign w6408 = ( ~w315 & w358 ) | ( ~w315 & w6405 ) | ( w358 & w6405 ) ;
  assign w6409 = w6407 | w6408 ;
  assign w6410 = ( w163 & w443 ) | ( w163 & ~w449 ) | ( w443 & ~w449 ) ;
  assign w6411 = w120 | w147 ;
  assign w6412 = ( ~w147 & w449 ) | ( ~w147 & w606 ) | ( w449 & w606 ) ;
  assign w6413 = w6411 | w6412 ;
  assign w6414 = w6410 | w6413 ;
  assign w6415 = ( w210 & w260 ) | ( w210 & ~w312 ) | ( w260 & ~w312 ) ;
  assign w6416 = w6312 | w6414 ;
  assign w6417 = ( w312 & w463 ) | ( w312 & ~w6414 ) | ( w463 & ~w6414 ) ;
  assign w6418 = w6416 | w6417 ;
  assign w6419 = w6415 | w6418 ;
  assign w6420 = ( w1881 & w2079 ) | ( w1881 & ~w2147 ) | ( w2079 & ~w2147 ) ;
  assign w6421 = w887 | w6419 ;
  assign w6422 = ( ~w887 & w2147 ) | ( ~w887 & w2872 ) | ( w2147 & w2872 ) ;
  assign w6423 = w6421 | w6422 ;
  assign w6424 = w6420 | w6423 ;
  assign w6425 = ( w415 & w608 ) | ( w415 & ~w726 ) | ( w608 & ~w726 ) ;
  assign w6426 = w384 | w6424 ;
  assign w6427 = ( ~w384 & w726 ) | ( ~w384 & w897 ) | ( w726 & w897 ) ;
  assign w6428 = w6426 | w6427 ;
  assign w6429 = w6425 | w6428 ;
  assign w6430 = w625 | w1153 ;
  assign w6431 = ( ~w625 & w637 ) | ( ~w625 & w1566 ) | ( w637 & w1566 ) ;
  assign w6432 = w6430 | w6431 ;
  assign w6433 = ( ~w533 & w1629 ) | ( ~w533 & w6432 ) | ( w1629 & w6432 ) ;
  assign w6434 = w2183 & ~w4229 ;
  assign w6435 = ( w533 & w663 ) | ( w533 & w2183 ) | ( w663 & w2183 ) ;
  assign w6436 = w6434 & ~w6435 ;
  assign w6437 = ~w6433 & w6436 ;
  assign w6438 = ( w270 & ~w510 ) | ( w270 & w6409 ) | ( ~w510 & w6409 ) ;
  assign w6439 = ~w6429 & w6437 ;
  assign w6440 = ( w510 & w1713 ) | ( w510 & ~w6429 ) | ( w1713 & ~w6429 ) ;
  assign w6441 = w6439 & ~w6440 ;
  assign w6442 = ~w6438 & w6441 ;
  assign w6443 = ( w201 & w221 ) | ( w201 & ~w232 ) | ( w221 & ~w232 ) ;
  assign w6444 = ~w822 & w6442 ;
  assign w6445 = ( w232 & w623 ) | ( w232 & ~w822 ) | ( w623 & ~w822 ) ;
  assign w6446 = w6444 & ~w6445 ;
  assign w6447 = ~w6443 & w6446 ;
  assign w6448 = ( w214 & w230 ) | ( w214 & ~w271 ) | ( w230 & ~w271 ) ;
  assign w6449 = ~w178 & w6447 ;
  assign w6450 = ( ~w178 & w271 ) | ( ~w178 & w511 ) | ( w271 & w511 ) ;
  assign w6451 = w6449 & ~w6450 ;
  assign w6452 = ~w6448 & w6451 ;
  assign w6453 = w224 | w787 ;
  assign w6454 = ( w224 & ~w353 ) | ( w224 & w6452 ) | ( ~w353 & w6452 ) ;
  assign w6455 = ~w6453 & w6454 ;
  assign w6456 = ~w2871 & w2973 ;
  assign w6457 = w2805 ^ w6456 ;
  assign w6458 = \pi31 & ~w2973 ;
  assign w6459 = w2805 ^ w6458 ;
  assign w6460 = ( \pi29 & \pi30 ) | ( \pi29 & w6459 ) | ( \pi30 & w6459 ) ;
  assign w6461 = \pi31 ^ w6460 ;
  assign w6462 = \pi30 & \pi31 ;
  assign w6463 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w2973 ) | ( \pi30 & w2973 ) ;
  assign w6464 = w6462 & ~w6463 ;
  assign w6465 = ( ~w2871 & w6461 ) | ( ~w2871 & w6464 ) | ( w6461 & w6464 ) ;
  assign w6466 = w36 & w2805 ;
  assign w6467 = ( w2871 & w6464 ) | ( w2871 & w6466 ) | ( w6464 & w6466 ) ;
  assign w6468 = w6465 | w6467 ;
  assign w6469 = ~w6455 & w6468 ;
  assign w6470 = w2694 ^ w2805 ;
  assign w6471 = w2805 & ~w2871 ;
  assign w6472 = ( w2871 & w2973 ) | ( w2871 & ~w6471 ) | ( w2973 & ~w6471 ) ;
  assign w6473 = w6470 ^ w6472 ;
  assign w6474 = ( \pi30 & \pi31 ) | ( \pi30 & w2805 ) | ( \pi31 & w2805 ) ;
  assign w6475 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w6474 ) | ( \pi30 & w6474 ) ;
  assign w6476 = ( \pi29 & ~\pi30 ) | ( \pi29 & w6474 ) | ( ~\pi30 & w6474 ) ;
  assign w6477 = ( \pi30 & w2871 ) | ( \pi30 & ~w6476 ) | ( w2871 & ~w6476 ) ;
  assign w6478 = ( ~w2694 & w6476 ) | ( ~w2694 & w6477 ) | ( w6476 & w6477 ) ;
  assign w6479 = ~\pi31 & w6478 ;
  assign w6480 = ( w6475 & ~w6477 ) | ( w6475 & w6479 ) | ( ~w6477 & w6479 ) ;
  assign w6481 = ( w37 & w6473 ) | ( w37 & w6480 ) | ( w6473 & w6480 ) ;
  assign w6482 = w6480 | w6481 ;
  assign w6483 = ( ~w6401 & w6469 ) | ( ~w6401 & w6482 ) | ( w6469 & w6482 ) ;
  assign w6484 = ( w6333 & w6346 ) | ( w6333 & w6483 ) | ( w6346 & w6483 ) ;
  assign w6485 = ( ~w6280 & w6290 ) | ( ~w6280 & w6484 ) | ( w6290 & w6484 ) ;
  assign w6486 = ( w6217 & w6227 ) | ( w6217 & w6485 ) | ( w6227 & w6485 ) ;
  assign w6487 = ( w6162 & w6172 ) | ( w6162 & w6486 ) | ( w6172 & w6486 ) ;
  assign w6488 = w2130 | w3717 ;
  assign w6489 = ~w2235 & w3649 ;
  assign w6490 = ( ~w2130 & w6488 ) | ( ~w2130 & w6489 ) | ( w6488 & w6489 ) ;
  assign w6491 = w2059 | w3549 ;
  assign w6492 = w5896 & ~w6490 ;
  assign w6493 = ( w3448 & w6490 ) | ( w3448 & ~w6492 ) | ( w6490 & ~w6492 ) ;
  assign w6494 = ( ~w2059 & w6491 ) | ( ~w2059 & w6493 ) | ( w6491 & w6493 ) ;
  assign w6495 = \pi29 ^ w6494 ;
  assign w6496 = ( w6116 & w6487 ) | ( w6116 & w6495 ) | ( w6487 & w6495 ) ;
  assign w6497 = ( w6104 & w6114 ) | ( w6104 & w6496 ) | ( w6114 & w6496 ) ;
  assign w6498 = ( ~w6092 & w6102 ) | ( ~w6092 & w6497 ) | ( w6102 & w6497 ) ;
  assign w6499 = w1939 | w3717 ;
  assign w6500 = w1976 & w3649 ;
  assign w6501 = ( ~w1939 & w6499 ) | ( ~w1939 & w6500 ) | ( w6499 & w6500 ) ;
  assign w6502 = w1834 | w3549 ;
  assign w6503 = w5659 & ~w6501 ;
  assign w6504 = ( w3448 & w6501 ) | ( w3448 & ~w6503 ) | ( w6501 & ~w6503 ) ;
  assign w6505 = ( ~w1834 & w6502 ) | ( ~w1834 & w6504 ) | ( w6502 & w6504 ) ;
  assign w6506 = \pi29 ^ w6505 ;
  assign w6507 = ( w6090 & w6498 ) | ( w6090 & w6506 ) | ( w6498 & w6506 ) ;
  assign w6508 = w5758 ^ w5914 ;
  assign w6509 = w5906 ^ w6508 ;
  assign w6510 = w1614 & ~w4052 ;
  assign w6511 = ~w1510 & w4143 ;
  assign w6512 = ( w1614 & ~w6510 ) | ( w1614 & w6511 ) | ( ~w6510 & w6511 ) ;
  assign w6513 = w4147 | w5069 ;
  assign w6514 = w1399 | w6512 ;
  assign w6515 = ( w3964 & w6512 ) | ( w3964 & w6514 ) | ( w6512 & w6514 ) ;
  assign w6516 = ( ~w5069 & w6513 ) | ( ~w5069 & w6515 ) | ( w6513 & w6515 ) ;
  assign w6517 = \pi26 ^ w6516 ;
  assign w6518 = ( w6507 & ~w6509 ) | ( w6507 & w6517 ) | ( ~w6509 & w6517 ) ;
  assign w6519 = w1085 & ~w4651 ;
  assign w6520 = w1205 & w4606 ;
  assign w6521 = ( w1085 & ~w6519 ) | ( w1085 & w6520 ) | ( ~w6519 & w6520 ) ;
  assign w6522 = w979 & ~w4706 ;
  assign w6523 = w4666 | w6521 ;
  assign w6524 = ( w4609 & w6521 ) | ( w4609 & w6523 ) | ( w6521 & w6523 ) ;
  assign w6525 = ( w979 & ~w6522 ) | ( w979 & w6524 ) | ( ~w6522 & w6524 ) ;
  assign w6526 = \pi23 ^ w6525 ;
  assign w6527 = ( w6088 & w6518 ) | ( w6088 & w6526 ) | ( w6518 & w6526 ) ;
  assign w6528 = ( w6084 & w6086 ) | ( w6084 & w6527 ) | ( w6086 & w6527 ) ;
  assign w6529 = w381 | w5343 ;
  assign w6530 = w592 & w4905 ;
  assign w6531 = ( ~w381 & w6529 ) | ( ~w381 & w6530 ) | ( w6529 & w6530 ) ;
  assign w6532 = w3094 | w5395 ;
  assign w6533 = w3096 | w6531 ;
  assign w6534 = ( w4908 & w6531 ) | ( w4908 & w6533 ) | ( w6531 & w6533 ) ;
  assign w6535 = ( ~w3094 & w6532 ) | ( ~w3094 & w6534 ) | ( w6532 & w6534 ) ;
  assign w6536 = \pi20 ^ w6535 ;
  assign w6537 = ( w6076 & w6528 ) | ( w6076 & w6536 ) | ( w6528 & w6536 ) ;
  assign w6538 = w3548 | w5710 ;
  assign w6539 = w3715 & w5494 ;
  assign w6540 = ( ~w3548 & w6538 ) | ( ~w3548 & w6539 ) | ( w6538 & w6539 ) ;
  assign w6541 = w3907 & ~w5948 ;
  assign w6542 = w3913 & ~w6540 ;
  assign w6543 = ( w5497 & w6540 ) | ( w5497 & ~w6542 ) | ( w6540 & ~w6542 ) ;
  assign w6544 = ( w3907 & ~w6541 ) | ( w3907 & w6543 ) | ( ~w6541 & w6543 ) ;
  assign w6545 = \pi17 ^ w6544 ;
  assign w6546 = ( w6074 & w6537 ) | ( w6074 & w6545 ) | ( w6537 & w6545 ) ;
  assign w6547 = ( w6070 & w6072 ) | ( w6070 & w6546 ) | ( w6072 & w6546 ) ;
  assign w6548 = ( \pi11 & \pi12 ) | ( \pi11 & \pi13 ) | ( \pi12 & \pi13 ) ;
  assign w6549 = \pi13 ^ w6548 ;
  assign w6550 = ~w4600 & w6549 ;
  assign w6551 = ( w3962 & w4600 ) | ( w3962 & ~w4601 ) | ( w4600 & ~w4601 ) ;
  assign w6552 = ( w3962 & w6045 ) | ( w3962 & w6551 ) | ( w6045 & w6551 ) ;
  assign w6553 = w3962 | w6048 ;
  assign w6554 = ( ~w3962 & w6552 ) | ( ~w3962 & w6553 ) | ( w6552 & w6553 ) ;
  assign w6555 = w3962 & w6551 ;
  assign w6556 = ( w6550 & w6554 ) | ( w6550 & ~w6555 ) | ( w6554 & ~w6555 ) ;
  assign w6557 = w5970 ^ w6041 ;
  assign w6558 = w6033 ^ w6557 ;
  assign w6559 = \pi14 ^ w6556 ;
  assign w6560 = ( w6547 & w6558 ) | ( w6547 & w6559 ) | ( w6558 & w6559 ) ;
  assign w6561 = w6074 ^ w6545 ;
  assign w6562 = w6537 ^ w6561 ;
  assign w6563 = w6076 ^ w6536 ;
  assign w6564 = w6528 ^ w6563 ;
  assign w6565 = w6084 ^ w6527 ;
  assign w6566 = w6086 ^ w6565 ;
  assign w6567 = w592 & ~w5343 ;
  assign w6568 = w721 & w4905 ;
  assign w6569 = ( w592 & ~w6567 ) | ( w592 & w6568 ) | ( ~w6567 & w6568 ) ;
  assign w6570 = w381 | w5395 ;
  assign w6571 = w3435 & ~w6569 ;
  assign w6572 = ( w4908 & w6569 ) | ( w4908 & ~w6571 ) | ( w6569 & ~w6571 ) ;
  assign w6573 = ( ~w381 & w6570 ) | ( ~w381 & w6572 ) | ( w6570 & w6572 ) ;
  assign w6574 = \pi20 ^ w6573 ;
  assign w6575 = w6088 ^ w6526 ;
  assign w6576 = w6518 ^ w6575 ;
  assign w6577 = w6509 ^ w6517 ;
  assign w6578 = w6507 ^ w6577 ;
  assign w6579 = w6498 ^ w6506 ;
  assign w6580 = w6090 ^ w6579 ;
  assign w6581 = w1614 & ~w4143 ;
  assign w6582 = w1711 & w4052 ;
  assign w6583 = ( w1614 & ~w6581 ) | ( w1614 & w6582 ) | ( ~w6581 & w6582 ) ;
  assign w6584 = w4147 | w5085 ;
  assign w6585 = w1510 & ~w6583 ;
  assign w6586 = ( w3964 & w6583 ) | ( w3964 & ~w6585 ) | ( w6583 & ~w6585 ) ;
  assign w6587 = ( ~w5085 & w6584 ) | ( ~w5085 & w6586 ) | ( w6584 & w6586 ) ;
  assign w6588 = \pi26 ^ w6587 ;
  assign w6589 = w6092 ^ w6497 ;
  assign w6590 = w6102 ^ w6589 ;
  assign w6591 = w2059 | w3649 ;
  assign w6592 = w1976 & w3717 ;
  assign w6593 = ( ~w2059 & w6591 ) | ( ~w2059 & w6592 ) | ( w6591 & w6592 ) ;
  assign w6594 = w1939 | w3549 ;
  assign w6595 = w5748 | w6593 ;
  assign w6596 = ( w3448 & w6593 ) | ( w3448 & w6595 ) | ( w6593 & w6595 ) ;
  assign w6597 = ( ~w1939 & w6594 ) | ( ~w1939 & w6596 ) | ( w6594 & w6596 ) ;
  assign w6598 = \pi29 ^ w6597 ;
  assign w6599 = w1711 & ~w4143 ;
  assign w6600 = ~w1834 & w4052 ;
  assign w6601 = ( w1711 & ~w6599 ) | ( w1711 & w6600 ) | ( ~w6599 & w6600 ) ;
  assign w6602 = w4147 | w5433 ;
  assign w6603 = w1614 | w6601 ;
  assign w6604 = ( w3964 & w6601 ) | ( w3964 & w6603 ) | ( w6601 & w6603 ) ;
  assign w6605 = ( ~w5433 & w6602 ) | ( ~w5433 & w6604 ) | ( w6602 & w6604 ) ;
  assign w6606 = \pi26 ^ w6605 ;
  assign w6607 = ( ~w6590 & w6598 ) | ( ~w6590 & w6606 ) | ( w6598 & w6606 ) ;
  assign w6608 = ( w6580 & w6588 ) | ( w6580 & w6607 ) | ( w6588 & w6607 ) ;
  assign w6609 = w1264 | w4606 ;
  assign w6610 = w1205 & w4651 ;
  assign w6611 = ( ~w1264 & w6609 ) | ( ~w1264 & w6610 ) | ( w6609 & w6610 ) ;
  assign w6612 = w1085 & ~w4706 ;
  assign w6613 = w4533 | w6611 ;
  assign w6614 = ( w4609 & w6611 ) | ( w4609 & w6613 ) | ( w6611 & w6613 ) ;
  assign w6615 = ( w1085 & ~w6612 ) | ( w1085 & w6614 ) | ( ~w6612 & w6614 ) ;
  assign w6616 = \pi23 ^ w6615 ;
  assign w6617 = ( ~w6578 & w6608 ) | ( ~w6578 & w6616 ) | ( w6608 & w6616 ) ;
  assign w6618 = w883 | w4905 ;
  assign w6619 = w721 & w5343 ;
  assign w6620 = ( ~w883 & w6618 ) | ( ~w883 & w6619 ) | ( w6618 & w6619 ) ;
  assign w6621 = w592 & ~w5395 ;
  assign w6622 = w3421 | w6620 ;
  assign w6623 = ( w4908 & w6620 ) | ( w4908 & w6622 ) | ( w6620 & w6622 ) ;
  assign w6624 = ( w592 & ~w6621 ) | ( w592 & w6623 ) | ( ~w6621 & w6623 ) ;
  assign w6625 = \pi20 ^ w6624 ;
  assign w6626 = ( w6576 & w6617 ) | ( w6576 & w6625 ) | ( w6617 & w6625 ) ;
  assign w6627 = ( w6566 & w6574 ) | ( w6566 & w6626 ) | ( w6574 & w6626 ) ;
  assign w6628 = w3647 & ~w5494 ;
  assign w6629 = w3715 & w5710 ;
  assign w6630 = ( w3647 & ~w6628 ) | ( w3647 & w6629 ) | ( ~w6628 & w6629 ) ;
  assign w6631 = w3548 | w5948 ;
  assign w6632 = w3725 & ~w6630 ;
  assign w6633 = ( w5497 & w6630 ) | ( w5497 & ~w6632 ) | ( w6630 & ~w6632 ) ;
  assign w6634 = ( ~w3548 & w6631 ) | ( ~w3548 & w6633 ) | ( w6631 & w6633 ) ;
  assign w6635 = \pi17 ^ w6634 ;
  assign w6636 = ( w6564 & w6627 ) | ( w6564 & w6635 ) | ( w6627 & w6635 ) ;
  assign w6637 = ~w6043 & w6044 ;
  assign w6638 = w4049 | w6048 ;
  assign w6639 = ~w4142 & w6549 ;
  assign w6640 = ( ~w4049 & w6638 ) | ( ~w4049 & w6639 ) | ( w6638 & w6639 ) ;
  assign w6641 = w3962 | w6637 ;
  assign w6642 = w4152 & ~w6640 ;
  assign w6643 = ( w6045 & w6640 ) | ( w6045 & ~w6642 ) | ( w6640 & ~w6642 ) ;
  assign w6644 = ( ~w3962 & w6641 ) | ( ~w3962 & w6643 ) | ( w6641 & w6643 ) ;
  assign w6645 = \pi14 ^ w6644 ;
  assign w6646 = ( w6562 & w6636 ) | ( w6562 & w6645 ) | ( w6636 & w6645 ) ;
  assign w6647 = ~w4142 & w6048 ;
  assign w6648 = ( ~w4600 & w6637 ) | ( ~w4600 & w6647 ) | ( w6637 & w6647 ) ;
  assign w6649 = w6549 | w6648 ;
  assign w6650 = ( ~w3962 & w6648 ) | ( ~w3962 & w6649 ) | ( w6648 & w6649 ) ;
  assign w6651 = w6647 | w6650 ;
  assign w6652 = w6070 ^ w6546 ;
  assign w6653 = w6072 ^ w6652 ;
  assign w6654 = w4722 & ~w6651 ;
  assign w6655 = ( w6045 & w6651 ) | ( w6045 & ~w6654 ) | ( w6651 & ~w6654 ) ;
  assign w6656 = \pi14 ^ w6655 ;
  assign w6657 = ( w6646 & w6653 ) | ( w6646 & w6656 ) | ( w6653 & w6656 ) ;
  assign w6658 = \pi14 ^ w6547 ;
  assign w6659 = w6556 ^ w6658 ;
  assign w6660 = w6558 ^ w6659 ;
  assign w6661 = w6564 ^ w6635 ;
  assign w6662 = w6627 ^ w6661 ;
  assign w6663 = w3647 & ~w5710 ;
  assign w6664 = ~w3094 & w5494 ;
  assign w6665 = ( w3647 & ~w6663 ) | ( w3647 & w6664 ) | ( ~w6663 & w6664 ) ;
  assign w6666 = w3715 & ~w5948 ;
  assign w6667 = w4164 & ~w6665 ;
  assign w6668 = ( w5497 & w6665 ) | ( w5497 & ~w6667 ) | ( w6665 & ~w6667 ) ;
  assign w6669 = ( w3715 & ~w6666 ) | ( w3715 & w6668 ) | ( ~w6666 & w6668 ) ;
  assign w6670 = \pi17 ^ w6669 ;
  assign w6671 = w6574 ^ w6626 ;
  assign w6672 = w6566 ^ w6671 ;
  assign w6673 = w6576 ^ w6625 ;
  assign w6674 = w6617 ^ w6673 ;
  assign w6675 = w6578 ^ w6616 ;
  assign w6676 = w6608 ^ w6675 ;
  assign w6677 = w1264 | w4651 ;
  assign w6678 = w1399 & w4606 ;
  assign w6679 = ( ~w1264 & w6677 ) | ( ~w1264 & w6678 ) | ( w6677 & w6678 ) ;
  assign w6680 = w1205 & ~w4706 ;
  assign w6681 = w4864 & ~w6679 ;
  assign w6682 = ( w4609 & w6679 ) | ( w4609 & ~w6681 ) | ( w6679 & ~w6681 ) ;
  assign w6683 = ( w1205 & ~w6680 ) | ( w1205 & w6682 ) | ( ~w6680 & w6682 ) ;
  assign w6684 = \pi23 ^ w6683 ;
  assign w6685 = w6588 ^ w6607 ;
  assign w6686 = w6580 ^ w6685 ;
  assign w6687 = w6590 ^ w6606 ;
  assign w6688 = w6598 ^ w6687 ;
  assign w6689 = w6104 ^ w6496 ;
  assign w6690 = w6114 ^ w6689 ;
  assign w6691 = w2059 | w3717 ;
  assign w6692 = ~w2130 & w3649 ;
  assign w6693 = ( ~w2059 & w6691 ) | ( ~w2059 & w6692 ) | ( w6691 & w6692 ) ;
  assign w6694 = w1976 & ~w3549 ;
  assign w6695 = w5646 | w6693 ;
  assign w6696 = ( w3448 & w6693 ) | ( w3448 & w6695 ) | ( w6693 & w6695 ) ;
  assign w6697 = ( w1976 & ~w6694 ) | ( w1976 & w6696 ) | ( ~w6694 & w6696 ) ;
  assign w6698 = \pi29 ^ w6697 ;
  assign w6699 = w1939 | w4052 ;
  assign w6700 = ~w1834 & w4143 ;
  assign w6701 = ( ~w1939 & w6699 ) | ( ~w1939 & w6700 ) | ( w6699 & w6700 ) ;
  assign w6702 = ~w4147 & w5296 ;
  assign w6703 = w1711 | w6701 ;
  assign w6704 = ( w3964 & w6701 ) | ( w3964 & w6703 ) | ( w6701 & w6703 ) ;
  assign w6705 = ( w5296 & ~w6702 ) | ( w5296 & w6704 ) | ( ~w6702 & w6704 ) ;
  assign w6706 = \pi26 ^ w6705 ;
  assign w6707 = ( w6690 & w6698 ) | ( w6690 & w6706 ) | ( w6698 & w6706 ) ;
  assign w6708 = w1399 & ~w4651 ;
  assign w6709 = ~w1510 & w4606 ;
  assign w6710 = ( w1399 & ~w6708 ) | ( w1399 & w6709 ) | ( ~w6708 & w6709 ) ;
  assign w6711 = w1264 | w4706 ;
  assign w6712 = w4852 & ~w6710 ;
  assign w6713 = ( w4609 & w6710 ) | ( w4609 & ~w6712 ) | ( w6710 & ~w6712 ) ;
  assign w6714 = ( ~w1264 & w6711 ) | ( ~w1264 & w6713 ) | ( w6711 & w6713 ) ;
  assign w6715 = \pi23 ^ w6714 ;
  assign w6716 = ( ~w6688 & w6707 ) | ( ~w6688 & w6715 ) | ( w6707 & w6715 ) ;
  assign w6717 = ( w6684 & w6686 ) | ( w6684 & w6716 ) | ( w6686 & w6716 ) ;
  assign w6718 = w883 | w5343 ;
  assign w6719 = w979 & w4905 ;
  assign w6720 = ( ~w883 & w6718 ) | ( ~w883 & w6719 ) | ( w6718 & w6719 ) ;
  assign w6721 = w721 & ~w5395 ;
  assign w6722 = w4257 & ~w6720 ;
  assign w6723 = ( w4908 & w6720 ) | ( w4908 & ~w6722 ) | ( w6720 & ~w6722 ) ;
  assign w6724 = ( w721 & ~w6721 ) | ( w721 & w6723 ) | ( ~w6721 & w6723 ) ;
  assign w6725 = \pi20 ^ w6724 ;
  assign w6726 = ( ~w6676 & w6717 ) | ( ~w6676 & w6725 ) | ( w6717 & w6725 ) ;
  assign w6727 = w381 | w5494 ;
  assign w6728 = ~w3094 & w5710 ;
  assign w6729 = ( ~w381 & w6727 ) | ( ~w381 & w6728 ) | ( w6727 & w6728 ) ;
  assign w6730 = w3647 & ~w5948 ;
  assign w6731 = w3810 | w6729 ;
  assign w6732 = ( w5497 & w6729 ) | ( w5497 & w6731 ) | ( w6729 & w6731 ) ;
  assign w6733 = ( w3647 & ~w6730 ) | ( w3647 & w6732 ) | ( ~w6730 & w6732 ) ;
  assign w6734 = \pi17 ^ w6733 ;
  assign w6735 = ( w6674 & w6726 ) | ( w6674 & w6734 ) | ( w6726 & w6734 ) ;
  assign w6736 = ( w6670 & w6672 ) | ( w6670 & w6735 ) | ( w6672 & w6735 ) ;
  assign w6737 = w4049 | w6549 ;
  assign w6738 = w3907 & w6048 ;
  assign w6739 = ( ~w4049 & w6737 ) | ( ~w4049 & w6738 ) | ( w6737 & w6738 ) ;
  assign w6740 = w4142 | w6637 ;
  assign w6741 = w4563 | w6739 ;
  assign w6742 = ( w6045 & w6739 ) | ( w6045 & w6741 ) | ( w6739 & w6741 ) ;
  assign w6743 = ( ~w4142 & w6740 ) | ( ~w4142 & w6742 ) | ( w6740 & w6742 ) ;
  assign w6744 = \pi14 ^ w6743 ;
  assign w6745 = ( w6662 & w6736 ) | ( w6662 & w6744 ) | ( w6736 & w6744 ) ;
  assign w6746 = ( \pi09 & ~\pi10 ) | ( \pi09 & \pi11 ) | ( ~\pi10 & \pi11 ) ;
  assign w6747 = ( \pi08 & \pi09 ) | ( \pi08 & w6746 ) | ( \pi09 & w6746 ) ;
  assign w6748 = w6746 ^ w6747 ;
  assign w6749 = \pi10 ^ \pi11 ;
  assign w6750 = \pi08 ^ \pi09 ;
  assign w6751 = w6749 & w6750 ;
  assign w6752 = ~w4600 & w6748 ;
  assign w6753 = w6751 | w6752 ;
  assign w6754 = ( ~w4603 & w6752 ) | ( ~w4603 & w6753 ) | ( w6752 & w6753 ) ;
  assign w6755 = \pi11 ^ w6754 ;
  assign w6756 = w6562 ^ w6645 ;
  assign w6757 = w6636 ^ w6756 ;
  assign w6758 = ( w6745 & w6755 ) | ( w6745 & w6757 ) | ( w6755 & w6757 ) ;
  assign w6759 = w4722 & w6045 ;
  assign w6760 = ( w6045 & w6651 ) | ( w6045 & ~w6759 ) | ( w6651 & ~w6759 ) ;
  assign w6761 = w6646 ^ w6760 ;
  assign w6762 = \pi14 ^ w6653 ;
  assign w6763 = w6761 ^ w6762 ;
  assign w6764 = w6755 ^ w6757 ;
  assign w6765 = w6745 ^ w6764 ;
  assign w6766 = w6670 ^ w6735 ;
  assign w6767 = w6672 ^ w6766 ;
  assign w6768 = w3548 | w6048 ;
  assign w6769 = w3907 & w6549 ;
  assign w6770 = ( ~w3548 & w6768 ) | ( ~w3548 & w6769 ) | ( w6768 & w6769 ) ;
  assign w6771 = w4049 | w6637 ;
  assign w6772 = w4622 & ~w6770 ;
  assign w6773 = ( w6045 & w6770 ) | ( w6045 & ~w6772 ) | ( w6770 & ~w6772 ) ;
  assign w6774 = ( ~w4049 & w6771 ) | ( ~w4049 & w6773 ) | ( w6771 & w6773 ) ;
  assign w6775 = \pi14 ^ w6774 ;
  assign w6776 = w6674 ^ w6734 ;
  assign w6777 = w6726 ^ w6776 ;
  assign w6778 = w6676 ^ w6725 ;
  assign w6779 = w6717 ^ w6778 ;
  assign w6780 = w6684 ^ w6716 ;
  assign w6781 = w6686 ^ w6780 ;
  assign w6782 = w979 & ~w5343 ;
  assign w6783 = w1085 & w4905 ;
  assign w6784 = ( w979 & ~w6782 ) | ( w979 & w6783 ) | ( ~w6782 & w6783 ) ;
  assign w6785 = w883 | w5395 ;
  assign w6786 = w4273 & ~w6784 ;
  assign w6787 = ( w4908 & w6784 ) | ( w4908 & ~w6786 ) | ( w6784 & ~w6786 ) ;
  assign w6788 = ( ~w883 & w6785 ) | ( ~w883 & w6787 ) | ( w6785 & w6787 ) ;
  assign w6789 = \pi20 ^ w6788 ;
  assign w6790 = w6688 ^ w6715 ;
  assign w6791 = w6707 ^ w6790 ;
  assign w6792 = w6690 ^ w6706 ;
  assign w6793 = w6698 ^ w6792 ;
  assign w6794 = w6172 ^ w6486 ;
  assign w6795 = w6162 ^ w6794 ;
  assign w6796 = w2273 & ~w3649 ;
  assign w6797 = ~w2235 & w3717 ;
  assign w6798 = ( w2273 & ~w6796 ) | ( w2273 & w6797 ) | ( ~w6796 & w6797 ) ;
  assign w6799 = w2130 | w3549 ;
  assign w6800 = w6094 | w6798 ;
  assign w6801 = ( w3448 & w6798 ) | ( w3448 & w6800 ) | ( w6798 & w6800 ) ;
  assign w6802 = ( ~w2130 & w6799 ) | ( ~w2130 & w6801 ) | ( w6799 & w6801 ) ;
  assign w6803 = \pi29 ^ w6802 ;
  assign w6804 = w6227 ^ w6485 ;
  assign w6805 = w6217 ^ w6804 ;
  assign w6806 = w2273 & ~w3717 ;
  assign w6807 = w2391 & w3649 ;
  assign w6808 = ( w2273 & ~w6806 ) | ( w2273 & w6807 ) | ( ~w6806 & w6807 ) ;
  assign w6809 = w2235 | w3549 ;
  assign w6810 = w6106 & ~w6808 ;
  assign w6811 = ( w3448 & w6808 ) | ( w3448 & ~w6810 ) | ( w6808 & ~w6810 ) ;
  assign w6812 = ( ~w2235 & w6809 ) | ( ~w2235 & w6811 ) | ( w6809 & w6811 ) ;
  assign w6813 = \pi29 ^ w6812 ;
  assign w6814 = w2391 & ~w3717 ;
  assign w6815 = w2500 & w3649 ;
  assign w6816 = ( w2391 & ~w6814 ) | ( w2391 & w6815 ) | ( ~w6814 & w6815 ) ;
  assign w6817 = w2273 & ~w3549 ;
  assign w6818 = w5880 | w6816 ;
  assign w6819 = ( w3448 & w6816 ) | ( w3448 & w6818 ) | ( w6816 & w6818 ) ;
  assign w6820 = ( w2273 & ~w6817 ) | ( w2273 & w6819 ) | ( ~w6817 & w6819 ) ;
  assign w6821 = \pi29 ^ w6820 ;
  assign w6822 = w6290 ^ w6484 ;
  assign w6823 = w6280 ^ w6822 ;
  assign w6824 = w2578 | w3649 ;
  assign w6825 = w2500 & w3717 ;
  assign w6826 = ( ~w2578 & w6824 ) | ( ~w2578 & w6825 ) | ( w6824 & w6825 ) ;
  assign w6827 = w2391 & ~w3549 ;
  assign w6828 = w6164 & ~w6826 ;
  assign w6829 = ( w3448 & w6826 ) | ( w3448 & ~w6828 ) | ( w6826 & ~w6828 ) ;
  assign w6830 = ( w2391 & ~w6827 ) | ( w2391 & w6829 ) | ( ~w6827 & w6829 ) ;
  assign w6831 = \pi29 ^ w6830 ;
  assign w6832 = w6346 ^ w6483 ;
  assign w6833 = w6333 ^ w6832 ;
  assign w6834 = w2578 | w3717 ;
  assign w6835 = ~w2653 & w3649 ;
  assign w6836 = ( ~w2578 & w6834 ) | ( ~w2578 & w6835 ) | ( w6834 & w6835 ) ;
  assign w6837 = w2500 & ~w3549 ;
  assign w6838 = w6219 | w6836 ;
  assign w6839 = ( w3448 & w6836 ) | ( w3448 & w6838 ) | ( w6836 & w6838 ) ;
  assign w6840 = ( w2500 & ~w6837 ) | ( w2500 & w6839 ) | ( ~w6837 & w6839 ) ;
  assign w6841 = \pi29 ^ w6840 ;
  assign w6842 = w6469 ^ w6482 ;
  assign w6843 = w6401 ^ w6842 ;
  assign w6844 = w2694 | w3649 ;
  assign w6845 = ~w2653 & w3717 ;
  assign w6846 = ( ~w2694 & w6844 ) | ( ~w2694 & w6845 ) | ( w6844 & w6845 ) ;
  assign w6847 = w2578 | w3549 ;
  assign w6848 = w6282 & ~w6846 ;
  assign w6849 = ( w3448 & w6846 ) | ( w3448 & ~w6848 ) | ( w6846 & ~w6848 ) ;
  assign w6850 = ( ~w2578 & w6847 ) | ( ~w2578 & w6849 ) | ( w6847 & w6849 ) ;
  assign w6851 = \pi29 ^ w6850 ;
  assign w6852 = w6455 ^ w6468 ;
  assign w6853 = w2805 & ~w3649 ;
  assign w6854 = ~w2694 & w3717 ;
  assign w6855 = ( w2805 & ~w6853 ) | ( w2805 & w6854 ) | ( ~w6853 & w6854 ) ;
  assign w6856 = w2653 | w3549 ;
  assign w6857 = w6338 & ~w6855 ;
  assign w6858 = ( w3448 & w6855 ) | ( w3448 & ~w6857 ) | ( w6855 & ~w6857 ) ;
  assign w6859 = ( ~w2653 & w6856 ) | ( ~w2653 & w6858 ) | ( w6856 & w6858 ) ;
  assign w6860 = \pi29 ^ w6859 ;
  assign w6861 = ( \pi29 & \pi30 ) | ( \pi29 & ~w2871 ) | ( \pi30 & ~w2871 ) ;
  assign w6862 = \pi29 & \pi30 ;
  assign w6863 = \pi31 ^ w2973 ;
  assign w6864 = ( \pi31 & w6862 ) | ( \pi31 & w6863 ) | ( w6862 & w6863 ) ;
  assign w6865 = w6861 ^ w6864 ;
  assign w6866 = ( \pi26 & \pi27 ) | ( \pi26 & ~\pi29 ) | ( \pi27 & ~\pi29 ) ;
  assign w6867 = \pi29 & w2973 ;
  assign w6868 = w2871 & w6867 ;
  assign w6869 = ( \pi26 & \pi27 ) | ( \pi26 & ~w6868 ) | ( \pi27 & ~w6868 ) ;
  assign w6870 = ( \pi28 & \pi29 ) | ( \pi28 & ~w6869 ) | ( \pi29 & ~w6869 ) ;
  assign w6871 = ( \pi28 & ~w6867 ) | ( \pi28 & w6869 ) | ( ~w6867 & w6869 ) ;
  assign w6872 = ( w6866 & w6870 ) | ( w6866 & ~w6871 ) | ( w6870 & ~w6871 ) ;
  assign w6873 = w2973 | w3649 ;
  assign w6874 = ~w2871 & w3717 ;
  assign w6875 = ( ~w2973 & w6873 ) | ( ~w2973 & w6874 ) | ( w6873 & w6874 ) ;
  assign w6876 = w2805 & ~w3549 ;
  assign w6877 = w6457 | w6875 ;
  assign w6878 = ( w3448 & w6875 ) | ( w3448 & w6877 ) | ( w6875 & w6877 ) ;
  assign w6879 = ( w2805 & ~w6876 ) | ( w2805 & w6878 ) | ( ~w6876 & w6878 ) ;
  assign w6880 = \pi29 ^ w6879 ;
  assign w6881 = w6872 & w6880 ;
  assign w6882 = w2805 & ~w3717 ;
  assign w6883 = ~w2871 & w3649 ;
  assign w6884 = ( w2805 & ~w6882 ) | ( w2805 & w6883 ) | ( ~w6882 & w6883 ) ;
  assign w6885 = w2694 | w3549 ;
  assign w6886 = w6473 | w6884 ;
  assign w6887 = ( w3448 & w6884 ) | ( w3448 & w6886 ) | ( w6884 & w6886 ) ;
  assign w6888 = ( ~w2694 & w6885 ) | ( ~w2694 & w6887 ) | ( w6885 & w6887 ) ;
  assign w6889 = \pi29 ^ w6888 ;
  assign w6890 = w36 & ~w2973 ;
  assign w6891 = ( w6881 & w6889 ) | ( w6881 & w6890 ) | ( w6889 & w6890 ) ;
  assign w6892 = ( w6860 & w6865 ) | ( w6860 & w6891 ) | ( w6865 & w6891 ) ;
  assign w6893 = ( w6851 & ~w6852 ) | ( w6851 & w6892 ) | ( ~w6852 & w6892 ) ;
  assign w6894 = ( w6841 & ~w6843 ) | ( w6841 & w6893 ) | ( ~w6843 & w6893 ) ;
  assign w6895 = ( w6831 & w6833 ) | ( w6831 & w6894 ) | ( w6833 & w6894 ) ;
  assign w6896 = ( w6821 & ~w6823 ) | ( w6821 & w6895 ) | ( ~w6823 & w6895 ) ;
  assign w6897 = ( w6805 & w6813 ) | ( w6805 & w6896 ) | ( w6813 & w6896 ) ;
  assign w6898 = ( w6795 & w6803 ) | ( w6795 & w6897 ) | ( w6803 & w6897 ) ;
  assign w6899 = w6116 ^ w6495 ;
  assign w6900 = w6487 ^ w6899 ;
  assign w6901 = w1939 | w4143 ;
  assign w6902 = w1976 & w4052 ;
  assign w6903 = ( ~w1939 & w6901 ) | ( ~w1939 & w6902 ) | ( w6901 & w6902 ) ;
  assign w6904 = w4147 | w5659 ;
  assign w6905 = w1834 & ~w6903 ;
  assign w6906 = ( w3964 & w6903 ) | ( w3964 & ~w6905 ) | ( w6903 & ~w6905 ) ;
  assign w6907 = ( ~w5659 & w6904 ) | ( ~w5659 & w6906 ) | ( w6904 & w6906 ) ;
  assign w6908 = \pi26 ^ w6907 ;
  assign w6909 = ( w6898 & w6900 ) | ( w6898 & w6908 ) | ( w6900 & w6908 ) ;
  assign w6910 = w1614 & ~w4606 ;
  assign w6911 = ~w1510 & w4651 ;
  assign w6912 = ( w1614 & ~w6910 ) | ( w1614 & w6911 ) | ( ~w6910 & w6911 ) ;
  assign w6913 = w1399 & ~w4706 ;
  assign w6914 = w5069 & ~w6912 ;
  assign w6915 = ( w4609 & w6912 ) | ( w4609 & ~w6914 ) | ( w6912 & ~w6914 ) ;
  assign w6916 = ( w1399 & ~w6913 ) | ( w1399 & w6915 ) | ( ~w6913 & w6915 ) ;
  assign w6917 = \pi23 ^ w6916 ;
  assign w6918 = ( w6793 & w6909 ) | ( w6793 & w6917 ) | ( w6909 & w6917 ) ;
  assign w6919 = w1085 & ~w5343 ;
  assign w6920 = w1205 & w4905 ;
  assign w6921 = ( w1085 & ~w6919 ) | ( w1085 & w6920 ) | ( ~w6919 & w6920 ) ;
  assign w6922 = w979 & ~w5395 ;
  assign w6923 = w4666 | w6921 ;
  assign w6924 = ( w4908 & w6921 ) | ( w4908 & w6923 ) | ( w6921 & w6923 ) ;
  assign w6925 = ( w979 & ~w6922 ) | ( w979 & w6924 ) | ( ~w6922 & w6924 ) ;
  assign w6926 = \pi20 ^ w6925 ;
  assign w6927 = ( ~w6791 & w6918 ) | ( ~w6791 & w6926 ) | ( w6918 & w6926 ) ;
  assign w6928 = ( w6781 & w6789 ) | ( w6781 & w6927 ) | ( w6789 & w6927 ) ;
  assign w6929 = w381 | w5710 ;
  assign w6930 = w592 & w5494 ;
  assign w6931 = ( ~w381 & w6929 ) | ( ~w381 & w6930 ) | ( w6929 & w6930 ) ;
  assign w6932 = w3094 | w5948 ;
  assign w6933 = w3096 | w6931 ;
  assign w6934 = ( w5497 & w6931 ) | ( w5497 & w6933 ) | ( w6931 & w6933 ) ;
  assign w6935 = ( ~w3094 & w6932 ) | ( ~w3094 & w6934 ) | ( w6932 & w6934 ) ;
  assign w6936 = \pi17 ^ w6935 ;
  assign w6937 = ( ~w6779 & w6928 ) | ( ~w6779 & w6936 ) | ( w6928 & w6936 ) ;
  assign w6938 = w3548 | w6549 ;
  assign w6939 = w3715 & w6048 ;
  assign w6940 = ( ~w3548 & w6938 ) | ( ~w3548 & w6939 ) | ( w6938 & w6939 ) ;
  assign w6941 = w3907 & ~w6637 ;
  assign w6942 = w3913 & ~w6940 ;
  assign w6943 = ( w6045 & w6940 ) | ( w6045 & ~w6942 ) | ( w6940 & ~w6942 ) ;
  assign w6944 = ( w3907 & ~w6941 ) | ( w3907 & w6943 ) | ( ~w6941 & w6943 ) ;
  assign w6945 = \pi14 ^ w6944 ;
  assign w6946 = ( w6777 & w6937 ) | ( w6777 & w6945 ) | ( w6937 & w6945 ) ;
  assign w6947 = ( w6767 & w6775 ) | ( w6767 & w6946 ) | ( w6775 & w6946 ) ;
  assign w6948 = ( \pi08 & \pi09 ) | ( \pi08 & \pi10 ) | ( \pi09 & \pi10 ) ;
  assign w6949 = \pi10 ^ w6948 ;
  assign w6950 = ~w4600 & w6949 ;
  assign w6951 = ( w3962 & w6551 ) | ( w3962 & w6751 ) | ( w6551 & w6751 ) ;
  assign w6952 = w3962 | w6748 ;
  assign w6953 = ( ~w3962 & w6951 ) | ( ~w3962 & w6952 ) | ( w6951 & w6952 ) ;
  assign w6954 = ( ~w6555 & w6950 ) | ( ~w6555 & w6953 ) | ( w6950 & w6953 ) ;
  assign w6955 = w6662 ^ w6744 ;
  assign w6956 = w6736 ^ w6955 ;
  assign w6957 = \pi11 ^ w6954 ;
  assign w6958 = ( w6947 & w6956 ) | ( w6947 & w6957 ) | ( w6956 & w6957 ) ;
  assign w6959 = w6777 ^ w6945 ;
  assign w6960 = w6937 ^ w6959 ;
  assign w6961 = w6779 ^ w6936 ;
  assign w6962 = w6928 ^ w6961 ;
  assign w6963 = w592 & ~w5710 ;
  assign w6964 = w721 & w5494 ;
  assign w6965 = ( w592 & ~w6963 ) | ( w592 & w6964 ) | ( ~w6963 & w6964 ) ;
  assign w6966 = w381 | w5948 ;
  assign w6967 = w3435 & ~w6965 ;
  assign w6968 = ( w5497 & w6965 ) | ( w5497 & ~w6967 ) | ( w6965 & ~w6967 ) ;
  assign w6969 = ( ~w381 & w6966 ) | ( ~w381 & w6968 ) | ( w6966 & w6968 ) ;
  assign w6970 = \pi17 ^ w6969 ;
  assign w6971 = w6789 ^ w6927 ;
  assign w6972 = w6781 ^ w6971 ;
  assign w6973 = w6791 ^ w6926 ;
  assign w6974 = w6918 ^ w6973 ;
  assign w6975 = w6793 ^ w6917 ;
  assign w6976 = w6909 ^ w6975 ;
  assign w6977 = w6803 ^ w6897 ;
  assign w6978 = w6795 ^ w6977 ;
  assign w6979 = w2059 | w4052 ;
  assign w6980 = w1976 & w4143 ;
  assign w6981 = ( ~w2059 & w6979 ) | ( ~w2059 & w6980 ) | ( w6979 & w6980 ) ;
  assign w6982 = ~w4147 & w5748 ;
  assign w6983 = w1939 & ~w6981 ;
  assign w6984 = ( w3964 & w6981 ) | ( w3964 & ~w6983 ) | ( w6981 & ~w6983 ) ;
  assign w6985 = ( w5748 & ~w6982 ) | ( w5748 & w6984 ) | ( ~w6982 & w6984 ) ;
  assign w6986 = \pi26 ^ w6985 ;
  assign w6987 = w6813 ^ w6896 ;
  assign w6988 = w6805 ^ w6987 ;
  assign w6989 = w2059 | w4143 ;
  assign w6990 = ~w2130 & w4052 ;
  assign w6991 = ( ~w2059 & w6989 ) | ( ~w2059 & w6990 ) | ( w6989 & w6990 ) ;
  assign w6992 = ~w4147 & w5646 ;
  assign w6993 = w1976 | w6991 ;
  assign w6994 = ( w3964 & w6991 ) | ( w3964 & w6993 ) | ( w6991 & w6993 ) ;
  assign w6995 = ( w5646 & ~w6992 ) | ( w5646 & w6994 ) | ( ~w6992 & w6994 ) ;
  assign w6996 = \pi26 ^ w6995 ;
  assign w6997 = w6821 ^ w6895 ;
  assign w6998 = w6823 ^ w6997 ;
  assign w6999 = w2130 | w4143 ;
  assign w7000 = ~w2235 & w4052 ;
  assign w7001 = ( ~w2130 & w6999 ) | ( ~w2130 & w7000 ) | ( w6999 & w7000 ) ;
  assign w7002 = w4147 | w5896 ;
  assign w7003 = w2059 & ~w7001 ;
  assign w7004 = ( w3964 & w7001 ) | ( w3964 & ~w7003 ) | ( w7001 & ~w7003 ) ;
  assign w7005 = ( ~w5896 & w7002 ) | ( ~w5896 & w7004 ) | ( w7002 & w7004 ) ;
  assign w7006 = \pi26 ^ w7005 ;
  assign w7007 = w6831 ^ w6894 ;
  assign w7008 = w6833 ^ w7007 ;
  assign w7009 = w2273 & ~w4052 ;
  assign w7010 = ~w2235 & w4143 ;
  assign w7011 = ( w2273 & ~w7009 ) | ( w2273 & w7010 ) | ( ~w7009 & w7010 ) ;
  assign w7012 = ~w4147 & w6094 ;
  assign w7013 = w2130 & ~w7011 ;
  assign w7014 = ( w3964 & w7011 ) | ( w3964 & ~w7013 ) | ( w7011 & ~w7013 ) ;
  assign w7015 = ( w6094 & ~w7012 ) | ( w6094 & w7014 ) | ( ~w7012 & w7014 ) ;
  assign w7016 = \pi26 ^ w7015 ;
  assign w7017 = w6841 ^ w6893 ;
  assign w7018 = w6843 ^ w7017 ;
  assign w7019 = w2273 & ~w4143 ;
  assign w7020 = w2391 & w4052 ;
  assign w7021 = ( w2273 & ~w7019 ) | ( w2273 & w7020 ) | ( ~w7019 & w7020 ) ;
  assign w7022 = w4147 | w6106 ;
  assign w7023 = w2235 & ~w7021 ;
  assign w7024 = ( w3964 & w7021 ) | ( w3964 & ~w7023 ) | ( w7021 & ~w7023 ) ;
  assign w7025 = ( ~w6106 & w7022 ) | ( ~w6106 & w7024 ) | ( w7022 & w7024 ) ;
  assign w7026 = \pi26 ^ w7025 ;
  assign w7027 = w6851 ^ w6892 ;
  assign w7028 = w6852 ^ w7027 ;
  assign w7029 = w2391 & ~w4143 ;
  assign w7030 = w2500 & w4052 ;
  assign w7031 = ( w2391 & ~w7029 ) | ( w2391 & w7030 ) | ( ~w7029 & w7030 ) ;
  assign w7032 = ~w4147 & w5880 ;
  assign w7033 = w2273 | w7031 ;
  assign w7034 = ( w3964 & w7031 ) | ( w3964 & w7033 ) | ( w7031 & w7033 ) ;
  assign w7035 = ( w5880 & ~w7032 ) | ( w5880 & w7034 ) | ( ~w7032 & w7034 ) ;
  assign w7036 = \pi26 ^ w7035 ;
  assign w7037 = w6860 ^ w6891 ;
  assign w7038 = w6865 ^ w7037 ;
  assign w7039 = w2578 | w4052 ;
  assign w7040 = w2500 & w4143 ;
  assign w7041 = ( ~w2578 & w7039 ) | ( ~w2578 & w7040 ) | ( w7039 & w7040 ) ;
  assign w7042 = w4147 | w6164 ;
  assign w7043 = w2391 | w7041 ;
  assign w7044 = ( w3964 & w7041 ) | ( w3964 & w7043 ) | ( w7041 & w7043 ) ;
  assign w7045 = ( ~w6164 & w7042 ) | ( ~w6164 & w7044 ) | ( w7042 & w7044 ) ;
  assign w7046 = \pi26 ^ w7045 ;
  assign w7047 = w2578 | w4143 ;
  assign w7048 = ~w2653 & w4052 ;
  assign w7049 = ( ~w2578 & w7047 ) | ( ~w2578 & w7048 ) | ( w7047 & w7048 ) ;
  assign w7050 = ~w4147 & w6219 ;
  assign w7051 = w2500 | w7049 ;
  assign w7052 = ( w3964 & w7049 ) | ( w3964 & w7051 ) | ( w7049 & w7051 ) ;
  assign w7053 = ( w6219 & ~w7050 ) | ( w6219 & w7052 ) | ( ~w7050 & w7052 ) ;
  assign w7054 = \pi26 ^ w7053 ;
  assign w7055 = w6881 ^ w6889 ;
  assign w7056 = w6890 ^ w7055 ;
  assign w7057 = w2694 | w4052 ;
  assign w7058 = ~w2653 & w4143 ;
  assign w7059 = ( ~w2694 & w7057 ) | ( ~w2694 & w7058 ) | ( w7057 & w7058 ) ;
  assign w7060 = w4147 | w6282 ;
  assign w7061 = w2578 & ~w7059 ;
  assign w7062 = ( w3964 & w7059 ) | ( w3964 & ~w7061 ) | ( w7059 & ~w7061 ) ;
  assign w7063 = ( ~w6282 & w7060 ) | ( ~w6282 & w7062 ) | ( w7060 & w7062 ) ;
  assign w7064 = \pi26 ^ w7063 ;
  assign w7065 = w6872 ^ w6880 ;
  assign w7066 = ( \pi26 & \pi27 ) | ( \pi26 & ~w2871 ) | ( \pi27 & ~w2871 ) ;
  assign w7067 = \pi26 & \pi27 ;
  assign w7068 = w2973 ^ w7067 ;
  assign w7069 = ( \pi28 & w7067 ) | ( \pi28 & ~w7068 ) | ( w7067 & ~w7068 ) ;
  assign w7070 = w7066 ^ w7069 ;
  assign w7071 = w2805 & ~w4052 ;
  assign w7072 = ~w2694 & w4143 ;
  assign w7073 = ( w2805 & ~w7071 ) | ( w2805 & w7072 ) | ( ~w7071 & w7072 ) ;
  assign w7074 = w4147 | w6338 ;
  assign w7075 = w2653 & ~w7073 ;
  assign w7076 = ( w3964 & w7073 ) | ( w3964 & ~w7075 ) | ( w7073 & ~w7075 ) ;
  assign w7077 = ( ~w6338 & w7074 ) | ( ~w6338 & w7076 ) | ( w7074 & w7076 ) ;
  assign w7078 = \pi26 ^ w7077 ;
  assign w7079 = ( \pi23 & \pi24 ) | ( \pi23 & ~\pi26 ) | ( \pi24 & ~\pi26 ) ;
  assign w7080 = \pi26 & w2973 ;
  assign w7081 = w2871 & w7080 ;
  assign w7082 = ( \pi23 & \pi24 ) | ( \pi23 & ~w7081 ) | ( \pi24 & ~w7081 ) ;
  assign w7083 = ( \pi25 & \pi26 ) | ( \pi25 & ~w7082 ) | ( \pi26 & ~w7082 ) ;
  assign w7084 = ( \pi25 & ~w7080 ) | ( \pi25 & w7082 ) | ( ~w7080 & w7082 ) ;
  assign w7085 = ( w7079 & w7083 ) | ( w7079 & ~w7084 ) | ( w7083 & ~w7084 ) ;
  assign w7086 = w2973 | w4052 ;
  assign w7087 = ~w2871 & w4143 ;
  assign w7088 = ( ~w2973 & w7086 ) | ( ~w2973 & w7087 ) | ( w7086 & w7087 ) ;
  assign w7089 = ~w4147 & w6457 ;
  assign w7090 = w2805 | w7088 ;
  assign w7091 = ( w3964 & w7088 ) | ( w3964 & w7090 ) | ( w7088 & w7090 ) ;
  assign w7092 = ( w6457 & ~w7089 ) | ( w6457 & w7091 ) | ( ~w7089 & w7091 ) ;
  assign w7093 = \pi26 ^ w7092 ;
  assign w7094 = w7085 & w7093 ;
  assign w7095 = w2805 & ~w4143 ;
  assign w7096 = ~w2871 & w4052 ;
  assign w7097 = ( w2805 & ~w7095 ) | ( w2805 & w7096 ) | ( ~w7095 & w7096 ) ;
  assign w7098 = ~w4147 & w6473 ;
  assign w7099 = w2694 & ~w7097 ;
  assign w7100 = ( w3964 & w7097 ) | ( w3964 & ~w7099 ) | ( w7097 & ~w7099 ) ;
  assign w7101 = ( w6473 & ~w7098 ) | ( w6473 & w7100 ) | ( ~w7098 & w7100 ) ;
  assign w7102 = \pi26 ^ w7101 ;
  assign w7103 = ~w2973 & w3447 ;
  assign w7104 = ( w7094 & w7102 ) | ( w7094 & w7103 ) | ( w7102 & w7103 ) ;
  assign w7105 = ( w7070 & w7078 ) | ( w7070 & w7104 ) | ( w7078 & w7104 ) ;
  assign w7106 = ( w7064 & w7065 ) | ( w7064 & w7105 ) | ( w7065 & w7105 ) ;
  assign w7107 = ( w7054 & w7056 ) | ( w7054 & w7106 ) | ( w7056 & w7106 ) ;
  assign w7108 = ( w7038 & w7046 ) | ( w7038 & w7107 ) | ( w7046 & w7107 ) ;
  assign w7109 = ( ~w7028 & w7036 ) | ( ~w7028 & w7108 ) | ( w7036 & w7108 ) ;
  assign w7110 = ( ~w7018 & w7026 ) | ( ~w7018 & w7109 ) | ( w7026 & w7109 ) ;
  assign w7111 = ( w7008 & w7016 ) | ( w7008 & w7110 ) | ( w7016 & w7110 ) ;
  assign w7112 = ( ~w6998 & w7006 ) | ( ~w6998 & w7111 ) | ( w7006 & w7111 ) ;
  assign w7113 = ( w6988 & w6996 ) | ( w6988 & w7112 ) | ( w6996 & w7112 ) ;
  assign w7114 = ( w6978 & w6986 ) | ( w6978 & w7113 ) | ( w6986 & w7113 ) ;
  assign w7115 = w6898 ^ w6908 ;
  assign w7116 = w6900 ^ w7115 ;
  assign w7117 = w1614 & ~w4651 ;
  assign w7118 = w1711 & w4606 ;
  assign w7119 = ( w1614 & ~w7117 ) | ( w1614 & w7118 ) | ( ~w7117 & w7118 ) ;
  assign w7120 = w1510 | w4706 ;
  assign w7121 = w5085 & ~w7119 ;
  assign w7122 = ( w4609 & w7119 ) | ( w4609 & ~w7121 ) | ( w7119 & ~w7121 ) ;
  assign w7123 = ( ~w1510 & w7120 ) | ( ~w1510 & w7122 ) | ( w7120 & w7122 ) ;
  assign w7124 = \pi23 ^ w7123 ;
  assign w7125 = ( w7114 & w7116 ) | ( w7114 & w7124 ) | ( w7116 & w7124 ) ;
  assign w7126 = w1264 | w4905 ;
  assign w7127 = w1205 & w5343 ;
  assign w7128 = ( ~w1264 & w7126 ) | ( ~w1264 & w7127 ) | ( w7126 & w7127 ) ;
  assign w7129 = w1085 & ~w5395 ;
  assign w7130 = w4533 | w7128 ;
  assign w7131 = ( w4908 & w7128 ) | ( w4908 & w7130 ) | ( w7128 & w7130 ) ;
  assign w7132 = ( w1085 & ~w7129 ) | ( w1085 & w7131 ) | ( ~w7129 & w7131 ) ;
  assign w7133 = \pi20 ^ w7132 ;
  assign w7134 = ( w6976 & w7125 ) | ( w6976 & w7133 ) | ( w7125 & w7133 ) ;
  assign w7135 = w883 | w5494 ;
  assign w7136 = w721 & w5710 ;
  assign w7137 = ( ~w883 & w7135 ) | ( ~w883 & w7136 ) | ( w7135 & w7136 ) ;
  assign w7138 = w592 & ~w5948 ;
  assign w7139 = w3421 | w7137 ;
  assign w7140 = ( w5497 & w7137 ) | ( w5497 & w7139 ) | ( w7137 & w7139 ) ;
  assign w7141 = ( w592 & ~w7138 ) | ( w592 & w7140 ) | ( ~w7138 & w7140 ) ;
  assign w7142 = \pi17 ^ w7141 ;
  assign w7143 = ( ~w6974 & w7134 ) | ( ~w6974 & w7142 ) | ( w7134 & w7142 ) ;
  assign w7144 = ( w6970 & w6972 ) | ( w6970 & w7143 ) | ( w6972 & w7143 ) ;
  assign w7145 = w3647 & ~w6048 ;
  assign w7146 = w3715 & w6549 ;
  assign w7147 = ( w3647 & ~w7145 ) | ( w3647 & w7146 ) | ( ~w7145 & w7146 ) ;
  assign w7148 = w3548 | w6637 ;
  assign w7149 = w3725 & ~w7147 ;
  assign w7150 = ( w6045 & w7147 ) | ( w6045 & ~w7149 ) | ( w7147 & ~w7149 ) ;
  assign w7151 = ( ~w3548 & w7148 ) | ( ~w3548 & w7150 ) | ( w7148 & w7150 ) ;
  assign w7152 = \pi14 ^ w7151 ;
  assign w7153 = ( ~w6962 & w7144 ) | ( ~w6962 & w7152 ) | ( w7144 & w7152 ) ;
  assign w7154 = ~w6749 & w6750 ;
  assign w7155 = w4049 | w6748 ;
  assign w7156 = ~w4142 & w6949 ;
  assign w7157 = ( ~w4049 & w7155 ) | ( ~w4049 & w7156 ) | ( w7155 & w7156 ) ;
  assign w7158 = w3962 | w7154 ;
  assign w7159 = w4152 & ~w7157 ;
  assign w7160 = ( w6751 & w7157 ) | ( w6751 & ~w7159 ) | ( w7157 & ~w7159 ) ;
  assign w7161 = ( ~w3962 & w7158 ) | ( ~w3962 & w7160 ) | ( w7158 & w7160 ) ;
  assign w7162 = \pi11 ^ w7161 ;
  assign w7163 = ( w6960 & w7153 ) | ( w6960 & w7162 ) | ( w7153 & w7162 ) ;
  assign w7164 = ~w4142 & w6748 ;
  assign w7165 = ( ~w4600 & w7154 ) | ( ~w4600 & w7164 ) | ( w7154 & w7164 ) ;
  assign w7166 = w6949 | w7165 ;
  assign w7167 = ( ~w3962 & w7165 ) | ( ~w3962 & w7166 ) | ( w7165 & w7166 ) ;
  assign w7168 = w7164 | w7167 ;
  assign w7169 = w6775 ^ w6946 ;
  assign w7170 = w6767 ^ w7169 ;
  assign w7171 = w4722 & ~w7168 ;
  assign w7172 = ( w6751 & w7168 ) | ( w6751 & ~w7171 ) | ( w7168 & ~w7171 ) ;
  assign w7173 = \pi11 ^ w7172 ;
  assign w7174 = ( w7163 & w7170 ) | ( w7163 & w7173 ) | ( w7170 & w7173 ) ;
  assign w7175 = \pi11 ^ w6947 ;
  assign w7176 = w6954 ^ w7175 ;
  assign w7177 = w6956 ^ w7176 ;
  assign w7178 = w4722 & w6751 ;
  assign w7179 = ( w6751 & w7168 ) | ( w6751 & ~w7178 ) | ( w7168 & ~w7178 ) ;
  assign w7180 = w7163 ^ w7179 ;
  assign w7181 = \pi11 ^ w7170 ;
  assign w7182 = w7180 ^ w7181 ;
  assign w7183 = w6962 ^ w7152 ;
  assign w7184 = w7144 ^ w7183 ;
  assign w7185 = w6970 ^ w7143 ;
  assign w7186 = w6972 ^ w7185 ;
  assign w7187 = w3647 & ~w6549 ;
  assign w7188 = ~w3094 & w6048 ;
  assign w7189 = ( w3647 & ~w7187 ) | ( w3647 & w7188 ) | ( ~w7187 & w7188 ) ;
  assign w7190 = w3715 & ~w6637 ;
  assign w7191 = w4164 & ~w7189 ;
  assign w7192 = ( w6045 & w7189 ) | ( w6045 & ~w7191 ) | ( w7189 & ~w7191 ) ;
  assign w7193 = ( w3715 & ~w7190 ) | ( w3715 & w7192 ) | ( ~w7190 & w7192 ) ;
  assign w7194 = \pi14 ^ w7193 ;
  assign w7195 = w6974 ^ w7142 ;
  assign w7196 = w7134 ^ w7195 ;
  assign w7197 = w6976 ^ w7133 ;
  assign w7198 = w7125 ^ w7197 ;
  assign w7199 = w1711 & ~w4651 ;
  assign w7200 = ~w1834 & w4606 ;
  assign w7201 = ( w1711 & ~w7199 ) | ( w1711 & w7200 ) | ( ~w7199 & w7200 ) ;
  assign w7202 = w1614 & ~w4706 ;
  assign w7203 = w5433 & ~w7201 ;
  assign w7204 = ( w4609 & w7201 ) | ( w4609 & ~w7203 ) | ( w7201 & ~w7203 ) ;
  assign w7205 = ( w1614 & ~w7202 ) | ( w1614 & w7204 ) | ( ~w7202 & w7204 ) ;
  assign w7206 = \pi23 ^ w7205 ;
  assign w7207 = w6978 ^ w7113 ;
  assign w7208 = w6986 ^ w7207 ;
  assign w7209 = w1939 | w4606 ;
  assign w7210 = ~w1834 & w4651 ;
  assign w7211 = ( ~w1939 & w7209 ) | ( ~w1939 & w7210 ) | ( w7209 & w7210 ) ;
  assign w7212 = w1711 & ~w4706 ;
  assign w7213 = w5296 | w7211 ;
  assign w7214 = ( w4609 & w7211 ) | ( w4609 & w7213 ) | ( w7211 & w7213 ) ;
  assign w7215 = ( w1711 & ~w7212 ) | ( w1711 & w7214 ) | ( ~w7212 & w7214 ) ;
  assign w7216 = \pi23 ^ w7215 ;
  assign w7217 = w6988 ^ w7112 ;
  assign w7218 = w6996 ^ w7217 ;
  assign w7219 = w1939 | w4651 ;
  assign w7220 = w1976 & w4606 ;
  assign w7221 = ( ~w1939 & w7219 ) | ( ~w1939 & w7220 ) | ( w7219 & w7220 ) ;
  assign w7222 = w1834 | w4706 ;
  assign w7223 = w5659 & ~w7221 ;
  assign w7224 = ( w4609 & w7221 ) | ( w4609 & ~w7223 ) | ( w7221 & ~w7223 ) ;
  assign w7225 = ( ~w1834 & w7222 ) | ( ~w1834 & w7224 ) | ( w7222 & w7224 ) ;
  assign w7226 = \pi23 ^ w7225 ;
  assign w7227 = w6998 ^ w7111 ;
  assign w7228 = w7006 ^ w7227 ;
  assign w7229 = w2059 | w4606 ;
  assign w7230 = w1976 & w4651 ;
  assign w7231 = ( ~w2059 & w7229 ) | ( ~w2059 & w7230 ) | ( w7229 & w7230 ) ;
  assign w7232 = w1939 | w4706 ;
  assign w7233 = w5748 | w7231 ;
  assign w7234 = ( w4609 & w7231 ) | ( w4609 & w7233 ) | ( w7231 & w7233 ) ;
  assign w7235 = ( ~w1939 & w7232 ) | ( ~w1939 & w7234 ) | ( w7232 & w7234 ) ;
  assign w7236 = \pi23 ^ w7235 ;
  assign w7237 = w7008 ^ w7110 ;
  assign w7238 = w7016 ^ w7237 ;
  assign w7239 = w2059 | w4651 ;
  assign w7240 = ~w2130 & w4606 ;
  assign w7241 = ( ~w2059 & w7239 ) | ( ~w2059 & w7240 ) | ( w7239 & w7240 ) ;
  assign w7242 = w1976 & ~w4706 ;
  assign w7243 = w5646 | w7241 ;
  assign w7244 = ( w4609 & w7241 ) | ( w4609 & w7243 ) | ( w7241 & w7243 ) ;
  assign w7245 = ( w1976 & ~w7242 ) | ( w1976 & w7244 ) | ( ~w7242 & w7244 ) ;
  assign w7246 = \pi23 ^ w7245 ;
  assign w7247 = w7018 ^ w7109 ;
  assign w7248 = w7026 ^ w7247 ;
  assign w7249 = w2130 | w4651 ;
  assign w7250 = ~w2235 & w4606 ;
  assign w7251 = ( ~w2130 & w7249 ) | ( ~w2130 & w7250 ) | ( w7249 & w7250 ) ;
  assign w7252 = w2059 | w4706 ;
  assign w7253 = w5896 & ~w7251 ;
  assign w7254 = ( w4609 & w7251 ) | ( w4609 & ~w7253 ) | ( w7251 & ~w7253 ) ;
  assign w7255 = ( ~w2059 & w7252 ) | ( ~w2059 & w7254 ) | ( w7252 & w7254 ) ;
  assign w7256 = \pi23 ^ w7255 ;
  assign w7257 = w7028 ^ w7108 ;
  assign w7258 = w7036 ^ w7257 ;
  assign w7259 = w2273 & ~w4606 ;
  assign w7260 = ~w2235 & w4651 ;
  assign w7261 = ( w2273 & ~w7259 ) | ( w2273 & w7260 ) | ( ~w7259 & w7260 ) ;
  assign w7262 = w2130 | w4706 ;
  assign w7263 = w6094 | w7261 ;
  assign w7264 = ( w4609 & w7261 ) | ( w4609 & w7263 ) | ( w7261 & w7263 ) ;
  assign w7265 = ( ~w2130 & w7262 ) | ( ~w2130 & w7264 ) | ( w7262 & w7264 ) ;
  assign w7266 = \pi23 ^ w7265 ;
  assign w7267 = w7038 ^ w7107 ;
  assign w7268 = w7046 ^ w7267 ;
  assign w7269 = w7054 ^ w7106 ;
  assign w7270 = w7056 ^ w7269 ;
  assign w7271 = w2273 & ~w4651 ;
  assign w7272 = w2391 & w4606 ;
  assign w7273 = ( w2273 & ~w7271 ) | ( w2273 & w7272 ) | ( ~w7271 & w7272 ) ;
  assign w7274 = w2235 | w4706 ;
  assign w7275 = w6106 & ~w7273 ;
  assign w7276 = ( w4609 & w7273 ) | ( w4609 & ~w7275 ) | ( w7273 & ~w7275 ) ;
  assign w7277 = ( ~w2235 & w7274 ) | ( ~w2235 & w7276 ) | ( w7274 & w7276 ) ;
  assign w7278 = \pi23 ^ w7277 ;
  assign w7279 = w7064 ^ w7105 ;
  assign w7280 = w7065 ^ w7279 ;
  assign w7281 = w2391 & ~w4651 ;
  assign w7282 = w2500 & w4606 ;
  assign w7283 = ( w2391 & ~w7281 ) | ( w2391 & w7282 ) | ( ~w7281 & w7282 ) ;
  assign w7284 = w2273 & ~w4706 ;
  assign w7285 = w5880 | w7283 ;
  assign w7286 = ( w4609 & w7283 ) | ( w4609 & w7285 ) | ( w7283 & w7285 ) ;
  assign w7287 = ( w2273 & ~w7284 ) | ( w2273 & w7286 ) | ( ~w7284 & w7286 ) ;
  assign w7288 = \pi23 ^ w7287 ;
  assign w7289 = w2578 | w4606 ;
  assign w7290 = w2500 & w4651 ;
  assign w7291 = ( ~w2578 & w7289 ) | ( ~w2578 & w7290 ) | ( w7289 & w7290 ) ;
  assign w7292 = w2391 & ~w4706 ;
  assign w7293 = w6164 & ~w7291 ;
  assign w7294 = ( w4609 & w7291 ) | ( w4609 & ~w7293 ) | ( w7291 & ~w7293 ) ;
  assign w7295 = ( w2391 & ~w7292 ) | ( w2391 & w7294 ) | ( ~w7292 & w7294 ) ;
  assign w7296 = \pi23 ^ w7295 ;
  assign w7297 = w7078 ^ w7104 ;
  assign w7298 = w7070 ^ w7297 ;
  assign w7299 = w7094 ^ w7102 ;
  assign w7300 = w7103 ^ w7299 ;
  assign w7301 = w2578 | w4651 ;
  assign w7302 = ~w2653 & w4606 ;
  assign w7303 = ( ~w2578 & w7301 ) | ( ~w2578 & w7302 ) | ( w7301 & w7302 ) ;
  assign w7304 = w2500 & ~w4706 ;
  assign w7305 = w6219 | w7303 ;
  assign w7306 = ( w4609 & w7303 ) | ( w4609 & w7305 ) | ( w7303 & w7305 ) ;
  assign w7307 = ( w2500 & ~w7304 ) | ( w2500 & w7306 ) | ( ~w7304 & w7306 ) ;
  assign w7308 = \pi23 ^ w7307 ;
  assign w7309 = w2694 | w4606 ;
  assign w7310 = ~w2653 & w4651 ;
  assign w7311 = ( ~w2694 & w7309 ) | ( ~w2694 & w7310 ) | ( w7309 & w7310 ) ;
  assign w7312 = w2578 | w4706 ;
  assign w7313 = w6282 & ~w7311 ;
  assign w7314 = ( w4609 & w7311 ) | ( w4609 & ~w7313 ) | ( w7311 & ~w7313 ) ;
  assign w7315 = ( ~w2578 & w7312 ) | ( ~w2578 & w7314 ) | ( w7312 & w7314 ) ;
  assign w7316 = \pi23 ^ w7315 ;
  assign w7317 = w7085 ^ w7093 ;
  assign w7318 = ( \pi23 & \pi24 ) | ( \pi23 & ~w2871 ) | ( \pi24 & ~w2871 ) ;
  assign w7319 = \pi23 & \pi24 ;
  assign w7320 = w2973 ^ w7319 ;
  assign w7321 = ( \pi25 & w7319 ) | ( \pi25 & ~w7320 ) | ( w7319 & ~w7320 ) ;
  assign w7322 = w7318 ^ w7321 ;
  assign w7323 = w2805 & ~w4606 ;
  assign w7324 = ~w2694 & w4651 ;
  assign w7325 = ( w2805 & ~w7323 ) | ( w2805 & w7324 ) | ( ~w7323 & w7324 ) ;
  assign w7326 = w2653 | w4706 ;
  assign w7327 = w6338 & ~w7325 ;
  assign w7328 = ( w4609 & w7325 ) | ( w4609 & ~w7327 ) | ( w7325 & ~w7327 ) ;
  assign w7329 = ( ~w2653 & w7326 ) | ( ~w2653 & w7328 ) | ( w7326 & w7328 ) ;
  assign w7330 = \pi23 ^ w7329 ;
  assign w7331 = ( \pi20 & \pi21 ) | ( \pi20 & ~\pi23 ) | ( \pi21 & ~\pi23 ) ;
  assign w7332 = \pi23 & w2973 ;
  assign w7333 = w2871 & w7332 ;
  assign w7334 = ( \pi20 & \pi21 ) | ( \pi20 & ~w7333 ) | ( \pi21 & ~w7333 ) ;
  assign w7335 = ( \pi22 & \pi23 ) | ( \pi22 & ~w7334 ) | ( \pi23 & ~w7334 ) ;
  assign w7336 = ( \pi22 & ~w7332 ) | ( \pi22 & w7334 ) | ( ~w7332 & w7334 ) ;
  assign w7337 = ( w7331 & w7335 ) | ( w7331 & ~w7336 ) | ( w7335 & ~w7336 ) ;
  assign w7338 = w2973 | w4606 ;
  assign w7339 = ~w2871 & w4651 ;
  assign w7340 = ( ~w2973 & w7338 ) | ( ~w2973 & w7339 ) | ( w7338 & w7339 ) ;
  assign w7341 = w2805 & ~w4706 ;
  assign w7342 = w6457 | w7340 ;
  assign w7343 = ( w4609 & w7340 ) | ( w4609 & w7342 ) | ( w7340 & w7342 ) ;
  assign w7344 = ( w2805 & ~w7341 ) | ( w2805 & w7343 ) | ( ~w7341 & w7343 ) ;
  assign w7345 = \pi23 ^ w7344 ;
  assign w7346 = w7337 & w7345 ;
  assign w7347 = w2805 & ~w4651 ;
  assign w7348 = ~w2871 & w4606 ;
  assign w7349 = ( w2805 & ~w7347 ) | ( w2805 & w7348 ) | ( ~w7347 & w7348 ) ;
  assign w7350 = w2694 | w4706 ;
  assign w7351 = w6473 | w7349 ;
  assign w7352 = ( w4609 & w7349 ) | ( w4609 & w7351 ) | ( w7349 & w7351 ) ;
  assign w7353 = ( ~w2694 & w7350 ) | ( ~w2694 & w7352 ) | ( w7350 & w7352 ) ;
  assign w7354 = \pi23 ^ w7353 ;
  assign w7355 = w2832 & ~w2973 ;
  assign w7356 = ( w7346 & w7354 ) | ( w7346 & w7355 ) | ( w7354 & w7355 ) ;
  assign w7357 = ( w7322 & w7330 ) | ( w7322 & w7356 ) | ( w7330 & w7356 ) ;
  assign w7358 = ( w7316 & w7317 ) | ( w7316 & w7357 ) | ( w7317 & w7357 ) ;
  assign w7359 = ( w7300 & w7308 ) | ( w7300 & w7358 ) | ( w7308 & w7358 ) ;
  assign w7360 = ( w7296 & w7298 ) | ( w7296 & w7359 ) | ( w7298 & w7359 ) ;
  assign w7361 = ( w7280 & w7288 ) | ( w7280 & w7360 ) | ( w7288 & w7360 ) ;
  assign w7362 = ( w7270 & w7278 ) | ( w7270 & w7361 ) | ( w7278 & w7361 ) ;
  assign w7363 = ( w7266 & w7268 ) | ( w7266 & w7362 ) | ( w7268 & w7362 ) ;
  assign w7364 = ( w7256 & ~w7258 ) | ( w7256 & w7363 ) | ( ~w7258 & w7363 ) ;
  assign w7365 = ( w7246 & ~w7248 ) | ( w7246 & w7364 ) | ( ~w7248 & w7364 ) ;
  assign w7366 = ( w7236 & w7238 ) | ( w7236 & w7365 ) | ( w7238 & w7365 ) ;
  assign w7367 = ( w7226 & ~w7228 ) | ( w7226 & w7366 ) | ( ~w7228 & w7366 ) ;
  assign w7368 = ( w7216 & w7218 ) | ( w7216 & w7367 ) | ( w7218 & w7367 ) ;
  assign w7369 = ( w7206 & w7208 ) | ( w7206 & w7368 ) | ( w7208 & w7368 ) ;
  assign w7370 = w7114 ^ w7124 ;
  assign w7371 = w7116 ^ w7370 ;
  assign w7372 = w1264 | w5343 ;
  assign w7373 = w1399 & w4905 ;
  assign w7374 = ( ~w1264 & w7372 ) | ( ~w1264 & w7373 ) | ( w7372 & w7373 ) ;
  assign w7375 = w1205 & ~w5395 ;
  assign w7376 = w4864 & ~w7374 ;
  assign w7377 = ( w4908 & w7374 ) | ( w4908 & ~w7376 ) | ( w7374 & ~w7376 ) ;
  assign w7378 = ( w1205 & ~w7375 ) | ( w1205 & w7377 ) | ( ~w7375 & w7377 ) ;
  assign w7379 = \pi20 ^ w7378 ;
  assign w7380 = ( w7369 & w7371 ) | ( w7369 & w7379 ) | ( w7371 & w7379 ) ;
  assign w7381 = w883 | w5710 ;
  assign w7382 = w979 & w5494 ;
  assign w7383 = ( ~w883 & w7381 ) | ( ~w883 & w7382 ) | ( w7381 & w7382 ) ;
  assign w7384 = w721 & ~w5948 ;
  assign w7385 = w4257 & ~w7383 ;
  assign w7386 = ( w5497 & w7383 ) | ( w5497 & ~w7385 ) | ( w7383 & ~w7385 ) ;
  assign w7387 = ( w721 & ~w7384 ) | ( w721 & w7386 ) | ( ~w7384 & w7386 ) ;
  assign w7388 = \pi17 ^ w7387 ;
  assign w7389 = ( w7198 & w7380 ) | ( w7198 & w7388 ) | ( w7380 & w7388 ) ;
  assign w7390 = w381 | w6048 ;
  assign w7391 = ~w3094 & w6549 ;
  assign w7392 = ( ~w381 & w7390 ) | ( ~w381 & w7391 ) | ( w7390 & w7391 ) ;
  assign w7393 = w3647 & ~w6637 ;
  assign w7394 = w3810 | w7392 ;
  assign w7395 = ( w6045 & w7392 ) | ( w6045 & w7394 ) | ( w7392 & w7394 ) ;
  assign w7396 = ( w3647 & ~w7393 ) | ( w3647 & w7395 ) | ( ~w7393 & w7395 ) ;
  assign w7397 = \pi14 ^ w7396 ;
  assign w7398 = ( ~w7196 & w7389 ) | ( ~w7196 & w7397 ) | ( w7389 & w7397 ) ;
  assign w7399 = ( w7186 & w7194 ) | ( w7186 & w7398 ) | ( w7194 & w7398 ) ;
  assign w7400 = w4049 | w6949 ;
  assign w7401 = w3907 & w6748 ;
  assign w7402 = ( ~w4049 & w7400 ) | ( ~w4049 & w7401 ) | ( w7400 & w7401 ) ;
  assign w7403 = w4142 | w7154 ;
  assign w7404 = w4563 | w7402 ;
  assign w7405 = ( w6751 & w7402 ) | ( w6751 & w7404 ) | ( w7402 & w7404 ) ;
  assign w7406 = ( ~w4142 & w7403 ) | ( ~w4142 & w7405 ) | ( w7403 & w7405 ) ;
  assign w7407 = \pi11 ^ w7406 ;
  assign w7408 = ( ~w7184 & w7399 ) | ( ~w7184 & w7407 ) | ( w7399 & w7407 ) ;
  assign w7409 = ( \pi06 & ~\pi07 ) | ( \pi06 & \pi08 ) | ( ~\pi07 & \pi08 ) ;
  assign w7410 = ( \pi05 & \pi06 ) | ( \pi05 & w7409 ) | ( \pi06 & w7409 ) ;
  assign w7411 = w7409 ^ w7410 ;
  assign w7412 = \pi07 ^ \pi08 ;
  assign w7413 = \pi05 ^ \pi06 ;
  assign w7414 = w7412 & w7413 ;
  assign w7415 = ~w4600 & w7411 ;
  assign w7416 = w7414 | w7415 ;
  assign w7417 = ( ~w4603 & w7415 ) | ( ~w4603 & w7416 ) | ( w7415 & w7416 ) ;
  assign w7418 = \pi08 ^ w7417 ;
  assign w7419 = w6960 ^ w7162 ;
  assign w7420 = w7153 ^ w7419 ;
  assign w7421 = ( w7408 & w7418 ) | ( w7408 & w7420 ) | ( w7418 & w7420 ) ;
  assign w7422 = w7418 ^ w7420 ;
  assign w7423 = w7408 ^ w7422 ;
  assign w7424 = w7196 ^ w7397 ;
  assign w7425 = w7389 ^ w7424 ;
  assign w7426 = w7198 ^ w7388 ;
  assign w7427 = w7380 ^ w7426 ;
  assign w7428 = w7206 ^ w7368 ;
  assign w7429 = w7208 ^ w7428 ;
  assign w7430 = w1399 & ~w5343 ;
  assign w7431 = ~w1510 & w4905 ;
  assign w7432 = ( w1399 & ~w7430 ) | ( w1399 & w7431 ) | ( ~w7430 & w7431 ) ;
  assign w7433 = w1264 | w5395 ;
  assign w7434 = w4852 & ~w7432 ;
  assign w7435 = ( w4908 & w7432 ) | ( w4908 & ~w7434 ) | ( w7432 & ~w7434 ) ;
  assign w7436 = ( ~w1264 & w7433 ) | ( ~w1264 & w7435 ) | ( w7433 & w7435 ) ;
  assign w7437 = \pi20 ^ w7436 ;
  assign w7438 = w7216 ^ w7367 ;
  assign w7439 = w7218 ^ w7438 ;
  assign w7440 = w1614 & ~w4905 ;
  assign w7441 = ~w1510 & w5343 ;
  assign w7442 = ( w1614 & ~w7440 ) | ( w1614 & w7441 ) | ( ~w7440 & w7441 ) ;
  assign w7443 = w1399 & ~w5395 ;
  assign w7444 = w5069 & ~w7442 ;
  assign w7445 = ( w4908 & w7442 ) | ( w4908 & ~w7444 ) | ( w7442 & ~w7444 ) ;
  assign w7446 = ( w1399 & ~w7443 ) | ( w1399 & w7445 ) | ( ~w7443 & w7445 ) ;
  assign w7447 = \pi20 ^ w7446 ;
  assign w7448 = w7226 ^ w7366 ;
  assign w7449 = w7228 ^ w7448 ;
  assign w7450 = w1614 & ~w5343 ;
  assign w7451 = w1711 & w4905 ;
  assign w7452 = ( w1614 & ~w7450 ) | ( w1614 & w7451 ) | ( ~w7450 & w7451 ) ;
  assign w7453 = w1510 | w5395 ;
  assign w7454 = w5085 & ~w7452 ;
  assign w7455 = ( w4908 & w7452 ) | ( w4908 & ~w7454 ) | ( w7452 & ~w7454 ) ;
  assign w7456 = ( ~w1510 & w7453 ) | ( ~w1510 & w7455 ) | ( w7453 & w7455 ) ;
  assign w7457 = \pi20 ^ w7456 ;
  assign w7458 = w7236 ^ w7365 ;
  assign w7459 = w7238 ^ w7458 ;
  assign w7460 = w1711 & ~w5343 ;
  assign w7461 = ~w1834 & w4905 ;
  assign w7462 = ( w1711 & ~w7460 ) | ( w1711 & w7461 ) | ( ~w7460 & w7461 ) ;
  assign w7463 = w1614 & ~w5395 ;
  assign w7464 = w5433 & ~w7462 ;
  assign w7465 = ( w4908 & w7462 ) | ( w4908 & ~w7464 ) | ( w7462 & ~w7464 ) ;
  assign w7466 = ( w1614 & ~w7463 ) | ( w1614 & w7465 ) | ( ~w7463 & w7465 ) ;
  assign w7467 = \pi20 ^ w7466 ;
  assign w7468 = w7246 ^ w7364 ;
  assign w7469 = w7248 ^ w7468 ;
  assign w7470 = w1939 | w4905 ;
  assign w7471 = ~w1834 & w5343 ;
  assign w7472 = ( ~w1939 & w7470 ) | ( ~w1939 & w7471 ) | ( w7470 & w7471 ) ;
  assign w7473 = w1711 & ~w5395 ;
  assign w7474 = w5296 | w7472 ;
  assign w7475 = ( w4908 & w7472 ) | ( w4908 & w7474 ) | ( w7472 & w7474 ) ;
  assign w7476 = ( w1711 & ~w7473 ) | ( w1711 & w7475 ) | ( ~w7473 & w7475 ) ;
  assign w7477 = \pi20 ^ w7476 ;
  assign w7478 = w7256 ^ w7363 ;
  assign w7479 = w7258 ^ w7478 ;
  assign w7480 = w1939 | w5343 ;
  assign w7481 = w1976 & w4905 ;
  assign w7482 = ( ~w1939 & w7480 ) | ( ~w1939 & w7481 ) | ( w7480 & w7481 ) ;
  assign w7483 = w1834 | w5395 ;
  assign w7484 = w5659 & ~w7482 ;
  assign w7485 = ( w4908 & w7482 ) | ( w4908 & ~w7484 ) | ( w7482 & ~w7484 ) ;
  assign w7486 = ( ~w1834 & w7483 ) | ( ~w1834 & w7485 ) | ( w7483 & w7485 ) ;
  assign w7487 = \pi20 ^ w7486 ;
  assign w7488 = w7266 ^ w7362 ;
  assign w7489 = w7268 ^ w7488 ;
  assign w7490 = w2059 | w4905 ;
  assign w7491 = w1976 & w5343 ;
  assign w7492 = ( ~w2059 & w7490 ) | ( ~w2059 & w7491 ) | ( w7490 & w7491 ) ;
  assign w7493 = w1939 | w5395 ;
  assign w7494 = w5748 | w7492 ;
  assign w7495 = ( w4908 & w7492 ) | ( w4908 & w7494 ) | ( w7492 & w7494 ) ;
  assign w7496 = ( ~w1939 & w7493 ) | ( ~w1939 & w7495 ) | ( w7493 & w7495 ) ;
  assign w7497 = \pi20 ^ w7496 ;
  assign w7498 = w2059 | w5343 ;
  assign w7499 = ~w2130 & w4905 ;
  assign w7500 = ( ~w2059 & w7498 ) | ( ~w2059 & w7499 ) | ( w7498 & w7499 ) ;
  assign w7501 = w1976 & ~w5395 ;
  assign w7502 = w5646 | w7500 ;
  assign w7503 = ( w4908 & w7500 ) | ( w4908 & w7502 ) | ( w7500 & w7502 ) ;
  assign w7504 = ( w1976 & ~w7501 ) | ( w1976 & w7503 ) | ( ~w7501 & w7503 ) ;
  assign w7505 = \pi20 ^ w7504 ;
  assign w7506 = w7270 ^ w7361 ;
  assign w7507 = w7278 ^ w7506 ;
  assign w7508 = w2130 | w5343 ;
  assign w7509 = ~w2235 & w4905 ;
  assign w7510 = ( ~w2130 & w7508 ) | ( ~w2130 & w7509 ) | ( w7508 & w7509 ) ;
  assign w7511 = w2059 | w5395 ;
  assign w7512 = w5896 & ~w7510 ;
  assign w7513 = ( w4908 & w7510 ) | ( w4908 & ~w7512 ) | ( w7510 & ~w7512 ) ;
  assign w7514 = ( ~w2059 & w7511 ) | ( ~w2059 & w7513 ) | ( w7511 & w7513 ) ;
  assign w7515 = \pi20 ^ w7514 ;
  assign w7516 = w7280 ^ w7360 ;
  assign w7517 = w7288 ^ w7516 ;
  assign w7518 = w7296 ^ w7359 ;
  assign w7519 = w7298 ^ w7518 ;
  assign w7520 = w2273 & ~w4905 ;
  assign w7521 = ~w2235 & w5343 ;
  assign w7522 = ( w2273 & ~w7520 ) | ( w2273 & w7521 ) | ( ~w7520 & w7521 ) ;
  assign w7523 = w2130 | w5395 ;
  assign w7524 = w6094 | w7522 ;
  assign w7525 = ( w4908 & w7522 ) | ( w4908 & w7524 ) | ( w7522 & w7524 ) ;
  assign w7526 = ( ~w2130 & w7523 ) | ( ~w2130 & w7525 ) | ( w7523 & w7525 ) ;
  assign w7527 = \pi20 ^ w7526 ;
  assign w7528 = w7300 ^ w7358 ;
  assign w7529 = w7308 ^ w7528 ;
  assign w7530 = w2273 & ~w5343 ;
  assign w7531 = w2391 & w4905 ;
  assign w7532 = ( w2273 & ~w7530 ) | ( w2273 & w7531 ) | ( ~w7530 & w7531 ) ;
  assign w7533 = w2235 | w5395 ;
  assign w7534 = w6106 & ~w7532 ;
  assign w7535 = ( w4908 & w7532 ) | ( w4908 & ~w7534 ) | ( w7532 & ~w7534 ) ;
  assign w7536 = ( ~w2235 & w7533 ) | ( ~w2235 & w7535 ) | ( w7533 & w7535 ) ;
  assign w7537 = \pi20 ^ w7536 ;
  assign w7538 = w7316 ^ w7357 ;
  assign w7539 = w7317 ^ w7538 ;
  assign w7540 = w2391 & ~w5343 ;
  assign w7541 = w2500 & w4905 ;
  assign w7542 = ( w2391 & ~w7540 ) | ( w2391 & w7541 ) | ( ~w7540 & w7541 ) ;
  assign w7543 = w2273 & ~w5395 ;
  assign w7544 = w5880 | w7542 ;
  assign w7545 = ( w4908 & w7542 ) | ( w4908 & w7544 ) | ( w7542 & w7544 ) ;
  assign w7546 = ( w2273 & ~w7543 ) | ( w2273 & w7545 ) | ( ~w7543 & w7545 ) ;
  assign w7547 = \pi20 ^ w7546 ;
  assign w7548 = w2578 | w4905 ;
  assign w7549 = w2500 & w5343 ;
  assign w7550 = ( ~w2578 & w7548 ) | ( ~w2578 & w7549 ) | ( w7548 & w7549 ) ;
  assign w7551 = w2391 & ~w5395 ;
  assign w7552 = w6164 & ~w7550 ;
  assign w7553 = ( w4908 & w7550 ) | ( w4908 & ~w7552 ) | ( w7550 & ~w7552 ) ;
  assign w7554 = ( w2391 & ~w7551 ) | ( w2391 & w7553 ) | ( ~w7551 & w7553 ) ;
  assign w7555 = \pi20 ^ w7554 ;
  assign w7556 = w7330 ^ w7356 ;
  assign w7557 = w7322 ^ w7556 ;
  assign w7558 = w7346 ^ w7354 ;
  assign w7559 = w7355 ^ w7558 ;
  assign w7560 = w2578 | w5343 ;
  assign w7561 = ~w2653 & w4905 ;
  assign w7562 = ( ~w2578 & w7560 ) | ( ~w2578 & w7561 ) | ( w7560 & w7561 ) ;
  assign w7563 = w2500 & ~w5395 ;
  assign w7564 = w6219 | w7562 ;
  assign w7565 = ( w4908 & w7562 ) | ( w4908 & w7564 ) | ( w7562 & w7564 ) ;
  assign w7566 = ( w2500 & ~w7563 ) | ( w2500 & w7565 ) | ( ~w7563 & w7565 ) ;
  assign w7567 = \pi20 ^ w7566 ;
  assign w7568 = w2694 | w4905 ;
  assign w7569 = ~w2653 & w5343 ;
  assign w7570 = ( ~w2694 & w7568 ) | ( ~w2694 & w7569 ) | ( w7568 & w7569 ) ;
  assign w7571 = w2578 | w5395 ;
  assign w7572 = w6282 & ~w7570 ;
  assign w7573 = ( w4908 & w7570 ) | ( w4908 & ~w7572 ) | ( w7570 & ~w7572 ) ;
  assign w7574 = ( ~w2578 & w7571 ) | ( ~w2578 & w7573 ) | ( w7571 & w7573 ) ;
  assign w7575 = \pi20 ^ w7574 ;
  assign w7576 = w7337 ^ w7345 ;
  assign w7577 = ( \pi20 & \pi21 ) | ( \pi20 & ~w2871 ) | ( \pi21 & ~w2871 ) ;
  assign w7578 = \pi20 & \pi21 ;
  assign w7579 = w2973 ^ w7578 ;
  assign w7580 = ( \pi22 & w7578 ) | ( \pi22 & ~w7579 ) | ( w7578 & ~w7579 ) ;
  assign w7581 = w7577 ^ w7580 ;
  assign w7582 = w2805 & ~w4905 ;
  assign w7583 = ~w2694 & w5343 ;
  assign w7584 = ( w2805 & ~w7582 ) | ( w2805 & w7583 ) | ( ~w7582 & w7583 ) ;
  assign w7585 = w2653 | w5395 ;
  assign w7586 = w6338 & ~w7584 ;
  assign w7587 = ( w4908 & w7584 ) | ( w4908 & ~w7586 ) | ( w7584 & ~w7586 ) ;
  assign w7588 = ( ~w2653 & w7585 ) | ( ~w2653 & w7587 ) | ( w7585 & w7587 ) ;
  assign w7589 = \pi20 ^ w7588 ;
  assign w7590 = ( \pi17 & \pi18 ) | ( \pi17 & ~\pi20 ) | ( \pi18 & ~\pi20 ) ;
  assign w7591 = \pi20 & w2973 ;
  assign w7592 = w2871 & w7591 ;
  assign w7593 = ( \pi17 & \pi18 ) | ( \pi17 & ~w7592 ) | ( \pi18 & ~w7592 ) ;
  assign w7594 = ( \pi19 & \pi20 ) | ( \pi19 & ~w7593 ) | ( \pi20 & ~w7593 ) ;
  assign w7595 = ( \pi19 & ~w7591 ) | ( \pi19 & w7593 ) | ( ~w7591 & w7593 ) ;
  assign w7596 = ( w7590 & w7594 ) | ( w7590 & ~w7595 ) | ( w7594 & ~w7595 ) ;
  assign w7597 = w2973 | w4905 ;
  assign w7598 = ~w2871 & w5343 ;
  assign w7599 = ( ~w2973 & w7597 ) | ( ~w2973 & w7598 ) | ( w7597 & w7598 ) ;
  assign w7600 = w2805 & ~w5395 ;
  assign w7601 = w6457 | w7599 ;
  assign w7602 = ( w4908 & w7599 ) | ( w4908 & w7601 ) | ( w7599 & w7601 ) ;
  assign w7603 = ( w2805 & ~w7600 ) | ( w2805 & w7602 ) | ( ~w7600 & w7602 ) ;
  assign w7604 = \pi20 ^ w7603 ;
  assign w7605 = w7596 & w7604 ;
  assign w7606 = w2805 & ~w5343 ;
  assign w7607 = ~w2871 & w4905 ;
  assign w7608 = ( w2805 & ~w7606 ) | ( w2805 & w7607 ) | ( ~w7606 & w7607 ) ;
  assign w7609 = w2694 | w5395 ;
  assign w7610 = w6473 | w7608 ;
  assign w7611 = ( w4908 & w7608 ) | ( w4908 & w7610 ) | ( w7608 & w7610 ) ;
  assign w7612 = ( ~w2694 & w7609 ) | ( ~w2694 & w7611 ) | ( w7609 & w7611 ) ;
  assign w7613 = \pi20 ^ w7612 ;
  assign w7614 = ~w2973 & w4608 ;
  assign w7615 = ( w7605 & w7613 ) | ( w7605 & w7614 ) | ( w7613 & w7614 ) ;
  assign w7616 = ( w7581 & w7589 ) | ( w7581 & w7615 ) | ( w7589 & w7615 ) ;
  assign w7617 = ( w7575 & w7576 ) | ( w7575 & w7616 ) | ( w7576 & w7616 ) ;
  assign w7618 = ( w7559 & w7567 ) | ( w7559 & w7617 ) | ( w7567 & w7617 ) ;
  assign w7619 = ( w7555 & w7557 ) | ( w7555 & w7618 ) | ( w7557 & w7618 ) ;
  assign w7620 = ( w7539 & w7547 ) | ( w7539 & w7619 ) | ( w7547 & w7619 ) ;
  assign w7621 = ( w7529 & w7537 ) | ( w7529 & w7620 ) | ( w7537 & w7620 ) ;
  assign w7622 = ( w7519 & w7527 ) | ( w7519 & w7621 ) | ( w7527 & w7621 ) ;
  assign w7623 = ( w7515 & w7517 ) | ( w7515 & w7622 ) | ( w7517 & w7622 ) ;
  assign w7624 = ( w7505 & w7507 ) | ( w7505 & w7623 ) | ( w7507 & w7623 ) ;
  assign w7625 = ( w7489 & w7497 ) | ( w7489 & w7624 ) | ( w7497 & w7624 ) ;
  assign w7626 = ( ~w7479 & w7487 ) | ( ~w7479 & w7625 ) | ( w7487 & w7625 ) ;
  assign w7627 = ( ~w7469 & w7477 ) | ( ~w7469 & w7626 ) | ( w7477 & w7626 ) ;
  assign w7628 = ( w7459 & w7467 ) | ( w7459 & w7627 ) | ( w7467 & w7627 ) ;
  assign w7629 = ( ~w7449 & w7457 ) | ( ~w7449 & w7628 ) | ( w7457 & w7628 ) ;
  assign w7630 = ( w7439 & w7447 ) | ( w7439 & w7629 ) | ( w7447 & w7629 ) ;
  assign w7631 = ( w7429 & w7437 ) | ( w7429 & w7630 ) | ( w7437 & w7630 ) ;
  assign w7632 = w7369 ^ w7379 ;
  assign w7633 = w7371 ^ w7632 ;
  assign w7634 = w979 & ~w5710 ;
  assign w7635 = w1085 & w5494 ;
  assign w7636 = ( w979 & ~w7634 ) | ( w979 & w7635 ) | ( ~w7634 & w7635 ) ;
  assign w7637 = w883 | w5948 ;
  assign w7638 = w4273 & ~w7636 ;
  assign w7639 = ( w5497 & w7636 ) | ( w5497 & ~w7638 ) | ( w7636 & ~w7638 ) ;
  assign w7640 = ( ~w883 & w7637 ) | ( ~w883 & w7639 ) | ( w7637 & w7639 ) ;
  assign w7641 = \pi17 ^ w7640 ;
  assign w7642 = ( w7631 & w7633 ) | ( w7631 & w7641 ) | ( w7633 & w7641 ) ;
  assign w7643 = w381 | w6549 ;
  assign w7644 = w592 & w6048 ;
  assign w7645 = ( ~w381 & w7643 ) | ( ~w381 & w7644 ) | ( w7643 & w7644 ) ;
  assign w7646 = w3094 | w6637 ;
  assign w7647 = w3096 | w7645 ;
  assign w7648 = ( w6045 & w7645 ) | ( w6045 & w7647 ) | ( w7645 & w7647 ) ;
  assign w7649 = ( ~w3094 & w7646 ) | ( ~w3094 & w7648 ) | ( w7646 & w7648 ) ;
  assign w7650 = \pi14 ^ w7649 ;
  assign w7651 = ( w7427 & w7642 ) | ( w7427 & w7650 ) | ( w7642 & w7650 ) ;
  assign w7652 = w3548 | w6949 ;
  assign w7653 = w3715 & w6748 ;
  assign w7654 = ( ~w3548 & w7652 ) | ( ~w3548 & w7653 ) | ( w7652 & w7653 ) ;
  assign w7655 = w3907 & ~w7154 ;
  assign w7656 = w3913 & ~w7654 ;
  assign w7657 = ( w6751 & w7654 ) | ( w6751 & ~w7656 ) | ( w7654 & ~w7656 ) ;
  assign w7658 = ( w3907 & ~w7655 ) | ( w3907 & w7657 ) | ( ~w7655 & w7657 ) ;
  assign w7659 = \pi11 ^ w7658 ;
  assign w7660 = ( ~w7425 & w7651 ) | ( ~w7425 & w7659 ) | ( w7651 & w7659 ) ;
  assign w7661 = w3548 | w6748 ;
  assign w7662 = w3907 & w6949 ;
  assign w7663 = ( ~w3548 & w7661 ) | ( ~w3548 & w7662 ) | ( w7661 & w7662 ) ;
  assign w7664 = w4049 | w7154 ;
  assign w7665 = w4622 & ~w7663 ;
  assign w7666 = ( w6751 & w7663 ) | ( w6751 & ~w7665 ) | ( w7663 & ~w7665 ) ;
  assign w7667 = ( ~w4049 & w7664 ) | ( ~w4049 & w7666 ) | ( w7664 & w7666 ) ;
  assign w7668 = \pi11 ^ w7667 ;
  assign w7669 = w7194 ^ w7398 ;
  assign w7670 = w7186 ^ w7669 ;
  assign w7671 = ( w7660 & w7668 ) | ( w7660 & w7670 ) | ( w7668 & w7670 ) ;
  assign w7672 = ( \pi05 & \pi06 ) | ( \pi05 & \pi07 ) | ( \pi06 & \pi07 ) ;
  assign w7673 = \pi07 ^ w7672 ;
  assign w7674 = ~w4600 & w7673 ;
  assign w7675 = ( w3962 & w6551 ) | ( w3962 & w7414 ) | ( w6551 & w7414 ) ;
  assign w7676 = w3962 | w7411 ;
  assign w7677 = ( ~w3962 & w7675 ) | ( ~w3962 & w7676 ) | ( w7675 & w7676 ) ;
  assign w7678 = ( ~w6555 & w7674 ) | ( ~w6555 & w7677 ) | ( w7674 & w7677 ) ;
  assign w7679 = w7184 ^ w7407 ;
  assign w7680 = w7399 ^ w7679 ;
  assign w7681 = \pi08 ^ w7678 ;
  assign w7682 = ( w7671 & ~w7680 ) | ( w7671 & w7681 ) | ( ~w7680 & w7681 ) ;
  assign w7683 = w7425 ^ w7659 ;
  assign w7684 = w7651 ^ w7683 ;
  assign w7685 = w7427 ^ w7650 ;
  assign w7686 = w7642 ^ w7685 ;
  assign w7687 = w1085 & ~w5710 ;
  assign w7688 = w1205 & w5494 ;
  assign w7689 = ( w1085 & ~w7687 ) | ( w1085 & w7688 ) | ( ~w7687 & w7688 ) ;
  assign w7690 = w979 & ~w5948 ;
  assign w7691 = w4666 | w7689 ;
  assign w7692 = ( w5497 & w7689 ) | ( w5497 & w7691 ) | ( w7689 & w7691 ) ;
  assign w7693 = ( w979 & ~w7690 ) | ( w979 & w7692 ) | ( ~w7690 & w7692 ) ;
  assign w7694 = \pi17 ^ w7693 ;
  assign w7695 = w7429 ^ w7630 ;
  assign w7696 = w7437 ^ w7695 ;
  assign w7697 = w1264 | w5494 ;
  assign w7698 = w1205 & w5710 ;
  assign w7699 = ( ~w1264 & w7697 ) | ( ~w1264 & w7698 ) | ( w7697 & w7698 ) ;
  assign w7700 = w1085 & ~w5948 ;
  assign w7701 = w4533 | w7699 ;
  assign w7702 = ( w5497 & w7699 ) | ( w5497 & w7701 ) | ( w7699 & w7701 ) ;
  assign w7703 = ( w1085 & ~w7700 ) | ( w1085 & w7702 ) | ( ~w7700 & w7702 ) ;
  assign w7704 = \pi17 ^ w7703 ;
  assign w7705 = w7439 ^ w7629 ;
  assign w7706 = w7447 ^ w7705 ;
  assign w7707 = w1264 | w5710 ;
  assign w7708 = w1399 & w5494 ;
  assign w7709 = ( ~w1264 & w7707 ) | ( ~w1264 & w7708 ) | ( w7707 & w7708 ) ;
  assign w7710 = w1205 & ~w5948 ;
  assign w7711 = w4864 & ~w7709 ;
  assign w7712 = ( w5497 & w7709 ) | ( w5497 & ~w7711 ) | ( w7709 & ~w7711 ) ;
  assign w7713 = ( w1205 & ~w7710 ) | ( w1205 & w7712 ) | ( ~w7710 & w7712 ) ;
  assign w7714 = \pi17 ^ w7713 ;
  assign w7715 = w7449 ^ w7628 ;
  assign w7716 = w7457 ^ w7715 ;
  assign w7717 = w1399 & ~w5710 ;
  assign w7718 = ~w1510 & w5494 ;
  assign w7719 = ( w1399 & ~w7717 ) | ( w1399 & w7718 ) | ( ~w7717 & w7718 ) ;
  assign w7720 = w1264 | w5948 ;
  assign w7721 = w4852 & ~w7719 ;
  assign w7722 = ( w5497 & w7719 ) | ( w5497 & ~w7721 ) | ( w7719 & ~w7721 ) ;
  assign w7723 = ( ~w1264 & w7720 ) | ( ~w1264 & w7722 ) | ( w7720 & w7722 ) ;
  assign w7724 = \pi17 ^ w7723 ;
  assign w7725 = w7459 ^ w7627 ;
  assign w7726 = w7467 ^ w7725 ;
  assign w7727 = w1614 & ~w5494 ;
  assign w7728 = ~w1510 & w5710 ;
  assign w7729 = ( w1614 & ~w7727 ) | ( w1614 & w7728 ) | ( ~w7727 & w7728 ) ;
  assign w7730 = w1399 & ~w5948 ;
  assign w7731 = w5069 & ~w7729 ;
  assign w7732 = ( w5497 & w7729 ) | ( w5497 & ~w7731 ) | ( w7729 & ~w7731 ) ;
  assign w7733 = ( w1399 & ~w7730 ) | ( w1399 & w7732 ) | ( ~w7730 & w7732 ) ;
  assign w7734 = \pi17 ^ w7733 ;
  assign w7735 = w7469 ^ w7626 ;
  assign w7736 = w7477 ^ w7735 ;
  assign w7737 = w1614 & ~w5710 ;
  assign w7738 = w1711 & w5494 ;
  assign w7739 = ( w1614 & ~w7737 ) | ( w1614 & w7738 ) | ( ~w7737 & w7738 ) ;
  assign w7740 = w1510 | w5948 ;
  assign w7741 = w5085 & ~w7739 ;
  assign w7742 = ( w5497 & w7739 ) | ( w5497 & ~w7741 ) | ( w7739 & ~w7741 ) ;
  assign w7743 = ( ~w1510 & w7740 ) | ( ~w1510 & w7742 ) | ( w7740 & w7742 ) ;
  assign w7744 = \pi17 ^ w7743 ;
  assign w7745 = w7479 ^ w7625 ;
  assign w7746 = w7487 ^ w7745 ;
  assign w7747 = w1711 & ~w5710 ;
  assign w7748 = ~w1834 & w5494 ;
  assign w7749 = ( w1711 & ~w7747 ) | ( w1711 & w7748 ) | ( ~w7747 & w7748 ) ;
  assign w7750 = w1614 & ~w5948 ;
  assign w7751 = w5433 & ~w7749 ;
  assign w7752 = ( w5497 & w7749 ) | ( w5497 & ~w7751 ) | ( w7749 & ~w7751 ) ;
  assign w7753 = ( w1614 & ~w7750 ) | ( w1614 & w7752 ) | ( ~w7750 & w7752 ) ;
  assign w7754 = \pi17 ^ w7753 ;
  assign w7755 = w7489 ^ w7624 ;
  assign w7756 = w7497 ^ w7755 ;
  assign w7757 = w7505 ^ w7623 ;
  assign w7758 = w7507 ^ w7757 ;
  assign w7759 = w1939 | w5494 ;
  assign w7760 = ~w1834 & w5710 ;
  assign w7761 = ( ~w1939 & w7759 ) | ( ~w1939 & w7760 ) | ( w7759 & w7760 ) ;
  assign w7762 = w1711 & ~w5948 ;
  assign w7763 = w5296 | w7761 ;
  assign w7764 = ( w5497 & w7761 ) | ( w5497 & w7763 ) | ( w7761 & w7763 ) ;
  assign w7765 = ( w1711 & ~w7762 ) | ( w1711 & w7764 ) | ( ~w7762 & w7764 ) ;
  assign w7766 = \pi17 ^ w7765 ;
  assign w7767 = w7515 ^ w7622 ;
  assign w7768 = w7517 ^ w7767 ;
  assign w7769 = w1939 | w5710 ;
  assign w7770 = w1976 & w5494 ;
  assign w7771 = ( ~w1939 & w7769 ) | ( ~w1939 & w7770 ) | ( w7769 & w7770 ) ;
  assign w7772 = w1834 | w5948 ;
  assign w7773 = w5659 & ~w7771 ;
  assign w7774 = ( w5497 & w7771 ) | ( w5497 & ~w7773 ) | ( w7771 & ~w7773 ) ;
  assign w7775 = ( ~w1834 & w7772 ) | ( ~w1834 & w7774 ) | ( w7772 & w7774 ) ;
  assign w7776 = \pi17 ^ w7775 ;
  assign w7777 = w2059 | w5494 ;
  assign w7778 = w1976 & w5710 ;
  assign w7779 = ( ~w2059 & w7777 ) | ( ~w2059 & w7778 ) | ( w7777 & w7778 ) ;
  assign w7780 = w1939 | w5948 ;
  assign w7781 = w5748 | w7779 ;
  assign w7782 = ( w5497 & w7779 ) | ( w5497 & w7781 ) | ( w7779 & w7781 ) ;
  assign w7783 = ( ~w1939 & w7780 ) | ( ~w1939 & w7782 ) | ( w7780 & w7782 ) ;
  assign w7784 = \pi17 ^ w7783 ;
  assign w7785 = w7519 ^ w7621 ;
  assign w7786 = w7527 ^ w7785 ;
  assign w7787 = w2059 | w5710 ;
  assign w7788 = ~w2130 & w5494 ;
  assign w7789 = ( ~w2059 & w7787 ) | ( ~w2059 & w7788 ) | ( w7787 & w7788 ) ;
  assign w7790 = w1976 & ~w5948 ;
  assign w7791 = w5646 | w7789 ;
  assign w7792 = ( w5497 & w7789 ) | ( w5497 & w7791 ) | ( w7789 & w7791 ) ;
  assign w7793 = ( w1976 & ~w7790 ) | ( w1976 & w7792 ) | ( ~w7790 & w7792 ) ;
  assign w7794 = \pi17 ^ w7793 ;
  assign w7795 = w7529 ^ w7620 ;
  assign w7796 = w7537 ^ w7795 ;
  assign w7797 = w2130 | w5710 ;
  assign w7798 = ~w2235 & w5494 ;
  assign w7799 = ( ~w2130 & w7797 ) | ( ~w2130 & w7798 ) | ( w7797 & w7798 ) ;
  assign w7800 = w2059 | w5948 ;
  assign w7801 = w5896 & ~w7799 ;
  assign w7802 = ( w5497 & w7799 ) | ( w5497 & ~w7801 ) | ( w7799 & ~w7801 ) ;
  assign w7803 = ( ~w2059 & w7800 ) | ( ~w2059 & w7802 ) | ( w7800 & w7802 ) ;
  assign w7804 = \pi17 ^ w7803 ;
  assign w7805 = w7539 ^ w7619 ;
  assign w7806 = w7547 ^ w7805 ;
  assign w7807 = w7555 ^ w7618 ;
  assign w7808 = w7557 ^ w7807 ;
  assign w7809 = w2273 & ~w5494 ;
  assign w7810 = ~w2235 & w5710 ;
  assign w7811 = ( w2273 & ~w7809 ) | ( w2273 & w7810 ) | ( ~w7809 & w7810 ) ;
  assign w7812 = w2130 | w5948 ;
  assign w7813 = w6094 | w7811 ;
  assign w7814 = ( w5497 & w7811 ) | ( w5497 & w7813 ) | ( w7811 & w7813 ) ;
  assign w7815 = ( ~w2130 & w7812 ) | ( ~w2130 & w7814 ) | ( w7812 & w7814 ) ;
  assign w7816 = \pi17 ^ w7815 ;
  assign w7817 = w7559 ^ w7617 ;
  assign w7818 = w7567 ^ w7817 ;
  assign w7819 = w2273 & ~w5710 ;
  assign w7820 = w2391 & w5494 ;
  assign w7821 = ( w2273 & ~w7819 ) | ( w2273 & w7820 ) | ( ~w7819 & w7820 ) ;
  assign w7822 = w2235 | w5948 ;
  assign w7823 = w6106 & ~w7821 ;
  assign w7824 = ( w5497 & w7821 ) | ( w5497 & ~w7823 ) | ( w7821 & ~w7823 ) ;
  assign w7825 = ( ~w2235 & w7822 ) | ( ~w2235 & w7824 ) | ( w7822 & w7824 ) ;
  assign w7826 = \pi17 ^ w7825 ;
  assign w7827 = w7575 ^ w7616 ;
  assign w7828 = w7576 ^ w7827 ;
  assign w7829 = w2391 & ~w5710 ;
  assign w7830 = w2500 & w5494 ;
  assign w7831 = ( w2391 & ~w7829 ) | ( w2391 & w7830 ) | ( ~w7829 & w7830 ) ;
  assign w7832 = w2273 & ~w5948 ;
  assign w7833 = w5880 | w7831 ;
  assign w7834 = ( w5497 & w7831 ) | ( w5497 & w7833 ) | ( w7831 & w7833 ) ;
  assign w7835 = ( w2273 & ~w7832 ) | ( w2273 & w7834 ) | ( ~w7832 & w7834 ) ;
  assign w7836 = \pi17 ^ w7835 ;
  assign w7837 = w2578 | w5494 ;
  assign w7838 = w2500 & w5710 ;
  assign w7839 = ( ~w2578 & w7837 ) | ( ~w2578 & w7838 ) | ( w7837 & w7838 ) ;
  assign w7840 = w2391 & ~w5948 ;
  assign w7841 = w6164 & ~w7839 ;
  assign w7842 = ( w5497 & w7839 ) | ( w5497 & ~w7841 ) | ( w7839 & ~w7841 ) ;
  assign w7843 = ( w2391 & ~w7840 ) | ( w2391 & w7842 ) | ( ~w7840 & w7842 ) ;
  assign w7844 = \pi17 ^ w7843 ;
  assign w7845 = w7589 ^ w7615 ;
  assign w7846 = w7581 ^ w7845 ;
  assign w7847 = w7605 ^ w7613 ;
  assign w7848 = w7614 ^ w7847 ;
  assign w7849 = w2578 | w5710 ;
  assign w7850 = ~w2653 & w5494 ;
  assign w7851 = ( ~w2578 & w7849 ) | ( ~w2578 & w7850 ) | ( w7849 & w7850 ) ;
  assign w7852 = w2500 & ~w5948 ;
  assign w7853 = w6219 | w7851 ;
  assign w7854 = ( w5497 & w7851 ) | ( w5497 & w7853 ) | ( w7851 & w7853 ) ;
  assign w7855 = ( w2500 & ~w7852 ) | ( w2500 & w7854 ) | ( ~w7852 & w7854 ) ;
  assign w7856 = \pi17 ^ w7855 ;
  assign w7857 = w2694 | w5494 ;
  assign w7858 = ~w2653 & w5710 ;
  assign w7859 = ( ~w2694 & w7857 ) | ( ~w2694 & w7858 ) | ( w7857 & w7858 ) ;
  assign w7860 = w2578 | w5948 ;
  assign w7861 = w6282 & ~w7859 ;
  assign w7862 = ( w5497 & w7859 ) | ( w5497 & ~w7861 ) | ( w7859 & ~w7861 ) ;
  assign w7863 = ( ~w2578 & w7860 ) | ( ~w2578 & w7862 ) | ( w7860 & w7862 ) ;
  assign w7864 = \pi17 ^ w7863 ;
  assign w7865 = w7596 ^ w7604 ;
  assign w7866 = ( \pi17 & \pi18 ) | ( \pi17 & ~w2871 ) | ( \pi18 & ~w2871 ) ;
  assign w7867 = \pi17 & \pi18 ;
  assign w7868 = w2973 ^ w7867 ;
  assign w7869 = ( \pi19 & w7867 ) | ( \pi19 & ~w7868 ) | ( w7867 & ~w7868 ) ;
  assign w7870 = w7866 ^ w7869 ;
  assign w7871 = w2805 & ~w5494 ;
  assign w7872 = ~w2694 & w5710 ;
  assign w7873 = ( w2805 & ~w7871 ) | ( w2805 & w7872 ) | ( ~w7871 & w7872 ) ;
  assign w7874 = w2653 | w5948 ;
  assign w7875 = w6338 & ~w7873 ;
  assign w7876 = ( w5497 & w7873 ) | ( w5497 & ~w7875 ) | ( w7873 & ~w7875 ) ;
  assign w7877 = ( ~w2653 & w7874 ) | ( ~w2653 & w7876 ) | ( w7874 & w7876 ) ;
  assign w7878 = \pi17 ^ w7877 ;
  assign w7879 = ( \pi14 & \pi15 ) | ( \pi14 & ~\pi17 ) | ( \pi15 & ~\pi17 ) ;
  assign w7880 = \pi17 & w2973 ;
  assign w7881 = w2871 & w7880 ;
  assign w7882 = ( \pi14 & \pi15 ) | ( \pi14 & ~w7881 ) | ( \pi15 & ~w7881 ) ;
  assign w7883 = ( \pi16 & \pi17 ) | ( \pi16 & ~w7882 ) | ( \pi17 & ~w7882 ) ;
  assign w7884 = ( \pi16 & ~w7880 ) | ( \pi16 & w7882 ) | ( ~w7880 & w7882 ) ;
  assign w7885 = ( w7879 & w7883 ) | ( w7879 & ~w7884 ) | ( w7883 & ~w7884 ) ;
  assign w7886 = w2973 | w5494 ;
  assign w7887 = ~w2871 & w5710 ;
  assign w7888 = ( ~w2973 & w7886 ) | ( ~w2973 & w7887 ) | ( w7886 & w7887 ) ;
  assign w7889 = w2805 & ~w5948 ;
  assign w7890 = w6457 | w7888 ;
  assign w7891 = ( w5497 & w7888 ) | ( w5497 & w7890 ) | ( w7888 & w7890 ) ;
  assign w7892 = ( w2805 & ~w7889 ) | ( w2805 & w7891 ) | ( ~w7889 & w7891 ) ;
  assign w7893 = \pi17 ^ w7892 ;
  assign w7894 = w7885 & w7893 ;
  assign w7895 = w2805 & ~w5710 ;
  assign w7896 = ~w2871 & w5494 ;
  assign w7897 = ( w2805 & ~w7895 ) | ( w2805 & w7896 ) | ( ~w7895 & w7896 ) ;
  assign w7898 = w2694 | w5948 ;
  assign w7899 = w6473 | w7897 ;
  assign w7900 = ( w5497 & w7897 ) | ( w5497 & w7899 ) | ( w7897 & w7899 ) ;
  assign w7901 = ( ~w2694 & w7898 ) | ( ~w2694 & w7900 ) | ( w7898 & w7900 ) ;
  assign w7902 = \pi17 ^ w7901 ;
  assign w7903 = ~w2973 & w4907 ;
  assign w7904 = ( w7894 & w7902 ) | ( w7894 & w7903 ) | ( w7902 & w7903 ) ;
  assign w7905 = ( w7870 & w7878 ) | ( w7870 & w7904 ) | ( w7878 & w7904 ) ;
  assign w7906 = ( w7864 & w7865 ) | ( w7864 & w7905 ) | ( w7865 & w7905 ) ;
  assign w7907 = ( w7848 & w7856 ) | ( w7848 & w7906 ) | ( w7856 & w7906 ) ;
  assign w7908 = ( w7844 & w7846 ) | ( w7844 & w7907 ) | ( w7846 & w7907 ) ;
  assign w7909 = ( w7828 & w7836 ) | ( w7828 & w7908 ) | ( w7836 & w7908 ) ;
  assign w7910 = ( w7818 & w7826 ) | ( w7818 & w7909 ) | ( w7826 & w7909 ) ;
  assign w7911 = ( w7808 & w7816 ) | ( w7808 & w7910 ) | ( w7816 & w7910 ) ;
  assign w7912 = ( w7804 & w7806 ) | ( w7804 & w7911 ) | ( w7806 & w7911 ) ;
  assign w7913 = ( w7794 & w7796 ) | ( w7794 & w7912 ) | ( w7796 & w7912 ) ;
  assign w7914 = ( w7784 & w7786 ) | ( w7784 & w7913 ) | ( w7786 & w7913 ) ;
  assign w7915 = ( w7768 & w7776 ) | ( w7768 & w7914 ) | ( w7776 & w7914 ) ;
  assign w7916 = ( w7758 & w7766 ) | ( w7758 & w7915 ) | ( w7766 & w7915 ) ;
  assign w7917 = ( w7754 & w7756 ) | ( w7754 & w7916 ) | ( w7756 & w7916 ) ;
  assign w7918 = ( w7744 & ~w7746 ) | ( w7744 & w7917 ) | ( ~w7746 & w7917 ) ;
  assign w7919 = ( w7734 & ~w7736 ) | ( w7734 & w7918 ) | ( ~w7736 & w7918 ) ;
  assign w7920 = ( w7724 & w7726 ) | ( w7724 & w7919 ) | ( w7726 & w7919 ) ;
  assign w7921 = ( w7714 & ~w7716 ) | ( w7714 & w7920 ) | ( ~w7716 & w7920 ) ;
  assign w7922 = ( w7704 & w7706 ) | ( w7704 & w7921 ) | ( w7706 & w7921 ) ;
  assign w7923 = ( w7694 & w7696 ) | ( w7694 & w7922 ) | ( w7696 & w7922 ) ;
  assign w7924 = w7631 ^ w7641 ;
  assign w7925 = w7633 ^ w7924 ;
  assign w7926 = w592 & ~w6549 ;
  assign w7927 = w721 & w6048 ;
  assign w7928 = ( w592 & ~w7926 ) | ( w592 & w7927 ) | ( ~w7926 & w7927 ) ;
  assign w7929 = w381 | w6637 ;
  assign w7930 = w3435 & ~w7928 ;
  assign w7931 = ( w6045 & w7928 ) | ( w6045 & ~w7930 ) | ( w7928 & ~w7930 ) ;
  assign w7932 = ( ~w381 & w7929 ) | ( ~w381 & w7931 ) | ( w7929 & w7931 ) ;
  assign w7933 = \pi14 ^ w7932 ;
  assign w7934 = ( w7923 & w7925 ) | ( w7923 & w7933 ) | ( w7925 & w7933 ) ;
  assign w7935 = w3647 & ~w6748 ;
  assign w7936 = w3715 & w6949 ;
  assign w7937 = ( w3647 & ~w7935 ) | ( w3647 & w7936 ) | ( ~w7935 & w7936 ) ;
  assign w7938 = w3548 | w7154 ;
  assign w7939 = w3725 & ~w7937 ;
  assign w7940 = ( w6751 & w7937 ) | ( w6751 & ~w7939 ) | ( w7937 & ~w7939 ) ;
  assign w7941 = ( ~w3548 & w7938 ) | ( ~w3548 & w7940 ) | ( w7938 & w7940 ) ;
  assign w7942 = \pi11 ^ w7941 ;
  assign w7943 = ( w7686 & w7934 ) | ( w7686 & w7942 ) | ( w7934 & w7942 ) ;
  assign w7944 = ~w7412 & w7413 ;
  assign w7945 = w4049 | w7411 ;
  assign w7946 = ~w4142 & w7673 ;
  assign w7947 = ( ~w4049 & w7945 ) | ( ~w4049 & w7946 ) | ( w7945 & w7946 ) ;
  assign w7948 = w3962 | w7944 ;
  assign w7949 = w4152 & ~w7947 ;
  assign w7950 = ( w7414 & w7947 ) | ( w7414 & ~w7949 ) | ( w7947 & ~w7949 ) ;
  assign w7951 = ( ~w3962 & w7948 ) | ( ~w3962 & w7950 ) | ( w7948 & w7950 ) ;
  assign w7952 = \pi08 ^ w7951 ;
  assign w7953 = ( ~w7684 & w7943 ) | ( ~w7684 & w7952 ) | ( w7943 & w7952 ) ;
  assign w7954 = ~w4142 & w7411 ;
  assign w7955 = ( ~w4600 & w7944 ) | ( ~w4600 & w7954 ) | ( w7944 & w7954 ) ;
  assign w7956 = w7673 | w7955 ;
  assign w7957 = ( ~w3962 & w7955 ) | ( ~w3962 & w7956 ) | ( w7955 & w7956 ) ;
  assign w7958 = w7954 | w7957 ;
  assign w7959 = w7660 ^ w7668 ;
  assign w7960 = w7670 ^ w7959 ;
  assign w7961 = w4722 & ~w7958 ;
  assign w7962 = ( w7414 & w7958 ) | ( w7414 & ~w7961 ) | ( w7958 & ~w7961 ) ;
  assign w7963 = \pi08 ^ w7962 ;
  assign w7964 = ( w7953 & w7960 ) | ( w7953 & w7963 ) | ( w7960 & w7963 ) ;
  assign w7965 = \pi08 ^ w7671 ;
  assign w7966 = w7678 ^ w7965 ;
  assign w7967 = w7680 ^ w7966 ;
  assign w7968 = w7686 ^ w7942 ;
  assign w7969 = w7934 ^ w7968 ;
  assign w7970 = w7694 ^ w7922 ;
  assign w7971 = w7696 ^ w7970 ;
  assign w7972 = w883 | w6048 ;
  assign w7973 = w721 & w6549 ;
  assign w7974 = ( ~w883 & w7972 ) | ( ~w883 & w7973 ) | ( w7972 & w7973 ) ;
  assign w7975 = w592 & ~w6637 ;
  assign w7976 = w3421 | w7974 ;
  assign w7977 = ( w6045 & w7974 ) | ( w6045 & w7976 ) | ( w7974 & w7976 ) ;
  assign w7978 = ( w592 & ~w7975 ) | ( w592 & w7977 ) | ( ~w7975 & w7977 ) ;
  assign w7979 = \pi14 ^ w7978 ;
  assign w7980 = w7704 ^ w7921 ;
  assign w7981 = w7706 ^ w7980 ;
  assign w7982 = w883 | w6549 ;
  assign w7983 = w979 & w6048 ;
  assign w7984 = ( ~w883 & w7982 ) | ( ~w883 & w7983 ) | ( w7982 & w7983 ) ;
  assign w7985 = w721 & ~w6637 ;
  assign w7986 = w4257 & ~w7984 ;
  assign w7987 = ( w6045 & w7984 ) | ( w6045 & ~w7986 ) | ( w7984 & ~w7986 ) ;
  assign w7988 = ( w721 & ~w7985 ) | ( w721 & w7987 ) | ( ~w7985 & w7987 ) ;
  assign w7989 = \pi14 ^ w7988 ;
  assign w7990 = w7714 ^ w7920 ;
  assign w7991 = w7716 ^ w7990 ;
  assign w7992 = w979 & ~w6549 ;
  assign w7993 = w1085 & w6048 ;
  assign w7994 = ( w979 & ~w7992 ) | ( w979 & w7993 ) | ( ~w7992 & w7993 ) ;
  assign w7995 = w883 | w6637 ;
  assign w7996 = w4273 & ~w7994 ;
  assign w7997 = ( w6045 & w7994 ) | ( w6045 & ~w7996 ) | ( w7994 & ~w7996 ) ;
  assign w7998 = ( ~w883 & w7995 ) | ( ~w883 & w7997 ) | ( w7995 & w7997 ) ;
  assign w7999 = \pi14 ^ w7998 ;
  assign w8000 = w7724 ^ w7919 ;
  assign w8001 = w7726 ^ w8000 ;
  assign w8002 = w1085 & ~w6549 ;
  assign w8003 = w1205 & w6048 ;
  assign w8004 = ( w1085 & ~w8002 ) | ( w1085 & w8003 ) | ( ~w8002 & w8003 ) ;
  assign w8005 = w979 & ~w6637 ;
  assign w8006 = w4666 | w8004 ;
  assign w8007 = ( w6045 & w8004 ) | ( w6045 & w8006 ) | ( w8004 & w8006 ) ;
  assign w8008 = ( w979 & ~w8005 ) | ( w979 & w8007 ) | ( ~w8005 & w8007 ) ;
  assign w8009 = \pi14 ^ w8008 ;
  assign w8010 = w7734 ^ w7918 ;
  assign w8011 = w7736 ^ w8010 ;
  assign w8012 = w1264 | w6048 ;
  assign w8013 = w1205 & w6549 ;
  assign w8014 = ( ~w1264 & w8012 ) | ( ~w1264 & w8013 ) | ( w8012 & w8013 ) ;
  assign w8015 = w1085 & ~w6637 ;
  assign w8016 = w4533 | w8014 ;
  assign w8017 = ( w6045 & w8014 ) | ( w6045 & w8016 ) | ( w8014 & w8016 ) ;
  assign w8018 = ( w1085 & ~w8015 ) | ( w1085 & w8017 ) | ( ~w8015 & w8017 ) ;
  assign w8019 = \pi14 ^ w8018 ;
  assign w8020 = w7744 ^ w7917 ;
  assign w8021 = w7746 ^ w8020 ;
  assign w8022 = w1264 | w6549 ;
  assign w8023 = w1399 & w6048 ;
  assign w8024 = ( ~w1264 & w8022 ) | ( ~w1264 & w8023 ) | ( w8022 & w8023 ) ;
  assign w8025 = w1205 & ~w6637 ;
  assign w8026 = w4864 & ~w8024 ;
  assign w8027 = ( w6045 & w8024 ) | ( w6045 & ~w8026 ) | ( w8024 & ~w8026 ) ;
  assign w8028 = ( w1205 & ~w8025 ) | ( w1205 & w8027 ) | ( ~w8025 & w8027 ) ;
  assign w8029 = \pi14 ^ w8028 ;
  assign w8030 = w7754 ^ w7916 ;
  assign w8031 = w7756 ^ w8030 ;
  assign w8032 = w1399 & ~w6549 ;
  assign w8033 = ~w1510 & w6048 ;
  assign w8034 = ( w1399 & ~w8032 ) | ( w1399 & w8033 ) | ( ~w8032 & w8033 ) ;
  assign w8035 = w1264 | w6637 ;
  assign w8036 = w4852 & ~w8034 ;
  assign w8037 = ( w6045 & w8034 ) | ( w6045 & ~w8036 ) | ( w8034 & ~w8036 ) ;
  assign w8038 = ( ~w1264 & w8035 ) | ( ~w1264 & w8037 ) | ( w8035 & w8037 ) ;
  assign w8039 = \pi14 ^ w8038 ;
  assign w8040 = w1614 & ~w6048 ;
  assign w8041 = ~w1510 & w6549 ;
  assign w8042 = ( w1614 & ~w8040 ) | ( w1614 & w8041 ) | ( ~w8040 & w8041 ) ;
  assign w8043 = w1399 & ~w6637 ;
  assign w8044 = w5069 & ~w8042 ;
  assign w8045 = ( w6045 & w8042 ) | ( w6045 & ~w8044 ) | ( w8042 & ~w8044 ) ;
  assign w8046 = ( w1399 & ~w8043 ) | ( w1399 & w8045 ) | ( ~w8043 & w8045 ) ;
  assign w8047 = \pi14 ^ w8046 ;
  assign w8048 = w7758 ^ w7915 ;
  assign w8049 = w7766 ^ w8048 ;
  assign w8050 = w1614 & ~w6549 ;
  assign w8051 = w1711 & w6048 ;
  assign w8052 = ( w1614 & ~w8050 ) | ( w1614 & w8051 ) | ( ~w8050 & w8051 ) ;
  assign w8053 = w1510 | w6637 ;
  assign w8054 = w5085 & ~w8052 ;
  assign w8055 = ( w6045 & w8052 ) | ( w6045 & ~w8054 ) | ( w8052 & ~w8054 ) ;
  assign w8056 = ( ~w1510 & w8053 ) | ( ~w1510 & w8055 ) | ( w8053 & w8055 ) ;
  assign w8057 = \pi14 ^ w8056 ;
  assign w8058 = w7768 ^ w7914 ;
  assign w8059 = w7776 ^ w8058 ;
  assign w8060 = w7784 ^ w7913 ;
  assign w8061 = w7786 ^ w8060 ;
  assign w8062 = w1711 & ~w6549 ;
  assign w8063 = ~w1834 & w6048 ;
  assign w8064 = ( w1711 & ~w8062 ) | ( w1711 & w8063 ) | ( ~w8062 & w8063 ) ;
  assign w8065 = w1614 & ~w6637 ;
  assign w8066 = w5433 & ~w8064 ;
  assign w8067 = ( w6045 & w8064 ) | ( w6045 & ~w8066 ) | ( w8064 & ~w8066 ) ;
  assign w8068 = ( w1614 & ~w8065 ) | ( w1614 & w8067 ) | ( ~w8065 & w8067 ) ;
  assign w8069 = \pi14 ^ w8068 ;
  assign w8070 = w7794 ^ w7912 ;
  assign w8071 = w7796 ^ w8070 ;
  assign w8072 = w1939 | w6048 ;
  assign w8073 = ~w1834 & w6549 ;
  assign w8074 = ( ~w1939 & w8072 ) | ( ~w1939 & w8073 ) | ( w8072 & w8073 ) ;
  assign w8075 = w1711 & ~w6637 ;
  assign w8076 = w5296 | w8074 ;
  assign w8077 = ( w6045 & w8074 ) | ( w6045 & w8076 ) | ( w8074 & w8076 ) ;
  assign w8078 = ( w1711 & ~w8075 ) | ( w1711 & w8077 ) | ( ~w8075 & w8077 ) ;
  assign w8079 = \pi14 ^ w8078 ;
  assign w8080 = w7804 ^ w7911 ;
  assign w8081 = w7806 ^ w8080 ;
  assign w8082 = w1939 | w6549 ;
  assign w8083 = w1976 & w6048 ;
  assign w8084 = ( ~w1939 & w8082 ) | ( ~w1939 & w8083 ) | ( w8082 & w8083 ) ;
  assign w8085 = w1834 | w6637 ;
  assign w8086 = w5659 & ~w8084 ;
  assign w8087 = ( w6045 & w8084 ) | ( w6045 & ~w8086 ) | ( w8084 & ~w8086 ) ;
  assign w8088 = ( ~w1834 & w8085 ) | ( ~w1834 & w8087 ) | ( w8085 & w8087 ) ;
  assign w8089 = \pi14 ^ w8088 ;
  assign w8090 = w2059 | w6048 ;
  assign w8091 = w1976 & w6549 ;
  assign w8092 = ( ~w2059 & w8090 ) | ( ~w2059 & w8091 ) | ( w8090 & w8091 ) ;
  assign w8093 = w1939 | w6637 ;
  assign w8094 = w5748 | w8092 ;
  assign w8095 = ( w6045 & w8092 ) | ( w6045 & w8094 ) | ( w8092 & w8094 ) ;
  assign w8096 = ( ~w1939 & w8093 ) | ( ~w1939 & w8095 ) | ( w8093 & w8095 ) ;
  assign w8097 = \pi14 ^ w8096 ;
  assign w8098 = w7808 ^ w7910 ;
  assign w8099 = w7816 ^ w8098 ;
  assign w8100 = w2059 | w6549 ;
  assign w8101 = ~w2130 & w6048 ;
  assign w8102 = ( ~w2059 & w8100 ) | ( ~w2059 & w8101 ) | ( w8100 & w8101 ) ;
  assign w8103 = w1976 & ~w6637 ;
  assign w8104 = w5646 | w8102 ;
  assign w8105 = ( w6045 & w8102 ) | ( w6045 & w8104 ) | ( w8102 & w8104 ) ;
  assign w8106 = ( w1976 & ~w8103 ) | ( w1976 & w8105 ) | ( ~w8103 & w8105 ) ;
  assign w8107 = \pi14 ^ w8106 ;
  assign w8108 = w7818 ^ w7909 ;
  assign w8109 = w7826 ^ w8108 ;
  assign w8110 = w2130 | w6549 ;
  assign w8111 = ~w2235 & w6048 ;
  assign w8112 = ( ~w2130 & w8110 ) | ( ~w2130 & w8111 ) | ( w8110 & w8111 ) ;
  assign w8113 = w2059 | w6637 ;
  assign w8114 = w5896 & ~w8112 ;
  assign w8115 = ( w6045 & w8112 ) | ( w6045 & ~w8114 ) | ( w8112 & ~w8114 ) ;
  assign w8116 = ( ~w2059 & w8113 ) | ( ~w2059 & w8115 ) | ( w8113 & w8115 ) ;
  assign w8117 = \pi14 ^ w8116 ;
  assign w8118 = w7828 ^ w7908 ;
  assign w8119 = w7836 ^ w8118 ;
  assign w8120 = w7844 ^ w7907 ;
  assign w8121 = w7846 ^ w8120 ;
  assign w8122 = w2273 & ~w6048 ;
  assign w8123 = ~w2235 & w6549 ;
  assign w8124 = ( w2273 & ~w8122 ) | ( w2273 & w8123 ) | ( ~w8122 & w8123 ) ;
  assign w8125 = w2130 | w6637 ;
  assign w8126 = w6094 | w8124 ;
  assign w8127 = ( w6045 & w8124 ) | ( w6045 & w8126 ) | ( w8124 & w8126 ) ;
  assign w8128 = ( ~w2130 & w8125 ) | ( ~w2130 & w8127 ) | ( w8125 & w8127 ) ;
  assign w8129 = \pi14 ^ w8128 ;
  assign w8130 = w7848 ^ w7906 ;
  assign w8131 = w7856 ^ w8130 ;
  assign w8132 = w2273 & ~w6549 ;
  assign w8133 = w2391 & w6048 ;
  assign w8134 = ( w2273 & ~w8132 ) | ( w2273 & w8133 ) | ( ~w8132 & w8133 ) ;
  assign w8135 = w2235 | w6637 ;
  assign w8136 = w6106 & ~w8134 ;
  assign w8137 = ( w6045 & w8134 ) | ( w6045 & ~w8136 ) | ( w8134 & ~w8136 ) ;
  assign w8138 = ( ~w2235 & w8135 ) | ( ~w2235 & w8137 ) | ( w8135 & w8137 ) ;
  assign w8139 = \pi14 ^ w8138 ;
  assign w8140 = w7864 ^ w7905 ;
  assign w8141 = w7865 ^ w8140 ;
  assign w8142 = w2391 & ~w6549 ;
  assign w8143 = w2500 & w6048 ;
  assign w8144 = ( w2391 & ~w8142 ) | ( w2391 & w8143 ) | ( ~w8142 & w8143 ) ;
  assign w8145 = w2273 & ~w6637 ;
  assign w8146 = w5880 | w8144 ;
  assign w8147 = ( w6045 & w8144 ) | ( w6045 & w8146 ) | ( w8144 & w8146 ) ;
  assign w8148 = ( w2273 & ~w8145 ) | ( w2273 & w8147 ) | ( ~w8145 & w8147 ) ;
  assign w8149 = \pi14 ^ w8148 ;
  assign w8150 = w2578 | w6048 ;
  assign w8151 = w2500 & w6549 ;
  assign w8152 = ( ~w2578 & w8150 ) | ( ~w2578 & w8151 ) | ( w8150 & w8151 ) ;
  assign w8153 = w2391 & ~w6637 ;
  assign w8154 = w6164 & ~w8152 ;
  assign w8155 = ( w6045 & w8152 ) | ( w6045 & ~w8154 ) | ( w8152 & ~w8154 ) ;
  assign w8156 = ( w2391 & ~w8153 ) | ( w2391 & w8155 ) | ( ~w8153 & w8155 ) ;
  assign w8157 = \pi14 ^ w8156 ;
  assign w8158 = w7878 ^ w7904 ;
  assign w8159 = w7870 ^ w8158 ;
  assign w8160 = w7894 ^ w7902 ;
  assign w8161 = w7903 ^ w8160 ;
  assign w8162 = w2578 | w6549 ;
  assign w8163 = ~w2653 & w6048 ;
  assign w8164 = ( ~w2578 & w8162 ) | ( ~w2578 & w8163 ) | ( w8162 & w8163 ) ;
  assign w8165 = w2500 & ~w6637 ;
  assign w8166 = w6219 | w8164 ;
  assign w8167 = ( w6045 & w8164 ) | ( w6045 & w8166 ) | ( w8164 & w8166 ) ;
  assign w8168 = ( w2500 & ~w8165 ) | ( w2500 & w8167 ) | ( ~w8165 & w8167 ) ;
  assign w8169 = \pi14 ^ w8168 ;
  assign w8170 = w2694 | w6048 ;
  assign w8171 = ~w2653 & w6549 ;
  assign w8172 = ( ~w2694 & w8170 ) | ( ~w2694 & w8171 ) | ( w8170 & w8171 ) ;
  assign w8173 = w2578 | w6637 ;
  assign w8174 = w6282 & ~w8172 ;
  assign w8175 = ( w6045 & w8172 ) | ( w6045 & ~w8174 ) | ( w8172 & ~w8174 ) ;
  assign w8176 = ( ~w2578 & w8173 ) | ( ~w2578 & w8175 ) | ( w8173 & w8175 ) ;
  assign w8177 = \pi14 ^ w8176 ;
  assign w8178 = w7885 ^ w7893 ;
  assign w8179 = ( \pi14 & \pi15 ) | ( \pi14 & ~w2871 ) | ( \pi15 & ~w2871 ) ;
  assign w8180 = \pi14 & \pi15 ;
  assign w8181 = w2973 ^ w8180 ;
  assign w8182 = ( \pi16 & w8180 ) | ( \pi16 & ~w8181 ) | ( w8180 & ~w8181 ) ;
  assign w8183 = w8179 ^ w8182 ;
  assign w8184 = w2805 & ~w6048 ;
  assign w8185 = ~w2694 & w6549 ;
  assign w8186 = ( w2805 & ~w8184 ) | ( w2805 & w8185 ) | ( ~w8184 & w8185 ) ;
  assign w8187 = w2653 | w6637 ;
  assign w8188 = w6338 & ~w8186 ;
  assign w8189 = ( w6045 & w8186 ) | ( w6045 & ~w8188 ) | ( w8186 & ~w8188 ) ;
  assign w8190 = ( ~w2653 & w8187 ) | ( ~w2653 & w8189 ) | ( w8187 & w8189 ) ;
  assign w8191 = \pi14 ^ w8190 ;
  assign w8192 = ( \pi11 & \pi12 ) | ( \pi11 & ~\pi14 ) | ( \pi12 & ~\pi14 ) ;
  assign w8193 = \pi14 & w2973 ;
  assign w8194 = w2871 & w8193 ;
  assign w8195 = ( \pi11 & \pi12 ) | ( \pi11 & ~w8194 ) | ( \pi12 & ~w8194 ) ;
  assign w8196 = ( \pi13 & \pi14 ) | ( \pi13 & ~w8195 ) | ( \pi14 & ~w8195 ) ;
  assign w8197 = ( \pi13 & ~w8193 ) | ( \pi13 & w8195 ) | ( ~w8193 & w8195 ) ;
  assign w8198 = ( w8192 & w8196 ) | ( w8192 & ~w8197 ) | ( w8196 & ~w8197 ) ;
  assign w8199 = w2973 | w6048 ;
  assign w8200 = ~w2871 & w6549 ;
  assign w8201 = ( ~w2973 & w8199 ) | ( ~w2973 & w8200 ) | ( w8199 & w8200 ) ;
  assign w8202 = w2805 & ~w6637 ;
  assign w8203 = w6457 | w8201 ;
  assign w8204 = ( w6045 & w8201 ) | ( w6045 & w8203 ) | ( w8201 & w8203 ) ;
  assign w8205 = ( w2805 & ~w8202 ) | ( w2805 & w8204 ) | ( ~w8202 & w8204 ) ;
  assign w8206 = \pi14 ^ w8205 ;
  assign w8207 = w8198 & w8206 ;
  assign w8208 = w2805 & ~w6549 ;
  assign w8209 = ~w2871 & w6048 ;
  assign w8210 = ( w2805 & ~w8208 ) | ( w2805 & w8209 ) | ( ~w8208 & w8209 ) ;
  assign w8211 = w2694 | w6637 ;
  assign w8212 = w6473 | w8210 ;
  assign w8213 = ( w6045 & w8210 ) | ( w6045 & w8212 ) | ( w8210 & w8212 ) ;
  assign w8214 = ( ~w2694 & w8211 ) | ( ~w2694 & w8213 ) | ( w8211 & w8213 ) ;
  assign w8215 = \pi14 ^ w8214 ;
  assign w8216 = ~w2973 & w5496 ;
  assign w8217 = ( w8207 & w8215 ) | ( w8207 & w8216 ) | ( w8215 & w8216 ) ;
  assign w8218 = ( w8183 & w8191 ) | ( w8183 & w8217 ) | ( w8191 & w8217 ) ;
  assign w8219 = ( w8177 & w8178 ) | ( w8177 & w8218 ) | ( w8178 & w8218 ) ;
  assign w8220 = ( w8161 & w8169 ) | ( w8161 & w8219 ) | ( w8169 & w8219 ) ;
  assign w8221 = ( w8157 & w8159 ) | ( w8157 & w8220 ) | ( w8159 & w8220 ) ;
  assign w8222 = ( w8141 & w8149 ) | ( w8141 & w8221 ) | ( w8149 & w8221 ) ;
  assign w8223 = ( w8131 & w8139 ) | ( w8131 & w8222 ) | ( w8139 & w8222 ) ;
  assign w8224 = ( w8121 & w8129 ) | ( w8121 & w8223 ) | ( w8129 & w8223 ) ;
  assign w8225 = ( w8117 & w8119 ) | ( w8117 & w8224 ) | ( w8119 & w8224 ) ;
  assign w8226 = ( w8107 & w8109 ) | ( w8107 & w8225 ) | ( w8109 & w8225 ) ;
  assign w8227 = ( w8097 & w8099 ) | ( w8097 & w8226 ) | ( w8099 & w8226 ) ;
  assign w8228 = ( w8081 & w8089 ) | ( w8081 & w8227 ) | ( w8089 & w8227 ) ;
  assign w8229 = ( w8071 & w8079 ) | ( w8071 & w8228 ) | ( w8079 & w8228 ) ;
  assign w8230 = ( w8061 & w8069 ) | ( w8061 & w8229 ) | ( w8069 & w8229 ) ;
  assign w8231 = ( w8057 & w8059 ) | ( w8057 & w8230 ) | ( w8059 & w8230 ) ;
  assign w8232 = ( w8047 & w8049 ) | ( w8047 & w8231 ) | ( w8049 & w8231 ) ;
  assign w8233 = ( w8031 & w8039 ) | ( w8031 & w8232 ) | ( w8039 & w8232 ) ;
  assign w8234 = ( ~w8021 & w8029 ) | ( ~w8021 & w8233 ) | ( w8029 & w8233 ) ;
  assign w8235 = ( ~w8011 & w8019 ) | ( ~w8011 & w8234 ) | ( w8019 & w8234 ) ;
  assign w8236 = ( w8001 & w8009 ) | ( w8001 & w8235 ) | ( w8009 & w8235 ) ;
  assign w8237 = ( ~w7991 & w7999 ) | ( ~w7991 & w8236 ) | ( w7999 & w8236 ) ;
  assign w8238 = ( w7981 & w7989 ) | ( w7981 & w8237 ) | ( w7989 & w8237 ) ;
  assign w8239 = ( w7971 & w7979 ) | ( w7971 & w8238 ) | ( w7979 & w8238 ) ;
  assign w8240 = w7923 ^ w7933 ;
  assign w8241 = w7925 ^ w8240 ;
  assign w8242 = w3647 & ~w6949 ;
  assign w8243 = ~w3094 & w6748 ;
  assign w8244 = ( w3647 & ~w8242 ) | ( w3647 & w8243 ) | ( ~w8242 & w8243 ) ;
  assign w8245 = w3715 & ~w7154 ;
  assign w8246 = w4164 & ~w8244 ;
  assign w8247 = ( w6751 & w8244 ) | ( w6751 & ~w8246 ) | ( w8244 & ~w8246 ) ;
  assign w8248 = ( w3715 & ~w8245 ) | ( w3715 & w8247 ) | ( ~w8245 & w8247 ) ;
  assign w8249 = \pi11 ^ w8248 ;
  assign w8250 = ( w8239 & w8241 ) | ( w8239 & w8249 ) | ( w8241 & w8249 ) ;
  assign w8251 = w4049 | w7673 ;
  assign w8252 = w3907 & w7411 ;
  assign w8253 = ( ~w4049 & w8251 ) | ( ~w4049 & w8252 ) | ( w8251 & w8252 ) ;
  assign w8254 = w4142 | w7944 ;
  assign w8255 = w4563 | w8253 ;
  assign w8256 = ( w7414 & w8253 ) | ( w7414 & w8255 ) | ( w8253 & w8255 ) ;
  assign w8257 = ( ~w4142 & w8254 ) | ( ~w4142 & w8256 ) | ( w8254 & w8256 ) ;
  assign w8258 = \pi08 ^ w8257 ;
  assign w8259 = ( w7969 & w8250 ) | ( w7969 & w8258 ) | ( w8250 & w8258 ) ;
  assign w8260 = ( \pi03 & ~\pi04 ) | ( \pi03 & \pi05 ) | ( ~\pi04 & \pi05 ) ;
  assign w8261 = ( \pi02 & \pi03 ) | ( \pi02 & w8260 ) | ( \pi03 & w8260 ) ;
  assign w8262 = w8260 ^ w8261 ;
  assign w8263 = w33 & w34 ;
  assign w8264 = ~w4600 & w8262 ;
  assign w8265 = w8263 | w8264 ;
  assign w8266 = ( ~w4603 & w8264 ) | ( ~w4603 & w8265 ) | ( w8264 & w8265 ) ;
  assign w8267 = \pi05 ^ w8266 ;
  assign w8268 = w7684 ^ w7952 ;
  assign w8269 = w7943 ^ w8268 ;
  assign w8270 = ( w8259 & w8267 ) | ( w8259 & ~w8269 ) | ( w8267 & ~w8269 ) ;
  assign w8271 = w4722 & w7414 ;
  assign w8272 = ( w7414 & w7958 ) | ( w7414 & ~w8271 ) | ( w7958 & ~w8271 ) ;
  assign w8273 = w7953 ^ w8272 ;
  assign w8274 = \pi08 ^ w7960 ;
  assign w8275 = w8273 ^ w8274 ;
  assign w8276 = w8267 ^ w8269 ;
  assign w8277 = w8259 ^ w8276 ;
  assign w8278 = w381 | w6748 ;
  assign w8279 = ~w3094 & w6949 ;
  assign w8280 = ( ~w381 & w8278 ) | ( ~w381 & w8279 ) | ( w8278 & w8279 ) ;
  assign w8281 = w3647 & ~w7154 ;
  assign w8282 = w3810 | w8280 ;
  assign w8283 = ( w6751 & w8280 ) | ( w6751 & w8282 ) | ( w8280 & w8282 ) ;
  assign w8284 = ( w3647 & ~w8281 ) | ( w3647 & w8283 ) | ( ~w8281 & w8283 ) ;
  assign w8285 = \pi11 ^ w8284 ;
  assign w8286 = w7971 ^ w8238 ;
  assign w8287 = w7979 ^ w8286 ;
  assign w8288 = w381 | w6949 ;
  assign w8289 = w592 & w6748 ;
  assign w8290 = ( ~w381 & w8288 ) | ( ~w381 & w8289 ) | ( w8288 & w8289 ) ;
  assign w8291 = w3094 | w7154 ;
  assign w8292 = w3096 | w8290 ;
  assign w8293 = ( w6751 & w8290 ) | ( w6751 & w8292 ) | ( w8290 & w8292 ) ;
  assign w8294 = ( ~w3094 & w8291 ) | ( ~w3094 & w8293 ) | ( w8291 & w8293 ) ;
  assign w8295 = \pi11 ^ w8294 ;
  assign w8296 = w7981 ^ w8237 ;
  assign w8297 = w7989 ^ w8296 ;
  assign w8298 = w592 & ~w6949 ;
  assign w8299 = w721 & w6748 ;
  assign w8300 = ( w592 & ~w8298 ) | ( w592 & w8299 ) | ( ~w8298 & w8299 ) ;
  assign w8301 = w381 | w7154 ;
  assign w8302 = w3435 & ~w8300 ;
  assign w8303 = ( w6751 & w8300 ) | ( w6751 & ~w8302 ) | ( w8300 & ~w8302 ) ;
  assign w8304 = ( ~w381 & w8301 ) | ( ~w381 & w8303 ) | ( w8301 & w8303 ) ;
  assign w8305 = \pi11 ^ w8304 ;
  assign w8306 = w7991 ^ w8236 ;
  assign w8307 = w7999 ^ w8306 ;
  assign w8308 = w883 | w6748 ;
  assign w8309 = w721 & w6949 ;
  assign w8310 = ( ~w883 & w8308 ) | ( ~w883 & w8309 ) | ( w8308 & w8309 ) ;
  assign w8311 = w592 & ~w7154 ;
  assign w8312 = w3421 | w8310 ;
  assign w8313 = ( w6751 & w8310 ) | ( w6751 & w8312 ) | ( w8310 & w8312 ) ;
  assign w8314 = ( w592 & ~w8311 ) | ( w592 & w8313 ) | ( ~w8311 & w8313 ) ;
  assign w8315 = \pi11 ^ w8314 ;
  assign w8316 = w8001 ^ w8235 ;
  assign w8317 = w8009 ^ w8316 ;
  assign w8318 = w883 | w6949 ;
  assign w8319 = w979 & w6748 ;
  assign w8320 = ( ~w883 & w8318 ) | ( ~w883 & w8319 ) | ( w8318 & w8319 ) ;
  assign w8321 = w721 & ~w7154 ;
  assign w8322 = w4257 & ~w8320 ;
  assign w8323 = ( w6751 & w8320 ) | ( w6751 & ~w8322 ) | ( w8320 & ~w8322 ) ;
  assign w8324 = ( w721 & ~w8321 ) | ( w721 & w8323 ) | ( ~w8321 & w8323 ) ;
  assign w8325 = \pi11 ^ w8324 ;
  assign w8326 = w8011 ^ w8234 ;
  assign w8327 = w8019 ^ w8326 ;
  assign w8328 = w979 & ~w6949 ;
  assign w8329 = w1085 & w6748 ;
  assign w8330 = ( w979 & ~w8328 ) | ( w979 & w8329 ) | ( ~w8328 & w8329 ) ;
  assign w8331 = w883 | w7154 ;
  assign w8332 = w4273 & ~w8330 ;
  assign w8333 = ( w6751 & w8330 ) | ( w6751 & ~w8332 ) | ( w8330 & ~w8332 ) ;
  assign w8334 = ( ~w883 & w8331 ) | ( ~w883 & w8333 ) | ( w8331 & w8333 ) ;
  assign w8335 = \pi11 ^ w8334 ;
  assign w8336 = w8021 ^ w8233 ;
  assign w8337 = w8029 ^ w8336 ;
  assign w8338 = w1085 & ~w6949 ;
  assign w8339 = w1205 & w6748 ;
  assign w8340 = ( w1085 & ~w8338 ) | ( w1085 & w8339 ) | ( ~w8338 & w8339 ) ;
  assign w8341 = w979 & ~w7154 ;
  assign w8342 = w4666 | w8340 ;
  assign w8343 = ( w6751 & w8340 ) | ( w6751 & w8342 ) | ( w8340 & w8342 ) ;
  assign w8344 = ( w979 & ~w8341 ) | ( w979 & w8343 ) | ( ~w8341 & w8343 ) ;
  assign w8345 = \pi11 ^ w8344 ;
  assign w8346 = w8031 ^ w8232 ;
  assign w8347 = w8039 ^ w8346 ;
  assign w8348 = w8047 ^ w8231 ;
  assign w8349 = w8049 ^ w8348 ;
  assign w8350 = w1264 | w6748 ;
  assign w8351 = w1205 & w6949 ;
  assign w8352 = ( ~w1264 & w8350 ) | ( ~w1264 & w8351 ) | ( w8350 & w8351 ) ;
  assign w8353 = w1085 & ~w7154 ;
  assign w8354 = w4533 | w8352 ;
  assign w8355 = ( w6751 & w8352 ) | ( w6751 & w8354 ) | ( w8352 & w8354 ) ;
  assign w8356 = ( w1085 & ~w8353 ) | ( w1085 & w8355 ) | ( ~w8353 & w8355 ) ;
  assign w8357 = \pi11 ^ w8356 ;
  assign w8358 = w8057 ^ w8230 ;
  assign w8359 = w8059 ^ w8358 ;
  assign w8360 = w1264 | w6949 ;
  assign w8361 = w1399 & w6748 ;
  assign w8362 = ( ~w1264 & w8360 ) | ( ~w1264 & w8361 ) | ( w8360 & w8361 ) ;
  assign w8363 = w1205 & ~w7154 ;
  assign w8364 = w4864 & ~w8362 ;
  assign w8365 = ( w6751 & w8362 ) | ( w6751 & ~w8364 ) | ( w8362 & ~w8364 ) ;
  assign w8366 = ( w1205 & ~w8363 ) | ( w1205 & w8365 ) | ( ~w8363 & w8365 ) ;
  assign w8367 = \pi11 ^ w8366 ;
  assign w8368 = w1399 & ~w6949 ;
  assign w8369 = ~w1510 & w6748 ;
  assign w8370 = ( w1399 & ~w8368 ) | ( w1399 & w8369 ) | ( ~w8368 & w8369 ) ;
  assign w8371 = w1264 | w7154 ;
  assign w8372 = w4852 & ~w8370 ;
  assign w8373 = ( w6751 & w8370 ) | ( w6751 & ~w8372 ) | ( w8370 & ~w8372 ) ;
  assign w8374 = ( ~w1264 & w8371 ) | ( ~w1264 & w8373 ) | ( w8371 & w8373 ) ;
  assign w8375 = \pi11 ^ w8374 ;
  assign w8376 = w8061 ^ w8229 ;
  assign w8377 = w8069 ^ w8376 ;
  assign w8378 = w1614 & ~w6748 ;
  assign w8379 = ~w1510 & w6949 ;
  assign w8380 = ( w1614 & ~w8378 ) | ( w1614 & w8379 ) | ( ~w8378 & w8379 ) ;
  assign w8381 = w1399 & ~w7154 ;
  assign w8382 = w5069 & ~w8380 ;
  assign w8383 = ( w6751 & w8380 ) | ( w6751 & ~w8382 ) | ( w8380 & ~w8382 ) ;
  assign w8384 = ( w1399 & ~w8381 ) | ( w1399 & w8383 ) | ( ~w8381 & w8383 ) ;
  assign w8385 = \pi11 ^ w8384 ;
  assign w8386 = w8071 ^ w8228 ;
  assign w8387 = w8079 ^ w8386 ;
  assign w8388 = w1614 & ~w6949 ;
  assign w8389 = w1711 & w6748 ;
  assign w8390 = ( w1614 & ~w8388 ) | ( w1614 & w8389 ) | ( ~w8388 & w8389 ) ;
  assign w8391 = w1510 | w7154 ;
  assign w8392 = w5085 & ~w8390 ;
  assign w8393 = ( w6751 & w8390 ) | ( w6751 & ~w8392 ) | ( w8390 & ~w8392 ) ;
  assign w8394 = ( ~w1510 & w8391 ) | ( ~w1510 & w8393 ) | ( w8391 & w8393 ) ;
  assign w8395 = \pi11 ^ w8394 ;
  assign w8396 = w8081 ^ w8227 ;
  assign w8397 = w8089 ^ w8396 ;
  assign w8398 = w8097 ^ w8226 ;
  assign w8399 = w8099 ^ w8398 ;
  assign w8400 = w1711 & ~w6949 ;
  assign w8401 = ~w1834 & w6748 ;
  assign w8402 = ( w1711 & ~w8400 ) | ( w1711 & w8401 ) | ( ~w8400 & w8401 ) ;
  assign w8403 = w1614 & ~w7154 ;
  assign w8404 = w5433 & ~w8402 ;
  assign w8405 = ( w6751 & w8402 ) | ( w6751 & ~w8404 ) | ( w8402 & ~w8404 ) ;
  assign w8406 = ( w1614 & ~w8403 ) | ( w1614 & w8405 ) | ( ~w8403 & w8405 ) ;
  assign w8407 = \pi11 ^ w8406 ;
  assign w8408 = w8107 ^ w8225 ;
  assign w8409 = w8109 ^ w8408 ;
  assign w8410 = w1939 | w6748 ;
  assign w8411 = ~w1834 & w6949 ;
  assign w8412 = ( ~w1939 & w8410 ) | ( ~w1939 & w8411 ) | ( w8410 & w8411 ) ;
  assign w8413 = w1711 & ~w7154 ;
  assign w8414 = w5296 | w8412 ;
  assign w8415 = ( w6751 & w8412 ) | ( w6751 & w8414 ) | ( w8412 & w8414 ) ;
  assign w8416 = ( w1711 & ~w8413 ) | ( w1711 & w8415 ) | ( ~w8413 & w8415 ) ;
  assign w8417 = \pi11 ^ w8416 ;
  assign w8418 = w8117 ^ w8224 ;
  assign w8419 = w8119 ^ w8418 ;
  assign w8420 = w1939 | w6949 ;
  assign w8421 = w1976 & w6748 ;
  assign w8422 = ( ~w1939 & w8420 ) | ( ~w1939 & w8421 ) | ( w8420 & w8421 ) ;
  assign w8423 = w1834 | w7154 ;
  assign w8424 = w5659 & ~w8422 ;
  assign w8425 = ( w6751 & w8422 ) | ( w6751 & ~w8424 ) | ( w8422 & ~w8424 ) ;
  assign w8426 = ( ~w1834 & w8423 ) | ( ~w1834 & w8425 ) | ( w8423 & w8425 ) ;
  assign w8427 = \pi11 ^ w8426 ;
  assign w8428 = w2059 | w6748 ;
  assign w8429 = w1976 & w6949 ;
  assign w8430 = ( ~w2059 & w8428 ) | ( ~w2059 & w8429 ) | ( w8428 & w8429 ) ;
  assign w8431 = w1939 | w7154 ;
  assign w8432 = w5748 | w8430 ;
  assign w8433 = ( w6751 & w8430 ) | ( w6751 & w8432 ) | ( w8430 & w8432 ) ;
  assign w8434 = ( ~w1939 & w8431 ) | ( ~w1939 & w8433 ) | ( w8431 & w8433 ) ;
  assign w8435 = \pi11 ^ w8434 ;
  assign w8436 = w8121 ^ w8223 ;
  assign w8437 = w8129 ^ w8436 ;
  assign w8438 = w2059 | w6949 ;
  assign w8439 = ~w2130 & w6748 ;
  assign w8440 = ( ~w2059 & w8438 ) | ( ~w2059 & w8439 ) | ( w8438 & w8439 ) ;
  assign w8441 = w1976 & ~w7154 ;
  assign w8442 = w5646 | w8440 ;
  assign w8443 = ( w6751 & w8440 ) | ( w6751 & w8442 ) | ( w8440 & w8442 ) ;
  assign w8444 = ( w1976 & ~w8441 ) | ( w1976 & w8443 ) | ( ~w8441 & w8443 ) ;
  assign w8445 = \pi11 ^ w8444 ;
  assign w8446 = w8131 ^ w8222 ;
  assign w8447 = w8139 ^ w8446 ;
  assign w8448 = w2130 | w6949 ;
  assign w8449 = ~w2235 & w6748 ;
  assign w8450 = ( ~w2130 & w8448 ) | ( ~w2130 & w8449 ) | ( w8448 & w8449 ) ;
  assign w8451 = w2059 | w7154 ;
  assign w8452 = w5896 & ~w8450 ;
  assign w8453 = ( w6751 & w8450 ) | ( w6751 & ~w8452 ) | ( w8450 & ~w8452 ) ;
  assign w8454 = ( ~w2059 & w8451 ) | ( ~w2059 & w8453 ) | ( w8451 & w8453 ) ;
  assign w8455 = \pi11 ^ w8454 ;
  assign w8456 = w8141 ^ w8221 ;
  assign w8457 = w8149 ^ w8456 ;
  assign w8458 = w8157 ^ w8220 ;
  assign w8459 = w8159 ^ w8458 ;
  assign w8460 = w2273 & ~w6748 ;
  assign w8461 = ~w2235 & w6949 ;
  assign w8462 = ( w2273 & ~w8460 ) | ( w2273 & w8461 ) | ( ~w8460 & w8461 ) ;
  assign w8463 = w2130 | w7154 ;
  assign w8464 = w6094 | w8462 ;
  assign w8465 = ( w6751 & w8462 ) | ( w6751 & w8464 ) | ( w8462 & w8464 ) ;
  assign w8466 = ( ~w2130 & w8463 ) | ( ~w2130 & w8465 ) | ( w8463 & w8465 ) ;
  assign w8467 = \pi11 ^ w8466 ;
  assign w8468 = w8161 ^ w8219 ;
  assign w8469 = w8169 ^ w8468 ;
  assign w8470 = w2273 & ~w6949 ;
  assign w8471 = w2391 & w6748 ;
  assign w8472 = ( w2273 & ~w8470 ) | ( w2273 & w8471 ) | ( ~w8470 & w8471 ) ;
  assign w8473 = w2235 | w7154 ;
  assign w8474 = w6106 & ~w8472 ;
  assign w8475 = ( w6751 & w8472 ) | ( w6751 & ~w8474 ) | ( w8472 & ~w8474 ) ;
  assign w8476 = ( ~w2235 & w8473 ) | ( ~w2235 & w8475 ) | ( w8473 & w8475 ) ;
  assign w8477 = \pi11 ^ w8476 ;
  assign w8478 = w8177 ^ w8218 ;
  assign w8479 = w8178 ^ w8478 ;
  assign w8480 = w2391 & ~w6949 ;
  assign w8481 = w2500 & w6748 ;
  assign w8482 = ( w2391 & ~w8480 ) | ( w2391 & w8481 ) | ( ~w8480 & w8481 ) ;
  assign w8483 = w2273 & ~w7154 ;
  assign w8484 = w5880 | w8482 ;
  assign w8485 = ( w6751 & w8482 ) | ( w6751 & w8484 ) | ( w8482 & w8484 ) ;
  assign w8486 = ( w2273 & ~w8483 ) | ( w2273 & w8485 ) | ( ~w8483 & w8485 ) ;
  assign w8487 = \pi11 ^ w8486 ;
  assign w8488 = w2578 | w6748 ;
  assign w8489 = w2500 & w6949 ;
  assign w8490 = ( ~w2578 & w8488 ) | ( ~w2578 & w8489 ) | ( w8488 & w8489 ) ;
  assign w8491 = w2391 & ~w7154 ;
  assign w8492 = w6164 & ~w8490 ;
  assign w8493 = ( w6751 & w8490 ) | ( w6751 & ~w8492 ) | ( w8490 & ~w8492 ) ;
  assign w8494 = ( w2391 & ~w8491 ) | ( w2391 & w8493 ) | ( ~w8491 & w8493 ) ;
  assign w8495 = \pi11 ^ w8494 ;
  assign w8496 = w8191 ^ w8217 ;
  assign w8497 = w8183 ^ w8496 ;
  assign w8498 = w8207 ^ w8215 ;
  assign w8499 = w8216 ^ w8498 ;
  assign w8500 = w2578 | w6949 ;
  assign w8501 = ~w2653 & w6748 ;
  assign w8502 = ( ~w2578 & w8500 ) | ( ~w2578 & w8501 ) | ( w8500 & w8501 ) ;
  assign w8503 = w2500 & ~w7154 ;
  assign w8504 = w6219 | w8502 ;
  assign w8505 = ( w6751 & w8502 ) | ( w6751 & w8504 ) | ( w8502 & w8504 ) ;
  assign w8506 = ( w2500 & ~w8503 ) | ( w2500 & w8505 ) | ( ~w8503 & w8505 ) ;
  assign w8507 = \pi11 ^ w8506 ;
  assign w8508 = w2694 | w6748 ;
  assign w8509 = ~w2653 & w6949 ;
  assign w8510 = ( ~w2694 & w8508 ) | ( ~w2694 & w8509 ) | ( w8508 & w8509 ) ;
  assign w8511 = w2578 | w7154 ;
  assign w8512 = w6282 & ~w8510 ;
  assign w8513 = ( w6751 & w8510 ) | ( w6751 & ~w8512 ) | ( w8510 & ~w8512 ) ;
  assign w8514 = ( ~w2578 & w8511 ) | ( ~w2578 & w8513 ) | ( w8511 & w8513 ) ;
  assign w8515 = \pi11 ^ w8514 ;
  assign w8516 = w8198 ^ w8206 ;
  assign w8517 = ( \pi11 & \pi12 ) | ( \pi11 & ~w2871 ) | ( \pi12 & ~w2871 ) ;
  assign w8518 = \pi11 & \pi12 ;
  assign w8519 = w2973 ^ w8518 ;
  assign w8520 = ( \pi13 & w8518 ) | ( \pi13 & ~w8519 ) | ( w8518 & ~w8519 ) ;
  assign w8521 = w8517 ^ w8520 ;
  assign w8522 = w2805 & ~w6748 ;
  assign w8523 = ~w2694 & w6949 ;
  assign w8524 = ( w2805 & ~w8522 ) | ( w2805 & w8523 ) | ( ~w8522 & w8523 ) ;
  assign w8525 = w2653 | w7154 ;
  assign w8526 = w6338 & ~w8524 ;
  assign w8527 = ( w6751 & w8524 ) | ( w6751 & ~w8526 ) | ( w8524 & ~w8526 ) ;
  assign w8528 = ( ~w2653 & w8525 ) | ( ~w2653 & w8527 ) | ( w8525 & w8527 ) ;
  assign w8529 = \pi11 ^ w8528 ;
  assign w8530 = ( \pi08 & \pi09 ) | ( \pi08 & ~\pi11 ) | ( \pi09 & ~\pi11 ) ;
  assign w8531 = \pi11 & w2973 ;
  assign w8532 = w2871 & w8531 ;
  assign w8533 = ( \pi08 & \pi09 ) | ( \pi08 & ~w8532 ) | ( \pi09 & ~w8532 ) ;
  assign w8534 = ( \pi10 & \pi11 ) | ( \pi10 & ~w8533 ) | ( \pi11 & ~w8533 ) ;
  assign w8535 = ( \pi10 & ~w8531 ) | ( \pi10 & w8533 ) | ( ~w8531 & w8533 ) ;
  assign w8536 = ( w8530 & w8534 ) | ( w8530 & ~w8535 ) | ( w8534 & ~w8535 ) ;
  assign w8537 = w2973 | w6748 ;
  assign w8538 = ~w2871 & w6949 ;
  assign w8539 = ( ~w2973 & w8537 ) | ( ~w2973 & w8538 ) | ( w8537 & w8538 ) ;
  assign w8540 = w2805 & ~w7154 ;
  assign w8541 = w6457 | w8539 ;
  assign w8542 = ( w6751 & w8539 ) | ( w6751 & w8541 ) | ( w8539 & w8541 ) ;
  assign w8543 = ( w2805 & ~w8540 ) | ( w2805 & w8542 ) | ( ~w8540 & w8542 ) ;
  assign w8544 = \pi11 ^ w8543 ;
  assign w8545 = w8536 & w8544 ;
  assign w8546 = w2805 & ~w6949 ;
  assign w8547 = ~w2871 & w6748 ;
  assign w8548 = ( w2805 & ~w8546 ) | ( w2805 & w8547 ) | ( ~w8546 & w8547 ) ;
  assign w8549 = w2694 | w7154 ;
  assign w8550 = w6473 | w8548 ;
  assign w8551 = ( w6751 & w8548 ) | ( w6751 & w8550 ) | ( w8548 & w8550 ) ;
  assign w8552 = ( ~w2694 & w8549 ) | ( ~w2694 & w8551 ) | ( w8549 & w8551 ) ;
  assign w8553 = \pi11 ^ w8552 ;
  assign w8554 = ~w2973 & w6044 ;
  assign w8555 = ( w8545 & w8553 ) | ( w8545 & w8554 ) | ( w8553 & w8554 ) ;
  assign w8556 = ( w8521 & w8529 ) | ( w8521 & w8555 ) | ( w8529 & w8555 ) ;
  assign w8557 = ( w8515 & w8516 ) | ( w8515 & w8556 ) | ( w8516 & w8556 ) ;
  assign w8558 = ( w8499 & w8507 ) | ( w8499 & w8557 ) | ( w8507 & w8557 ) ;
  assign w8559 = ( w8495 & w8497 ) | ( w8495 & w8558 ) | ( w8497 & w8558 ) ;
  assign w8560 = ( w8479 & w8487 ) | ( w8479 & w8559 ) | ( w8487 & w8559 ) ;
  assign w8561 = ( w8469 & w8477 ) | ( w8469 & w8560 ) | ( w8477 & w8560 ) ;
  assign w8562 = ( w8459 & w8467 ) | ( w8459 & w8561 ) | ( w8467 & w8561 ) ;
  assign w8563 = ( w8455 & w8457 ) | ( w8455 & w8562 ) | ( w8457 & w8562 ) ;
  assign w8564 = ( w8445 & w8447 ) | ( w8445 & w8563 ) | ( w8447 & w8563 ) ;
  assign w8565 = ( w8435 & w8437 ) | ( w8435 & w8564 ) | ( w8437 & w8564 ) ;
  assign w8566 = ( w8419 & w8427 ) | ( w8419 & w8565 ) | ( w8427 & w8565 ) ;
  assign w8567 = ( w8409 & w8417 ) | ( w8409 & w8566 ) | ( w8417 & w8566 ) ;
  assign w8568 = ( w8399 & w8407 ) | ( w8399 & w8567 ) | ( w8407 & w8567 ) ;
  assign w8569 = ( w8395 & w8397 ) | ( w8395 & w8568 ) | ( w8397 & w8568 ) ;
  assign w8570 = ( w8385 & w8387 ) | ( w8385 & w8569 ) | ( w8387 & w8569 ) ;
  assign w8571 = ( w8375 & w8377 ) | ( w8375 & w8570 ) | ( w8377 & w8570 ) ;
  assign w8572 = ( w8359 & w8367 ) | ( w8359 & w8571 ) | ( w8367 & w8571 ) ;
  assign w8573 = ( w8349 & w8357 ) | ( w8349 & w8572 ) | ( w8357 & w8572 ) ;
  assign w8574 = ( w8345 & w8347 ) | ( w8345 & w8573 ) | ( w8347 & w8573 ) ;
  assign w8575 = ( w8335 & ~w8337 ) | ( w8335 & w8574 ) | ( ~w8337 & w8574 ) ;
  assign w8576 = ( w8325 & ~w8327 ) | ( w8325 & w8575 ) | ( ~w8327 & w8575 ) ;
  assign w8577 = ( w8315 & w8317 ) | ( w8315 & w8576 ) | ( w8317 & w8576 ) ;
  assign w8578 = ( w8305 & ~w8307 ) | ( w8305 & w8577 ) | ( ~w8307 & w8577 ) ;
  assign w8579 = ( w8295 & w8297 ) | ( w8295 & w8578 ) | ( w8297 & w8578 ) ;
  assign w8580 = ( w8285 & w8287 ) | ( w8285 & w8579 ) | ( w8287 & w8579 ) ;
  assign w8581 = w8239 ^ w8249 ;
  assign w8582 = w8241 ^ w8581 ;
  assign w8583 = w3548 | w7411 ;
  assign w8584 = w3907 & w7673 ;
  assign w8585 = ( ~w3548 & w8583 ) | ( ~w3548 & w8584 ) | ( w8583 & w8584 ) ;
  assign w8586 = w4049 | w7944 ;
  assign w8587 = w4622 & ~w8585 ;
  assign w8588 = ( w7414 & w8585 ) | ( w7414 & ~w8587 ) | ( w8585 & ~w8587 ) ;
  assign w8589 = ( ~w4049 & w8586 ) | ( ~w4049 & w8588 ) | ( w8586 & w8588 ) ;
  assign w8590 = \pi08 ^ w8589 ;
  assign w8591 = ( w8580 & w8582 ) | ( w8580 & w8590 ) | ( w8582 & w8590 ) ;
  assign w8592 = ( \pi02 & \pi03 ) | ( \pi02 & \pi04 ) | ( \pi03 & \pi04 ) ;
  assign w8593 = \pi04 ^ w8592 ;
  assign w8594 = ~w4600 & w8593 ;
  assign w8595 = ( w3962 & w6551 ) | ( w3962 & w8263 ) | ( w6551 & w8263 ) ;
  assign w8596 = w3962 | w8262 ;
  assign w8597 = ( ~w3962 & w8595 ) | ( ~w3962 & w8596 ) | ( w8595 & w8596 ) ;
  assign w8598 = ( ~w6555 & w8594 ) | ( ~w6555 & w8597 ) | ( w8594 & w8597 ) ;
  assign w8599 = w7969 ^ w8258 ;
  assign w8600 = w8250 ^ w8599 ;
  assign w8601 = \pi05 ^ w8598 ;
  assign w8602 = ( w8591 & w8600 ) | ( w8591 & w8601 ) | ( w8600 & w8601 ) ;
  assign w8603 = w8285 ^ w8579 ;
  assign w8604 = w8287 ^ w8603 ;
  assign w8605 = w3548 | w7673 ;
  assign w8606 = w3715 & w7411 ;
  assign w8607 = ( ~w3548 & w8605 ) | ( ~w3548 & w8606 ) | ( w8605 & w8606 ) ;
  assign w8608 = w3907 & ~w7944 ;
  assign w8609 = w3913 & ~w8607 ;
  assign w8610 = ( w7414 & w8607 ) | ( w7414 & ~w8609 ) | ( w8607 & ~w8609 ) ;
  assign w8611 = ( w3907 & ~w8608 ) | ( w3907 & w8610 ) | ( ~w8608 & w8610 ) ;
  assign w8612 = \pi08 ^ w8611 ;
  assign w8613 = w8295 ^ w8578 ;
  assign w8614 = w8297 ^ w8613 ;
  assign w8615 = w3647 & ~w7411 ;
  assign w8616 = w3715 & w7673 ;
  assign w8617 = ( w3647 & ~w8615 ) | ( w3647 & w8616 ) | ( ~w8615 & w8616 ) ;
  assign w8618 = w3548 | w7944 ;
  assign w8619 = w3725 & ~w8617 ;
  assign w8620 = ( w7414 & w8617 ) | ( w7414 & ~w8619 ) | ( w8617 & ~w8619 ) ;
  assign w8621 = ( ~w3548 & w8618 ) | ( ~w3548 & w8620 ) | ( w8618 & w8620 ) ;
  assign w8622 = \pi08 ^ w8621 ;
  assign w8623 = w8305 ^ w8577 ;
  assign w8624 = w8307 ^ w8623 ;
  assign w8625 = w3647 & ~w7673 ;
  assign w8626 = ~w3094 & w7411 ;
  assign w8627 = ( w3647 & ~w8625 ) | ( w3647 & w8626 ) | ( ~w8625 & w8626 ) ;
  assign w8628 = w3715 & ~w7944 ;
  assign w8629 = w4164 & ~w8627 ;
  assign w8630 = ( w7414 & w8627 ) | ( w7414 & ~w8629 ) | ( w8627 & ~w8629 ) ;
  assign w8631 = ( w3715 & ~w8628 ) | ( w3715 & w8630 ) | ( ~w8628 & w8630 ) ;
  assign w8632 = \pi08 ^ w8631 ;
  assign w8633 = w8315 ^ w8576 ;
  assign w8634 = w8317 ^ w8633 ;
  assign w8635 = w381 | w7411 ;
  assign w8636 = ~w3094 & w7673 ;
  assign w8637 = ( ~w381 & w8635 ) | ( ~w381 & w8636 ) | ( w8635 & w8636 ) ;
  assign w8638 = w3647 & ~w7944 ;
  assign w8639 = w3810 | w8637 ;
  assign w8640 = ( w7414 & w8637 ) | ( w7414 & w8639 ) | ( w8637 & w8639 ) ;
  assign w8641 = ( w3647 & ~w8638 ) | ( w3647 & w8640 ) | ( ~w8638 & w8640 ) ;
  assign w8642 = \pi08 ^ w8641 ;
  assign w8643 = w8325 ^ w8575 ;
  assign w8644 = w8327 ^ w8643 ;
  assign w8645 = w381 | w7673 ;
  assign w8646 = w592 & w7411 ;
  assign w8647 = ( ~w381 & w8645 ) | ( ~w381 & w8646 ) | ( w8645 & w8646 ) ;
  assign w8648 = w3094 | w7944 ;
  assign w8649 = w3096 | w8647 ;
  assign w8650 = ( w7414 & w8647 ) | ( w7414 & w8649 ) | ( w8647 & w8649 ) ;
  assign w8651 = ( ~w3094 & w8648 ) | ( ~w3094 & w8650 ) | ( w8648 & w8650 ) ;
  assign w8652 = \pi08 ^ w8651 ;
  assign w8653 = w8335 ^ w8574 ;
  assign w8654 = w8337 ^ w8653 ;
  assign w8655 = w592 & ~w7673 ;
  assign w8656 = w721 & w7411 ;
  assign w8657 = ( w592 & ~w8655 ) | ( w592 & w8656 ) | ( ~w8655 & w8656 ) ;
  assign w8658 = w381 | w7944 ;
  assign w8659 = w3435 & ~w8657 ;
  assign w8660 = ( w7414 & w8657 ) | ( w7414 & ~w8659 ) | ( w8657 & ~w8659 ) ;
  assign w8661 = ( ~w381 & w8658 ) | ( ~w381 & w8660 ) | ( w8658 & w8660 ) ;
  assign w8662 = \pi08 ^ w8661 ;
  assign w8663 = w8345 ^ w8573 ;
  assign w8664 = w8347 ^ w8663 ;
  assign w8665 = w883 | w7411 ;
  assign w8666 = w721 & w7673 ;
  assign w8667 = ( ~w883 & w8665 ) | ( ~w883 & w8666 ) | ( w8665 & w8666 ) ;
  assign w8668 = w592 & ~w7944 ;
  assign w8669 = w3421 | w8667 ;
  assign w8670 = ( w7414 & w8667 ) | ( w7414 & w8669 ) | ( w8667 & w8669 ) ;
  assign w8671 = ( w592 & ~w8668 ) | ( w592 & w8670 ) | ( ~w8668 & w8670 ) ;
  assign w8672 = \pi08 ^ w8671 ;
  assign w8673 = w883 | w7673 ;
  assign w8674 = w979 & w7411 ;
  assign w8675 = ( ~w883 & w8673 ) | ( ~w883 & w8674 ) | ( w8673 & w8674 ) ;
  assign w8676 = w721 & ~w7944 ;
  assign w8677 = w4257 & ~w8675 ;
  assign w8678 = ( w7414 & w8675 ) | ( w7414 & ~w8677 ) | ( w8675 & ~w8677 ) ;
  assign w8679 = ( w721 & ~w8676 ) | ( w721 & w8678 ) | ( ~w8676 & w8678 ) ;
  assign w8680 = \pi08 ^ w8679 ;
  assign w8681 = w8349 ^ w8572 ;
  assign w8682 = w8357 ^ w8681 ;
  assign w8683 = w979 & ~w7673 ;
  assign w8684 = w1085 & w7411 ;
  assign w8685 = ( w979 & ~w8683 ) | ( w979 & w8684 ) | ( ~w8683 & w8684 ) ;
  assign w8686 = w883 | w7944 ;
  assign w8687 = w4273 & ~w8685 ;
  assign w8688 = ( w7414 & w8685 ) | ( w7414 & ~w8687 ) | ( w8685 & ~w8687 ) ;
  assign w8689 = ( ~w883 & w8686 ) | ( ~w883 & w8688 ) | ( w8686 & w8688 ) ;
  assign w8690 = \pi08 ^ w8689 ;
  assign w8691 = w8359 ^ w8571 ;
  assign w8692 = w8367 ^ w8691 ;
  assign w8693 = w8375 ^ w8570 ;
  assign w8694 = w8377 ^ w8693 ;
  assign w8695 = w1085 & ~w7673 ;
  assign w8696 = w1205 & w7411 ;
  assign w8697 = ( w1085 & ~w8695 ) | ( w1085 & w8696 ) | ( ~w8695 & w8696 ) ;
  assign w8698 = w979 & ~w7944 ;
  assign w8699 = w4666 | w8697 ;
  assign w8700 = ( w7414 & w8697 ) | ( w7414 & w8699 ) | ( w8697 & w8699 ) ;
  assign w8701 = ( w979 & ~w8698 ) | ( w979 & w8700 ) | ( ~w8698 & w8700 ) ;
  assign w8702 = \pi08 ^ w8701 ;
  assign w8703 = w8385 ^ w8569 ;
  assign w8704 = w8387 ^ w8703 ;
  assign w8705 = w1264 | w7411 ;
  assign w8706 = w1205 & w7673 ;
  assign w8707 = ( ~w1264 & w8705 ) | ( ~w1264 & w8706 ) | ( w8705 & w8706 ) ;
  assign w8708 = w1085 & ~w7944 ;
  assign w8709 = w4533 | w8707 ;
  assign w8710 = ( w7414 & w8707 ) | ( w7414 & w8709 ) | ( w8707 & w8709 ) ;
  assign w8711 = ( w1085 & ~w8708 ) | ( w1085 & w8710 ) | ( ~w8708 & w8710 ) ;
  assign w8712 = \pi08 ^ w8711 ;
  assign w8713 = w8395 ^ w8568 ;
  assign w8714 = w8397 ^ w8713 ;
  assign w8715 = w1264 | w7673 ;
  assign w8716 = w1399 & w7411 ;
  assign w8717 = ( ~w1264 & w8715 ) | ( ~w1264 & w8716 ) | ( w8715 & w8716 ) ;
  assign w8718 = w1205 & ~w7944 ;
  assign w8719 = w4864 & ~w8717 ;
  assign w8720 = ( w7414 & w8717 ) | ( w7414 & ~w8719 ) | ( w8717 & ~w8719 ) ;
  assign w8721 = ( w1205 & ~w8718 ) | ( w1205 & w8720 ) | ( ~w8718 & w8720 ) ;
  assign w8722 = \pi08 ^ w8721 ;
  assign w8723 = w1399 & ~w7673 ;
  assign w8724 = ~w1510 & w7411 ;
  assign w8725 = ( w1399 & ~w8723 ) | ( w1399 & w8724 ) | ( ~w8723 & w8724 ) ;
  assign w8726 = w1264 | w7944 ;
  assign w8727 = w4852 & ~w8725 ;
  assign w8728 = ( w7414 & w8725 ) | ( w7414 & ~w8727 ) | ( w8725 & ~w8727 ) ;
  assign w8729 = ( ~w1264 & w8726 ) | ( ~w1264 & w8728 ) | ( w8726 & w8728 ) ;
  assign w8730 = \pi08 ^ w8729 ;
  assign w8731 = w8399 ^ w8567 ;
  assign w8732 = w8407 ^ w8731 ;
  assign w8733 = w1614 & ~w7411 ;
  assign w8734 = ~w1510 & w7673 ;
  assign w8735 = ( w1614 & ~w8733 ) | ( w1614 & w8734 ) | ( ~w8733 & w8734 ) ;
  assign w8736 = w1399 & ~w7944 ;
  assign w8737 = w5069 & ~w8735 ;
  assign w8738 = ( w7414 & w8735 ) | ( w7414 & ~w8737 ) | ( w8735 & ~w8737 ) ;
  assign w8739 = ( w1399 & ~w8736 ) | ( w1399 & w8738 ) | ( ~w8736 & w8738 ) ;
  assign w8740 = \pi08 ^ w8739 ;
  assign w8741 = w8409 ^ w8566 ;
  assign w8742 = w8417 ^ w8741 ;
  assign w8743 = w1614 & ~w7673 ;
  assign w8744 = w1711 & w7411 ;
  assign w8745 = ( w1614 & ~w8743 ) | ( w1614 & w8744 ) | ( ~w8743 & w8744 ) ;
  assign w8746 = w1510 | w7944 ;
  assign w8747 = w5085 & ~w8745 ;
  assign w8748 = ( w7414 & w8745 ) | ( w7414 & ~w8747 ) | ( w8745 & ~w8747 ) ;
  assign w8749 = ( ~w1510 & w8746 ) | ( ~w1510 & w8748 ) | ( w8746 & w8748 ) ;
  assign w8750 = \pi08 ^ w8749 ;
  assign w8751 = w8419 ^ w8565 ;
  assign w8752 = w8427 ^ w8751 ;
  assign w8753 = w8435 ^ w8564 ;
  assign w8754 = w8437 ^ w8753 ;
  assign w8755 = w1711 & ~w7673 ;
  assign w8756 = ~w1834 & w7411 ;
  assign w8757 = ( w1711 & ~w8755 ) | ( w1711 & w8756 ) | ( ~w8755 & w8756 ) ;
  assign w8758 = w1614 & ~w7944 ;
  assign w8759 = w5433 & ~w8757 ;
  assign w8760 = ( w7414 & w8757 ) | ( w7414 & ~w8759 ) | ( w8757 & ~w8759 ) ;
  assign w8761 = ( w1614 & ~w8758 ) | ( w1614 & w8760 ) | ( ~w8758 & w8760 ) ;
  assign w8762 = \pi08 ^ w8761 ;
  assign w8763 = w8445 ^ w8563 ;
  assign w8764 = w8447 ^ w8763 ;
  assign w8765 = w1939 | w7411 ;
  assign w8766 = ~w1834 & w7673 ;
  assign w8767 = ( ~w1939 & w8765 ) | ( ~w1939 & w8766 ) | ( w8765 & w8766 ) ;
  assign w8768 = w1711 & ~w7944 ;
  assign w8769 = w5296 | w8767 ;
  assign w8770 = ( w7414 & w8767 ) | ( w7414 & w8769 ) | ( w8767 & w8769 ) ;
  assign w8771 = ( w1711 & ~w8768 ) | ( w1711 & w8770 ) | ( ~w8768 & w8770 ) ;
  assign w8772 = \pi08 ^ w8771 ;
  assign w8773 = w8455 ^ w8562 ;
  assign w8774 = w8457 ^ w8773 ;
  assign w8775 = w1939 | w7673 ;
  assign w8776 = w1976 & w7411 ;
  assign w8777 = ( ~w1939 & w8775 ) | ( ~w1939 & w8776 ) | ( w8775 & w8776 ) ;
  assign w8778 = w1834 | w7944 ;
  assign w8779 = w5659 & ~w8777 ;
  assign w8780 = ( w7414 & w8777 ) | ( w7414 & ~w8779 ) | ( w8777 & ~w8779 ) ;
  assign w8781 = ( ~w1834 & w8778 ) | ( ~w1834 & w8780 ) | ( w8778 & w8780 ) ;
  assign w8782 = \pi08 ^ w8781 ;
  assign w8783 = w2059 | w7411 ;
  assign w8784 = w1976 & w7673 ;
  assign w8785 = ( ~w2059 & w8783 ) | ( ~w2059 & w8784 ) | ( w8783 & w8784 ) ;
  assign w8786 = w1939 | w7944 ;
  assign w8787 = w5748 | w8785 ;
  assign w8788 = ( w7414 & w8785 ) | ( w7414 & w8787 ) | ( w8785 & w8787 ) ;
  assign w8789 = ( ~w1939 & w8786 ) | ( ~w1939 & w8788 ) | ( w8786 & w8788 ) ;
  assign w8790 = \pi08 ^ w8789 ;
  assign w8791 = w8459 ^ w8561 ;
  assign w8792 = w8467 ^ w8791 ;
  assign w8793 = w2059 | w7673 ;
  assign w8794 = ~w2130 & w7411 ;
  assign w8795 = ( ~w2059 & w8793 ) | ( ~w2059 & w8794 ) | ( w8793 & w8794 ) ;
  assign w8796 = w1976 & ~w7944 ;
  assign w8797 = w5646 | w8795 ;
  assign w8798 = ( w7414 & w8795 ) | ( w7414 & w8797 ) | ( w8795 & w8797 ) ;
  assign w8799 = ( w1976 & ~w8796 ) | ( w1976 & w8798 ) | ( ~w8796 & w8798 ) ;
  assign w8800 = \pi08 ^ w8799 ;
  assign w8801 = w8469 ^ w8560 ;
  assign w8802 = w8477 ^ w8801 ;
  assign w8803 = w2130 | w7673 ;
  assign w8804 = ~w2235 & w7411 ;
  assign w8805 = ( ~w2130 & w8803 ) | ( ~w2130 & w8804 ) | ( w8803 & w8804 ) ;
  assign w8806 = w2059 | w7944 ;
  assign w8807 = w5896 & ~w8805 ;
  assign w8808 = ( w7414 & w8805 ) | ( w7414 & ~w8807 ) | ( w8805 & ~w8807 ) ;
  assign w8809 = ( ~w2059 & w8806 ) | ( ~w2059 & w8808 ) | ( w8806 & w8808 ) ;
  assign w8810 = \pi08 ^ w8809 ;
  assign w8811 = w8479 ^ w8559 ;
  assign w8812 = w8487 ^ w8811 ;
  assign w8813 = w8495 ^ w8558 ;
  assign w8814 = w8497 ^ w8813 ;
  assign w8815 = w2273 & ~w7411 ;
  assign w8816 = ~w2235 & w7673 ;
  assign w8817 = ( w2273 & ~w8815 ) | ( w2273 & w8816 ) | ( ~w8815 & w8816 ) ;
  assign w8818 = w2130 | w7944 ;
  assign w8819 = w6094 | w8817 ;
  assign w8820 = ( w7414 & w8817 ) | ( w7414 & w8819 ) | ( w8817 & w8819 ) ;
  assign w8821 = ( ~w2130 & w8818 ) | ( ~w2130 & w8820 ) | ( w8818 & w8820 ) ;
  assign w8822 = \pi08 ^ w8821 ;
  assign w8823 = w8499 ^ w8557 ;
  assign w8824 = w8507 ^ w8823 ;
  assign w8825 = w2273 & ~w7673 ;
  assign w8826 = w2391 & w7411 ;
  assign w8827 = ( w2273 & ~w8825 ) | ( w2273 & w8826 ) | ( ~w8825 & w8826 ) ;
  assign w8828 = w2235 | w7944 ;
  assign w8829 = w6106 & ~w8827 ;
  assign w8830 = ( w7414 & w8827 ) | ( w7414 & ~w8829 ) | ( w8827 & ~w8829 ) ;
  assign w8831 = ( ~w2235 & w8828 ) | ( ~w2235 & w8830 ) | ( w8828 & w8830 ) ;
  assign w8832 = \pi08 ^ w8831 ;
  assign w8833 = w8515 ^ w8556 ;
  assign w8834 = w8516 ^ w8833 ;
  assign w8835 = w2391 & ~w7673 ;
  assign w8836 = w2500 & w7411 ;
  assign w8837 = ( w2391 & ~w8835 ) | ( w2391 & w8836 ) | ( ~w8835 & w8836 ) ;
  assign w8838 = w2273 & ~w7944 ;
  assign w8839 = w5880 | w8837 ;
  assign w8840 = ( w7414 & w8837 ) | ( w7414 & w8839 ) | ( w8837 & w8839 ) ;
  assign w8841 = ( w2273 & ~w8838 ) | ( w2273 & w8840 ) | ( ~w8838 & w8840 ) ;
  assign w8842 = \pi08 ^ w8841 ;
  assign w8843 = w2578 | w7411 ;
  assign w8844 = w2500 & w7673 ;
  assign w8845 = ( ~w2578 & w8843 ) | ( ~w2578 & w8844 ) | ( w8843 & w8844 ) ;
  assign w8846 = w2391 & ~w7944 ;
  assign w8847 = w6164 & ~w8845 ;
  assign w8848 = ( w7414 & w8845 ) | ( w7414 & ~w8847 ) | ( w8845 & ~w8847 ) ;
  assign w8849 = ( w2391 & ~w8846 ) | ( w2391 & w8848 ) | ( ~w8846 & w8848 ) ;
  assign w8850 = \pi08 ^ w8849 ;
  assign w8851 = w8529 ^ w8555 ;
  assign w8852 = w8521 ^ w8851 ;
  assign w8853 = w8545 ^ w8553 ;
  assign w8854 = w8554 ^ w8853 ;
  assign w8855 = w2578 | w7673 ;
  assign w8856 = ~w2653 & w7411 ;
  assign w8857 = ( ~w2578 & w8855 ) | ( ~w2578 & w8856 ) | ( w8855 & w8856 ) ;
  assign w8858 = w2500 & ~w7944 ;
  assign w8859 = w6219 | w8857 ;
  assign w8860 = ( w7414 & w8857 ) | ( w7414 & w8859 ) | ( w8857 & w8859 ) ;
  assign w8861 = ( w2500 & ~w8858 ) | ( w2500 & w8860 ) | ( ~w8858 & w8860 ) ;
  assign w8862 = \pi08 ^ w8861 ;
  assign w8863 = w2694 | w7411 ;
  assign w8864 = ~w2653 & w7673 ;
  assign w8865 = ( ~w2694 & w8863 ) | ( ~w2694 & w8864 ) | ( w8863 & w8864 ) ;
  assign w8866 = w2578 | w7944 ;
  assign w8867 = w6282 & ~w8865 ;
  assign w8868 = ( w7414 & w8865 ) | ( w7414 & ~w8867 ) | ( w8865 & ~w8867 ) ;
  assign w8869 = ( ~w2578 & w8866 ) | ( ~w2578 & w8868 ) | ( w8866 & w8868 ) ;
  assign w8870 = \pi08 ^ w8869 ;
  assign w8871 = w8536 ^ w8544 ;
  assign w8872 = ( \pi08 & \pi09 ) | ( \pi08 & ~w2871 ) | ( \pi09 & ~w2871 ) ;
  assign w8873 = \pi08 & \pi09 ;
  assign w8874 = w2973 ^ w8873 ;
  assign w8875 = ( \pi10 & w8873 ) | ( \pi10 & ~w8874 ) | ( w8873 & ~w8874 ) ;
  assign w8876 = w8872 ^ w8875 ;
  assign w8877 = w2805 & ~w7411 ;
  assign w8878 = ~w2694 & w7673 ;
  assign w8879 = ( w2805 & ~w8877 ) | ( w2805 & w8878 ) | ( ~w8877 & w8878 ) ;
  assign w8880 = w2653 | w7944 ;
  assign w8881 = w6338 & ~w8879 ;
  assign w8882 = ( w7414 & w8879 ) | ( w7414 & ~w8881 ) | ( w8879 & ~w8881 ) ;
  assign w8883 = ( ~w2653 & w8880 ) | ( ~w2653 & w8882 ) | ( w8880 & w8882 ) ;
  assign w8884 = \pi08 ^ w8883 ;
  assign w8885 = ( \pi05 & \pi06 ) | ( \pi05 & ~\pi08 ) | ( \pi06 & ~\pi08 ) ;
  assign w8886 = \pi08 & w2973 ;
  assign w8887 = w2871 & w8886 ;
  assign w8888 = ( \pi05 & \pi06 ) | ( \pi05 & ~w8887 ) | ( \pi06 & ~w8887 ) ;
  assign w8889 = ( \pi07 & \pi08 ) | ( \pi07 & ~w8888 ) | ( \pi08 & ~w8888 ) ;
  assign w8890 = ( \pi07 & ~w8886 ) | ( \pi07 & w8888 ) | ( ~w8886 & w8888 ) ;
  assign w8891 = ( w8885 & w8889 ) | ( w8885 & ~w8890 ) | ( w8889 & ~w8890 ) ;
  assign w8892 = w2973 | w7411 ;
  assign w8893 = ~w2871 & w7673 ;
  assign w8894 = ( ~w2973 & w8892 ) | ( ~w2973 & w8893 ) | ( w8892 & w8893 ) ;
  assign w8895 = w2805 & ~w7944 ;
  assign w8896 = w6457 | w8894 ;
  assign w8897 = ( w7414 & w8894 ) | ( w7414 & w8896 ) | ( w8894 & w8896 ) ;
  assign w8898 = ( w2805 & ~w8895 ) | ( w2805 & w8897 ) | ( ~w8895 & w8897 ) ;
  assign w8899 = \pi08 ^ w8898 ;
  assign w8900 = w8891 & w8899 ;
  assign w8901 = w2805 & ~w7673 ;
  assign w8902 = ~w2871 & w7411 ;
  assign w8903 = ( w2805 & ~w8901 ) | ( w2805 & w8902 ) | ( ~w8901 & w8902 ) ;
  assign w8904 = w2694 | w7944 ;
  assign w8905 = w6473 | w8903 ;
  assign w8906 = ( w7414 & w8903 ) | ( w7414 & w8905 ) | ( w8903 & w8905 ) ;
  assign w8907 = ( ~w2694 & w8904 ) | ( ~w2694 & w8906 ) | ( w8904 & w8906 ) ;
  assign w8908 = \pi08 ^ w8907 ;
  assign w8909 = ~w2973 & w6750 ;
  assign w8910 = ( w8900 & w8908 ) | ( w8900 & w8909 ) | ( w8908 & w8909 ) ;
  assign w8911 = ( w8876 & w8884 ) | ( w8876 & w8910 ) | ( w8884 & w8910 ) ;
  assign w8912 = ( w8870 & w8871 ) | ( w8870 & w8911 ) | ( w8871 & w8911 ) ;
  assign w8913 = ( w8854 & w8862 ) | ( w8854 & w8912 ) | ( w8862 & w8912 ) ;
  assign w8914 = ( w8850 & w8852 ) | ( w8850 & w8913 ) | ( w8852 & w8913 ) ;
  assign w8915 = ( w8834 & w8842 ) | ( w8834 & w8914 ) | ( w8842 & w8914 ) ;
  assign w8916 = ( w8824 & w8832 ) | ( w8824 & w8915 ) | ( w8832 & w8915 ) ;
  assign w8917 = ( w8814 & w8822 ) | ( w8814 & w8916 ) | ( w8822 & w8916 ) ;
  assign w8918 = ( w8810 & w8812 ) | ( w8810 & w8917 ) | ( w8812 & w8917 ) ;
  assign w8919 = ( w8800 & w8802 ) | ( w8800 & w8918 ) | ( w8802 & w8918 ) ;
  assign w8920 = ( w8790 & w8792 ) | ( w8790 & w8919 ) | ( w8792 & w8919 ) ;
  assign w8921 = ( w8774 & w8782 ) | ( w8774 & w8920 ) | ( w8782 & w8920 ) ;
  assign w8922 = ( w8764 & w8772 ) | ( w8764 & w8921 ) | ( w8772 & w8921 ) ;
  assign w8923 = ( w8754 & w8762 ) | ( w8754 & w8922 ) | ( w8762 & w8922 ) ;
  assign w8924 = ( w8750 & w8752 ) | ( w8750 & w8923 ) | ( w8752 & w8923 ) ;
  assign w8925 = ( w8740 & w8742 ) | ( w8740 & w8924 ) | ( w8742 & w8924 ) ;
  assign w8926 = ( w8730 & w8732 ) | ( w8730 & w8925 ) | ( w8732 & w8925 ) ;
  assign w8927 = ( w8714 & w8722 ) | ( w8714 & w8926 ) | ( w8722 & w8926 ) ;
  assign w8928 = ( w8704 & w8712 ) | ( w8704 & w8927 ) | ( w8712 & w8927 ) ;
  assign w8929 = ( w8694 & w8702 ) | ( w8694 & w8928 ) | ( w8702 & w8928 ) ;
  assign w8930 = ( w8690 & w8692 ) | ( w8690 & w8929 ) | ( w8692 & w8929 ) ;
  assign w8931 = ( w8680 & w8682 ) | ( w8680 & w8930 ) | ( w8682 & w8930 ) ;
  assign w8932 = ( w8664 & w8672 ) | ( w8664 & w8931 ) | ( w8672 & w8931 ) ;
  assign w8933 = ( ~w8654 & w8662 ) | ( ~w8654 & w8932 ) | ( w8662 & w8932 ) ;
  assign w8934 = ( ~w8644 & w8652 ) | ( ~w8644 & w8933 ) | ( w8652 & w8933 ) ;
  assign w8935 = ( w8634 & w8642 ) | ( w8634 & w8934 ) | ( w8642 & w8934 ) ;
  assign w8936 = ( ~w8624 & w8632 ) | ( ~w8624 & w8935 ) | ( w8632 & w8935 ) ;
  assign w8937 = ( w8614 & w8622 ) | ( w8614 & w8936 ) | ( w8622 & w8936 ) ;
  assign w8938 = ( w8604 & w8612 ) | ( w8604 & w8937 ) | ( w8612 & w8937 ) ;
  assign w8939 = w8580 ^ w8590 ;
  assign w8940 = w8582 ^ w8939 ;
  assign w8941 = w3962 | w8593 ;
  assign w8942 = ~w4142 & w8262 ;
  assign w8943 = ( ~w3962 & w8941 ) | ( ~w3962 & w8942 ) | ( w8941 & w8942 ) ;
  assign w8944 = w4722 | w8263 ;
  assign w8945 = w4600 & ~w8943 ;
  assign w8946 = ( w35 & w8943 ) | ( w35 & ~w8945 ) | ( w8943 & ~w8945 ) ;
  assign w8947 = ( ~w4722 & w8944 ) | ( ~w4722 & w8946 ) | ( w8944 & w8946 ) ;
  assign w8948 = \pi05 ^ w8947 ;
  assign w8949 = ( w8938 & w8940 ) | ( w8938 & w8948 ) | ( w8940 & w8948 ) ;
  assign w8950 = \pi05 ^ w8591 ;
  assign w8951 = w8598 ^ w8950 ;
  assign w8952 = w8600 ^ w8951 ;
  assign w8953 = \pi01 ^ \pi02 ;
  assign w8954 = \pi00 & w8953 ;
  assign w8955 = \pi02 & w4603 ;
  assign w8956 = ( \pi00 & \pi02 ) | ( \pi00 & ~w4603 ) | ( \pi02 & ~w4603 ) ;
  assign w8957 = \pi00 | w4600 ;
  assign w8958 = ( ~\pi00 & \pi01 ) | ( ~\pi00 & w8957 ) | ( \pi01 & w8957 ) ;
  assign w8959 = ( w8955 & w8956 ) | ( w8955 & w8958 ) | ( w8956 & w8958 ) ;
  assign w8960 = w4049 | w8262 ;
  assign w8961 = ~w4142 & w8593 ;
  assign w8962 = ( ~w4049 & w8960 ) | ( ~w4049 & w8961 ) | ( w8960 & w8961 ) ;
  assign w8963 = w4152 | w8263 ;
  assign w8964 = w3962 & ~w8962 ;
  assign w8965 = ( w35 & w8962 ) | ( w35 & ~w8964 ) | ( w8962 & ~w8964 ) ;
  assign w8966 = ( ~w4152 & w8963 ) | ( ~w4152 & w8965 ) | ( w8963 & w8965 ) ;
  assign w8967 = \pi05 ^ w8966 ;
  assign w8968 = w8604 ^ w8937 ;
  assign w8969 = w8612 ^ w8968 ;
  assign w8970 = ( w8959 & w8967 ) | ( w8959 & w8969 ) | ( w8967 & w8969 ) ;
  assign w8971 = w8938 ^ w8948 ;
  assign w8972 = w8940 ^ w8971 ;
  assign w8973 = w8959 ^ w8967 ;
  assign w8974 = w8969 ^ w8973 ;
  assign w8975 = w4049 | w8593 ;
  assign w8976 = w3907 & w8262 ;
  assign w8977 = ( ~w4049 & w8975 ) | ( ~w4049 & w8976 ) | ( w8975 & w8976 ) ;
  assign w8978 = w4563 & ~w8263 ;
  assign w8979 = w4142 & ~w8977 ;
  assign w8980 = ( w35 & w8977 ) | ( w35 & ~w8979 ) | ( w8977 & ~w8979 ) ;
  assign w8981 = ( w4563 & ~w8978 ) | ( w4563 & w8980 ) | ( ~w8978 & w8980 ) ;
  assign w8982 = \pi05 ^ w8981 ;
  assign w8983 = w8614 ^ w8936 ;
  assign w8984 = w8622 ^ w8983 ;
  assign w8985 = w3548 | w8262 ;
  assign w8986 = w3907 & w8593 ;
  assign w8987 = ( ~w3548 & w8985 ) | ( ~w3548 & w8986 ) | ( w8985 & w8986 ) ;
  assign w8988 = w4622 | w8263 ;
  assign w8989 = w4049 & ~w8987 ;
  assign w8990 = ( w35 & w8987 ) | ( w35 & ~w8989 ) | ( w8987 & ~w8989 ) ;
  assign w8991 = ( ~w4622 & w8988 ) | ( ~w4622 & w8990 ) | ( w8988 & w8990 ) ;
  assign w8992 = \pi05 ^ w8991 ;
  assign w8993 = w8624 ^ w8935 ;
  assign w8994 = w8632 ^ w8993 ;
  assign w8995 = w3548 | w8593 ;
  assign w8996 = w3715 & w8262 ;
  assign w8997 = ( ~w3548 & w8995 ) | ( ~w3548 & w8996 ) | ( w8995 & w8996 ) ;
  assign w8998 = w3913 | w8263 ;
  assign w8999 = w3907 | w8997 ;
  assign w9000 = ( w35 & w8997 ) | ( w35 & w8999 ) | ( w8997 & w8999 ) ;
  assign w9001 = ( ~w3913 & w8998 ) | ( ~w3913 & w9000 ) | ( w8998 & w9000 ) ;
  assign w9002 = \pi05 ^ w9001 ;
  assign w9003 = w8634 ^ w8934 ;
  assign w9004 = w8642 ^ w9003 ;
  assign w9005 = w3647 & ~w8262 ;
  assign w9006 = w3715 & w8593 ;
  assign w9007 = ( w3647 & ~w9005 ) | ( w3647 & w9006 ) | ( ~w9005 & w9006 ) ;
  assign w9008 = w3725 | w8263 ;
  assign w9009 = w3548 & ~w9007 ;
  assign w9010 = ( w35 & w9007 ) | ( w35 & ~w9009 ) | ( w9007 & ~w9009 ) ;
  assign w9011 = ( ~w3725 & w9008 ) | ( ~w3725 & w9010 ) | ( w9008 & w9010 ) ;
  assign w9012 = \pi05 ^ w9011 ;
  assign w9013 = w8644 ^ w8933 ;
  assign w9014 = w8652 ^ w9013 ;
  assign w9015 = w3647 & ~w8593 ;
  assign w9016 = ~w3094 & w8262 ;
  assign w9017 = ( w3647 & ~w9015 ) | ( w3647 & w9016 ) | ( ~w9015 & w9016 ) ;
  assign w9018 = w4164 | w8263 ;
  assign w9019 = w3715 | w9017 ;
  assign w9020 = ( w35 & w9017 ) | ( w35 & w9019 ) | ( w9017 & w9019 ) ;
  assign w9021 = ( ~w4164 & w9018 ) | ( ~w4164 & w9020 ) | ( w9018 & w9020 ) ;
  assign w9022 = \pi05 ^ w9021 ;
  assign w9023 = w8654 ^ w8932 ;
  assign w9024 = w8662 ^ w9023 ;
  assign w9025 = w381 | w8262 ;
  assign w9026 = ~w3094 & w8593 ;
  assign w9027 = ( ~w381 & w9025 ) | ( ~w381 & w9026 ) | ( w9025 & w9026 ) ;
  assign w9028 = w3810 & ~w8263 ;
  assign w9029 = w3647 | w9027 ;
  assign w9030 = ( w35 & w9027 ) | ( w35 & w9029 ) | ( w9027 & w9029 ) ;
  assign w9031 = ( w3810 & ~w9028 ) | ( w3810 & w9030 ) | ( ~w9028 & w9030 ) ;
  assign w9032 = \pi05 ^ w9031 ;
  assign w9033 = w8664 ^ w8931 ;
  assign w9034 = w8672 ^ w9033 ;
  assign w9035 = w8680 ^ w8930 ;
  assign w9036 = w8682 ^ w9035 ;
  assign w9037 = w381 | w8593 ;
  assign w9038 = w592 & w8262 ;
  assign w9039 = ( ~w381 & w9037 ) | ( ~w381 & w9038 ) | ( w9037 & w9038 ) ;
  assign w9040 = w3096 & ~w8263 ;
  assign w9041 = w3094 & ~w9039 ;
  assign w9042 = ( w35 & w9039 ) | ( w35 & ~w9041 ) | ( w9039 & ~w9041 ) ;
  assign w9043 = ( w3096 & ~w9040 ) | ( w3096 & w9042 ) | ( ~w9040 & w9042 ) ;
  assign w9044 = \pi05 ^ w9043 ;
  assign w9045 = w8690 ^ w8929 ;
  assign w9046 = w8692 ^ w9045 ;
  assign w9047 = w592 & ~w8593 ;
  assign w9048 = w721 & w8262 ;
  assign w9049 = ( w592 & ~w9047 ) | ( w592 & w9048 ) | ( ~w9047 & w9048 ) ;
  assign w9050 = w3435 | w8263 ;
  assign w9051 = w381 & ~w9049 ;
  assign w9052 = ( w35 & w9049 ) | ( w35 & ~w9051 ) | ( w9049 & ~w9051 ) ;
  assign w9053 = ( ~w3435 & w9050 ) | ( ~w3435 & w9052 ) | ( w9050 & w9052 ) ;
  assign w9054 = \pi05 ^ w9053 ;
  assign w9055 = w883 | w8262 ;
  assign w9056 = w721 & w8593 ;
  assign w9057 = ( ~w883 & w9055 ) | ( ~w883 & w9056 ) | ( w9055 & w9056 ) ;
  assign w9058 = w3421 & ~w8263 ;
  assign w9059 = w592 | w9057 ;
  assign w9060 = ( w35 & w9057 ) | ( w35 & w9059 ) | ( w9057 & w9059 ) ;
  assign w9061 = ( w3421 & ~w9058 ) | ( w3421 & w9060 ) | ( ~w9058 & w9060 ) ;
  assign w9062 = \pi05 ^ w9061 ;
  assign w9063 = w8694 ^ w8928 ;
  assign w9064 = w8702 ^ w9063 ;
  assign w9065 = w883 | w8593 ;
  assign w9066 = w979 & w8262 ;
  assign w9067 = ( ~w883 & w9065 ) | ( ~w883 & w9066 ) | ( w9065 & w9066 ) ;
  assign w9068 = w4257 | w8263 ;
  assign w9069 = w721 | w9067 ;
  assign w9070 = ( w35 & w9067 ) | ( w35 & w9069 ) | ( w9067 & w9069 ) ;
  assign w9071 = ( ~w4257 & w9068 ) | ( ~w4257 & w9070 ) | ( w9068 & w9070 ) ;
  assign w9072 = \pi05 ^ w9071 ;
  assign w9073 = w8704 ^ w8927 ;
  assign w9074 = w8712 ^ w9073 ;
  assign w9075 = w979 & ~w8593 ;
  assign w9076 = w1085 & w8262 ;
  assign w9077 = ( w979 & ~w9075 ) | ( w979 & w9076 ) | ( ~w9075 & w9076 ) ;
  assign w9078 = w4273 | w8263 ;
  assign w9079 = w883 & ~w9077 ;
  assign w9080 = ( w35 & w9077 ) | ( w35 & ~w9079 ) | ( w9077 & ~w9079 ) ;
  assign w9081 = ( ~w4273 & w9078 ) | ( ~w4273 & w9080 ) | ( w9078 & w9080 ) ;
  assign w9082 = \pi05 ^ w9081 ;
  assign w9083 = w8714 ^ w8926 ;
  assign w9084 = w8722 ^ w9083 ;
  assign w9085 = w8730 ^ w8925 ;
  assign w9086 = w8732 ^ w9085 ;
  assign w9087 = w1085 & ~w8593 ;
  assign w9088 = w1205 & w8262 ;
  assign w9089 = ( w1085 & ~w9087 ) | ( w1085 & w9088 ) | ( ~w9087 & w9088 ) ;
  assign w9090 = w4666 & ~w8263 ;
  assign w9091 = w979 | w9089 ;
  assign w9092 = ( w35 & w9089 ) | ( w35 & w9091 ) | ( w9089 & w9091 ) ;
  assign w9093 = ( w4666 & ~w9090 ) | ( w4666 & w9092 ) | ( ~w9090 & w9092 ) ;
  assign w9094 = \pi05 ^ w9093 ;
  assign w9095 = w8740 ^ w8924 ;
  assign w9096 = w8742 ^ w9095 ;
  assign w9097 = w1264 | w8262 ;
  assign w9098 = w1205 & w8593 ;
  assign w9099 = ( ~w1264 & w9097 ) | ( ~w1264 & w9098 ) | ( w9097 & w9098 ) ;
  assign w9100 = w4533 & ~w8263 ;
  assign w9101 = w1085 | w9099 ;
  assign w9102 = ( w35 & w9099 ) | ( w35 & w9101 ) | ( w9099 & w9101 ) ;
  assign w9103 = ( w4533 & ~w9100 ) | ( w4533 & w9102 ) | ( ~w9100 & w9102 ) ;
  assign w9104 = \pi05 ^ w9103 ;
  assign w9105 = w8750 ^ w8923 ;
  assign w9106 = w8752 ^ w9105 ;
  assign w9107 = w1264 | w8593 ;
  assign w9108 = w1399 & w8262 ;
  assign w9109 = ( ~w1264 & w9107 ) | ( ~w1264 & w9108 ) | ( w9107 & w9108 ) ;
  assign w9110 = w4864 | w8263 ;
  assign w9111 = w1205 | w9109 ;
  assign w9112 = ( w35 & w9109 ) | ( w35 & w9111 ) | ( w9109 & w9111 ) ;
  assign w9113 = ( ~w4864 & w9110 ) | ( ~w4864 & w9112 ) | ( w9110 & w9112 ) ;
  assign w9114 = \pi05 ^ w9113 ;
  assign w9115 = w1399 & ~w8593 ;
  assign w9116 = ~w1510 & w8262 ;
  assign w9117 = ( w1399 & ~w9115 ) | ( w1399 & w9116 ) | ( ~w9115 & w9116 ) ;
  assign w9118 = w4852 | w8263 ;
  assign w9119 = w1264 & ~w9117 ;
  assign w9120 = ( w35 & w9117 ) | ( w35 & ~w9119 ) | ( w9117 & ~w9119 ) ;
  assign w9121 = ( ~w4852 & w9118 ) | ( ~w4852 & w9120 ) | ( w9118 & w9120 ) ;
  assign w9122 = \pi05 ^ w9121 ;
  assign w9123 = w8754 ^ w8922 ;
  assign w9124 = w8762 ^ w9123 ;
  assign w9125 = w1614 & ~w8262 ;
  assign w9126 = ~w1510 & w8593 ;
  assign w9127 = ( w1614 & ~w9125 ) | ( w1614 & w9126 ) | ( ~w9125 & w9126 ) ;
  assign w9128 = w5069 | w8263 ;
  assign w9129 = w1399 | w9127 ;
  assign w9130 = ( w35 & w9127 ) | ( w35 & w9129 ) | ( w9127 & w9129 ) ;
  assign w9131 = ( ~w5069 & w9128 ) | ( ~w5069 & w9130 ) | ( w9128 & w9130 ) ;
  assign w9132 = \pi05 ^ w9131 ;
  assign w9133 = w8764 ^ w8921 ;
  assign w9134 = w8772 ^ w9133 ;
  assign w9135 = w1614 & ~w8593 ;
  assign w9136 = w1711 & w8262 ;
  assign w9137 = ( w1614 & ~w9135 ) | ( w1614 & w9136 ) | ( ~w9135 & w9136 ) ;
  assign w9138 = w5085 | w8263 ;
  assign w9139 = w1510 & ~w9137 ;
  assign w9140 = ( w35 & w9137 ) | ( w35 & ~w9139 ) | ( w9137 & ~w9139 ) ;
  assign w9141 = ( ~w5085 & w9138 ) | ( ~w5085 & w9140 ) | ( w9138 & w9140 ) ;
  assign w9142 = \pi05 ^ w9141 ;
  assign w9143 = w8774 ^ w8920 ;
  assign w9144 = w8782 ^ w9143 ;
  assign w9145 = w8790 ^ w8919 ;
  assign w9146 = w8792 ^ w9145 ;
  assign w9147 = w1711 & ~w8593 ;
  assign w9148 = ~w1834 & w8262 ;
  assign w9149 = ( w1711 & ~w9147 ) | ( w1711 & w9148 ) | ( ~w9147 & w9148 ) ;
  assign w9150 = w5433 | w8263 ;
  assign w9151 = w1614 | w9149 ;
  assign w9152 = ( w35 & w9149 ) | ( w35 & w9151 ) | ( w9149 & w9151 ) ;
  assign w9153 = ( ~w5433 & w9150 ) | ( ~w5433 & w9152 ) | ( w9150 & w9152 ) ;
  assign w9154 = \pi05 ^ w9153 ;
  assign w9155 = w8800 ^ w8918 ;
  assign w9156 = w8802 ^ w9155 ;
  assign w9157 = w1939 | w8262 ;
  assign w9158 = ~w1834 & w8593 ;
  assign w9159 = ( ~w1939 & w9157 ) | ( ~w1939 & w9158 ) | ( w9157 & w9158 ) ;
  assign w9160 = w5296 & ~w8263 ;
  assign w9161 = w1711 | w9159 ;
  assign w9162 = ( w35 & w9159 ) | ( w35 & w9161 ) | ( w9159 & w9161 ) ;
  assign w9163 = ( w5296 & ~w9160 ) | ( w5296 & w9162 ) | ( ~w9160 & w9162 ) ;
  assign w9164 = \pi05 ^ w9163 ;
  assign w9165 = w8810 ^ w8917 ;
  assign w9166 = w8812 ^ w9165 ;
  assign w9167 = w1939 | w8593 ;
  assign w9168 = w1976 & w8262 ;
  assign w9169 = ( ~w1939 & w9167 ) | ( ~w1939 & w9168 ) | ( w9167 & w9168 ) ;
  assign w9170 = w5659 | w8263 ;
  assign w9171 = w1834 & ~w9169 ;
  assign w9172 = ( w35 & w9169 ) | ( w35 & ~w9171 ) | ( w9169 & ~w9171 ) ;
  assign w9173 = ( ~w5659 & w9170 ) | ( ~w5659 & w9172 ) | ( w9170 & w9172 ) ;
  assign w9174 = \pi05 ^ w9173 ;
  assign w9175 = w2059 | w8262 ;
  assign w9176 = w1976 & w8593 ;
  assign w9177 = ( ~w2059 & w9175 ) | ( ~w2059 & w9176 ) | ( w9175 & w9176 ) ;
  assign w9178 = w5748 & ~w8263 ;
  assign w9179 = w1939 & ~w9177 ;
  assign w9180 = ( w35 & w9177 ) | ( w35 & ~w9179 ) | ( w9177 & ~w9179 ) ;
  assign w9181 = ( w5748 & ~w9178 ) | ( w5748 & w9180 ) | ( ~w9178 & w9180 ) ;
  assign w9182 = \pi05 ^ w9181 ;
  assign w9183 = w8814 ^ w8916 ;
  assign w9184 = w8822 ^ w9183 ;
  assign w9185 = w2059 | w8593 ;
  assign w9186 = ~w2130 & w8262 ;
  assign w9187 = ( ~w2059 & w9185 ) | ( ~w2059 & w9186 ) | ( w9185 & w9186 ) ;
  assign w9188 = w5646 & ~w8263 ;
  assign w9189 = w1976 | w9187 ;
  assign w9190 = ( w35 & w9187 ) | ( w35 & w9189 ) | ( w9187 & w9189 ) ;
  assign w9191 = ( w5646 & ~w9188 ) | ( w5646 & w9190 ) | ( ~w9188 & w9190 ) ;
  assign w9192 = \pi05 ^ w9191 ;
  assign w9193 = w8824 ^ w8915 ;
  assign w9194 = w8832 ^ w9193 ;
  assign w9195 = w2130 | w8593 ;
  assign w9196 = ~w2235 & w8262 ;
  assign w9197 = ( ~w2130 & w9195 ) | ( ~w2130 & w9196 ) | ( w9195 & w9196 ) ;
  assign w9198 = w5896 | w8263 ;
  assign w9199 = w2059 & ~w9197 ;
  assign w9200 = ( w35 & w9197 ) | ( w35 & ~w9199 ) | ( w9197 & ~w9199 ) ;
  assign w9201 = ( ~w5896 & w9198 ) | ( ~w5896 & w9200 ) | ( w9198 & w9200 ) ;
  assign w9202 = \pi05 ^ w9201 ;
  assign w9203 = w8834 ^ w8914 ;
  assign w9204 = w8842 ^ w9203 ;
  assign w9205 = w8850 ^ w8913 ;
  assign w9206 = w8852 ^ w9205 ;
  assign w9207 = w2273 & ~w8262 ;
  assign w9208 = ~w2235 & w8593 ;
  assign w9209 = ( w2273 & ~w9207 ) | ( w2273 & w9208 ) | ( ~w9207 & w9208 ) ;
  assign w9210 = w6094 & ~w8263 ;
  assign w9211 = w2130 & ~w9209 ;
  assign w9212 = ( w35 & w9209 ) | ( w35 & ~w9211 ) | ( w9209 & ~w9211 ) ;
  assign w9213 = ( w6094 & ~w9210 ) | ( w6094 & w9212 ) | ( ~w9210 & w9212 ) ;
  assign w9214 = \pi05 ^ w9213 ;
  assign w9215 = w8854 ^ w8912 ;
  assign w9216 = w8862 ^ w9215 ;
  assign w9217 = w2273 & ~w8593 ;
  assign w9218 = w2391 & w8262 ;
  assign w9219 = ( w2273 & ~w9217 ) | ( w2273 & w9218 ) | ( ~w9217 & w9218 ) ;
  assign w9220 = w6106 | w8263 ;
  assign w9221 = w2235 & ~w9219 ;
  assign w9222 = ( w35 & w9219 ) | ( w35 & ~w9221 ) | ( w9219 & ~w9221 ) ;
  assign w9223 = ( ~w6106 & w9220 ) | ( ~w6106 & w9222 ) | ( w9220 & w9222 ) ;
  assign w9224 = \pi05 ^ w9223 ;
  assign w9225 = w8870 ^ w8911 ;
  assign w9226 = w8871 ^ w9225 ;
  assign w9227 = w2391 & ~w8593 ;
  assign w9228 = w2500 & w8262 ;
  assign w9229 = ( w2391 & ~w9227 ) | ( w2391 & w9228 ) | ( ~w9227 & w9228 ) ;
  assign w9230 = w5880 & ~w8263 ;
  assign w9231 = w2273 | w9229 ;
  assign w9232 = ( w35 & w9229 ) | ( w35 & w9231 ) | ( w9229 & w9231 ) ;
  assign w9233 = ( w5880 & ~w9230 ) | ( w5880 & w9232 ) | ( ~w9230 & w9232 ) ;
  assign w9234 = \pi05 ^ w9233 ;
  assign w9235 = w2578 | w8262 ;
  assign w9236 = w2500 & w8593 ;
  assign w9237 = ( ~w2578 & w9235 ) | ( ~w2578 & w9236 ) | ( w9235 & w9236 ) ;
  assign w9238 = w6164 | w8263 ;
  assign w9239 = w2391 | w9237 ;
  assign w9240 = ( w35 & w9237 ) | ( w35 & w9239 ) | ( w9237 & w9239 ) ;
  assign w9241 = ( ~w6164 & w9238 ) | ( ~w6164 & w9240 ) | ( w9238 & w9240 ) ;
  assign w9242 = \pi05 ^ w9241 ;
  assign w9243 = w8884 ^ w8910 ;
  assign w9244 = w8876 ^ w9243 ;
  assign w9245 = w8900 ^ w8908 ;
  assign w9246 = w8909 ^ w9245 ;
  assign w9247 = w2578 | w8593 ;
  assign w9248 = ~w2653 & w8262 ;
  assign w9249 = ( ~w2578 & w9247 ) | ( ~w2578 & w9248 ) | ( w9247 & w9248 ) ;
  assign w9250 = w6219 & ~w8263 ;
  assign w9251 = w2500 | w9249 ;
  assign w9252 = ( w35 & w9249 ) | ( w35 & w9251 ) | ( w9249 & w9251 ) ;
  assign w9253 = ( w6219 & ~w9250 ) | ( w6219 & w9252 ) | ( ~w9250 & w9252 ) ;
  assign w9254 = \pi05 ^ w9253 ;
  assign w9255 = w2694 | w8262 ;
  assign w9256 = ~w2653 & w8593 ;
  assign w9257 = ( ~w2694 & w9255 ) | ( ~w2694 & w9256 ) | ( w9255 & w9256 ) ;
  assign w9258 = w6282 | w8263 ;
  assign w9259 = w2578 & ~w9257 ;
  assign w9260 = ( w35 & w9257 ) | ( w35 & ~w9259 ) | ( w9257 & ~w9259 ) ;
  assign w9261 = ( ~w6282 & w9258 ) | ( ~w6282 & w9260 ) | ( w9258 & w9260 ) ;
  assign w9262 = \pi05 ^ w9261 ;
  assign w9263 = w8891 ^ w8899 ;
  assign w9264 = ( \pi05 & \pi06 ) | ( \pi05 & ~w2871 ) | ( \pi06 & ~w2871 ) ;
  assign w9265 = \pi05 & \pi06 ;
  assign w9266 = w2973 ^ w9265 ;
  assign w9267 = ( \pi07 & w9265 ) | ( \pi07 & ~w9266 ) | ( w9265 & ~w9266 ) ;
  assign w9268 = w9264 ^ w9267 ;
  assign w9269 = w2805 & ~w8262 ;
  assign w9270 = ~w2694 & w8593 ;
  assign w9271 = ( w2805 & ~w9269 ) | ( w2805 & w9270 ) | ( ~w9269 & w9270 ) ;
  assign w9272 = w6338 | w8263 ;
  assign w9273 = w2653 & ~w9271 ;
  assign w9274 = ( w35 & w9271 ) | ( w35 & ~w9273 ) | ( w9271 & ~w9273 ) ;
  assign w9275 = ( ~w6338 & w9272 ) | ( ~w6338 & w9274 ) | ( w9272 & w9274 ) ;
  assign w9276 = \pi05 ^ w9275 ;
  assign w9277 = ( \pi02 & \pi03 ) | ( \pi02 & ~\pi05 ) | ( \pi03 & ~\pi05 ) ;
  assign w9278 = \pi05 & w2973 ;
  assign w9279 = w2871 & w9278 ;
  assign w9280 = ( \pi02 & \pi03 ) | ( \pi02 & ~w9279 ) | ( \pi03 & ~w9279 ) ;
  assign w9281 = ( \pi04 & \pi05 ) | ( \pi04 & ~w9280 ) | ( \pi05 & ~w9280 ) ;
  assign w9282 = ( \pi04 & ~w9278 ) | ( \pi04 & w9280 ) | ( ~w9278 & w9280 ) ;
  assign w9283 = ( w9277 & w9281 ) | ( w9277 & ~w9282 ) | ( w9281 & ~w9282 ) ;
  assign w9284 = w2973 | w8262 ;
  assign w9285 = ~w2871 & w8593 ;
  assign w9286 = ( ~w2973 & w9284 ) | ( ~w2973 & w9285 ) | ( w9284 & w9285 ) ;
  assign w9287 = w6457 & ~w8263 ;
  assign w9288 = w2805 | w9286 ;
  assign w9289 = ( w35 & w9286 ) | ( w35 & w9288 ) | ( w9286 & w9288 ) ;
  assign w9290 = ( w6457 & ~w9287 ) | ( w6457 & w9289 ) | ( ~w9287 & w9289 ) ;
  assign w9291 = \pi05 ^ w9290 ;
  assign w9292 = w9283 & w9291 ;
  assign w9293 = ~w2973 & w7413 ;
  assign w9294 = w9292 ^ w9293 ;
  assign w9295 = w2805 & ~w8593 ;
  assign w9296 = ~w2871 & w8262 ;
  assign w9297 = ( w2805 & ~w9295 ) | ( w2805 & w9296 ) | ( ~w9295 & w9296 ) ;
  assign w9298 = w6473 & ~w8263 ;
  assign w9299 = w2694 & ~w9297 ;
  assign w9300 = ( w35 & w9297 ) | ( w35 & ~w9299 ) | ( w9297 & ~w9299 ) ;
  assign w9301 = ( w6473 & ~w9298 ) | ( w6473 & w9300 ) | ( ~w9298 & w9300 ) ;
  assign w9302 = \pi05 ^ w9301 ;
  assign w9303 = ( w9292 & w9293 ) | ( w9292 & w9302 ) | ( w9293 & w9302 ) ;
  assign w9304 = ( w9268 & w9276 ) | ( w9268 & w9303 ) | ( w9276 & w9303 ) ;
  assign w9305 = ( w9262 & w9263 ) | ( w9262 & w9304 ) | ( w9263 & w9304 ) ;
  assign w9306 = ( w9246 & w9254 ) | ( w9246 & w9305 ) | ( w9254 & w9305 ) ;
  assign w9307 = ( w9242 & w9244 ) | ( w9242 & w9306 ) | ( w9244 & w9306 ) ;
  assign w9308 = ( w9226 & w9234 ) | ( w9226 & w9307 ) | ( w9234 & w9307 ) ;
  assign w9309 = ( w9216 & w9224 ) | ( w9216 & w9308 ) | ( w9224 & w9308 ) ;
  assign w9310 = ( w9206 & w9214 ) | ( w9206 & w9309 ) | ( w9214 & w9309 ) ;
  assign w9311 = ( w9202 & w9204 ) | ( w9202 & w9310 ) | ( w9204 & w9310 ) ;
  assign w9312 = ( w9192 & w9194 ) | ( w9192 & w9311 ) | ( w9194 & w9311 ) ;
  assign w9313 = ( w9182 & w9184 ) | ( w9182 & w9312 ) | ( w9184 & w9312 ) ;
  assign w9314 = ( w9166 & w9174 ) | ( w9166 & w9313 ) | ( w9174 & w9313 ) ;
  assign w9315 = ( w9156 & w9164 ) | ( w9156 & w9314 ) | ( w9164 & w9314 ) ;
  assign w9316 = ( w9146 & w9154 ) | ( w9146 & w9315 ) | ( w9154 & w9315 ) ;
  assign w9317 = ( w9142 & w9144 ) | ( w9142 & w9316 ) | ( w9144 & w9316 ) ;
  assign w9318 = ( w9132 & w9134 ) | ( w9132 & w9317 ) | ( w9134 & w9317 ) ;
  assign w9319 = ( w9122 & w9124 ) | ( w9122 & w9318 ) | ( w9124 & w9318 ) ;
  assign w9320 = ( w9106 & w9114 ) | ( w9106 & w9319 ) | ( w9114 & w9319 ) ;
  assign w9321 = ( w9096 & w9104 ) | ( w9096 & w9320 ) | ( w9104 & w9320 ) ;
  assign w9322 = ( w9086 & w9094 ) | ( w9086 & w9321 ) | ( w9094 & w9321 ) ;
  assign w9323 = ( w9082 & w9084 ) | ( w9082 & w9322 ) | ( w9084 & w9322 ) ;
  assign w9324 = ( w9072 & w9074 ) | ( w9072 & w9323 ) | ( w9074 & w9323 ) ;
  assign w9325 = ( w9062 & w9064 ) | ( w9062 & w9324 ) | ( w9064 & w9324 ) ;
  assign w9326 = ( w9046 & w9054 ) | ( w9046 & w9325 ) | ( w9054 & w9325 ) ;
  assign w9327 = ( w9036 & w9044 ) | ( w9036 & w9326 ) | ( w9044 & w9326 ) ;
  assign w9328 = ( w9032 & w9034 ) | ( w9032 & w9327 ) | ( w9034 & w9327 ) ;
  assign w9329 = ( w9022 & ~w9024 ) | ( w9022 & w9328 ) | ( ~w9024 & w9328 ) ;
  assign w9330 = ( w9012 & ~w9014 ) | ( w9012 & w9329 ) | ( ~w9014 & w9329 ) ;
  assign w9331 = ( w9002 & w9004 ) | ( w9002 & w9330 ) | ( w9004 & w9330 ) ;
  assign w9332 = ( w8992 & ~w8994 ) | ( w8992 & w9331 ) | ( ~w8994 & w9331 ) ;
  assign w9333 = ( w8982 & w8984 ) | ( w8982 & w9332 ) | ( w8984 & w9332 ) ;
  assign w9334 = w8982 ^ w9332 ;
  assign w9335 = w8984 ^ w9334 ;
  assign w9336 = \pi00 & \pi02 ;
  assign w9337 = \pi00 & ~w4602 ;
  assign w9338 = w4600 ^ w9337 ;
  assign w9339 = ~\pi02 & w9338 ;
  assign w9340 = \pi01 & ~w9339 ;
  assign w9341 = ( \pi02 & ~w4600 ) | ( \pi02 & w9336 ) | ( ~w4600 & w9336 ) ;
  assign w9342 = ( w9336 & w9340 ) | ( w9336 & ~w9341 ) | ( w9340 & ~w9341 ) ;
  assign w9343 = ~\pi01 & \pi02 ;
  assign w9344 = \pi00 & ~w6551 ;
  assign w9345 = w3962 ^ w9344 ;
  assign w9346 = w9343 & w9345 ;
  assign w9347 = w9342 | w9346 ;
  assign w9348 = w8992 ^ w9331 ;
  assign w9349 = w8994 ^ w9348 ;
  assign w9350 = ( \pi02 & w3962 ) | ( \pi02 & w4600 ) | ( w3962 & w4600 ) ;
  assign w9351 = \pi00 ^ w9350 ;
  assign w9352 = ( \pi02 & ~w4600 ) | ( \pi02 & w9351 ) | ( ~w4600 & w9351 ) ;
  assign w9353 = ( ~\pi02 & w3962 ) | ( ~\pi02 & w9351 ) | ( w3962 & w9351 ) ;
  assign w9354 = \pi01 & ~w9353 ;
  assign w9355 = ( \pi00 & w4142 ) | ( \pi00 & ~w9354 ) | ( w4142 & ~w9354 ) ;
  assign w9356 = ( \pi01 & \pi02 ) | ( \pi01 & w9355 ) | ( \pi02 & w9355 ) ;
  assign w9357 = ( w9352 & w9354 ) | ( w9352 & ~w9356 ) | ( w9354 & ~w9356 ) ;
  assign w9358 = w9002 ^ w9330 ;
  assign w9359 = w9004 ^ w9358 ;
  assign w9360 = ( \pi02 & w3962 ) | ( \pi02 & w4142 ) | ( w3962 & w4142 ) ;
  assign w9361 = \pi00 ^ w9360 ;
  assign w9362 = ( \pi02 & ~w3962 ) | ( \pi02 & w9361 ) | ( ~w3962 & w9361 ) ;
  assign w9363 = ( ~\pi02 & w4142 ) | ( ~\pi02 & w9361 ) | ( w4142 & w9361 ) ;
  assign w9364 = \pi01 & ~w9363 ;
  assign w9365 = ( \pi00 & w4049 ) | ( \pi00 & ~w9364 ) | ( w4049 & ~w9364 ) ;
  assign w9366 = ( \pi01 & \pi02 ) | ( \pi01 & w9365 ) | ( \pi02 & w9365 ) ;
  assign w9367 = ( w9362 & w9364 ) | ( w9362 & ~w9366 ) | ( w9364 & ~w9366 ) ;
  assign w9368 = w9012 ^ w9329 ;
  assign w9369 = w9014 ^ w9368 ;
  assign w9370 = ( \pi02 & w4049 ) | ( \pi02 & w4142 ) | ( w4049 & w4142 ) ;
  assign w9371 = \pi00 ^ w9370 ;
  assign w9372 = ( \pi02 & ~w4142 ) | ( \pi02 & w9371 ) | ( ~w4142 & w9371 ) ;
  assign w9373 = ( ~\pi02 & w4049 ) | ( ~\pi02 & w9371 ) | ( w4049 & w9371 ) ;
  assign w9374 = \pi01 & ~w9373 ;
  assign w9375 = ( ~\pi00 & w3907 ) | ( ~\pi00 & w9374 ) | ( w3907 & w9374 ) ;
  assign w9376 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9375 ) | ( \pi02 & ~w9375 ) ;
  assign w9377 = ( w9372 & w9374 ) | ( w9372 & ~w9376 ) | ( w9374 & ~w9376 ) ;
  assign w9378 = w9022 ^ w9328 ;
  assign w9379 = w9024 ^ w9378 ;
  assign w9380 = ( \pi02 & ~w3907 ) | ( \pi02 & w4049 ) | ( ~w3907 & w4049 ) ;
  assign w9381 = \pi00 ^ w9380 ;
  assign w9382 = ( \pi02 & ~w4049 ) | ( \pi02 & w9381 ) | ( ~w4049 & w9381 ) ;
  assign w9383 = ( \pi02 & w3907 ) | ( \pi02 & ~w9381 ) | ( w3907 & ~w9381 ) ;
  assign w9384 = \pi01 & w9383 ;
  assign w9385 = ( \pi00 & w3548 ) | ( \pi00 & ~w9384 ) | ( w3548 & ~w9384 ) ;
  assign w9386 = ( \pi01 & \pi02 ) | ( \pi01 & w9385 ) | ( \pi02 & w9385 ) ;
  assign w9387 = ( w9382 & w9384 ) | ( w9382 & ~w9386 ) | ( w9384 & ~w9386 ) ;
  assign w9388 = w9036 ^ w9326 ;
  assign w9389 = w9044 ^ w9388 ;
  assign w9390 = w9086 ^ w9321 ;
  assign w9391 = w9094 ^ w9390 ;
  assign w9392 = w9146 ^ w9315 ;
  assign w9393 = w9154 ^ w9392 ;
  assign w9394 = w9206 ^ w9309 ;
  assign w9395 = w9214 ^ w9394 ;
  assign w9396 = \pi00 ^ w2805 ;
  assign w9397 = ( \pi01 & w2805 ) | ( \pi01 & ~w9396 ) | ( w2805 & ~w9396 ) ;
  assign w9398 = ( \pi00 & ~w2871 ) | ( \pi00 & w9397 ) | ( ~w2871 & w9397 ) ;
  assign w9399 = ( \pi02 & ~w2973 ) | ( \pi02 & w9398 ) | ( ~w2973 & w9398 ) ;
  assign w9400 = \pi02 & ~w9399 ;
  assign w9401 = ( \pi02 & w2694 ) | ( \pi02 & ~w2805 ) | ( w2694 & ~w2805 ) ;
  assign w9402 = \pi00 ^ w9401 ;
  assign w9403 = ( \pi02 & ~w2694 ) | ( \pi02 & w9402 ) | ( ~w2694 & w9402 ) ;
  assign w9404 = ( \pi02 & w2805 ) | ( \pi02 & ~w9402 ) | ( w2805 & ~w9402 ) ;
  assign w9405 = \pi01 & w9404 ;
  assign w9406 = ( \pi00 & w2871 ) | ( \pi00 & ~w9405 ) | ( w2871 & ~w9405 ) ;
  assign w9407 = ( \pi01 & \pi02 ) | ( \pi01 & w9406 ) | ( \pi02 & w9406 ) ;
  assign w9408 = ( w9403 & w9405 ) | ( w9403 & ~w9407 ) | ( w9405 & ~w9407 ) ;
  assign w9409 = ( w6473 & w8954 ) | ( w6473 & w9408 ) | ( w8954 & w9408 ) ;
  assign w9410 = w9408 | w9409 ;
  assign w9411 = \pi02 ^ w9410 ;
  assign w9412 = w34 & ~w2973 ;
  assign w9413 = ( w9400 & w9411 ) | ( w9400 & w9412 ) | ( w9411 & w9412 ) ;
  assign w9414 = ( \pi02 & w2653 ) | ( \pi02 & w2694 ) | ( w2653 & w2694 ) ;
  assign w9415 = \pi00 ^ w9414 ;
  assign w9416 = ( \pi02 & ~w2653 ) | ( \pi02 & w9415 ) | ( ~w2653 & w9415 ) ;
  assign w9417 = ( ~\pi02 & w2694 ) | ( ~\pi02 & w9415 ) | ( w2694 & w9415 ) ;
  assign w9418 = \pi01 & ~w9417 ;
  assign w9419 = ( ~\pi00 & w2805 ) | ( ~\pi00 & w9418 ) | ( w2805 & w9418 ) ;
  assign w9420 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9419 ) | ( \pi02 & ~w9419 ) ;
  assign w9421 = ( w9416 & w9418 ) | ( w9416 & ~w9420 ) | ( w9418 & ~w9420 ) ;
  assign w9422 = ( \pi02 & \pi03 ) | ( \pi02 & ~w2871 ) | ( \pi03 & ~w2871 ) ;
  assign w9423 = \pi02 & \pi03 ;
  assign w9424 = w2973 ^ w9423 ;
  assign w9425 = ( \pi04 & w9423 ) | ( \pi04 & ~w9424 ) | ( w9423 & ~w9424 ) ;
  assign w9426 = w9422 ^ w9425 ;
  assign w9427 = w6338 & ~w9421 ;
  assign w9428 = ( w8954 & w9421 ) | ( w8954 & ~w9427 ) | ( w9421 & ~w9427 ) ;
  assign w9429 = \pi02 ^ w9428 ;
  assign w9430 = ( w9413 & w9426 ) | ( w9413 & w9429 ) | ( w9426 & w9429 ) ;
  assign w9431 = ( \pi02 & w2578 ) | ( \pi02 & w2653 ) | ( w2578 & w2653 ) ;
  assign w9432 = \pi00 ^ w9431 ;
  assign w9433 = ( \pi02 & ~w2578 ) | ( \pi02 & w9432 ) | ( ~w2578 & w9432 ) ;
  assign w9434 = ( ~\pi02 & w2653 ) | ( ~\pi02 & w9432 ) | ( w2653 & w9432 ) ;
  assign w9435 = \pi01 & ~w9434 ;
  assign w9436 = ( \pi00 & w2694 ) | ( \pi00 & ~w9435 ) | ( w2694 & ~w9435 ) ;
  assign w9437 = ( \pi01 & \pi02 ) | ( \pi01 & w9436 ) | ( \pi02 & w9436 ) ;
  assign w9438 = ( w9433 & w9435 ) | ( w9433 & ~w9437 ) | ( w9435 & ~w9437 ) ;
  assign w9439 = w6282 | w8954 ;
  assign w9440 = ( ~w6282 & w9438 ) | ( ~w6282 & w9439 ) | ( w9438 & w9439 ) ;
  assign w9441 = \pi02 ^ w9440 ;
  assign w9442 = w9283 ^ w9291 ;
  assign w9443 = ( w9430 & w9441 ) | ( w9430 & w9442 ) | ( w9441 & w9442 ) ;
  assign w9444 = ( \pi02 & ~w2500 ) | ( \pi02 & w2578 ) | ( ~w2500 & w2578 ) ;
  assign w9445 = \pi00 ^ w9444 ;
  assign w9446 = ( \pi02 & w2500 ) | ( \pi02 & w9445 ) | ( w2500 & w9445 ) ;
  assign w9447 = ( ~\pi02 & w2578 ) | ( ~\pi02 & w9445 ) | ( w2578 & w9445 ) ;
  assign w9448 = \pi01 & ~w9447 ;
  assign w9449 = ( \pi00 & w2653 ) | ( \pi00 & ~w9448 ) | ( w2653 & ~w9448 ) ;
  assign w9450 = ( \pi01 & \pi02 ) | ( \pi01 & w9449 ) | ( \pi02 & w9449 ) ;
  assign w9451 = ( w9446 & w9448 ) | ( w9446 & ~w9450 ) | ( w9448 & ~w9450 ) ;
  assign w9452 = w6219 & ~w8954 ;
  assign w9453 = ( w6219 & w9451 ) | ( w6219 & ~w9452 ) | ( w9451 & ~w9452 ) ;
  assign w9454 = \pi02 ^ w9453 ;
  assign w9455 = w9294 ^ w9302 ;
  assign w9456 = ( w9443 & w9454 ) | ( w9443 & w9455 ) | ( w9454 & w9455 ) ;
  assign w9457 = ( ~\pi02 & w2391 ) | ( ~\pi02 & w2500 ) | ( w2391 & w2500 ) ;
  assign w9458 = \pi00 ^ w9457 ;
  assign w9459 = ( \pi02 & w2391 ) | ( \pi02 & ~w9458 ) | ( w2391 & ~w9458 ) ;
  assign w9460 = ( \pi02 & w2500 ) | ( \pi02 & w9458 ) | ( w2500 & w9458 ) ;
  assign w9461 = \pi01 & w9460 ;
  assign w9462 = ( \pi00 & w2578 ) | ( \pi00 & ~w9461 ) | ( w2578 & ~w9461 ) ;
  assign w9463 = ( \pi01 & \pi02 ) | ( \pi01 & w9462 ) | ( \pi02 & w9462 ) ;
  assign w9464 = ( w9459 & w9461 ) | ( w9459 & ~w9463 ) | ( w9461 & ~w9463 ) ;
  assign w9465 = w6164 | w8954 ;
  assign w9466 = ( ~w6164 & w9464 ) | ( ~w6164 & w9465 ) | ( w9464 & w9465 ) ;
  assign w9467 = \pi02 ^ w9466 ;
  assign w9468 = w9276 ^ w9303 ;
  assign w9469 = w9268 ^ w9468 ;
  assign w9470 = ( w9456 & w9467 ) | ( w9456 & w9469 ) | ( w9467 & w9469 ) ;
  assign w9471 = ( ~\pi02 & w2273 ) | ( ~\pi02 & w2391 ) | ( w2273 & w2391 ) ;
  assign w9472 = \pi00 ^ w9471 ;
  assign w9473 = ( \pi02 & w2273 ) | ( \pi02 & ~w9472 ) | ( w2273 & ~w9472 ) ;
  assign w9474 = ( \pi02 & w2391 ) | ( \pi02 & w9472 ) | ( w2391 & w9472 ) ;
  assign w9475 = \pi01 & w9474 ;
  assign w9476 = ( ~\pi00 & w2500 ) | ( ~\pi00 & w9475 ) | ( w2500 & w9475 ) ;
  assign w9477 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9476 ) | ( \pi02 & ~w9476 ) ;
  assign w9478 = ( w9473 & w9475 ) | ( w9473 & ~w9477 ) | ( w9475 & ~w9477 ) ;
  assign w9479 = w5880 & ~w8954 ;
  assign w9480 = ( w5880 & w9478 ) | ( w5880 & ~w9479 ) | ( w9478 & ~w9479 ) ;
  assign w9481 = \pi02 ^ w9480 ;
  assign w9482 = w9262 ^ w9304 ;
  assign w9483 = w9263 ^ w9482 ;
  assign w9484 = ( w9470 & w9481 ) | ( w9470 & w9483 ) | ( w9481 & w9483 ) ;
  assign w9485 = ( \pi02 & w2235 ) | ( \pi02 & ~w2273 ) | ( w2235 & ~w2273 ) ;
  assign w9486 = \pi00 ^ w9485 ;
  assign w9487 = ( \pi02 & ~w2235 ) | ( \pi02 & w9486 ) | ( ~w2235 & w9486 ) ;
  assign w9488 = ( \pi02 & w2273 ) | ( \pi02 & ~w9486 ) | ( w2273 & ~w9486 ) ;
  assign w9489 = \pi01 & w9488 ;
  assign w9490 = ( ~\pi00 & w2391 ) | ( ~\pi00 & w9489 ) | ( w2391 & w9489 ) ;
  assign w9491 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9490 ) | ( \pi02 & ~w9490 ) ;
  assign w9492 = ( w9487 & w9489 ) | ( w9487 & ~w9491 ) | ( w9489 & ~w9491 ) ;
  assign w9493 = w6106 | w8954 ;
  assign w9494 = ( ~w6106 & w9492 ) | ( ~w6106 & w9493 ) | ( w9492 & w9493 ) ;
  assign w9495 = \pi02 ^ w9494 ;
  assign w9496 = w9246 ^ w9305 ;
  assign w9497 = w9254 ^ w9496 ;
  assign w9498 = ( w9484 & w9495 ) | ( w9484 & w9497 ) | ( w9495 & w9497 ) ;
  assign w9499 = ( \pi02 & w2130 ) | ( \pi02 & w2235 ) | ( w2130 & w2235 ) ;
  assign w9500 = \pi00 ^ w9499 ;
  assign w9501 = ( \pi02 & ~w2130 ) | ( \pi02 & w9500 ) | ( ~w2130 & w9500 ) ;
  assign w9502 = ( ~\pi02 & w2235 ) | ( ~\pi02 & w9500 ) | ( w2235 & w9500 ) ;
  assign w9503 = \pi01 & ~w9502 ;
  assign w9504 = ( ~\pi00 & w2273 ) | ( ~\pi00 & w9503 ) | ( w2273 & w9503 ) ;
  assign w9505 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9504 ) | ( \pi02 & ~w9504 ) ;
  assign w9506 = ( w9501 & w9503 ) | ( w9501 & ~w9505 ) | ( w9503 & ~w9505 ) ;
  assign w9507 = w6094 & ~w8954 ;
  assign w9508 = ( w6094 & w9506 ) | ( w6094 & ~w9507 ) | ( w9506 & ~w9507 ) ;
  assign w9509 = \pi02 ^ w9508 ;
  assign w9510 = w9242 ^ w9306 ;
  assign w9511 = w9244 ^ w9510 ;
  assign w9512 = ( w9498 & w9509 ) | ( w9498 & w9511 ) | ( w9509 & w9511 ) ;
  assign w9513 = w9226 ^ w9307 ;
  assign w9514 = w9234 ^ w9513 ;
  assign w9515 = ( \pi02 & w2059 ) | ( \pi02 & w2130 ) | ( w2059 & w2130 ) ;
  assign w9516 = \pi00 ^ w9515 ;
  assign w9517 = ( \pi02 & ~w2059 ) | ( \pi02 & w9516 ) | ( ~w2059 & w9516 ) ;
  assign w9518 = ( ~\pi02 & w2130 ) | ( ~\pi02 & w9516 ) | ( w2130 & w9516 ) ;
  assign w9519 = \pi01 & ~w9518 ;
  assign w9520 = ( \pi00 & w2235 ) | ( \pi00 & ~w9519 ) | ( w2235 & ~w9519 ) ;
  assign w9521 = ( \pi01 & \pi02 ) | ( \pi01 & w9520 ) | ( \pi02 & w9520 ) ;
  assign w9522 = ( w9517 & w9519 ) | ( w9517 & ~w9521 ) | ( w9519 & ~w9521 ) ;
  assign w9523 = ( ~w5896 & w8954 ) | ( ~w5896 & w9522 ) | ( w8954 & w9522 ) ;
  assign w9524 = w9522 | w9523 ;
  assign w9525 = w9216 ^ w9308 ;
  assign w9526 = w9224 ^ w9525 ;
  assign w9527 = ( \pi02 & ~w1976 ) | ( \pi02 & w2059 ) | ( ~w1976 & w2059 ) ;
  assign w9528 = \pi00 ^ w9527 ;
  assign w9529 = ( \pi02 & w1976 ) | ( \pi02 & w9528 ) | ( w1976 & w9528 ) ;
  assign w9530 = ( ~\pi02 & w2059 ) | ( ~\pi02 & w9528 ) | ( w2059 & w9528 ) ;
  assign w9531 = \pi01 & ~w9530 ;
  assign w9532 = ( \pi00 & w2130 ) | ( \pi00 & ~w9531 ) | ( w2130 & ~w9531 ) ;
  assign w9533 = ( \pi01 & \pi02 ) | ( \pi01 & w9532 ) | ( \pi02 & w9532 ) ;
  assign w9534 = ( w9529 & w9531 ) | ( w9529 & ~w9533 ) | ( w9531 & ~w9533 ) ;
  assign w9535 = ( w5646 & w8954 ) | ( w5646 & w9534 ) | ( w8954 & w9534 ) ;
  assign w9536 = w9534 | w9535 ;
  assign w9537 = \pi02 ^ w9524 ;
  assign w9538 = ( w9512 & w9514 ) | ( w9512 & w9537 ) | ( w9514 & w9537 ) ;
  assign w9539 = \pi02 ^ w9536 ;
  assign w9540 = ( w9526 & w9538 ) | ( w9526 & w9539 ) | ( w9538 & w9539 ) ;
  assign w9541 = ( \pi02 & w1939 ) | ( \pi02 & ~w1976 ) | ( w1939 & ~w1976 ) ;
  assign w9542 = \pi00 ^ w9541 ;
  assign w9543 = ( \pi02 & ~w1939 ) | ( \pi02 & w9542 ) | ( ~w1939 & w9542 ) ;
  assign w9544 = ( \pi02 & w1976 ) | ( \pi02 & ~w9542 ) | ( w1976 & ~w9542 ) ;
  assign w9545 = \pi01 & w9544 ;
  assign w9546 = ( \pi00 & w2059 ) | ( \pi00 & ~w9545 ) | ( w2059 & ~w9545 ) ;
  assign w9547 = ( \pi01 & \pi02 ) | ( \pi01 & w9546 ) | ( \pi02 & w9546 ) ;
  assign w9548 = ( w9543 & w9545 ) | ( w9543 & ~w9547 ) | ( w9545 & ~w9547 ) ;
  assign w9549 = ( w5748 & w8954 ) | ( w5748 & w9548 ) | ( w8954 & w9548 ) ;
  assign w9550 = w9548 | w9549 ;
  assign w9551 = ( \pi02 & w1834 ) | ( \pi02 & w1939 ) | ( w1834 & w1939 ) ;
  assign w9552 = \pi00 ^ w9551 ;
  assign w9553 = ( \pi02 & ~w1834 ) | ( \pi02 & w9552 ) | ( ~w1834 & w9552 ) ;
  assign w9554 = ( ~\pi02 & w1939 ) | ( ~\pi02 & w9552 ) | ( w1939 & w9552 ) ;
  assign w9555 = \pi01 & ~w9554 ;
  assign w9556 = ( ~\pi00 & w1976 ) | ( ~\pi00 & w9555 ) | ( w1976 & w9555 ) ;
  assign w9557 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9556 ) | ( \pi02 & ~w9556 ) ;
  assign w9558 = ( w9553 & w9555 ) | ( w9553 & ~w9557 ) | ( w9555 & ~w9557 ) ;
  assign w9559 = ( ~w5659 & w8954 ) | ( ~w5659 & w9558 ) | ( w8954 & w9558 ) ;
  assign w9560 = w9558 | w9559 ;
  assign w9561 = w9202 ^ w9310 ;
  assign w9562 = w9204 ^ w9561 ;
  assign w9563 = \pi02 ^ w9550 ;
  assign w9564 = ( w9395 & w9540 ) | ( w9395 & w9563 ) | ( w9540 & w9563 ) ;
  assign w9565 = \pi02 ^ w9560 ;
  assign w9566 = ( w9562 & w9564 ) | ( w9562 & w9565 ) | ( w9564 & w9565 ) ;
  assign w9567 = ( \pi02 & ~w1711 ) | ( \pi02 & w1834 ) | ( ~w1711 & w1834 ) ;
  assign w9568 = \pi00 ^ w9567 ;
  assign w9569 = ( \pi02 & w1711 ) | ( \pi02 & w9568 ) | ( w1711 & w9568 ) ;
  assign w9570 = ( ~\pi02 & w1834 ) | ( ~\pi02 & w9568 ) | ( w1834 & w9568 ) ;
  assign w9571 = \pi01 & ~w9570 ;
  assign w9572 = ( \pi00 & w1939 ) | ( \pi00 & ~w9571 ) | ( w1939 & ~w9571 ) ;
  assign w9573 = ( \pi01 & \pi02 ) | ( \pi01 & w9572 ) | ( \pi02 & w9572 ) ;
  assign w9574 = ( w9569 & w9571 ) | ( w9569 & ~w9573 ) | ( w9571 & ~w9573 ) ;
  assign w9575 = w5296 & ~w8954 ;
  assign w9576 = ( w5296 & w9574 ) | ( w5296 & ~w9575 ) | ( w9574 & ~w9575 ) ;
  assign w9577 = \pi02 ^ w9576 ;
  assign w9578 = w9192 ^ w9311 ;
  assign w9579 = w9194 ^ w9578 ;
  assign w9580 = ( w9566 & w9577 ) | ( w9566 & w9579 ) | ( w9577 & w9579 ) ;
  assign w9581 = ( ~\pi02 & w1614 ) | ( ~\pi02 & w1711 ) | ( w1614 & w1711 ) ;
  assign w9582 = \pi00 ^ w9581 ;
  assign w9583 = ( \pi02 & w1614 ) | ( \pi02 & ~w9582 ) | ( w1614 & ~w9582 ) ;
  assign w9584 = ( \pi02 & w1711 ) | ( \pi02 & w9582 ) | ( w1711 & w9582 ) ;
  assign w9585 = \pi01 & w9584 ;
  assign w9586 = ( \pi00 & w1834 ) | ( \pi00 & ~w9585 ) | ( w1834 & ~w9585 ) ;
  assign w9587 = ( \pi01 & \pi02 ) | ( \pi01 & w9586 ) | ( \pi02 & w9586 ) ;
  assign w9588 = ( w9583 & w9585 ) | ( w9583 & ~w9587 ) | ( w9585 & ~w9587 ) ;
  assign w9589 = w5433 | w8954 ;
  assign w9590 = ( ~w5433 & w9588 ) | ( ~w5433 & w9589 ) | ( w9588 & w9589 ) ;
  assign w9591 = \pi02 ^ w9590 ;
  assign w9592 = w9182 ^ w9312 ;
  assign w9593 = w9184 ^ w9592 ;
  assign w9594 = ( w9580 & w9591 ) | ( w9580 & w9593 ) | ( w9591 & w9593 ) ;
  assign w9595 = w9166 ^ w9313 ;
  assign w9596 = w9174 ^ w9595 ;
  assign w9597 = ( \pi02 & w1510 ) | ( \pi02 & ~w1614 ) | ( w1510 & ~w1614 ) ;
  assign w9598 = \pi00 ^ w9597 ;
  assign w9599 = ( \pi02 & ~w1510 ) | ( \pi02 & w9598 ) | ( ~w1510 & w9598 ) ;
  assign w9600 = ( \pi02 & w1614 ) | ( \pi02 & ~w9598 ) | ( w1614 & ~w9598 ) ;
  assign w9601 = \pi01 & w9600 ;
  assign w9602 = ( ~\pi00 & w1711 ) | ( ~\pi00 & w9601 ) | ( w1711 & w9601 ) ;
  assign w9603 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9602 ) | ( \pi02 & ~w9602 ) ;
  assign w9604 = ( w9599 & w9601 ) | ( w9599 & ~w9603 ) | ( w9601 & ~w9603 ) ;
  assign w9605 = ( ~w5085 & w8954 ) | ( ~w5085 & w9604 ) | ( w8954 & w9604 ) ;
  assign w9606 = w9604 | w9605 ;
  assign w9607 = w9156 ^ w9314 ;
  assign w9608 = w9164 ^ w9607 ;
  assign w9609 = ( \pi02 & ~w1399 ) | ( \pi02 & w1510 ) | ( ~w1399 & w1510 ) ;
  assign w9610 = \pi00 ^ w9609 ;
  assign w9611 = ( \pi02 & w1399 ) | ( \pi02 & w9610 ) | ( w1399 & w9610 ) ;
  assign w9612 = ( ~\pi02 & w1510 ) | ( ~\pi02 & w9610 ) | ( w1510 & w9610 ) ;
  assign w9613 = \pi01 & ~w9612 ;
  assign w9614 = ( ~\pi00 & w1614 ) | ( ~\pi00 & w9613 ) | ( w1614 & w9613 ) ;
  assign w9615 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9614 ) | ( \pi02 & ~w9614 ) ;
  assign w9616 = ( w9611 & w9613 ) | ( w9611 & ~w9615 ) | ( w9613 & ~w9615 ) ;
  assign w9617 = ( ~w5069 & w8954 ) | ( ~w5069 & w9616 ) | ( w8954 & w9616 ) ;
  assign w9618 = w9616 | w9617 ;
  assign w9619 = \pi02 ^ w9606 ;
  assign w9620 = ( w9594 & w9596 ) | ( w9594 & w9619 ) | ( w9596 & w9619 ) ;
  assign w9621 = \pi02 ^ w9618 ;
  assign w9622 = ( w9608 & w9620 ) | ( w9608 & w9621 ) | ( w9620 & w9621 ) ;
  assign w9623 = ( \pi02 & w1264 ) | ( \pi02 & ~w1399 ) | ( w1264 & ~w1399 ) ;
  assign w9624 = \pi00 ^ w9623 ;
  assign w9625 = ( \pi02 & ~w1264 ) | ( \pi02 & w9624 ) | ( ~w1264 & w9624 ) ;
  assign w9626 = ( \pi02 & w1399 ) | ( \pi02 & ~w9624 ) | ( w1399 & ~w9624 ) ;
  assign w9627 = \pi01 & w9626 ;
  assign w9628 = ( \pi00 & w1510 ) | ( \pi00 & ~w9627 ) | ( w1510 & ~w9627 ) ;
  assign w9629 = ( \pi01 & \pi02 ) | ( \pi01 & w9628 ) | ( \pi02 & w9628 ) ;
  assign w9630 = ( w9625 & w9627 ) | ( w9625 & ~w9629 ) | ( w9627 & ~w9629 ) ;
  assign w9631 = ( ~w4852 & w8954 ) | ( ~w4852 & w9630 ) | ( w8954 & w9630 ) ;
  assign w9632 = w9630 | w9631 ;
  assign w9633 = ( \pi02 & ~w1205 ) | ( \pi02 & w1264 ) | ( ~w1205 & w1264 ) ;
  assign w9634 = \pi00 ^ w9633 ;
  assign w9635 = ( \pi02 & w1205 ) | ( \pi02 & w9634 ) | ( w1205 & w9634 ) ;
  assign w9636 = ( ~\pi02 & w1264 ) | ( ~\pi02 & w9634 ) | ( w1264 & w9634 ) ;
  assign w9637 = \pi01 & ~w9636 ;
  assign w9638 = ( ~\pi00 & w1399 ) | ( ~\pi00 & w9637 ) | ( w1399 & w9637 ) ;
  assign w9639 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9638 ) | ( \pi02 & ~w9638 ) ;
  assign w9640 = ( w9635 & w9637 ) | ( w9635 & ~w9639 ) | ( w9637 & ~w9639 ) ;
  assign w9641 = ( ~w4864 & w8954 ) | ( ~w4864 & w9640 ) | ( w8954 & w9640 ) ;
  assign w9642 = w9640 | w9641 ;
  assign w9643 = w9142 ^ w9316 ;
  assign w9644 = w9144 ^ w9643 ;
  assign w9645 = \pi02 ^ w9632 ;
  assign w9646 = ( w9393 & w9622 ) | ( w9393 & w9645 ) | ( w9622 & w9645 ) ;
  assign w9647 = \pi02 ^ w9642 ;
  assign w9648 = ( w9644 & w9646 ) | ( w9644 & w9647 ) | ( w9646 & w9647 ) ;
  assign w9649 = ( ~\pi02 & w1085 ) | ( ~\pi02 & w1205 ) | ( w1085 & w1205 ) ;
  assign w9650 = \pi00 ^ w9649 ;
  assign w9651 = ( \pi02 & w1085 ) | ( \pi02 & ~w9650 ) | ( w1085 & ~w9650 ) ;
  assign w9652 = ( \pi02 & w1205 ) | ( \pi02 & w9650 ) | ( w1205 & w9650 ) ;
  assign w9653 = \pi01 & w9652 ;
  assign w9654 = ( \pi00 & w1264 ) | ( \pi00 & ~w9653 ) | ( w1264 & ~w9653 ) ;
  assign w9655 = ( \pi01 & \pi02 ) | ( \pi01 & w9654 ) | ( \pi02 & w9654 ) ;
  assign w9656 = ( w9651 & w9653 ) | ( w9651 & ~w9655 ) | ( w9653 & ~w9655 ) ;
  assign w9657 = w4533 & ~w8954 ;
  assign w9658 = ( w4533 & w9656 ) | ( w4533 & ~w9657 ) | ( w9656 & ~w9657 ) ;
  assign w9659 = \pi02 ^ w9658 ;
  assign w9660 = w9132 ^ w9317 ;
  assign w9661 = w9134 ^ w9660 ;
  assign w9662 = ( w9648 & w9659 ) | ( w9648 & w9661 ) | ( w9659 & w9661 ) ;
  assign w9663 = ( ~\pi02 & w979 ) | ( ~\pi02 & w1085 ) | ( w979 & w1085 ) ;
  assign w9664 = \pi00 ^ w9663 ;
  assign w9665 = ( \pi02 & w979 ) | ( \pi02 & ~w9664 ) | ( w979 & ~w9664 ) ;
  assign w9666 = ( \pi02 & w1085 ) | ( \pi02 & w9664 ) | ( w1085 & w9664 ) ;
  assign w9667 = \pi01 & w9666 ;
  assign w9668 = ( ~\pi00 & w1205 ) | ( ~\pi00 & w9667 ) | ( w1205 & w9667 ) ;
  assign w9669 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9668 ) | ( \pi02 & ~w9668 ) ;
  assign w9670 = ( w9665 & w9667 ) | ( w9665 & ~w9669 ) | ( w9667 & ~w9669 ) ;
  assign w9671 = w4666 & ~w8954 ;
  assign w9672 = ( w4666 & w9670 ) | ( w4666 & ~w9671 ) | ( w9670 & ~w9671 ) ;
  assign w9673 = \pi02 ^ w9672 ;
  assign w9674 = w9122 ^ w9318 ;
  assign w9675 = w9124 ^ w9674 ;
  assign w9676 = ( w9662 & w9673 ) | ( w9662 & w9675 ) | ( w9673 & w9675 ) ;
  assign w9677 = w9106 ^ w9319 ;
  assign w9678 = w9114 ^ w9677 ;
  assign w9679 = ( \pi02 & w883 ) | ( \pi02 & ~w979 ) | ( w883 & ~w979 ) ;
  assign w9680 = \pi00 ^ w9679 ;
  assign w9681 = ( \pi02 & ~w883 ) | ( \pi02 & w9680 ) | ( ~w883 & w9680 ) ;
  assign w9682 = ( \pi02 & w979 ) | ( \pi02 & ~w9680 ) | ( w979 & ~w9680 ) ;
  assign w9683 = \pi01 & w9682 ;
  assign w9684 = ( ~\pi00 & w1085 ) | ( ~\pi00 & w9683 ) | ( w1085 & w9683 ) ;
  assign w9685 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9684 ) | ( \pi02 & ~w9684 ) ;
  assign w9686 = ( w9681 & w9683 ) | ( w9681 & ~w9685 ) | ( w9683 & ~w9685 ) ;
  assign w9687 = ( ~w4273 & w8954 ) | ( ~w4273 & w9686 ) | ( w8954 & w9686 ) ;
  assign w9688 = w9686 | w9687 ;
  assign w9689 = w9096 ^ w9320 ;
  assign w9690 = w9104 ^ w9689 ;
  assign w9691 = ( \pi02 & ~w721 ) | ( \pi02 & w883 ) | ( ~w721 & w883 ) ;
  assign w9692 = \pi00 ^ w9691 ;
  assign w9693 = ( \pi02 & w721 ) | ( \pi02 & w9692 ) | ( w721 & w9692 ) ;
  assign w9694 = ( ~\pi02 & w883 ) | ( ~\pi02 & w9692 ) | ( w883 & w9692 ) ;
  assign w9695 = \pi01 & ~w9694 ;
  assign w9696 = ( ~\pi00 & w979 ) | ( ~\pi00 & w9695 ) | ( w979 & w9695 ) ;
  assign w9697 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9696 ) | ( \pi02 & ~w9696 ) ;
  assign w9698 = ( w9693 & w9695 ) | ( w9693 & ~w9697 ) | ( w9695 & ~w9697 ) ;
  assign w9699 = ( ~w4257 & w8954 ) | ( ~w4257 & w9698 ) | ( w8954 & w9698 ) ;
  assign w9700 = w9698 | w9699 ;
  assign w9701 = \pi02 ^ w9688 ;
  assign w9702 = ( w9676 & w9678 ) | ( w9676 & w9701 ) | ( w9678 & w9701 ) ;
  assign w9703 = \pi02 ^ w9700 ;
  assign w9704 = ( w9690 & w9702 ) | ( w9690 & w9703 ) | ( w9702 & w9703 ) ;
  assign w9705 = ( ~\pi02 & w592 ) | ( ~\pi02 & w721 ) | ( w592 & w721 ) ;
  assign w9706 = \pi00 ^ w9705 ;
  assign w9707 = ( \pi02 & w592 ) | ( \pi02 & ~w9706 ) | ( w592 & ~w9706 ) ;
  assign w9708 = ( \pi02 & w721 ) | ( \pi02 & w9706 ) | ( w721 & w9706 ) ;
  assign w9709 = \pi01 & w9708 ;
  assign w9710 = ( \pi00 & w883 ) | ( \pi00 & ~w9709 ) | ( w883 & ~w9709 ) ;
  assign w9711 = ( \pi01 & \pi02 ) | ( \pi01 & w9710 ) | ( \pi02 & w9710 ) ;
  assign w9712 = ( w9707 & w9709 ) | ( w9707 & ~w9711 ) | ( w9709 & ~w9711 ) ;
  assign w9713 = ( w3421 & w8954 ) | ( w3421 & w9712 ) | ( w8954 & w9712 ) ;
  assign w9714 = w9712 | w9713 ;
  assign w9715 = ( \pi02 & w381 ) | ( \pi02 & ~w592 ) | ( w381 & ~w592 ) ;
  assign w9716 = \pi00 ^ w9715 ;
  assign w9717 = ( \pi02 & ~w381 ) | ( \pi02 & w9716 ) | ( ~w381 & w9716 ) ;
  assign w9718 = ( \pi02 & w592 ) | ( \pi02 & ~w9716 ) | ( w592 & ~w9716 ) ;
  assign w9719 = \pi01 & w9718 ;
  assign w9720 = ( ~\pi00 & w721 ) | ( ~\pi00 & w9719 ) | ( w721 & w9719 ) ;
  assign w9721 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9720 ) | ( \pi02 & ~w9720 ) ;
  assign w9722 = ( w9717 & w9719 ) | ( w9717 & ~w9721 ) | ( w9719 & ~w9721 ) ;
  assign w9723 = ( ~w3435 & w8954 ) | ( ~w3435 & w9722 ) | ( w8954 & w9722 ) ;
  assign w9724 = w9722 | w9723 ;
  assign w9725 = w9082 ^ w9322 ;
  assign w9726 = w9084 ^ w9725 ;
  assign w9727 = \pi02 ^ w9714 ;
  assign w9728 = ( w9391 & w9704 ) | ( w9391 & w9727 ) | ( w9704 & w9727 ) ;
  assign w9729 = \pi02 ^ w9724 ;
  assign w9730 = ( w9726 & w9728 ) | ( w9726 & w9729 ) | ( w9728 & w9729 ) ;
  assign w9731 = ( \pi02 & w381 ) | ( \pi02 & w3094 ) | ( w381 & w3094 ) ;
  assign w9732 = \pi00 ^ w9731 ;
  assign w9733 = ( \pi02 & ~w3094 ) | ( \pi02 & w9732 ) | ( ~w3094 & w9732 ) ;
  assign w9734 = ( ~\pi02 & w381 ) | ( ~\pi02 & w9732 ) | ( w381 & w9732 ) ;
  assign w9735 = \pi01 & ~w9734 ;
  assign w9736 = ( ~\pi00 & w592 ) | ( ~\pi00 & w9735 ) | ( w592 & w9735 ) ;
  assign w9737 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9736 ) | ( \pi02 & ~w9736 ) ;
  assign w9738 = ( w9733 & w9735 ) | ( w9733 & ~w9737 ) | ( w9735 & ~w9737 ) ;
  assign w9739 = w3096 & ~w8954 ;
  assign w9740 = ( w3096 & w9738 ) | ( w3096 & ~w9739 ) | ( w9738 & ~w9739 ) ;
  assign w9741 = \pi02 ^ w9740 ;
  assign w9742 = w9072 ^ w9323 ;
  assign w9743 = w9074 ^ w9742 ;
  assign w9744 = ( w9730 & w9741 ) | ( w9730 & w9743 ) | ( w9741 & w9743 ) ;
  assign w9745 = ( \pi02 & w3094 ) | ( \pi02 & ~w3647 ) | ( w3094 & ~w3647 ) ;
  assign w9746 = \pi00 ^ w9745 ;
  assign w9747 = ( \pi02 & w3647 ) | ( \pi02 & w9746 ) | ( w3647 & w9746 ) ;
  assign w9748 = ( ~\pi02 & w3094 ) | ( ~\pi02 & w9746 ) | ( w3094 & w9746 ) ;
  assign w9749 = \pi01 & ~w9748 ;
  assign w9750 = ( \pi00 & w381 ) | ( \pi00 & ~w9749 ) | ( w381 & ~w9749 ) ;
  assign w9751 = ( \pi01 & \pi02 ) | ( \pi01 & w9750 ) | ( \pi02 & w9750 ) ;
  assign w9752 = ( w9747 & w9749 ) | ( w9747 & ~w9751 ) | ( w9749 & ~w9751 ) ;
  assign w9753 = w3810 & ~w8954 ;
  assign w9754 = ( w3810 & w9752 ) | ( w3810 & ~w9753 ) | ( w9752 & ~w9753 ) ;
  assign w9755 = \pi02 ^ w9754 ;
  assign w9756 = w9062 ^ w9324 ;
  assign w9757 = w9064 ^ w9756 ;
  assign w9758 = ( w9744 & w9755 ) | ( w9744 & w9757 ) | ( w9755 & w9757 ) ;
  assign w9759 = w9046 ^ w9325 ;
  assign w9760 = w9054 ^ w9759 ;
  assign w9761 = ( ~\pi02 & w3647 ) | ( ~\pi02 & w3715 ) | ( w3647 & w3715 ) ;
  assign w9762 = \pi00 ^ w9761 ;
  assign w9763 = ( \pi02 & w3715 ) | ( \pi02 & ~w9762 ) | ( w3715 & ~w9762 ) ;
  assign w9764 = ( \pi02 & w3647 ) | ( \pi02 & w9762 ) | ( w3647 & w9762 ) ;
  assign w9765 = \pi01 & w9764 ;
  assign w9766 = ( \pi00 & w3094 ) | ( \pi00 & ~w9765 ) | ( w3094 & ~w9765 ) ;
  assign w9767 = ( \pi01 & \pi02 ) | ( \pi01 & w9766 ) | ( \pi02 & w9766 ) ;
  assign w9768 = ( w9763 & w9765 ) | ( w9763 & ~w9767 ) | ( w9765 & ~w9767 ) ;
  assign w9769 = ( ~w4164 & w8954 ) | ( ~w4164 & w9768 ) | ( w8954 & w9768 ) ;
  assign w9770 = w9768 | w9769 ;
  assign w9771 = ( \pi02 & w3548 ) | ( \pi02 & ~w3715 ) | ( w3548 & ~w3715 ) ;
  assign w9772 = \pi00 ^ w9771 ;
  assign w9773 = ( \pi02 & ~w3548 ) | ( \pi02 & w9772 ) | ( ~w3548 & w9772 ) ;
  assign w9774 = ( \pi02 & w3715 ) | ( \pi02 & ~w9772 ) | ( w3715 & ~w9772 ) ;
  assign w9775 = \pi01 & w9774 ;
  assign w9776 = ( ~\pi00 & w3647 ) | ( ~\pi00 & w9775 ) | ( w3647 & w9775 ) ;
  assign w9777 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9776 ) | ( \pi02 & ~w9776 ) ;
  assign w9778 = ( w9773 & w9775 ) | ( w9773 & ~w9777 ) | ( w9775 & ~w9777 ) ;
  assign w9779 = ( ~w3725 & w8954 ) | ( ~w3725 & w9778 ) | ( w8954 & w9778 ) ;
  assign w9780 = w9778 | w9779 ;
  assign w9781 = \pi02 ^ w9770 ;
  assign w9782 = ( w9758 & w9760 ) | ( w9758 & w9781 ) | ( w9760 & w9781 ) ;
  assign w9783 = \pi02 ^ w9780 ;
  assign w9784 = ( w9389 & w9782 ) | ( w9389 & w9783 ) | ( w9782 & w9783 ) ;
  assign w9785 = ( \pi02 & w3548 ) | ( \pi02 & ~w3907 ) | ( w3548 & ~w3907 ) ;
  assign w9786 = \pi00 ^ w9785 ;
  assign w9787 = ( \pi02 & w3907 ) | ( \pi02 & w9786 ) | ( w3907 & w9786 ) ;
  assign w9788 = ( ~\pi02 & w3548 ) | ( ~\pi02 & w9786 ) | ( w3548 & w9786 ) ;
  assign w9789 = \pi01 & ~w9788 ;
  assign w9790 = ( ~\pi00 & w3715 ) | ( ~\pi00 & w9789 ) | ( w3715 & w9789 ) ;
  assign w9791 = ( \pi01 & \pi02 ) | ( \pi01 & ~w9790 ) | ( \pi02 & ~w9790 ) ;
  assign w9792 = ( w9787 & w9789 ) | ( w9787 & ~w9791 ) | ( w9789 & ~w9791 ) ;
  assign w9793 = w3913 | w8954 ;
  assign w9794 = ( ~w3913 & w9792 ) | ( ~w3913 & w9793 ) | ( w9792 & w9793 ) ;
  assign w9795 = \pi02 ^ w9794 ;
  assign w9796 = w9032 ^ w9327 ;
  assign w9797 = w9034 ^ w9796 ;
  assign w9798 = ( w9784 & w9795 ) | ( w9784 & w9797 ) | ( w9795 & w9797 ) ;
  assign w9799 = w4622 & ~w9387 ;
  assign w9800 = ( w8954 & w9387 ) | ( w8954 & ~w9799 ) | ( w9387 & ~w9799 ) ;
  assign w9801 = \pi02 ^ w9800 ;
  assign w9802 = ( ~w9379 & w9798 ) | ( ~w9379 & w9801 ) | ( w9798 & w9801 ) ;
  assign w9803 = w4563 | w9377 ;
  assign w9804 = ( w8954 & w9377 ) | ( w8954 & w9803 ) | ( w9377 & w9803 ) ;
  assign w9805 = \pi02 ^ w9804 ;
  assign w9806 = ( ~w9369 & w9802 ) | ( ~w9369 & w9805 ) | ( w9802 & w9805 ) ;
  assign w9807 = w4152 & ~w9367 ;
  assign w9808 = ( w8954 & w9367 ) | ( w8954 & ~w9807 ) | ( w9367 & ~w9807 ) ;
  assign w9809 = \pi02 ^ w9808 ;
  assign w9810 = ( w9359 & w9806 ) | ( w9359 & w9809 ) | ( w9806 & w9809 ) ;
  assign w9811 = w4722 & ~w9357 ;
  assign w9812 = ( w8954 & w9357 ) | ( w8954 & ~w9811 ) | ( w9357 & ~w9811 ) ;
  assign w9813 = \pi02 ^ w9812 ;
  assign w9814 = ( ~w9349 & w9810 ) | ( ~w9349 & w9813 ) | ( w9810 & w9813 ) ;
  assign w9815 = ( w9335 & w9347 ) | ( w9335 & w9814 ) | ( w9347 & w9814 ) ;
  assign w9816 = ( w8974 & w9333 ) | ( w8974 & w9815 ) | ( w9333 & w9815 ) ;
  assign w9817 = ( w8970 & w8972 ) | ( w8970 & w9816 ) | ( w8972 & w9816 ) ;
  assign w9818 = ( w8949 & w8952 ) | ( w8949 & w9817 ) | ( w8952 & w9817 ) ;
  assign w9819 = ( ~w8277 & w8602 ) | ( ~w8277 & w9818 ) | ( w8602 & w9818 ) ;
  assign w9820 = ( w8270 & w8275 ) | ( w8270 & w9819 ) | ( w8275 & w9819 ) ;
  assign w9821 = ( w7964 & ~w7967 ) | ( w7964 & w9820 ) | ( ~w7967 & w9820 ) ;
  assign w9822 = ( w7423 & w7682 ) | ( w7423 & w9821 ) | ( w7682 & w9821 ) ;
  assign w9823 = ( w7182 & w7421 ) | ( w7182 & w9822 ) | ( w7421 & w9822 ) ;
  assign w9824 = ( w7174 & w7177 ) | ( w7174 & w9823 ) | ( w7177 & w9823 ) ;
  assign w9825 = ( w6765 & w6958 ) | ( w6765 & w9824 ) | ( w6958 & w9824 ) ;
  assign w9826 = ( w6758 & w6763 ) | ( w6758 & w9825 ) | ( w6763 & w9825 ) ;
  assign w9827 = ( w6657 & w6660 ) | ( w6657 & w9826 ) | ( w6660 & w9826 ) ;
  assign w9828 = ( w6062 & w6560 ) | ( w6062 & w9827 ) | ( w6560 & w9827 ) ;
  assign w9829 = ( w6055 & ~w6060 ) | ( w6055 & w9828 ) | ( ~w6060 & w9828 ) ;
  assign w9830 = w5708 ^ w5716 ;
  assign w9831 = \pi17 ^ w9830 ;
  assign w9832 = ( w5968 & w9829 ) | ( w5968 & w9831 ) | ( w9829 & w9831 ) ;
  assign w9833 = ( ~w5511 & w5718 ) | ( ~w5511 & w9832 ) | ( w5718 & w9832 ) ;
  assign w9834 = ( w5504 & w5509 ) | ( w5504 & w9833 ) | ( w5509 & w9833 ) ;
  assign w9835 = w5341 ^ w5349 ;
  assign w9836 = \pi20 ^ w9835 ;
  assign w9837 = ( w5415 & w9834 ) | ( w5415 & w9836 ) | ( w9834 & w9836 ) ;
  assign w9838 = ( ~w4917 & w5351 ) | ( ~w4917 & w9837 ) | ( w5351 & w9837 ) ;
  assign w9839 = ( w4736 & w4915 ) | ( w4736 & w9838 ) | ( w4915 & w9838 ) ;
  assign w9840 = ( w4728 & ~w4731 ) | ( w4728 & w9839 ) | ( ~w4731 & w9839 ) ;
  assign w9841 = w4615 ^ w9840 ;
  assign w9842 = w4660 ^ w9841 ;
  assign w9843 = ( w4615 & w4660 ) | ( w4615 & w9840 ) | ( w4660 & w9840 ) ;
  assign w9844 = ( w4159 & w4569 ) | ( w4159 & w4613 ) | ( w4569 & w4613 ) ;
  assign w9845 = w3548 | w3649 ;
  assign w9846 = w3717 & w3907 ;
  assign w9847 = ( ~w3548 & w9845 ) | ( ~w3548 & w9846 ) | ( w9845 & w9846 ) ;
  assign w9848 = w3549 | w4049 ;
  assign w9849 = w4622 & ~w9847 ;
  assign w9850 = ( w3448 & w9847 ) | ( w3448 & ~w9849 ) | ( w9847 & ~w9849 ) ;
  assign w9851 = ( ~w4049 & w9848 ) | ( ~w4049 & w9850 ) | ( w9848 & w9850 ) ;
  assign w9852 = \pi29 ^ w9851 ;
  assign w9853 = ( w3731 & w3808 ) | ( w3731 & w3818 ) | ( w3808 & w3818 ) ;
  assign w9854 = w208 | w2374 ;
  assign w9855 = ( w90 & w270 ) | ( w90 & ~w2374 ) | ( w270 & ~w2374 ) ;
  assign w9856 = w9854 | w9855 ;
  assign w9857 = w353 | w495 ;
  assign w9858 = w257 | w9857 ;
  assign w9859 = ( w179 & ~w257 ) | ( w179 & w317 ) | ( ~w257 & w317 ) ;
  assign w9860 = w9858 | w9859 ;
  assign w9861 = w389 | w465 ;
  assign w9862 = w2704 | w9861 ;
  assign w9863 = ( ~w2704 & w9856 ) | ( ~w2704 & w9860 ) | ( w9856 & w9860 ) ;
  assign w9864 = w9862 | w9863 ;
  assign w9865 = w88 | w143 ;
  assign w9866 = ( ~w88 & w133 ) | ( ~w88 & w9864 ) | ( w133 & w9864 ) ;
  assign w9867 = w9865 | w9866 ;
  assign w9868 = w390 | w1229 ;
  assign w9869 = w76 | w9868 ;
  assign w9870 = ( ~w76 & w271 ) | ( ~w76 & w1590 ) | ( w271 & w1590 ) ;
  assign w9871 = w9869 | w9870 ;
  assign w9872 = w467 | w951 ;
  assign w9873 = w253 | w9872 ;
  assign w9874 = ( ~w253 & w420 ) | ( ~w253 & w9871 ) | ( w420 & w9871 ) ;
  assign w9875 = w9873 | w9874 ;
  assign w9876 = ( w136 & w169 ) | ( w136 & ~w178 ) | ( w169 & ~w178 ) ;
  assign w9877 = w116 | w532 ;
  assign w9878 = ( ~w116 & w178 ) | ( ~w116 & w215 ) | ( w178 & w215 ) ;
  assign w9879 = w9877 | w9878 ;
  assign w9880 = w9876 | w9879 ;
  assign w9881 = w393 | w9880 ;
  assign w9882 = w272 | w447 ;
  assign w9883 = ( ~w272 & w287 ) | ( ~w272 & w2452 ) | ( w287 & w2452 ) ;
  assign w9884 = w9882 | w9883 ;
  assign w9885 = ( ~w205 & w3037 ) | ( ~w205 & w9884 ) | ( w3037 & w9884 ) ;
  assign w9886 = w1531 | w9881 ;
  assign w9887 = ( w205 & w787 ) | ( w205 & ~w1531 ) | ( w787 & ~w1531 ) ;
  assign w9888 = w9886 | w9887 ;
  assign w9889 = w9885 | w9888 ;
  assign w9890 = w266 | w785 ;
  assign w9891 = ( w119 & ~w785 ) | ( w119 & w9889 ) | ( ~w785 & w9889 ) ;
  assign w9892 = w9890 | w9891 ;
  assign w9893 = ( ~w258 & w1282 ) | ( ~w258 & w2060 ) | ( w1282 & w2060 ) ;
  assign w9894 = w900 | w9892 ;
  assign w9895 = ( w258 & w860 ) | ( w258 & ~w900 ) | ( w860 & ~w900 ) ;
  assign w9896 = w9894 | w9895 ;
  assign w9897 = w9893 | w9896 ;
  assign w9898 = ( w56 & w342 ) | ( w56 & ~w418 ) | ( w342 & ~w418 ) ;
  assign w9899 = w44 | w9897 ;
  assign w9900 = ( ~w44 & w418 ) | ( ~w44 & w445 ) | ( w418 & w445 ) ;
  assign w9901 = w9899 | w9900 ;
  assign w9902 = w9898 | w9901 ;
  assign w9903 = w283 | w637 ;
  assign w9904 = ( w111 & ~w283 ) | ( w111 & w568 ) | ( ~w283 & w568 ) ;
  assign w9905 = w9903 | w9904 ;
  assign w9906 = ( w227 & w229 ) | ( w227 & ~w361 ) | ( w229 & ~w361 ) ;
  assign w9907 = w125 | w1184 ;
  assign w9908 = ( ~w125 & w361 ) | ( ~w125 & w466 ) | ( w361 & w466 ) ;
  assign w9909 = w9907 | w9908 ;
  assign w9910 = w9906 | w9909 ;
  assign w9911 = ( w9867 & w9875 ) | ( w9867 & ~w9910 ) | ( w9875 & ~w9910 ) ;
  assign w9912 = w6429 | w9902 ;
  assign w9913 = ( ~w6429 & w9905 ) | ( ~w6429 & w9910 ) | ( w9905 & w9910 ) ;
  assign w9914 = w9912 | w9913 ;
  assign w9915 = w9911 | w9914 ;
  assign w9916 = ( w209 & w573 ) | ( w209 & ~w663 ) | ( w573 & ~w663 ) ;
  assign w9917 = w3251 | w9915 ;
  assign w9918 = ( w663 & w1340 ) | ( w663 & ~w3251 ) | ( w1340 & ~w3251 ) ;
  assign w9919 = w9917 | w9918 ;
  assign w9920 = w9916 | w9919 ;
  assign w9921 = ( w344 & w358 ) | ( w344 & ~w423 ) | ( w358 & ~w423 ) ;
  assign w9922 = w86 | w9920 ;
  assign w9923 = ( ~w86 & w423 ) | ( ~w86 & w571 ) | ( w423 & w571 ) ;
  assign w9924 = w9922 | w9923 ;
  assign w9925 = w9921 | w9924 ;
  assign w9926 = ( ~\pi23 & w3805 ) | ( ~\pi23 & w9925 ) | ( w3805 & w9925 ) ;
  assign w9927 = w3805 ^ w9925 ;
  assign w9928 = \pi23 ^ w9927 ;
  assign w9929 = w37 | w4164 ;
  assign w9930 = ~w3094 & w3098 ;
  assign w9931 = ( ~w4164 & w9929 ) | ( ~w4164 & w9930 ) | ( w9929 & w9930 ) ;
  assign w9932 = ( \pi29 & \pi30 ) | ( \pi29 & w3715 ) | ( \pi30 & w3715 ) ;
  assign w9933 = \pi31 | w9932 ;
  assign w9934 = ( \pi29 & ~\pi30 ) | ( \pi29 & w3647 ) | ( ~\pi30 & w3647 ) ;
  assign w9935 = ( \pi29 & \pi31 ) | ( \pi29 & ~w9934 ) | ( \pi31 & ~w9934 ) ;
  assign w9936 = ( w9931 & w9933 ) | ( w9931 & ~w9935 ) | ( w9933 & ~w9935 ) ;
  assign w9937 = w3806 ^ w9936 ;
  assign w9938 = w9928 ^ w9937 ;
  assign w9939 = w9852 ^ w9853 ;
  assign w9940 = w9938 ^ w9939 ;
  assign w9941 = ( w3820 & w3918 ) | ( w3820 & w4157 ) | ( w3918 & w4157 ) ;
  assign w9942 = w3964 & ~w4600 ;
  assign w9943 = ( ~w3962 & w4143 ) | ( ~w3962 & w9942 ) | ( w4143 & w9942 ) ;
  assign w9944 = w4052 | w9943 ;
  assign w9945 = ( ~w4142 & w9943 ) | ( ~w4142 & w9944 ) | ( w9943 & w9944 ) ;
  assign w9946 = w9942 | w9945 ;
  assign w9947 = w4147 & w4722 ;
  assign w9948 = ( w4147 & w9946 ) | ( w4147 & ~w9947 ) | ( w9946 & ~w9947 ) ;
  assign w9949 = w9941 ^ w9948 ;
  assign w9950 = \pi26 ^ w9940 ;
  assign w9951 = w9949 ^ w9950 ;
  assign w9952 = w9843 ^ w9844 ;
  assign w9953 = w9951 ^ w9952 ;
  assign w9954 = w4728 ^ w9839 ;
  assign w9955 = w4731 ^ w9954 ;
  assign w9956 = w4736 ^ w9838 ;
  assign w9957 = w4915 ^ w9956 ;
  assign w9958 = w5341 ^ w5415 ;
  assign w9959 = w5349 ^ w9834 ;
  assign w9960 = \pi20 ^ w9959 ;
  assign w9961 = w9958 ^ w9960 ;
  assign w9962 = w4917 ^ w9837 ;
  assign w9963 = w5351 ^ w9962 ;
  assign w9964 = w5504 ^ w9833 ;
  assign w9965 = w5509 ^ w9964 ;
  assign w9966 = w5511 ^ w9832 ;
  assign w9967 = w5718 ^ w9966 ;
  assign w9968 = w5708 ^ w5968 ;
  assign w9969 = w5716 ^ w9829 ;
  assign w9970 = \pi17 ^ w9969 ;
  assign w9971 = w9968 ^ w9970 ;
  assign w9972 = w6055 ^ w9828 ;
  assign w9973 = w6060 ^ w9972 ;
  assign w9974 = w6062 ^ w9827 ;
  assign w9975 = w6560 ^ w9974 ;
  assign w9976 = w6657 ^ w9826 ;
  assign w9977 = w6660 ^ w9976 ;
  assign w9978 = w6758 ^ w9825 ;
  assign w9979 = w6763 ^ w9978 ;
  assign w9980 = w6765 ^ w9824 ;
  assign w9981 = w6958 ^ w9980 ;
  assign w9982 = w7174 ^ w9823 ;
  assign w9983 = w7177 ^ w9982 ;
  assign w9984 = w7182 ^ w9822 ;
  assign w9985 = w7421 ^ w9984 ;
  assign w9986 = w7423 ^ w9821 ;
  assign w9987 = w7682 ^ w9986 ;
  assign w9988 = w7964 ^ w9820 ;
  assign w9989 = w7967 ^ w9988 ;
  assign w9990 = w8270 ^ w9819 ;
  assign w9991 = w8275 ^ w9990 ;
  assign w9992 = w8277 ^ w9818 ;
  assign w9993 = w8602 ^ w9992 ;
  assign w9994 = w8949 ^ w9817 ;
  assign w9995 = w8952 ^ w9994 ;
  assign w9996 = w8970 ^ w9816 ;
  assign w9997 = w8972 ^ w9996 ;
  assign w9998 = w8974 ^ w9815 ;
  assign w9999 = w9333 ^ w9998 ;
  assign w10000 = w9335 ^ w9814 ;
  assign w10001 = w9347 ^ w10000 ;
  assign w10002 = w4722 & w8954 ;
  assign w10003 = ( w8954 & w9357 ) | ( w8954 & ~w10002 ) | ( w9357 & ~w10002 ) ;
  assign w10004 = w9349 ^ w10003 ;
  assign w10005 = \pi02 ^ w9810 ;
  assign w10006 = w10004 ^ w10005 ;
  assign w10007 = w4152 & w8954 ;
  assign w10008 = ( w8954 & w9367 ) | ( w8954 & ~w10007 ) | ( w9367 & ~w10007 ) ;
  assign w10009 = w9359 ^ w10008 ;
  assign w10010 = \pi02 ^ w9806 ;
  assign w10011 = w10009 ^ w10010 ;
  assign w10012 = ~w4563 & w8954 ;
  assign w10013 = ( w8954 & w9377 ) | ( w8954 & ~w10012 ) | ( w9377 & ~w10012 ) ;
  assign w10014 = w9369 ^ w10013 ;
  assign w10015 = \pi02 ^ w9802 ;
  assign w10016 = w10014 ^ w10015 ;
  assign w10017 = w4622 & w8954 ;
  assign w10018 = ( w8954 & w9387 ) | ( w8954 & ~w10017 ) | ( w9387 & ~w10017 ) ;
  assign w10019 = w9379 ^ w10018 ;
  assign w10020 = \pi02 ^ w9798 ;
  assign w10021 = w10019 ^ w10020 ;
  assign w10022 = ( w9999 & w10001 ) | ( w9999 & ~w10006 ) | ( w10001 & ~w10006 ) ;
  assign w10023 = w10001 & ~w10016 ;
  assign w10024 = ( w10016 & w10021 ) | ( w10016 & ~w10023 ) | ( w10021 & ~w10023 ) ;
  assign w10025 = ( w10001 & ~w10011 ) | ( w10001 & w10024 ) | ( ~w10011 & w10024 ) ;
  assign w10026 = ( w10001 & w10022 ) | ( w10001 & ~w10025 ) | ( w10022 & ~w10025 ) ;
  assign w10027 = ( w9997 & w9999 ) | ( w9997 & w10026 ) | ( w9999 & w10026 ) ;
  assign w10028 = ( ~w9993 & w9995 ) | ( ~w9993 & w10027 ) | ( w9995 & w10027 ) ;
  assign w10029 = ( w9995 & w9997 ) | ( w9995 & w10028 ) | ( w9997 & w10028 ) ;
  assign w10030 = ( w9991 & ~w9993 ) | ( w9991 & w10029 ) | ( ~w9993 & w10029 ) ;
  assign w10031 = ( w9987 & ~w9989 ) | ( w9987 & w10030 ) | ( ~w9989 & w10030 ) ;
  assign w10032 = ( ~w9989 & w9991 ) | ( ~w9989 & w10031 ) | ( w9991 & w10031 ) ;
  assign w10033 = ( w9983 & w9985 ) | ( w9983 & w10032 ) | ( w9985 & w10032 ) ;
  assign w10034 = ( w9985 & w9987 ) | ( w9985 & w10033 ) | ( w9987 & w10033 ) ;
  assign w10035 = ( w9981 & w9983 ) | ( w9981 & w10034 ) | ( w9983 & w10034 ) ;
  assign w10036 = ( w9979 & w9981 ) | ( w9979 & w10035 ) | ( w9981 & w10035 ) ;
  assign w10037 = ( w9975 & w9977 ) | ( w9975 & w10036 ) | ( w9977 & w10036 ) ;
  assign w10038 = ( w9977 & w9979 ) | ( w9977 & w10037 ) | ( w9979 & w10037 ) ;
  assign w10039 = ( w9971 & ~w9973 ) | ( w9971 & w10038 ) | ( ~w9973 & w10038 ) ;
  assign w10040 = ( ~w9973 & w9975 ) | ( ~w9973 & w10039 ) | ( w9975 & w10039 ) ;
  assign w10041 = ( ~w9967 & w9971 ) | ( ~w9967 & w10040 ) | ( w9971 & w10040 ) ;
  assign w10042 = ( w9965 & ~w9967 ) | ( w9965 & w10041 ) | ( ~w9967 & w10041 ) ;
  assign w10043 = ( w9961 & w9965 ) | ( w9961 & w10042 ) | ( w9965 & w10042 ) ;
  assign w10044 = ( w9957 & ~w9963 ) | ( w9957 & w10043 ) | ( ~w9963 & w10043 ) ;
  assign w10045 = ( w9961 & ~w9963 ) | ( w9961 & w10044 ) | ( ~w9963 & w10044 ) ;
  assign w10046 = ( ~w9955 & w9957 ) | ( ~w9955 & w10045 ) | ( w9957 & w10045 ) ;
  assign w10047 = ( w9842 & ~w9955 ) | ( w9842 & w10046 ) | ( ~w9955 & w10046 ) ;
  assign w10048 = ( w9842 & w9953 ) | ( w9842 & w10047 ) | ( w9953 & w10047 ) ;
  assign w10049 = ( w9843 & w9844 ) | ( w9843 & w9951 ) | ( w9844 & w9951 ) ;
  assign w10050 = w4722 & ~w9946 ;
  assign w10051 = ( w4147 & w9946 ) | ( w4147 & ~w10050 ) | ( w9946 & ~w10050 ) ;
  assign w10052 = \pi26 ^ w10051 ;
  assign w10053 = ( w9940 & w9941 ) | ( w9940 & w10052 ) | ( w9941 & w10052 ) ;
  assign w10054 = w4143 & ~w4600 ;
  assign w10055 = ( ~w3962 & w4052 ) | ( ~w3962 & w10054 ) | ( w4052 & w10054 ) ;
  assign w10056 = ( ~w3962 & w4601 ) | ( ~w3962 & w10055 ) | ( w4601 & w10055 ) ;
  assign w10057 = ( w4147 & w4600 ) | ( w4147 & w4601 ) | ( w4600 & w4601 ) ;
  assign w10058 = ( w10054 & ~w10056 ) | ( w10054 & w10057 ) | ( ~w10056 & w10057 ) ;
  assign w10059 = ( ~w4657 & w10055 ) | ( ~w4657 & w10058 ) | ( w10055 & w10058 ) ;
  assign w10060 = ( w9852 & w9853 ) | ( w9852 & w9938 ) | ( w9853 & w9938 ) ;
  assign w10061 = ( \pi29 & \pi31 ) | ( \pi29 & w3715 ) | ( \pi31 & w3715 ) ;
  assign w10062 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10061 ) | ( ~\pi30 & w10061 ) ;
  assign w10063 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10061 ) | ( \pi30 & w10061 ) ;
  assign w10064 = ( ~\pi29 & w3647 ) | ( ~\pi29 & w10063 ) | ( w3647 & w10063 ) ;
  assign w10065 = ( w3548 & ~w10063 ) | ( w3548 & w10064 ) | ( ~w10063 & w10064 ) ;
  assign w10066 = \pi31 | w10065 ;
  assign w10067 = ( w10062 & w10064 ) | ( w10062 & ~w10066 ) | ( w10064 & ~w10066 ) ;
  assign w10068 = ( w37 & ~w3725 ) | ( w37 & w10067 ) | ( ~w3725 & w10067 ) ;
  assign w10069 = w10067 | w10068 ;
  assign w10070 = ( w384 & w411 ) | ( w384 & ~w817 ) | ( w411 & ~w817 ) ;
  assign w10071 = w141 | w169 ;
  assign w10072 = ( ~w169 & w817 ) | ( ~w169 & w1126 ) | ( w817 & w1126 ) ;
  assign w10073 = w10071 | w10072 ;
  assign w10074 = w10070 | w10073 ;
  assign w10075 = ( ~w131 & w664 ) | ( ~w131 & w10074 ) | ( w664 & w10074 ) ;
  assign w10076 = w131 | w10075 ;
  assign w10077 = w209 | w383 ;
  assign w10078 = w2470 | w10077 ;
  assign w10079 = ( w176 & w1940 ) | ( w176 & ~w2470 ) | ( w1940 & ~w2470 ) ;
  assign w10080 = w10078 | w10079 ;
  assign w10081 = ( ~w1618 & w5804 ) | ( ~w1618 & w10080 ) | ( w5804 & w10080 ) ;
  assign w10082 = w1589 | w5624 ;
  assign w10083 = ( w1618 & w2625 ) | ( w1618 & ~w5624 ) | ( w2625 & ~w5624 ) ;
  assign w10084 = w10082 | w10083 ;
  assign w10085 = w10081 | w10084 ;
  assign w10086 = w2695 | w4784 ;
  assign w10087 = w10076 | w10086 ;
  assign w10088 = ( w87 & ~w10076 ) | ( w87 & w10085 ) | ( ~w10076 & w10085 ) ;
  assign w10089 = w10087 | w10088 ;
  assign w10090 = ( w68 & ~w124 ) | ( w68 & w343 ) | ( ~w124 & w343 ) ;
  assign w10091 = w82 | w10089 ;
  assign w10092 = ( ~w82 & w124 ) | ( ~w82 & w725 ) | ( w124 & w725 ) ;
  assign w10093 = w10091 | w10092 ;
  assign w10094 = w10090 | w10093 ;
  assign w10095 = ( ~w252 & w259 ) | ( ~w252 & w10094 ) | ( w259 & w10094 ) ;
  assign w10096 = w252 | w10095 ;
  assign w10097 = w9926 ^ w10069 ;
  assign w10098 = w10096 ^ w10097 ;
  assign w10099 = ( w3806 & w9928 ) | ( w3806 & ~w9936 ) | ( w9928 & ~w9936 ) ;
  assign w10100 = w3717 | w4049 ;
  assign w10101 = w3649 & w3907 ;
  assign w10102 = ( ~w4049 & w10100 ) | ( ~w4049 & w10101 ) | ( w10100 & w10101 ) ;
  assign w10103 = w3549 | w4142 ;
  assign w10104 = w4563 | w10102 ;
  assign w10105 = ( w3448 & w10102 ) | ( w3448 & w10104 ) | ( w10102 & w10104 ) ;
  assign w10106 = ( ~w4142 & w10103 ) | ( ~w4142 & w10105 ) | ( w10103 & w10105 ) ;
  assign w10107 = \pi29 ^ w10106 ;
  assign w10108 = w10098 ^ w10107 ;
  assign w10109 = w10099 ^ w10108 ;
  assign w10110 = \pi26 ^ w10060 ;
  assign w10111 = w10059 ^ w10110 ;
  assign w10112 = w10109 ^ w10111 ;
  assign w10113 = w10049 ^ w10053 ;
  assign w10114 = w10112 ^ w10113 ;
  assign w10115 = ( w10049 & w10053 ) | ( w10049 & w10112 ) | ( w10053 & w10112 ) ;
  assign w10116 = \pi26 ^ w10059 ;
  assign w10117 = ( w10060 & w10109 ) | ( w10060 & w10116 ) | ( w10109 & w10116 ) ;
  assign w10118 = ( \pi30 & \pi31 ) | ( \pi30 & ~w3548 ) | ( \pi31 & ~w3548 ) ;
  assign w10119 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10118 ) | ( \pi30 & w10118 ) ;
  assign w10120 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10118 ) | ( ~\pi30 & w10118 ) ;
  assign w10121 = ( ~\pi30 & w3715 ) | ( ~\pi30 & w10120 ) | ( w3715 & w10120 ) ;
  assign w10122 = ( w3907 & w10120 ) | ( w3907 & ~w10121 ) | ( w10120 & ~w10121 ) ;
  assign w10123 = ~\pi31 & w10122 ;
  assign w10124 = ( w10119 & w10121 ) | ( w10119 & w10123 ) | ( w10121 & w10123 ) ;
  assign w10125 = ( w37 & ~w3913 ) | ( w37 & w10124 ) | ( ~w3913 & w10124 ) ;
  assign w10126 = w10124 | w10125 ;
  assign w10127 = ( w201 & ~w286 ) | ( w201 & w2704 ) | ( ~w286 & w2704 ) ;
  assign w10128 = w660 | w2695 ;
  assign w10129 = ( w286 & w724 ) | ( w286 & ~w2695 ) | ( w724 & ~w2695 ) ;
  assign w10130 = w10128 | w10129 ;
  assign w10131 = w10127 | w10130 ;
  assign w10132 = ( ~w258 & w456 ) | ( ~w258 & w10131 ) | ( w456 & w10131 ) ;
  assign w10133 = w258 | w10132 ;
  assign w10134 = ( w208 & w255 ) | ( w208 & ~w722 ) | ( w255 & ~w722 ) ;
  assign w10135 = w202 | w10133 ;
  assign w10136 = ( ~w202 & w722 ) | ( ~w202 & w951 ) | ( w722 & w951 ) ;
  assign w10137 = w10135 | w10136 ;
  assign w10138 = w10134 | w10137 ;
  assign w10139 = w316 | w5626 ;
  assign w10140 = ( w209 & w564 ) | ( w209 & ~w5626 ) | ( w564 & ~w5626 ) ;
  assign w10141 = w10139 | w10140 ;
  assign w10142 = w264 | w2253 ;
  assign w10143 = ( ~w264 & w988 ) | ( ~w264 & w10141 ) | ( w988 & w10141 ) ;
  assign w10144 = w10142 | w10143 ;
  assign w10145 = ( w180 & w530 ) | ( w180 & ~w681 ) | ( w530 & ~w681 ) ;
  assign w10146 = w1275 | w10144 ;
  assign w10147 = ( w681 & w1130 ) | ( w681 & ~w1275 ) | ( w1130 & ~w1275 ) ;
  assign w10148 = w10146 | w10147 ;
  assign w10149 = w10145 | w10148 ;
  assign w10150 = ( w445 & w459 ) | ( w445 & ~w674 ) | ( w459 & ~w674 ) ;
  assign w10151 = w92 | w120 ;
  assign w10152 = ( ~w120 & w674 ) | ( ~w120 & w1086 ) | ( w674 & w1086 ) ;
  assign w10153 = w10151 | w10152 ;
  assign w10154 = w10150 | w10153 ;
  assign w10155 = ( w393 & ~w506 ) | ( w393 & w10154 ) | ( ~w506 & w10154 ) ;
  assign w10156 = w1564 | w10149 ;
  assign w10157 = ( w506 & w605 ) | ( w506 & ~w1564 ) | ( w605 & ~w1564 ) ;
  assign w10158 = w10156 | w10157 ;
  assign w10159 = w10155 | w10158 ;
  assign w10160 = ( w164 & w177 ) | ( w164 & ~w218 ) | ( w177 & ~w218 ) ;
  assign w10161 = w4793 | w10159 ;
  assign w10162 = ( w218 & w232 ) | ( w218 & ~w4793 ) | ( w232 & ~w4793 ) ;
  assign w10163 = w10161 | w10162 ;
  assign w10164 = w10160 | w10163 ;
  assign w10165 = ( w221 & w269 ) | ( w221 & ~w284 ) | ( w269 & ~w284 ) ;
  assign w10166 = w88 | w10164 ;
  assign w10167 = ( ~w88 & w284 ) | ( ~w88 & w392 ) | ( w284 & w392 ) ;
  assign w10168 = w10166 | w10167 ;
  assign w10169 = w10165 | w10168 ;
  assign w10170 = w253 | w516 ;
  assign w10171 = ( ~w253 & w423 ) | ( ~w253 & w10169 ) | ( w423 & w10169 ) ;
  assign w10172 = w10170 | w10171 ;
  assign w10173 = ( w229 & ~w317 ) | ( w229 & w429 ) | ( ~w317 & w429 ) ;
  assign w10174 = w317 | w10173 ;
  assign w10175 = ( w268 & w277 ) | ( w268 & ~w385 ) | ( w277 & ~w385 ) ;
  assign w10176 = w10172 | w10174 ;
  assign w10177 = ( w385 & w431 ) | ( w385 & ~w10174 ) | ( w431 & ~w10174 ) ;
  assign w10178 = w10176 | w10177 ;
  assign w10179 = w10175 | w10178 ;
  assign w10180 = w1513 | w1712 ;
  assign w10181 = w10138 | w10180 ;
  assign w10182 = ( w129 & ~w10138 ) | ( w129 & w10179 ) | ( ~w10138 & w10179 ) ;
  assign w10183 = w10181 | w10182 ;
  assign w10184 = ( w165 & w266 ) | ( w165 & ~w447 ) | ( w266 & ~w447 ) ;
  assign w10185 = w572 | w10183 ;
  assign w10186 = ( w447 & w470 ) | ( w447 & ~w572 ) | ( w470 & ~w572 ) ;
  assign w10187 = w10185 | w10186 ;
  assign w10188 = w10184 | w10187 ;
  assign w10189 = ( ~w10096 & w10126 ) | ( ~w10096 & w10188 ) | ( w10126 & w10188 ) ;
  assign w10190 = w10096 ^ w10126 ;
  assign w10191 = w10188 ^ w10190 ;
  assign w10192 = ( w9926 & w10069 ) | ( w9926 & ~w10096 ) | ( w10069 & ~w10096 ) ;
  assign w10193 = ( w10098 & w10099 ) | ( w10098 & ~w10107 ) | ( w10099 & ~w10107 ) ;
  assign w10194 = w10191 ^ w10193 ;
  assign w10195 = w10192 ^ w10194 ;
  assign w10196 = w4052 & ~w4600 ;
  assign w10197 = w4147 | w10196 ;
  assign w10198 = ( ~w4603 & w10196 ) | ( ~w4603 & w10197 ) | ( w10196 & w10197 ) ;
  assign w10199 = \pi26 ^ w10198 ;
  assign w10200 = w3649 | w4049 ;
  assign w10201 = w3717 & ~w4142 ;
  assign w10202 = ( ~w4049 & w10200 ) | ( ~w4049 & w10201 ) | ( w10200 & w10201 ) ;
  assign w10203 = w3549 | w3962 ;
  assign w10204 = w4152 & ~w10202 ;
  assign w10205 = ( w3448 & w10202 ) | ( w3448 & ~w10204 ) | ( w10202 & ~w10204 ) ;
  assign w10206 = ( ~w3962 & w10203 ) | ( ~w3962 & w10205 ) | ( w10203 & w10205 ) ;
  assign w10207 = \pi29 ^ w10206 ;
  assign w10208 = w10195 ^ w10199 ;
  assign w10209 = w10207 ^ w10208 ;
  assign w10210 = w10115 ^ w10209 ;
  assign w10211 = w10117 ^ w10210 ;
  assign w10212 = ( ~w9953 & w10048 ) | ( ~w9953 & w10114 ) | ( w10048 & w10114 ) ;
  assign w10213 = w10048 ^ w10212 ;
  assign w10214 = w10211 ^ w10213 ;
  assign w10215 = ( \pi29 & \pi31 ) | ( \pi29 & w10114 ) | ( \pi31 & w10114 ) ;
  assign w10216 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10215 ) | ( ~\pi30 & w10215 ) ;
  assign w10217 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10215 ) | ( \pi30 & w10215 ) ;
  assign w10218 = ( ~\pi29 & w9953 ) | ( ~\pi29 & w10217 ) | ( w9953 & w10217 ) ;
  assign w10219 = ( w10211 & w10217 ) | ( w10211 & ~w10218 ) | ( w10217 & ~w10218 ) ;
  assign w10220 = ~\pi31 & w10219 ;
  assign w10221 = ( w10216 & w10218 ) | ( w10216 & w10220 ) | ( w10218 & w10220 ) ;
  assign w10222 = ( w37 & w10214 ) | ( w37 & w10221 ) | ( w10214 & w10221 ) ;
  assign w10223 = w10221 | w10222 ;
  assign w10224 = ( w164 & ~w258 ) | ( w164 & w674 ) | ( ~w258 & w674 ) ;
  assign w10225 = w258 | w10224 ;
  assign w10226 = ( w386 & w415 ) | ( w386 & ~w449 ) | ( w415 & ~w449 ) ;
  assign w10227 = w101 | w10225 ;
  assign w10228 = ( ~w101 & w449 ) | ( ~w101 & w1126 ) | ( w449 & w1126 ) ;
  assign w10229 = w10227 | w10228 ;
  assign w10230 = w10226 | w10229 ;
  assign w10231 = w206 | w287 ;
  assign w10232 = ( w205 & ~w206 ) | ( w205 & w254 ) | ( ~w206 & w254 ) ;
  assign w10233 = w10231 | w10232 ;
  assign w10234 = w637 | w1030 ;
  assign w10235 = w420 | w10234 ;
  assign w10236 = ( w256 & ~w420 ) | ( w256 & w491 ) | ( ~w420 & w491 ) ;
  assign w10237 = w10235 | w10236 ;
  assign w10238 = ( w125 & w10233 ) | ( w125 & ~w10237 ) | ( w10233 & ~w10237 ) ;
  assign w10239 = w10237 | w10238 ;
  assign w10240 = ( w320 & w392 ) | ( w320 & ~w897 ) | ( w392 & ~w897 ) ;
  assign w10241 = w161 | w10239 ;
  assign w10242 = ( ~w161 & w897 ) | ( ~w161 & w1130 ) | ( w897 & w1130 ) ;
  assign w10243 = w10241 | w10242 ;
  assign w10244 = w10240 | w10243 ;
  assign w10245 = ( w275 & w569 ) | ( w275 & ~w605 ) | ( w569 & ~w605 ) ;
  assign w10246 = w218 | w2170 ;
  assign w10247 = ( ~w218 & w605 ) | ( ~w218 & w837 ) | ( w605 & w837 ) ;
  assign w10248 = w10246 | w10247 ;
  assign w10249 = w10245 | w10248 ;
  assign w10250 = w76 | w220 ;
  assign w10251 = w2060 | w10250 ;
  assign w10252 = ( w1836 & ~w2060 ) | ( w1836 & w6142 ) | ( ~w2060 & w6142 ) ;
  assign w10253 = w10251 | w10252 ;
  assign w10254 = w311 | w385 ;
  assign w10255 = w51 | w10254 ;
  assign w10256 = ( ~w51 & w116 ) | ( ~w51 & w10253 ) | ( w116 & w10253 ) ;
  assign w10257 = w10255 | w10256 ;
  assign w10258 = ( w505 & ~w641 ) | ( w505 & w2518 ) | ( ~w641 & w2518 ) ;
  assign w10259 = w999 | w10257 ;
  assign w10260 = ( w641 & ~w999 ) | ( w641 & w1094 ) | ( ~w999 & w1094 ) ;
  assign w10261 = w10259 | w10260 ;
  assign w10262 = w10258 | w10261 ;
  assign w10263 = ( w104 & ~w345 ) | ( w104 & w2556 ) | ( ~w345 & w2556 ) ;
  assign w10264 = w10249 | w10262 ;
  assign w10265 = ( w345 & w901 ) | ( w345 & ~w10249 ) | ( w901 & ~w10249 ) ;
  assign w10266 = w10264 | w10265 ;
  assign w10267 = w10263 | w10266 ;
  assign w10268 = ( w143 & w342 ) | ( w143 & ~w568 ) | ( w342 & ~w568 ) ;
  assign w10269 = w360 & ~w1265 ;
  assign w10270 = ( w568 & w1031 ) | ( w568 & ~w1265 ) | ( w1031 & ~w1265 ) ;
  assign w10271 = w10269 & ~w10270 ;
  assign w10272 = ~w10268 & w10271 ;
  assign w10273 = w573 | w640 ;
  assign w10274 = w167 | w10273 ;
  assign w10275 = ( ~w167 & w227 ) | ( ~w167 & w2319 ) | ( w227 & w2319 ) ;
  assign w10276 = w10274 | w10275 ;
  assign w10277 = ( w352 & w10272 ) | ( w352 & ~w10276 ) | ( w10272 & ~w10276 ) ;
  assign w10278 = w2750 | w10267 ;
  assign w10279 = ( w352 & w697 ) | ( w352 & ~w10267 ) | ( w697 & ~w10267 ) ;
  assign w10280 = w10278 | w10279 ;
  assign w10281 = w10277 & ~w10280 ;
  assign w10282 = w1155 | w4381 ;
  assign w10283 = w10244 | w10282 ;
  assign w10284 = ( ~w10230 & w10244 ) | ( ~w10230 & w10281 ) | ( w10244 & w10281 ) ;
  assign w10285 = ~w10283 & w10284 ;
  assign w10286 = w274 | w314 ;
  assign w10287 = w56 | w10286 ;
  assign w10288 = ( w56 & ~w230 ) | ( w56 & w10285 ) | ( ~w230 & w10285 ) ;
  assign w10289 = ~w10287 & w10288 ;
  assign w10290 = w219 | w2814 ;
  assign w10291 = ( w51 & w528 ) | ( w51 & ~w2814 ) | ( w528 & ~w2814 ) ;
  assign w10292 = w10290 | w10291 ;
  assign w10293 = ( ~w467 & w1283 ) | ( ~w467 & w1884 ) | ( w1283 & w1884 ) ;
  assign w10294 = w1987 | w10292 ;
  assign w10295 = ( w467 & w674 ) | ( w467 & ~w10292 ) | ( w674 & ~w10292 ) ;
  assign w10296 = w10294 | w10295 ;
  assign w10297 = w10293 | w10296 ;
  assign w10298 = w625 | w860 ;
  assign w10299 = w1185 | w10298 ;
  assign w10300 = ( w125 & ~w1185 ) | ( w125 & w10297 ) | ( ~w1185 & w10297 ) ;
  assign w10301 = w10299 | w10300 ;
  assign w10302 = ( w316 & w384 ) | ( w316 & ~w640 ) | ( w384 & ~w640 ) ;
  assign w10303 = w202 | w10301 ;
  assign w10304 = ( ~w202 & w640 ) | ( ~w202 & w1001 ) | ( w640 & w1001 ) ;
  assign w10305 = w10303 | w10304 ;
  assign w10306 = w10302 | w10305 ;
  assign w10307 = w420 | w458 ;
  assign w10308 = w208 | w10307 ;
  assign w10309 = ( w163 & ~w208 ) | ( w163 & w263 ) | ( ~w208 & w263 ) ;
  assign w10310 = w10308 | w10309 ;
  assign w10311 = ( w272 & w325 ) | ( w272 & ~w509 ) | ( w325 & ~w509 ) ;
  assign w10312 = w167 | w10310 ;
  assign w10313 = ( ~w167 & w509 ) | ( ~w167 & w899 ) | ( w509 & w899 ) ;
  assign w10314 = w10312 | w10313 ;
  assign w10315 = w10311 | w10314 ;
  assign w10316 = w1242 | w10315 ;
  assign w10317 = w10306 | w10316 ;
  assign w10318 = ( ~w2035 & w5180 ) | ( ~w2035 & w10306 ) | ( w5180 & w10306 ) ;
  assign w10319 = ~w10317 & w10318 ;
  assign w10320 = w1560 | w2760 ;
  assign w10321 = ( w1560 & ~w1882 ) | ( w1560 & w10319 ) | ( ~w1882 & w10319 ) ;
  assign w10322 = ~w10320 & w10321 ;
  assign w10323 = ( w220 & w224 ) | ( w220 & ~w342 ) | ( w224 & ~w342 ) ;
  assign w10324 = ~w1281 & w10322 ;
  assign w10325 = ( w342 & w495 ) | ( w342 & ~w1281 ) | ( w495 & ~w1281 ) ;
  assign w10326 = w10324 & ~w10325 ;
  assign w10327 = ~w10323 & w10326 ;
  assign w10328 = ( w135 & w215 ) | ( w135 & ~w362 ) | ( w215 & ~w362 ) ;
  assign w10329 = ~w114 & w10327 ;
  assign w10330 = ( ~w114 & w362 ) | ( ~w114 & w568 ) | ( w362 & w568 ) ;
  assign w10331 = w10329 & ~w10330 ;
  assign w10332 = ~w10328 & w10331 ;
  assign w10333 = w10048 ^ w10114 ;
  assign w10334 = w9953 ^ w10333 ;
  assign w10335 = ( \pi29 & \pi31 ) | ( \pi29 & w9953 ) | ( \pi31 & w9953 ) ;
  assign w10336 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10335 ) | ( ~\pi30 & w10335 ) ;
  assign w10337 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10335 ) | ( \pi30 & w10335 ) ;
  assign w10338 = ( ~\pi29 & w9842 ) | ( ~\pi29 & w10337 ) | ( w9842 & w10337 ) ;
  assign w10339 = ( w10114 & w10337 ) | ( w10114 & ~w10338 ) | ( w10337 & ~w10338 ) ;
  assign w10340 = ~\pi31 & w10339 ;
  assign w10341 = ( w10336 & w10338 ) | ( w10336 & w10340 ) | ( w10338 & w10340 ) ;
  assign w10342 = ( w37 & w10334 ) | ( w37 & w10341 ) | ( w10334 & w10341 ) ;
  assign w10343 = w10341 | w10342 ;
  assign w10344 = ( w10289 & ~w10332 ) | ( w10289 & w10343 ) | ( ~w10332 & w10343 ) ;
  assign w10345 = w86 | w513 ;
  assign w10346 = ( ~w86 & w141 ) | ( ~w86 & w216 ) | ( w141 & w216 ) ;
  assign w10347 = w10345 | w10346 ;
  assign w10348 = ( w411 & w492 ) | ( w411 & ~w697 ) | ( w492 & ~w697 ) ;
  assign w10349 = w310 | w340 ;
  assign w10350 = ( ~w340 & w697 ) | ( ~w340 & w860 ) | ( w697 & w860 ) ;
  assign w10351 = w10349 | w10350 ;
  assign w10352 = w10348 | w10351 ;
  assign w10353 = ( ~w104 & w10347 ) | ( ~w104 & w10352 ) | ( w10347 & w10352 ) ;
  assign w10354 = w1548 | w10138 ;
  assign w10355 = ( w104 & w281 ) | ( w104 & ~w1548 ) | ( w281 & ~w1548 ) ;
  assign w10356 = w10354 | w10355 ;
  assign w10357 = w10353 | w10356 ;
  assign w10358 = ( w1276 & w1884 ) | ( w1276 & ~w2625 ) | ( w1884 & ~w2625 ) ;
  assign w10359 = w2922 | w10357 ;
  assign w10360 = ( w283 & w2625 ) | ( w283 & ~w2922 ) | ( w2625 & ~w2922 ) ;
  assign w10361 = w10359 | w10360 ;
  assign w10362 = w10358 | w10361 ;
  assign w10363 = ( w81 & w260 ) | ( w81 & ~w430 ) | ( w260 & ~w430 ) ;
  assign w10364 = w56 | w10362 ;
  assign w10365 = ( ~w56 & w430 ) | ( ~w56 & w504 ) | ( w430 & w504 ) ;
  assign w10366 = w10364 | w10365 ;
  assign w10367 = w10363 | w10366 ;
  assign w10368 = ( ~w98 & w352 ) | ( ~w98 & w4232 ) | ( w352 & w4232 ) ;
  assign w10369 = w98 | w10368 ;
  assign w10370 = w421 | w490 ;
  assign w10371 = w169 | w10370 ;
  assign w10372 = ( ~w169 & w322 ) | ( ~w169 & w10369 ) | ( w322 & w10369 ) ;
  assign w10373 = w10371 | w10372 ;
  assign w10374 = ( w409 & w525 ) | ( w409 & ~w596 ) | ( w525 & ~w596 ) ;
  assign w10375 = w136 | w10373 ;
  assign w10376 = ( ~w136 & w596 ) | ( ~w136 & w663 ) | ( w596 & w663 ) ;
  assign w10377 = w10375 | w10376 ;
  assign w10378 = w10374 | w10377 ;
  assign w10379 = ( ~w275 & w680 ) | ( ~w275 & w10378 ) | ( w680 & w10378 ) ;
  assign w10380 = w275 | w10379 ;
  assign w10381 = ( w345 & w422 ) | ( w345 & ~w515 ) | ( w422 & ~w515 ) ;
  assign w10382 = w205 | w2090 ;
  assign w10383 = ( ~w205 & w515 ) | ( ~w205 & w595 ) | ( w515 & w595 ) ;
  assign w10384 = w10382 | w10383 ;
  assign w10385 = w10381 | w10384 ;
  assign w10386 = ( w1559 & ~w6241 ) | ( w1559 & w10380 ) | ( ~w6241 & w10380 ) ;
  assign w10387 = w10172 | w10367 ;
  assign w10388 = ( w6241 & ~w10172 ) | ( w6241 & w10385 ) | ( ~w10172 & w10385 ) ;
  assign w10389 = w10387 | w10388 ;
  assign w10390 = w10386 | w10389 ;
  assign w10391 = ( ~w224 & w1051 ) | ( ~w224 & w1165 ) | ( w1051 & w1165 ) ;
  assign w10392 = w273 | w10390 ;
  assign w10393 = ( w224 & ~w273 ) | ( w224 & w413 ) | ( ~w273 & w413 ) ;
  assign w10394 = w10392 | w10393 ;
  assign w10395 = w10391 | w10394 ;
  assign w10396 = w1128 | w1153 ;
  assign w10397 = w326 | w10396 ;
  assign w10398 = ( ~w326 & w1421 ) | ( ~w326 & w10395 ) | ( w1421 & w10395 ) ;
  assign w10399 = w10397 | w10398 ;
  assign w10400 = w168 | w3923 ;
  assign w10401 = ( ~w168 & w447 ) | ( ~w168 & w10399 ) | ( w447 & w10399 ) ;
  assign w10402 = w10400 | w10401 ;
  assign w10403 = ( w226 & w443 ) | ( w226 & ~w593 ) | ( w443 & ~w593 ) ;
  assign w10404 = w63 | w1835 ;
  assign w10405 = ( ~w63 & w593 ) | ( ~w63 & w4073 ) | ( w593 & w4073 ) ;
  assign w10406 = w10404 | w10405 ;
  assign w10407 = w10403 | w10406 ;
  assign w10408 = ( ~w131 & w759 ) | ( ~w131 & w998 ) | ( w759 & w998 ) ;
  assign w10409 = w177 | w3690 ;
  assign w10410 = ( w131 & ~w177 ) | ( w131 & w680 ) | ( ~w177 & w680 ) ;
  assign w10411 = w10409 | w10410 ;
  assign w10412 = w10408 | w10411 ;
  assign w10413 = ( w3937 & ~w4586 ) | ( w3937 & w5191 ) | ( ~w4586 & w5191 ) ;
  assign w10414 = w4110 & ~w10412 ;
  assign w10415 = ( w4586 & w10407 ) | ( w4586 & ~w10412 ) | ( w10407 & ~w10412 ) ;
  assign w10416 = w10414 & ~w10415 ;
  assign w10417 = ~w10413 & w10416 ;
  assign w10418 = w220 | w515 ;
  assign w10419 = w2705 | w10418 ;
  assign w10420 = ( w2705 & ~w2872 ) | ( w2705 & w10417 ) | ( ~w2872 & w10417 ) ;
  assign w10421 = ~w10419 & w10420 ;
  assign w10422 = ( w759 & ~w998 ) | ( w759 & w3677 ) | ( ~w998 & w3677 ) ;
  assign w10423 = w998 | w10422 ;
  assign w10424 = w980 | w3953 ;
  assign w10425 = w10423 | w10424 ;
  assign w10426 = ( ~w280 & w4130 ) | ( ~w280 & w10423 ) | ( w4130 & w10423 ) ;
  assign w10427 = ~w10425 & w10426 ;
  assign w10428 = w312 | w569 ;
  assign w10429 = ( w312 & ~w533 ) | ( w312 & w10427 ) | ( ~w533 & w10427 ) ;
  assign w10430 = ~w10428 & w10429 ;
  assign w10431 = w10421 & w10430 ;
  assign w10432 = ~w43 & w62 ;
  assign w10433 = ( ~\pi23 & \pi24 ) | ( ~\pi23 & w43 ) | ( \pi24 & w43 ) ;
  assign w10434 = ( ~\pi24 & \pi25 ) | ( ~\pi24 & w10433 ) | ( \pi25 & w10433 ) ;
  assign w10435 = ( \pi25 & w10432 ) | ( \pi25 & ~w10434 ) | ( w10432 & ~w10434 ) ;
  assign w10436 = \pi26 ^ w62 ;
  assign w10437 = ( ~\pi23 & w62 ) | ( ~\pi23 & w10436 ) | ( w62 & w10436 ) ;
  assign w10438 = ( \pi24 & \pi26 ) | ( \pi24 & ~w10437 ) | ( \pi26 & ~w10437 ) ;
  assign w10439 = \pi25 | w10438 ;
  assign w10440 = \pi26 ^ w10439 ;
  assign w10441 = ~w10435 & w10440 ;
  assign w10442 = w359 & ~w10441 ;
  assign w10443 = ( w359 & w443 ) | ( w359 & w1514 ) | ( w443 & w1514 ) ;
  assign w10444 = w10442 & ~w10443 ;
  assign w10445 = ~w4573 & w10444 ;
  assign w10446 = ( w672 & w3945 ) | ( w672 & w10444 ) | ( w3945 & w10444 ) ;
  assign w10447 = w10445 & ~w10446 ;
  assign w10448 = w605 | w681 ;
  assign w10449 = w1814 | w10448 ;
  assign w10450 = ( ~w63 & w1814 ) | ( ~w63 & w10447 ) | ( w1814 & w10447 ) ;
  assign w10451 = ~w10449 & w10450 ;
  assign w10452 = w3098 & ~w4600 ;
  assign w10453 = ( w37 & ~w4603 ) | ( w37 & w10452 ) | ( ~w4603 & w10452 ) ;
  assign w10454 = w10452 | w10453 ;
  assign w10455 = ( w10421 & ~w10451 ) | ( w10421 & w10454 ) | ( ~w10451 & w10454 ) ;
  assign w10456 = w10421 ^ w10430 ;
  assign w10457 = w10421 ^ w10451 ;
  assign w10458 = w37 & w4603 ;
  assign w10459 = ( w37 & w10452 ) | ( w37 & ~w10458 ) | ( w10452 & ~w10458 ) ;
  assign w10460 = w10457 ^ w10459 ;
  assign w10461 = w1229 | w1340 ;
  assign w10462 = w265 | w10461 ;
  assign w10463 = ( w226 & ~w265 ) | ( w226 & w390 ) | ( ~w265 & w390 ) ;
  assign w10464 = w10462 | w10463 ;
  assign w10465 = ( w286 & w386 ) | ( w286 & ~w393 ) | ( w386 & ~w393 ) ;
  assign w10466 = w1978 | w10464 ;
  assign w10467 = ( w393 & w424 ) | ( w393 & ~w10464 ) | ( w424 & ~w10464 ) ;
  assign w10468 = w10466 | w10467 ;
  assign w10469 = w10465 | w10468 ;
  assign w10470 = w275 | w516 ;
  assign w10471 = w92 | w10470 ;
  assign w10472 = ( ~w92 & w224 ) | ( ~w92 & w10469 ) | ( w224 & w10469 ) ;
  assign w10473 = w10471 | w10472 ;
  assign w10474 = w422 | w2704 ;
  assign w10475 = ( w528 & ~w2704 ) | ( w528 & w2873 ) | ( ~w2704 & w2873 ) ;
  assign w10476 = w10474 | w10475 ;
  assign w10477 = ( w203 & w209 ) | ( w203 & ~w271 ) | ( w209 & ~w271 ) ;
  assign w10478 = w118 | w10476 ;
  assign w10479 = ( ~w118 & w271 ) | ( ~w118 & w490 ) | ( w271 & w490 ) ;
  assign w10480 = w10478 | w10479 ;
  assign w10481 = w10477 | w10480 ;
  assign w10482 = ( w127 & w496 ) | ( w127 & ~w628 ) | ( w496 & ~w628 ) ;
  assign w10483 = w51 | w10481 ;
  assign w10484 = ( ~w51 & w628 ) | ( ~w51 & w783 ) | ( w628 & w783 ) ;
  assign w10485 = w10483 | w10484 ;
  assign w10486 = w10482 | w10485 ;
  assign w10487 = w128 | w138 ;
  assign w10488 = ( ~w128 & w136 ) | ( ~w128 & w10486 ) | ( w136 & w10486 ) ;
  assign w10489 = w10487 | w10488 ;
  assign w10490 = ( w263 & w389 ) | ( w263 & ~w596 ) | ( w389 & ~w596 ) ;
  assign w10491 = w1185 | w10489 ;
  assign w10492 = ( w596 & w724 ) | ( w596 & ~w1185 ) | ( w724 & ~w1185 ) ;
  assign w10493 = w10491 | w10492 ;
  assign w10494 = w10490 | w10493 ;
  assign w10495 = w1787 | w10494 ;
  assign w10496 = ( w1400 & ~w2762 ) | ( w1400 & w10473 ) | ( ~w2762 & w10473 ) ;
  assign w10497 = w1228 & ~w10495 ;
  assign w10498 = ( w2762 & w5039 ) | ( w2762 & ~w10495 ) | ( w5039 & ~w10495 ) ;
  assign w10499 = w10497 & ~w10498 ;
  assign w10500 = ~w10496 & w10499 ;
  assign w10501 = w232 | w623 ;
  assign w10502 = w741 | w10501 ;
  assign w10503 = ( w741 & ~w1281 ) | ( w741 & w10500 ) | ( ~w1281 & w10500 ) ;
  assign w10504 = ~w10502 & w10503 ;
  assign w10505 = ( w90 & w266 ) | ( w90 & ~w353 ) | ( w266 & ~w353 ) ;
  assign w10506 = ~w998 & w10504 ;
  assign w10507 = ( w353 & w860 ) | ( w353 & ~w998 ) | ( w860 & ~w998 ) ;
  assign w10508 = w10506 & ~w10507 ;
  assign w10509 = ~w10505 & w10508 ;
  assign w10510 = w524 | w680 ;
  assign w10511 = w256 | w10510 ;
  assign w10512 = ( w256 & ~w274 ) | ( w256 & w10509 ) | ( ~w274 & w10509 ) ;
  assign w10513 = ~w10511 & w10512 ;
  assign w10514 = w202 | w726 ;
  assign w10515 = w900 | w10514 ;
  assign w10516 = ( w113 & ~w900 ) | ( w113 & w4015 ) | ( ~w900 & w4015 ) ;
  assign w10517 = w10515 | w10516 ;
  assign w10518 = ( w227 & w495 ) | ( w227 & ~w625 ) | ( w495 & ~w625 ) ;
  assign w10519 = w86 | w167 ;
  assign w10520 = ( ~w167 & w625 ) | ( ~w167 & w783 ) | ( w625 & w783 ) ;
  assign w10521 = w10519 | w10520 ;
  assign w10522 = w10518 | w10521 ;
  assign w10523 = w4032 | w10441 ;
  assign w10524 = w10407 | w10523 ;
  assign w10525 = ( ~w10407 & w10517 ) | ( ~w10407 & w10522 ) | ( w10517 & w10522 ) ;
  assign w10526 = w10524 | w10525 ;
  assign w10527 = ( w275 & w524 ) | ( w275 & ~w569 ) | ( w524 & ~w569 ) ;
  assign w10528 = w1069 | w10526 ;
  assign w10529 = ( w569 & ~w1069 ) | ( w569 & w4101 ) | ( ~w1069 & w4101 ) ;
  assign w10530 = w10528 | w10529 ;
  assign w10531 = w10527 | w10530 ;
  assign w10532 = ( \pi29 & w10513 ) | ( \pi29 & ~w10531 ) | ( w10513 & ~w10531 ) ;
  assign w10533 = w3962 ^ w6862 ;
  assign w10534 = ( ~w3962 & w4600 ) | ( ~w3962 & w10533 ) | ( w4600 & w10533 ) ;
  assign w10535 = ( w4601 & w10533 ) | ( w4601 & w10534 ) | ( w10533 & w10534 ) ;
  assign w10536 = ( \pi29 & \pi30 ) | ( \pi29 & ~w10535 ) | ( \pi30 & ~w10535 ) ;
  assign w10537 = w10534 ^ w10536 ;
  assign w10538 = \pi30 & ~w4600 ;
  assign w10539 = \pi29 & w10538 ;
  assign w10540 = \pi31 ^ w10539 ;
  assign w10541 = ( ~w10537 & w10539 ) | ( ~w10537 & w10540 ) | ( w10539 & w10540 ) ;
  assign w10542 = ( w10421 & ~w10532 ) | ( w10421 & w10541 ) | ( ~w10532 & w10541 ) ;
  assign w10543 = w10532 ^ w10541 ;
  assign w10544 = w10421 ^ w10543 ;
  assign w10545 = w10513 ^ w10531 ;
  assign w10546 = \pi29 ^ w10545 ;
  assign w10547 = ( w385 & w421 ) | ( w385 & ~w447 ) | ( w421 & ~w447 ) ;
  assign w10548 = w351 | w1164 ;
  assign w10549 = ( ~w351 & w447 ) | ( ~w351 & w488 ) | ( w447 & w488 ) ;
  assign w10550 = w10548 | w10549 ;
  assign w10551 = w10547 | w10550 ;
  assign w10552 = w147 | w205 ;
  assign w10553 = w270 | w10552 ;
  assign w10554 = ( ~w270 & w468 ) | ( ~w270 & w10551 ) | ( w468 & w10551 ) ;
  assign w10555 = w10553 | w10554 ;
  assign w10556 = w1064 | w4353 ;
  assign w10557 = ( w341 & ~w1064 ) | ( w341 & w10555 ) | ( ~w1064 & w10555 ) ;
  assign w10558 = w10556 | w10557 ;
  assign w10559 = ( w316 & w463 ) | ( w316 & ~w505 ) | ( w463 & ~w505 ) ;
  assign w10560 = w59 | w10558 ;
  assign w10561 = ( ~w59 & w505 ) | ( ~w59 & w980 ) | ( w505 & w980 ) ;
  assign w10562 = w10560 | w10561 ;
  assign w10563 = w10559 | w10562 ;
  assign w10564 = w253 | w413 ;
  assign w10565 = w86 | w10564 ;
  assign w10566 = ( ~w86 & w224 ) | ( ~w86 & w627 ) | ( w224 & w627 ) ;
  assign w10567 = w10565 | w10566 ;
  assign w10568 = ( w312 & w353 ) | ( w312 & ~w409 ) | ( w353 & ~w409 ) ;
  assign w10569 = w120 | w10567 ;
  assign w10570 = ( ~w120 & w409 ) | ( ~w120 & w723 ) | ( w409 & w723 ) ;
  assign w10571 = w10569 | w10570 ;
  assign w10572 = w10568 | w10571 ;
  assign w10573 = w175 | w662 ;
  assign w10574 = w56 | w10573 ;
  assign w10575 = ( ~w56 & w101 ) | ( ~w56 & w10572 ) | ( w101 & w10572 ) ;
  assign w10576 = w10574 | w10575 ;
  assign w10577 = w350 | w951 ;
  assign w10578 = ( ~w350 & w445 ) | ( ~w350 & w3196 ) | ( w445 & w3196 ) ;
  assign w10579 = w10577 | w10578 ;
  assign w10580 = w122 | w493 ;
  assign w10581 = ( w103 & ~w493 ) | ( w103 & w10579 ) | ( ~w493 & w10579 ) ;
  assign w10582 = w10580 | w10581 ;
  assign w10583 = ( w3067 & w10576 ) | ( w3067 & w10582 ) | ( w10576 & w10582 ) ;
  assign w10584 = w4311 | w10563 ;
  assign w10585 = ( w3067 & ~w6353 ) | ( w3067 & w10563 ) | ( ~w6353 & w10563 ) ;
  assign w10586 = ~w10584 & w10585 ;
  assign w10587 = ~w10583 & w10586 ;
  assign w10588 = w201 | w725 ;
  assign w10589 = w1283 | w10588 ;
  assign w10590 = ( w1283 & ~w1566 ) | ( w1283 & w10587 ) | ( ~w1566 & w10587 ) ;
  assign w10591 = ~w10589 & w10590 ;
  assign w10592 = ( w449 & w491 ) | ( w449 & ~w504 ) | ( w491 & ~w504 ) ;
  assign w10593 = ~w142 & w10591 ;
  assign w10594 = ( ~w142 & w504 ) | ( ~w142 & w570 ) | ( w504 & w570 ) ;
  assign w10595 = w10593 & ~w10594 ;
  assign w10596 = ~w10592 & w10595 ;
  assign w10597 = ( ~w1883 & w4796 ) | ( ~w1883 & w9884 ) | ( w4796 & w9884 ) ;
  assign w10598 = w1883 | w10597 ;
  assign w10599 = ( w113 & w309 ) | ( w113 & ~w339 ) | ( w309 & ~w339 ) ;
  assign w10600 = w410 | w10598 ;
  assign w10601 = ( w339 & ~w410 ) | ( w339 & w443 ) | ( ~w410 & w443 ) ;
  assign w10602 = w10600 | w10601 ;
  assign w10603 = w10599 | w10602 ;
  assign w10604 = ( w115 & w277 ) | ( w115 & ~w385 ) | ( w277 & ~w385 ) ;
  assign w10605 = ( ~w95 & w385 ) | ( ~w95 & w723 ) | ( w385 & w723 ) ;
  assign w10606 = w6144 | w10605 ;
  assign w10607 = w10604 | w10606 ;
  assign w10608 = ( w210 & w561 ) | ( w210 & ~w817 ) | ( w561 & ~w817 ) ;
  assign w10609 = w5837 | w10607 ;
  assign w10610 = ( w817 & w899 ) | ( w817 & ~w10607 ) | ( w899 & ~w10607 ) ;
  assign w10611 = w10609 | w10610 ;
  assign w10612 = w10608 | w10611 ;
  assign w10613 = w267 | w1882 ;
  assign w10614 = ( ~w267 & w1400 ) | ( ~w267 & w10612 ) | ( w1400 & w10612 ) ;
  assign w10615 = w10613 | w10614 ;
  assign w10616 = ( w269 & w490 ) | ( w269 & ~w1128 ) | ( w490 & ~w1128 ) ;
  assign w10617 = w214 | w10615 ;
  assign w10618 = ( ~w214 & w1128 ) | ( ~w214 & w1340 ) | ( w1128 & w1340 ) ;
  assign w10619 = w10617 | w10618 ;
  assign w10620 = w10616 | w10619 ;
  assign w10621 = w167 | w673 ;
  assign w10622 = ( ~w167 & w224 ) | ( ~w167 & w10620 ) | ( w224 & w10620 ) ;
  assign w10623 = w10621 | w10622 ;
  assign w10624 = w92 | w422 ;
  assign w10625 = ( ~w92 & w352 ) | ( ~w92 & w594 ) | ( w352 & w594 ) ;
  assign w10626 = w10624 | w10625 ;
  assign w10627 = w133 | w608 ;
  assign w10628 = w76 | w10627 ;
  assign w10629 = ( ~w76 & w101 ) | ( ~w76 & w4464 ) | ( w101 & w4464 ) ;
  assign w10630 = w10628 | w10629 ;
  assign w10631 = ( ~w253 & w10626 ) | ( ~w253 & w10630 ) | ( w10626 & w10630 ) ;
  assign w10632 = w2909 | w10623 ;
  assign w10633 = ( w253 & w459 ) | ( w253 & ~w10623 ) | ( w459 & ~w10623 ) ;
  assign w10634 = w10632 | w10633 ;
  assign w10635 = w10631 | w10634 ;
  assign w10636 = w2168 | w10603 ;
  assign w10637 = ( w1363 & ~w10603 ) | ( w1363 & w10635 ) | ( ~w10603 & w10635 ) ;
  assign w10638 = w10636 | w10637 ;
  assign w10639 = w259 | w260 ;
  assign w10640 = w126 | w10639 ;
  assign w10641 = ( ~w126 & w2518 ) | ( ~w126 & w10638 ) | ( w2518 & w10638 ) ;
  assign w10642 = w10640 | w10641 ;
  assign w10643 = w209 | w311 ;
  assign w10644 = w114 | w10643 ;
  assign w10645 = ( ~w114 & w136 ) | ( ~w114 & w10642 ) | ( w136 & w10642 ) ;
  assign w10646 = w10644 | w10645 ;
  assign w10647 = ( ~\pi26 & w10096 ) | ( ~\pi26 & w10646 ) | ( w10096 & w10646 ) ;
  assign w10648 = ( \pi30 & \pi31 ) | ( \pi30 & ~w4049 ) | ( \pi31 & ~w4049 ) ;
  assign w10649 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10648 ) | ( \pi30 & w10648 ) ;
  assign w10650 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10648 ) | ( ~\pi30 & w10648 ) ;
  assign w10651 = ( ~\pi30 & w3907 ) | ( ~\pi30 & w10650 ) | ( w3907 & w10650 ) ;
  assign w10652 = ( w4142 & ~w10650 ) | ( w4142 & w10651 ) | ( ~w10650 & w10651 ) ;
  assign w10653 = \pi31 | w10652 ;
  assign w10654 = ( w10649 & w10651 ) | ( w10649 & ~w10653 ) | ( w10651 & ~w10653 ) ;
  assign w10655 = ( w37 & w4563 ) | ( w37 & w10654 ) | ( w4563 & w10654 ) ;
  assign w10656 = w10654 | w10655 ;
  assign w10657 = ( w10596 & w10647 ) | ( w10596 & w10656 ) | ( w10647 & w10656 ) ;
  assign w10658 = ( w10513 & ~w10596 ) | ( w10513 & w10657 ) | ( ~w10596 & w10657 ) ;
  assign w10659 = ( \pi30 & \pi31 ) | ( \pi30 & ~w3962 ) | ( \pi31 & ~w3962 ) ;
  assign w10660 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10659 ) | ( \pi30 & w10659 ) ;
  assign w10661 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10659 ) | ( ~\pi30 & w10659 ) ;
  assign w10662 = ( \pi30 & w4142 ) | ( \pi30 & ~w10661 ) | ( w4142 & ~w10661 ) ;
  assign w10663 = ( ~w4600 & w10661 ) | ( ~w4600 & w10662 ) | ( w10661 & w10662 ) ;
  assign w10664 = ~\pi31 & w10663 ;
  assign w10665 = ( w10660 & ~w10662 ) | ( w10660 & w10664 ) | ( ~w10662 & w10664 ) ;
  assign w10666 = ( w37 & ~w4722 ) | ( w37 & w10665 ) | ( ~w4722 & w10665 ) ;
  assign w10667 = w10665 | w10666 ;
  assign w10668 = ( w10546 & w10658 ) | ( w10546 & w10667 ) | ( w10658 & w10667 ) ;
  assign w10669 = w3649 & ~w4600 ;
  assign w10670 = w3448 | w10669 ;
  assign w10671 = ( ~w4603 & w10669 ) | ( ~w4603 & w10670 ) | ( w10669 & w10670 ) ;
  assign w10672 = \pi29 ^ w10671 ;
  assign w10673 = ( \pi29 & \pi31 ) | ( \pi29 & ~w4142 ) | ( \pi31 & ~w4142 ) ;
  assign w10674 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10673 ) | ( ~\pi30 & w10673 ) ;
  assign w10675 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10673 ) | ( \pi30 & w10673 ) ;
  assign w10676 = ( \pi29 & w4049 ) | ( \pi29 & ~w10675 ) | ( w4049 & ~w10675 ) ;
  assign w10677 = ( ~w3962 & w10675 ) | ( ~w3962 & w10676 ) | ( w10675 & w10676 ) ;
  assign w10678 = ~\pi31 & w10677 ;
  assign w10679 = ( w10674 & ~w10676 ) | ( w10674 & w10678 ) | ( ~w10676 & w10678 ) ;
  assign w10680 = ( w37 & ~w4152 ) | ( w37 & w10679 ) | ( ~w4152 & w10679 ) ;
  assign w10681 = w10679 | w10680 ;
  assign w10682 = w10513 ^ w10657 ;
  assign w10683 = w10596 ^ w10682 ;
  assign w10684 = ( w10672 & w10681 ) | ( w10672 & ~w10683 ) | ( w10681 & ~w10683 ) ;
  assign w10685 = w10658 ^ w10667 ;
  assign w10686 = w10546 ^ w10685 ;
  assign w10687 = w10647 ^ w10656 ;
  assign w10688 = w10596 ^ w10687 ;
  assign w10689 = w10096 ^ w10646 ;
  assign w10690 = \pi26 ^ w10689 ;
  assign w10691 = ( \pi29 & \pi31 ) | ( \pi29 & w3907 ) | ( \pi31 & w3907 ) ;
  assign w10692 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10691 ) | ( ~\pi30 & w10691 ) ;
  assign w10693 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10691 ) | ( \pi30 & w10691 ) ;
  assign w10694 = ( \pi29 & w3548 ) | ( \pi29 & ~w10693 ) | ( w3548 & ~w10693 ) ;
  assign w10695 = ( ~w4049 & w10693 ) | ( ~w4049 & w10694 ) | ( w10693 & w10694 ) ;
  assign w10696 = ~\pi31 & w10695 ;
  assign w10697 = ( w10692 & ~w10694 ) | ( w10692 & w10696 ) | ( ~w10694 & w10696 ) ;
  assign w10698 = ( w37 & ~w4622 ) | ( w37 & w10697 ) | ( ~w4622 & w10697 ) ;
  assign w10699 = w10697 | w10698 ;
  assign w10700 = ( w10189 & ~w10690 ) | ( w10189 & w10699 ) | ( ~w10690 & w10699 ) ;
  assign w10701 = w10688 ^ w10700 ;
  assign w10702 = w3717 & ~w4600 ;
  assign w10703 = ( w3649 & ~w3962 ) | ( w3649 & w10702 ) | ( ~w3962 & w10702 ) ;
  assign w10704 = ( ~w3962 & w4601 ) | ( ~w3962 & w10703 ) | ( w4601 & w10703 ) ;
  assign w10705 = ( w3448 & w4600 ) | ( w3448 & w4601 ) | ( w4600 & w4601 ) ;
  assign w10706 = ( w10702 & ~w10704 ) | ( w10702 & w10705 ) | ( ~w10704 & w10705 ) ;
  assign w10707 = ( ~w4657 & w10703 ) | ( ~w4657 & w10706 ) | ( w10703 & w10706 ) ;
  assign w10708 = \pi29 ^ w10707 ;
  assign w10709 = ( w10688 & w10700 ) | ( w10688 & w10708 ) | ( w10700 & w10708 ) ;
  assign w10710 = w10672 ^ w10683 ;
  assign w10711 = w10681 ^ w10710 ;
  assign w10712 = ( w10191 & ~w10192 ) | ( w10191 & w10193 ) | ( ~w10192 & w10193 ) ;
  assign w10713 = w10189 ^ w10699 ;
  assign w10714 = w10690 ^ w10713 ;
  assign w10715 = w3717 | w3962 ;
  assign w10716 = w3649 & ~w4142 ;
  assign w10717 = ( ~w3962 & w10715 ) | ( ~w3962 & w10716 ) | ( w10715 & w10716 ) ;
  assign w10718 = w3549 | w4600 ;
  assign w10719 = w4722 & ~w10717 ;
  assign w10720 = ( w3448 & w10717 ) | ( w3448 & ~w10719 ) | ( w10717 & ~w10719 ) ;
  assign w10721 = ( ~w4600 & w10718 ) | ( ~w4600 & w10720 ) | ( w10718 & w10720 ) ;
  assign w10722 = \pi29 ^ w10721 ;
  assign w10723 = ( w10712 & w10714 ) | ( w10712 & ~w10722 ) | ( w10714 & ~w10722 ) ;
  assign w10724 = w10712 ^ w10722 ;
  assign w10725 = w10714 ^ w10724 ;
  assign w10726 = ( w10195 & w10199 ) | ( w10195 & w10207 ) | ( w10199 & w10207 ) ;
  assign w10727 = ( w10115 & w10117 ) | ( w10115 & w10209 ) | ( w10117 & w10209 ) ;
  assign w10728 = ( w10725 & w10726 ) | ( w10725 & w10727 ) | ( w10726 & w10727 ) ;
  assign w10729 = w10701 ^ w10707 ;
  assign w10730 = \pi29 ^ w10729 ;
  assign w10731 = ( ~w10723 & w10728 ) | ( ~w10723 & w10730 ) | ( w10728 & w10730 ) ;
  assign w10732 = ( w10709 & ~w10711 ) | ( w10709 & w10731 ) | ( ~w10711 & w10731 ) ;
  assign w10733 = ( w10684 & w10686 ) | ( w10684 & w10732 ) | ( w10686 & w10732 ) ;
  assign w10734 = ( ~w10544 & w10668 ) | ( ~w10544 & w10733 ) | ( w10668 & w10733 ) ;
  assign w10735 = ( ~w10460 & w10542 ) | ( ~w10460 & w10734 ) | ( w10542 & w10734 ) ;
  assign w10736 = ( w10455 & ~w10456 ) | ( w10455 & w10735 ) | ( ~w10456 & w10735 ) ;
  assign w10737 = ( w10402 & w10431 ) | ( w10402 & ~w10736 ) | ( w10431 & ~w10736 ) ;
  assign w10738 = w10402 & ~w10737 ;
  assign w10739 = ( \pi17 & \pi18 ) | ( \pi17 & ~\pi19 ) | ( \pi18 & ~\pi19 ) ;
  assign w10740 = ( \pi19 & ~\pi20 ) | ( \pi19 & w10739 ) | ( ~\pi20 & w10739 ) ;
  assign w10741 = w10738 ^ w10740 ;
  assign w10742 = ( \pi20 & w10740 ) | ( \pi20 & w10741 ) | ( w10740 & w10741 ) ;
  assign w10743 = ( w317 & w318 ) | ( w317 & ~w384 ) | ( w318 & ~w384 ) ;
  assign w10744 = w2715 | w3525 ;
  assign w10745 = ( w384 & w1086 ) | ( w384 & ~w3525 ) | ( w1086 & ~w3525 ) ;
  assign w10746 = w10744 | w10745 ;
  assign w10747 = w10743 | w10746 ;
  assign w10748 = w218 | w219 ;
  assign w10749 = w1273 | w10748 ;
  assign w10750 = ( ~w1273 & w1955 ) | ( ~w1273 & w10747 ) | ( w1955 & w10747 ) ;
  assign w10751 = w10749 | w10750 ;
  assign w10752 = w206 | w209 ;
  assign w10753 = w276 | w10752 ;
  assign w10754 = ( ~w276 & w1281 ) | ( ~w276 & w10751 ) | ( w1281 & w10751 ) ;
  assign w10755 = w10753 | w10754 ;
  assign w10756 = w266 | w722 ;
  assign w10757 = ( ~w266 & w565 ) | ( ~w266 & w10755 ) | ( w565 & w10755 ) ;
  assign w10758 = w10756 | w10757 ;
  assign w10759 = w230 | w1031 ;
  assign w10760 = w507 | w10759 ;
  assign w10761 = ( w114 & ~w507 ) | ( w114 & w2948 ) | ( ~w507 & w2948 ) ;
  assign w10762 = w10760 | w10761 ;
  assign w10763 = ( ~w495 & w1009 ) | ( ~w495 & w10762 ) | ( w1009 & w10762 ) ;
  assign w10764 = w1758 & ~w10758 ;
  assign w10765 = ( w495 & w513 ) | ( w495 & w1758 ) | ( w513 & w1758 ) ;
  assign w10766 = w10764 & ~w10765 ;
  assign w10767 = ~w10763 & w10766 ;
  assign w10768 = w201 | w221 ;
  assign w10769 = w444 | w10768 ;
  assign w10770 = ( w444 & ~w627 ) | ( w444 & w10767 ) | ( ~w627 & w10767 ) ;
  assign w10771 = ~w10769 & w10770 ;
  assign w10772 = ( w232 & w560 ) | ( w232 & ~w571 ) | ( w560 & ~w571 ) ;
  assign w10773 = ~w229 & w10771 ;
  assign w10774 = ( ~w229 & w571 ) | ( ~w229 & w897 ) | ( w571 & w897 ) ;
  assign w10775 = w10773 & ~w10774 ;
  assign w10776 = ~w10772 & w10775 ;
  assign w10777 = ( w783 & ~w889 ) | ( w783 & w10776 ) | ( ~w889 & w10776 ) ;
  assign w10778 = ~w783 & w10777 ;
  assign w10779 = w10289 ^ w10742 ;
  assign w10780 = w10778 ^ w10779 ;
  assign w10781 = ( w10223 & w10344 ) | ( w10223 & ~w10780 ) | ( w10344 & ~w10780 ) ;
  assign w10782 = ( w10289 & w10742 ) | ( w10289 & w10778 ) | ( w10742 & w10778 ) ;
  assign w10783 = w10725 ^ w10727 ;
  assign w10784 = w10726 ^ w10783 ;
  assign w10785 = ( w9953 & w10048 ) | ( w9953 & w10114 ) | ( w10048 & w10114 ) ;
  assign w10786 = ( w10114 & w10211 ) | ( w10114 & w10785 ) | ( w10211 & w10785 ) ;
  assign w10787 = ( w10211 & w10784 ) | ( w10211 & w10786 ) | ( w10784 & w10786 ) ;
  assign w10788 = w10784 ^ w10786 ;
  assign w10789 = w10211 ^ w10788 ;
  assign w10790 = ~w37 & w10789 ;
  assign w10791 = w3098 & w10114 ;
  assign w10792 = ( w10789 & ~w10790 ) | ( w10789 & w10791 ) | ( ~w10790 & w10791 ) ;
  assign w10793 = ( \pi29 & \pi30 ) | ( \pi29 & w10784 ) | ( \pi30 & w10784 ) ;
  assign w10794 = \pi31 | w10793 ;
  assign w10795 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10211 ) | ( ~\pi30 & w10211 ) ;
  assign w10796 = ( \pi29 & \pi31 ) | ( \pi29 & ~w10795 ) | ( \pi31 & ~w10795 ) ;
  assign w10797 = ( w10792 & w10794 ) | ( w10792 & ~w10796 ) | ( w10794 & ~w10796 ) ;
  assign w10798 = w10782 ^ w10797 ;
  assign w10799 = w10367 ^ w10798 ;
  assign w10800 = w10684 ^ w10732 ;
  assign w10801 = w10686 ^ w10800 ;
  assign w10802 = w10701 ^ w10723 ;
  assign w10803 = w10707 ^ w10728 ;
  assign w10804 = \pi29 ^ w10803 ;
  assign w10805 = w10802 ^ w10804 ;
  assign w10806 = w10711 ^ w10731 ;
  assign w10807 = w10709 ^ w10806 ;
  assign w10808 = w3717 | w10807 ;
  assign w10809 = w3649 & ~w10805 ;
  assign w10810 = ( ~w10807 & w10808 ) | ( ~w10807 & w10809 ) | ( w10808 & w10809 ) ;
  assign w10811 = ( w10784 & w10787 ) | ( w10784 & ~w10805 ) | ( w10787 & ~w10805 ) ;
  assign w10812 = ( w10805 & w10807 ) | ( w10805 & ~w10811 ) | ( w10807 & ~w10811 ) ;
  assign w10813 = w10801 ^ w10812 ;
  assign w10814 = w10807 ^ w10813 ;
  assign w10815 = ~w3549 & w10801 ;
  assign w10816 = w10810 | w10814 ;
  assign w10817 = ( w3448 & w10810 ) | ( w3448 & w10816 ) | ( w10810 & w10816 ) ;
  assign w10818 = ( w10801 & ~w10815 ) | ( w10801 & w10817 ) | ( ~w10815 & w10817 ) ;
  assign w10819 = \pi29 ^ w10818 ;
  assign w10820 = ( w10781 & w10799 ) | ( w10781 & w10819 ) | ( w10799 & w10819 ) ;
  assign w10821 = ( w10367 & w10782 ) | ( w10367 & ~w10797 ) | ( w10782 & ~w10797 ) ;
  assign w10822 = ( w285 & ~w362 ) | ( w285 & w3892 ) | ( ~w362 & w3892 ) ;
  assign w10823 = w1010 | w2480 ;
  assign w10824 = ( w362 & w511 ) | ( w362 & ~w2480 ) | ( w511 & ~w2480 ) ;
  assign w10825 = w10823 | w10824 ;
  assign w10826 = w10822 | w10825 ;
  assign w10827 = w389 | w899 ;
  assign w10828 = w267 | w10827 ;
  assign w10829 = ( w210 & ~w267 ) | ( w210 & w10826 ) | ( ~w267 & w10826 ) ;
  assign w10830 = w10828 | w10829 ;
  assign w10831 = ( w253 & w467 ) | ( w253 & ~w625 ) | ( w467 & ~w625 ) ;
  assign w10832 = w92 | w10830 ;
  assign w10833 = ( ~w92 & w625 ) | ( ~w92 & w1086 ) | ( w625 & w1086 ) ;
  assign w10834 = w10832 | w10833 ;
  assign w10835 = w10831 | w10834 ;
  assign w10836 = ( ~w203 & w5546 ) | ( ~w203 & w9860 ) | ( w5546 & w9860 ) ;
  assign w10837 = w3471 | w10267 ;
  assign w10838 = ( w203 & w1153 ) | ( w203 & ~w3471 ) | ( w1153 & ~w3471 ) ;
  assign w10839 = w10837 | w10838 ;
  assign w10840 = w10836 | w10839 ;
  assign w10841 = ( w911 & ~w2091 ) | ( w911 & w10835 ) | ( ~w2091 & w10835 ) ;
  assign w10842 = w4379 | w10840 ;
  assign w10843 = ( w2091 & w3965 ) | ( w2091 & ~w10840 ) | ( w3965 & ~w10840 ) ;
  assign w10844 = w10842 | w10843 ;
  assign w10845 = w10841 | w10844 ;
  assign w10846 = ( w268 & w354 ) | ( w268 & ~w567 ) | ( w354 & ~w567 ) ;
  assign w10847 = w147 | w10845 ;
  assign w10848 = ( ~w147 & w567 ) | ( ~w147 & w860 ) | ( w567 & w860 ) ;
  assign w10849 = w10847 | w10848 ;
  assign w10850 = w10846 | w10849 ;
  assign w10851 = ( ~w10367 & w10821 ) | ( ~w10367 & w10850 ) | ( w10821 & w10850 ) ;
  assign w10852 = w10367 ^ w10821 ;
  assign w10853 = w10850 ^ w10852 ;
  assign w10854 = w10787 ^ w10805 ;
  assign w10855 = w10784 ^ w10854 ;
  assign w10856 = ( \pi29 & \pi31 ) | ( \pi29 & w10784 ) | ( \pi31 & w10784 ) ;
  assign w10857 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10856 ) | ( ~\pi30 & w10856 ) ;
  assign w10858 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10856 ) | ( \pi30 & w10856 ) ;
  assign w10859 = ( ~\pi29 & w10211 ) | ( ~\pi29 & w10858 ) | ( w10211 & w10858 ) ;
  assign w10860 = ( w10805 & ~w10858 ) | ( w10805 & w10859 ) | ( ~w10858 & w10859 ) ;
  assign w10861 = \pi31 | w10860 ;
  assign w10862 = ( w10857 & w10859 ) | ( w10857 & ~w10861 ) | ( w10859 & ~w10861 ) ;
  assign w10863 = ( w37 & ~w10855 ) | ( w37 & w10862 ) | ( ~w10855 & w10862 ) ;
  assign w10864 = w10862 | w10863 ;
  assign w10865 = w10668 ^ w10733 ;
  assign w10866 = w10544 ^ w10865 ;
  assign w10867 = ~w3717 & w10801 ;
  assign w10868 = w3649 & ~w10807 ;
  assign w10869 = ( w10801 & ~w10867 ) | ( w10801 & w10868 ) | ( ~w10867 & w10868 ) ;
  assign w10870 = ( ~w10801 & w10812 ) | ( ~w10801 & w10866 ) | ( w10812 & w10866 ) ;
  assign w10871 = ( ~w10801 & w10807 ) | ( ~w10801 & w10870 ) | ( w10807 & w10870 ) ;
  assign w10872 = ( ~w10801 & w10807 ) | ( ~w10801 & w10812 ) | ( w10807 & w10812 ) ;
  assign w10873 = w10801 ^ w10872 ;
  assign w10874 = w10866 ^ w10873 ;
  assign w10875 = w3549 | w10866 ;
  assign w10876 = w10869 | w10874 ;
  assign w10877 = ( w3448 & w10869 ) | ( w3448 & w10876 ) | ( w10869 & w10876 ) ;
  assign w10878 = ( ~w10866 & w10875 ) | ( ~w10866 & w10877 ) | ( w10875 & w10877 ) ;
  assign w10879 = \pi29 ^ w10878 ;
  assign w10880 = w10853 ^ w10879 ;
  assign w10881 = w10864 ^ w10880 ;
  assign w10882 = w10402 ^ w10736 ;
  assign w10883 = w10431 ^ w10882 ;
  assign w10884 = w10460 ^ w10734 ;
  assign w10885 = w10542 ^ w10884 ;
  assign w10886 = w10455 ^ w10735 ;
  assign w10887 = w10456 ^ w10886 ;
  assign w10888 = w4143 | w10887 ;
  assign w10889 = w4052 & ~w10885 ;
  assign w10890 = ( ~w10887 & w10888 ) | ( ~w10887 & w10889 ) | ( w10888 & w10889 ) ;
  assign w10891 = ( w10866 & w10871 ) | ( w10866 & w10885 ) | ( w10871 & w10885 ) ;
  assign w10892 = ( w10885 & w10887 ) | ( w10885 & w10891 ) | ( w10887 & w10891 ) ;
  assign w10893 = ( ~w10883 & w10887 ) | ( ~w10883 & w10892 ) | ( w10887 & w10892 ) ;
  assign w10894 = w10883 ^ w10892 ;
  assign w10895 = w10887 ^ w10894 ;
  assign w10896 = ~w4147 & w10895 ;
  assign w10897 = w10883 | w10890 ;
  assign w10898 = ( w3964 & w10890 ) | ( w3964 & w10897 ) | ( w10890 & w10897 ) ;
  assign w10899 = ( w10895 & ~w10896 ) | ( w10895 & w10898 ) | ( ~w10896 & w10898 ) ;
  assign w10900 = \pi26 ^ w10899 ;
  assign w10901 = w10820 ^ w10881 ;
  assign w10902 = w10900 ^ w10901 ;
  assign w10903 = w10223 ^ w10780 ;
  assign w10904 = w10344 ^ w10903 ;
  assign w10905 = w10289 ^ w10343 ;
  assign w10906 = w10332 ^ w10905 ;
  assign w10907 = w860 | w1094 ;
  assign w10908 = w409 | w10907 ;
  assign w10909 = ( w409 & ~w560 ) | ( w409 & w2949 ) | ( ~w560 & w2949 ) ;
  assign w10910 = ~w10908 & w10909 ;
  assign w10911 = ( w179 & ~w570 ) | ( w179 & w10910 ) | ( ~w570 & w10910 ) ;
  assign w10912 = ~w179 & w10911 ;
  assign w10913 = ( w385 & w506 ) | ( w385 & ~w573 ) | ( w506 & ~w573 ) ;
  assign w10914 = w255 | w2603 ;
  assign w10915 = ( ~w255 & w573 ) | ( ~w255 & w837 ) | ( w573 & w837 ) ;
  assign w10916 = w10914 | w10915 ;
  assign w10917 = w10913 | w10916 ;
  assign w10918 = ( w445 & w10912 ) | ( w445 & ~w10917 ) | ( w10912 & ~w10917 ) ;
  assign w10919 = w2451 | w3190 ;
  assign w10920 = ( w445 & w783 ) | ( w445 & ~w2451 ) | ( w783 & ~w2451 ) ;
  assign w10921 = w10919 | w10920 ;
  assign w10922 = w10918 & ~w10921 ;
  assign w10923 = w2705 | w4784 ;
  assign w10924 = w5230 | w10923 ;
  assign w10925 = ( ~w1881 & w5230 ) | ( ~w1881 & w10922 ) | ( w5230 & w10922 ) ;
  assign w10926 = ~w10924 & w10925 ;
  assign w10927 = ( w232 & w314 ) | ( w232 & ~w339 ) | ( w314 & ~w339 ) ;
  assign w10928 = ~w163 & w10926 ;
  assign w10929 = ( ~w163 & w339 ) | ( ~w163 & w623 ) | ( w339 & w623 ) ;
  assign w10930 = w10928 & ~w10929 ;
  assign w10931 = ~w10927 & w10930 ;
  assign w10932 = ( w176 & w467 ) | ( w176 & ~w491 ) | ( w467 & ~w491 ) ;
  assign w10933 = ~w51 & w10931 ;
  assign w10934 = ( ~w51 & w491 ) | ( ~w51 & w663 ) | ( w491 & w663 ) ;
  assign w10935 = w10933 & ~w10934 ;
  assign w10936 = ~w10932 & w10935 ;
  assign w10937 = ( w414 & ~w595 ) | ( w414 & w641 ) | ( ~w595 & w641 ) ;
  assign w10938 = w595 | w10937 ;
  assign w10939 = ( w390 & ~w517 ) | ( w390 & w10938 ) | ( ~w517 & w10938 ) ;
  assign w10940 = w517 | w10939 ;
  assign w10941 = w6313 | w10940 ;
  assign w10942 = ( w609 & w10489 ) | ( w609 & ~w10940 ) | ( w10489 & ~w10940 ) ;
  assign w10943 = w10941 | w10942 ;
  assign w10944 = ( w114 & w488 ) | ( w114 & ~w663 ) | ( w488 & ~w663 ) ;
  assign w10945 = w10244 | w10943 ;
  assign w10946 = ( w663 & w821 ) | ( w663 & ~w10244 ) | ( w821 & ~w10244 ) ;
  assign w10947 = w10945 | w10946 ;
  assign w10948 = w10944 | w10947 ;
  assign w10949 = ( w177 & ~w1616 ) | ( w177 & w2729 ) | ( ~w1616 & w2729 ) ;
  assign w10950 = w4814 | w10948 ;
  assign w10951 = ( w1616 & w2518 ) | ( w1616 & ~w4814 ) | ( w2518 & ~w4814 ) ;
  assign w10952 = w10950 | w10951 ;
  assign w10953 = w10949 | w10952 ;
  assign w10954 = ( w104 & w252 ) | ( w104 & ~w311 ) | ( w252 & ~w311 ) ;
  assign w10955 = w1413 | w10953 ;
  assign w10956 = ( w311 & w383 ) | ( w311 & ~w1413 ) | ( w383 & ~w1413 ) ;
  assign w10957 = w10955 | w10956 ;
  assign w10958 = w10954 | w10957 ;
  assign w10959 = ( \pi14 & \pi15 ) | ( \pi14 & ~\pi16 ) | ( \pi15 & ~\pi16 ) ;
  assign w10960 = ( \pi16 & ~\pi17 ) | ( \pi16 & w10959 ) | ( ~\pi17 & w10959 ) ;
  assign w10961 = w10738 ^ w10960 ;
  assign w10962 = ( \pi17 & w10960 ) | ( \pi17 & w10961 ) | ( w10960 & w10961 ) ;
  assign w10963 = ( w10936 & ~w10958 ) | ( w10936 & w10962 ) | ( ~w10958 & w10962 ) ;
  assign w10964 = w9953 ^ w10047 ;
  assign w10965 = w9842 ^ w10964 ;
  assign w10966 = ~w37 & w10965 ;
  assign w10967 = w3098 & ~w9955 ;
  assign w10968 = ( w10965 & ~w10966 ) | ( w10965 & w10967 ) | ( ~w10966 & w10967 ) ;
  assign w10969 = ( \pi29 & \pi30 ) | ( \pi29 & w9953 ) | ( \pi30 & w9953 ) ;
  assign w10970 = \pi31 | w10969 ;
  assign w10971 = ( \pi29 & ~\pi30 ) | ( \pi29 & w9842 ) | ( ~\pi30 & w9842 ) ;
  assign w10972 = ( \pi29 & \pi31 ) | ( \pi29 & ~w10971 ) | ( \pi31 & ~w10971 ) ;
  assign w10973 = ( w10968 & w10970 ) | ( w10968 & ~w10972 ) | ( w10970 & ~w10972 ) ;
  assign w10974 = ( w10289 & ~w10963 ) | ( w10289 & w10973 ) | ( ~w10963 & w10973 ) ;
  assign w10975 = w9842 ^ w10046 ;
  assign w10976 = w9955 ^ w10975 ;
  assign w10977 = ( \pi29 & \pi31 ) | ( \pi29 & ~w9955 ) | ( \pi31 & ~w9955 ) ;
  assign w10978 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10977 ) | ( ~\pi30 & w10977 ) ;
  assign w10979 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10977 ) | ( \pi30 & w10977 ) ;
  assign w10980 = ( ~\pi29 & w9957 ) | ( ~\pi29 & w10979 ) | ( w9957 & w10979 ) ;
  assign w10981 = ( w9842 & w10979 ) | ( w9842 & ~w10980 ) | ( w10979 & ~w10980 ) ;
  assign w10982 = ~\pi31 & w10981 ;
  assign w10983 = ( w10978 & w10980 ) | ( w10978 & w10982 ) | ( w10980 & w10982 ) ;
  assign w10984 = ( w37 & ~w10976 ) | ( w37 & w10983 ) | ( ~w10976 & w10983 ) ;
  assign w10985 = w10983 | w10984 ;
  assign w10986 = w10936 ^ w10962 ;
  assign w10987 = w10958 ^ w10986 ;
  assign w10988 = w663 | w2168 ;
  assign w10989 = ( w317 & w1282 ) | ( w317 & ~w2168 ) | ( w1282 & ~w2168 ) ;
  assign w10990 = w10988 | w10989 ;
  assign w10991 = w318 | w421 ;
  assign w10992 = w216 | w10991 ;
  assign w10993 = ( ~w216 & w262 ) | ( ~w216 & w10990 ) | ( w262 & w10990 ) ;
  assign w10994 = w10992 | w10993 ;
  assign w10995 = w456 | w664 ;
  assign w10996 = w51 | w10995 ;
  assign w10997 = ( ~w51 & w218 ) | ( ~w51 & w10994 ) | ( w218 & w10994 ) ;
  assign w10998 = w10996 | w10997 ;
  assign w10999 = ( w606 & w623 ) | ( w606 & ~w764 ) | ( w623 & ~w764 ) ;
  assign w11000 = w268 | w531 ;
  assign w11001 = ( ~w531 & w764 ) | ( ~w531 & w1340 ) | ( w764 & w1340 ) ;
  assign w11002 = w11000 | w11001 ;
  assign w11003 = w10999 | w11002 ;
  assign w11004 = ( w98 & w113 ) | ( w98 & ~w309 ) | ( w113 & ~w309 ) ;
  assign w11005 = w4415 | w11003 ;
  assign w11006 = ( w309 & w817 ) | ( w309 & ~w11003 ) | ( w817 & ~w11003 ) ;
  assign w11007 = w11005 | w11006 ;
  assign w11008 = w11004 | w11007 ;
  assign w11009 = ( w209 & ~w495 ) | ( w209 & w1400 ) | ( ~w495 & w1400 ) ;
  assign w11010 = w5763 | w11008 ;
  assign w11011 = ( w495 & w674 ) | ( w495 & ~w5763 ) | ( w674 & ~w5763 ) ;
  assign w11012 = w11010 | w11011 ;
  assign w11013 = w11009 | w11012 ;
  assign w11014 = ( w225 & w254 ) | ( w225 & ~w429 ) | ( w254 & ~w429 ) ;
  assign w11015 = w56 | w11013 ;
  assign w11016 = ( ~w56 & w429 ) | ( ~w56 & w901 ) | ( w429 & w901 ) ;
  assign w11017 = w11015 | w11016 ;
  assign w11018 = w11014 | w11017 ;
  assign w11019 = w139 | w269 ;
  assign w11020 = ( ~w139 & w198 ) | ( ~w139 & w11018 ) | ( w198 & w11018 ) ;
  assign w11021 = w11019 | w11020 ;
  assign w11022 = ( w385 & ~w449 ) | ( w385 & w2005 ) | ( ~w449 & w2005 ) ;
  assign w11023 = w5608 | w11021 ;
  assign w11024 = ( w449 & w697 ) | ( w449 & ~w5608 ) | ( w697 & ~w5608 ) ;
  assign w11025 = w11023 | w11024 ;
  assign w11026 = w11022 | w11025 ;
  assign w11027 = ( ~w138 & w1616 ) | ( ~w138 & w10998 ) | ( w1616 & w10998 ) ;
  assign w11028 = w2938 | w11026 ;
  assign w11029 = ( w138 & w424 ) | ( w138 & ~w2938 ) | ( w424 & ~w2938 ) ;
  assign w11030 = w11028 | w11029 ;
  assign w11031 = w11027 | w11030 ;
  assign w11032 = w206 | w313 ;
  assign w11033 = w129 | w11032 ;
  assign w11034 = ( ~w129 & w1185 ) | ( ~w129 & w11031 ) | ( w1185 & w11031 ) ;
  assign w11035 = w11033 | w11034 ;
  assign w11036 = ( w340 & w569 ) | ( w340 & ~w641 ) | ( w569 & ~w641 ) ;
  assign w11037 = w285 | w11035 ;
  assign w11038 = ( ~w285 & w641 ) | ( ~w285 & w722 ) | ( w641 & w722 ) ;
  assign w11039 = w11037 | w11038 ;
  assign w11040 = w11036 | w11039 ;
  assign w11041 = ( ~w104 & w899 ) | ( ~w104 & w5036 ) | ( w899 & w5036 ) ;
  assign w11042 = w104 | w11041 ;
  assign w11043 = w422 | w512 ;
  assign w11044 = w177 | w11043 ;
  assign w11045 = ( ~w177 & w3115 ) | ( ~w177 & w11042 ) | ( w3115 & w11042 ) ;
  assign w11046 = w11044 | w11045 ;
  assign w11047 = w3590 | w4464 ;
  assign w11048 = ( w2850 & ~w3590 ) | ( w2850 & w11046 ) | ( ~w3590 & w11046 ) ;
  assign w11049 = w11047 | w11048 ;
  assign w11050 = w515 | w606 ;
  assign w11051 = w1104 | w11050 ;
  assign w11052 = ( w115 & ~w1104 ) | ( w115 & w11049 ) | ( ~w1104 & w11049 ) ;
  assign w11053 = w11051 | w11052 ;
  assign w11054 = ( w310 & w568 ) | ( w310 & ~w640 ) | ( w568 & ~w640 ) ;
  assign w11055 = w92 | w11053 ;
  assign w11056 = ( ~w92 & w640 ) | ( ~w92 & w681 ) | ( w640 & w681 ) ;
  assign w11057 = w11055 | w11056 ;
  assign w11058 = w11054 | w11057 ;
  assign w11059 = ( w120 & w198 ) | ( w120 & ~w362 ) | ( w198 & ~w362 ) ;
  assign w11060 = w416 | w1400 ;
  assign w11061 = ( w362 & w534 ) | ( w362 & ~w1400 ) | ( w534 & ~w1400 ) ;
  assign w11062 = w11060 | w11061 ;
  assign w11063 = w11059 | w11062 ;
  assign w11064 = ( ~w84 & w1565 ) | ( ~w84 & w4384 ) | ( w1565 & w4384 ) ;
  assign w11065 = w784 | w3143 ;
  assign w11066 = ( w84 & w341 ) | ( w84 & ~w784 ) | ( w341 & ~w784 ) ;
  assign w11067 = w11065 | w11066 ;
  assign w11068 = w11064 | w11067 ;
  assign w11069 = w428 | w11063 ;
  assign w11070 = w1870 & ~w11069 ;
  assign w11071 = ( w1870 & w6135 ) | ( w1870 & w11068 ) | ( w6135 & w11068 ) ;
  assign w11072 = w11070 & ~w11071 ;
  assign w11073 = w209 | w640 ;
  assign w11074 = w1896 | w11073 ;
  assign w11075 = ( ~w785 & w1896 ) | ( ~w785 & w11072 ) | ( w1896 & w11072 ) ;
  assign w11076 = ~w11074 & w11075 ;
  assign w11077 = ( w205 & w277 ) | ( w205 & ~w280 ) | ( w277 & ~w280 ) ;
  assign w11078 = ~w95 & w11076 ;
  assign w11079 = ( ~w95 & w280 ) | ( ~w95 & w284 ) | ( w280 & w284 ) ;
  assign w11080 = w11078 & ~w11079 ;
  assign w11081 = ~w11077 & w11080 ;
  assign w11082 = ( \pi11 & \pi12 ) | ( \pi11 & ~\pi13 ) | ( \pi12 & ~\pi13 ) ;
  assign w11083 = ( \pi13 & ~\pi14 ) | ( \pi13 & w11082 ) | ( ~\pi14 & w11082 ) ;
  assign w11084 = w10738 ^ w11083 ;
  assign w11085 = ( \pi14 & w11083 ) | ( \pi14 & w11084 ) | ( w11083 & w11084 ) ;
  assign w11086 = ( ~w11058 & w11081 ) | ( ~w11058 & w11085 ) | ( w11081 & w11085 ) ;
  assign w11087 = ( w9961 & ~w9963 ) | ( w9961 & w10043 ) | ( ~w9963 & w10043 ) ;
  assign w11088 = w9963 ^ w11087 ;
  assign w11089 = w9957 ^ w11088 ;
  assign w11090 = w37 | w11089 ;
  assign w11091 = w3098 & w9961 ;
  assign w11092 = ( ~w11089 & w11090 ) | ( ~w11089 & w11091 ) | ( w11090 & w11091 ) ;
  assign w11093 = ( \pi29 & \pi30 ) | ( \pi29 & w9957 ) | ( \pi30 & w9957 ) ;
  assign w11094 = \pi31 | w11093 ;
  assign w11095 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w9963 ) | ( \pi30 & w9963 ) ;
  assign w11096 = ( \pi29 & \pi31 ) | ( \pi29 & w11095 ) | ( \pi31 & w11095 ) ;
  assign w11097 = ( w11092 & w11094 ) | ( w11092 & ~w11096 ) | ( w11094 & ~w11096 ) ;
  assign w11098 = ( w11040 & w11086 ) | ( w11040 & ~w11097 ) | ( w11086 & ~w11097 ) ;
  assign w11099 = ( w10936 & w11040 ) | ( w10936 & ~w11098 ) | ( w11040 & ~w11098 ) ;
  assign w11100 = ( w10985 & w10987 ) | ( w10985 & w11099 ) | ( w10987 & w11099 ) ;
  assign w11101 = w10963 ^ w10973 ;
  assign w11102 = w10289 ^ w11101 ;
  assign w11103 = ~w3717 & w10211 ;
  assign w11104 = w3649 & w10114 ;
  assign w11105 = ( w10211 & ~w11103 ) | ( w10211 & w11104 ) | ( ~w11103 & w11104 ) ;
  assign w11106 = ~w3549 & w10784 ;
  assign w11107 = w10789 | w11105 ;
  assign w11108 = ( w3448 & w11105 ) | ( w3448 & w11107 ) | ( w11105 & w11107 ) ;
  assign w11109 = ( w10784 & ~w11106 ) | ( w10784 & w11108 ) | ( ~w11106 & w11108 ) ;
  assign w11110 = \pi29 ^ w11109 ;
  assign w11111 = ( w11100 & ~w11102 ) | ( w11100 & w11110 ) | ( ~w11102 & w11110 ) ;
  assign w11112 = ( ~w10906 & w10974 ) | ( ~w10906 & w11111 ) | ( w10974 & w11111 ) ;
  assign w11113 = w3717 | w10805 ;
  assign w11114 = w3649 & w10784 ;
  assign w11115 = ( ~w10805 & w11113 ) | ( ~w10805 & w11114 ) | ( w11113 & w11114 ) ;
  assign w11116 = w10807 ^ w10811 ;
  assign w11117 = w10805 ^ w11116 ;
  assign w11118 = w3549 | w10807 ;
  assign w11119 = w11115 | w11117 ;
  assign w11120 = ( w3448 & w11115 ) | ( w3448 & w11119 ) | ( w11115 & w11119 ) ;
  assign w11121 = ( ~w10807 & w11118 ) | ( ~w10807 & w11120 ) | ( w11118 & w11120 ) ;
  assign w11122 = \pi29 ^ w11121 ;
  assign w11123 = ( ~w10904 & w11112 ) | ( ~w10904 & w11122 ) | ( w11112 & w11122 ) ;
  assign w11124 = w10781 ^ w10799 ;
  assign w11125 = w10819 ^ w11124 ;
  assign w11126 = w4143 | w10885 ;
  assign w11127 = w4052 & ~w10866 ;
  assign w11128 = ( ~w10885 & w11126 ) | ( ~w10885 & w11127 ) | ( w11126 & w11127 ) ;
  assign w11129 = ( ~w10866 & w10871 ) | ( ~w10866 & w10885 ) | ( w10871 & w10885 ) ;
  assign w11130 = w10871 ^ w11129 ;
  assign w11131 = w10887 ^ w11130 ;
  assign w11132 = w4147 | w11131 ;
  assign w11133 = w10887 & ~w11128 ;
  assign w11134 = ( w3964 & w11128 ) | ( w3964 & ~w11133 ) | ( w11128 & ~w11133 ) ;
  assign w11135 = ( ~w11131 & w11132 ) | ( ~w11131 & w11134 ) | ( w11132 & w11134 ) ;
  assign w11136 = \pi26 ^ w11135 ;
  assign w11137 = ( w11123 & w11125 ) | ( w11123 & w11136 ) | ( w11125 & w11136 ) ;
  assign w11138 = ~w10402 & w10737 ;
  assign w11139 = w10738 | w11138 ;
  assign w11140 = ( w4606 & w4651 ) | ( w4606 & ~w11138 ) | ( w4651 & ~w11138 ) ;
  assign w11141 = w4651 & ~w11140 ;
  assign w11142 = ( w4706 & ~w11140 ) | ( w4706 & w11141 ) | ( ~w11140 & w11141 ) ;
  assign w11143 = ( ~w10738 & w11140 ) | ( ~w10738 & w11142 ) | ( w11140 & w11142 ) ;
  assign w11144 = ( ~w10883 & w10893 ) | ( ~w10883 & w11139 ) | ( w10893 & w11139 ) ;
  assign w11145 = w11138 ^ w11144 ;
  assign w11146 = ( w10738 & w11144 ) | ( w10738 & ~w11145 ) | ( w11144 & ~w11145 ) ;
  assign w11147 = w4609 & w11146 ;
  assign w11148 = ( w4609 & w11143 ) | ( w4609 & ~w11147 ) | ( w11143 & ~w11147 ) ;
  assign w11149 = w11137 ^ w11148 ;
  assign w11150 = \pi23 ^ w10902 ;
  assign w11151 = w11149 ^ w11150 ;
  assign w11152 = w11123 ^ w11125 ;
  assign w11153 = w11136 ^ w11152 ;
  assign w11154 = w10904 ^ w11112 ;
  assign w11155 = w11122 ^ w11154 ;
  assign w11156 = w4143 | w10866 ;
  assign w11157 = w4052 & w10801 ;
  assign w11158 = ( ~w10866 & w11156 ) | ( ~w10866 & w11157 ) | ( w11156 & w11157 ) ;
  assign w11159 = w10871 ^ w10885 ;
  assign w11160 = w10866 ^ w11159 ;
  assign w11161 = w4147 | w11160 ;
  assign w11162 = w10885 & ~w11158 ;
  assign w11163 = ( w3964 & w11158 ) | ( w3964 & ~w11162 ) | ( w11158 & ~w11162 ) ;
  assign w11164 = ( ~w11160 & w11161 ) | ( ~w11160 & w11163 ) | ( w11161 & w11163 ) ;
  assign w11165 = \pi26 ^ w11164 ;
  assign w11166 = w10974 ^ w11111 ;
  assign w11167 = w10906 ^ w11166 ;
  assign w11168 = ~w3717 & w10784 ;
  assign w11169 = w3649 & w10211 ;
  assign w11170 = ( w10784 & ~w11168 ) | ( w10784 & w11169 ) | ( ~w11168 & w11169 ) ;
  assign w11171 = w3549 | w10805 ;
  assign w11172 = w10855 & ~w11170 ;
  assign w11173 = ( w3448 & w11170 ) | ( w3448 & ~w11172 ) | ( w11170 & ~w11172 ) ;
  assign w11174 = ( ~w10805 & w11171 ) | ( ~w10805 & w11173 ) | ( w11171 & w11173 ) ;
  assign w11175 = \pi29 ^ w11174 ;
  assign w11176 = ~w4143 & w10801 ;
  assign w11177 = w4052 & ~w10807 ;
  assign w11178 = ( w10801 & ~w11176 ) | ( w10801 & w11177 ) | ( ~w11176 & w11177 ) ;
  assign w11179 = ~w4147 & w10874 ;
  assign w11180 = w10866 & ~w11178 ;
  assign w11181 = ( w3964 & w11178 ) | ( w3964 & ~w11180 ) | ( w11178 & ~w11180 ) ;
  assign w11182 = ( w10874 & ~w11179 ) | ( w10874 & w11181 ) | ( ~w11179 & w11181 ) ;
  assign w11183 = \pi26 ^ w11182 ;
  assign w11184 = ( ~w11167 & w11175 ) | ( ~w11167 & w11183 ) | ( w11175 & w11183 ) ;
  assign w11185 = ( ~w11155 & w11165 ) | ( ~w11155 & w11184 ) | ( w11165 & w11184 ) ;
  assign w11186 = w4651 | w11139 ;
  assign w11187 = w4606 & w10883 ;
  assign w11188 = ( ~w11139 & w11186 ) | ( ~w11139 & w11187 ) | ( w11186 & w11187 ) ;
  assign w11189 = w4706 | w10738 ;
  assign w11190 = w11145 & ~w11188 ;
  assign w11191 = ( w4609 & w11188 ) | ( w4609 & ~w11190 ) | ( w11188 & ~w11190 ) ;
  assign w11192 = ( ~w10738 & w11189 ) | ( ~w10738 & w11191 ) | ( w11189 & w11191 ) ;
  assign w11193 = \pi23 ^ w11192 ;
  assign w11194 = ( w11153 & w11185 ) | ( w11153 & w11193 ) | ( w11185 & w11193 ) ;
  assign w11195 = w11153 ^ w11185 ;
  assign w11196 = w11193 ^ w11195 ;
  assign w11197 = w11167 ^ w11183 ;
  assign w11198 = w11175 ^ w11197 ;
  assign w11199 = w11040 ^ w11098 ;
  assign w11200 = w10936 ^ w11199 ;
  assign w11201 = w9955 ^ w10045 ;
  assign w11202 = w9957 ^ w11201 ;
  assign w11203 = ( \pi29 & \pi31 ) | ( \pi29 & w9957 ) | ( \pi31 & w9957 ) ;
  assign w11204 = ( \pi29 & ~\pi30 ) | ( \pi29 & w11203 ) | ( ~\pi30 & w11203 ) ;
  assign w11205 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w11203 ) | ( \pi30 & w11203 ) ;
  assign w11206 = ( \pi29 & w9963 ) | ( \pi29 & ~w11205 ) | ( w9963 & ~w11205 ) ;
  assign w11207 = ( ~w9955 & w11205 ) | ( ~w9955 & w11206 ) | ( w11205 & w11206 ) ;
  assign w11208 = ~\pi31 & w11207 ;
  assign w11209 = ( w11204 & ~w11206 ) | ( w11204 & w11208 ) | ( ~w11206 & w11208 ) ;
  assign w11210 = ( w37 & ~w11202 ) | ( w37 & w11209 ) | ( ~w11202 & w11209 ) ;
  assign w11211 = w11209 | w11210 ;
  assign w11212 = ~w3717 & w9953 ;
  assign w11213 = w3649 & w9842 ;
  assign w11214 = ( w9953 & ~w11212 ) | ( w9953 & w11213 ) | ( ~w11212 & w11213 ) ;
  assign w11215 = ~w3549 & w10114 ;
  assign w11216 = w10334 | w11214 ;
  assign w11217 = ( w3448 & w11214 ) | ( w3448 & w11216 ) | ( w11214 & w11216 ) ;
  assign w11218 = ( w10114 & ~w11215 ) | ( w10114 & w11217 ) | ( ~w11215 & w11217 ) ;
  assign w11219 = \pi29 ^ w11218 ;
  assign w11220 = ( ~w11200 & w11211 ) | ( ~w11200 & w11219 ) | ( w11211 & w11219 ) ;
  assign w11221 = w10987 ^ w11099 ;
  assign w11222 = w10985 ^ w11221 ;
  assign w11223 = ~w3717 & w10114 ;
  assign w11224 = w3649 & w9953 ;
  assign w11225 = ( w10114 & ~w11223 ) | ( w10114 & w11224 ) | ( ~w11223 & w11224 ) ;
  assign w11226 = ~w3549 & w10211 ;
  assign w11227 = w10214 | w11225 ;
  assign w11228 = ( w3448 & w11225 ) | ( w3448 & w11227 ) | ( w11225 & w11227 ) ;
  assign w11229 = ( w10211 & ~w11226 ) | ( w10211 & w11228 ) | ( ~w11226 & w11228 ) ;
  assign w11230 = \pi29 ^ w11229 ;
  assign w11231 = ( w11220 & w11222 ) | ( w11220 & w11230 ) | ( w11222 & w11230 ) ;
  assign w11232 = w11100 ^ w11102 ;
  assign w11233 = w11110 ^ w11232 ;
  assign w11234 = w4143 | w10807 ;
  assign w11235 = w4052 & ~w10805 ;
  assign w11236 = ( ~w10807 & w11234 ) | ( ~w10807 & w11235 ) | ( w11234 & w11235 ) ;
  assign w11237 = ~w4147 & w10814 ;
  assign w11238 = w10801 | w11236 ;
  assign w11239 = ( w3964 & w11236 ) | ( w3964 & w11238 ) | ( w11236 & w11238 ) ;
  assign w11240 = ( w10814 & ~w11237 ) | ( w10814 & w11239 ) | ( ~w11237 & w11239 ) ;
  assign w11241 = \pi26 ^ w11240 ;
  assign w11242 = ( w11231 & ~w11233 ) | ( w11231 & w11241 ) | ( ~w11233 & w11241 ) ;
  assign w11243 = w4651 | w10887 ;
  assign w11244 = w4606 & ~w10885 ;
  assign w11245 = ( ~w10887 & w11243 ) | ( ~w10887 & w11244 ) | ( w11243 & w11244 ) ;
  assign w11246 = ~w4706 & w10883 ;
  assign w11247 = w10895 | w11245 ;
  assign w11248 = ( w4609 & w11245 ) | ( w4609 & w11247 ) | ( w11245 & w11247 ) ;
  assign w11249 = ( w10883 & ~w11246 ) | ( w10883 & w11248 ) | ( ~w11246 & w11248 ) ;
  assign w11250 = \pi23 ^ w11249 ;
  assign w11251 = ( ~w11198 & w11242 ) | ( ~w11198 & w11250 ) | ( w11242 & w11250 ) ;
  assign w11252 = ~w4651 & w10883 ;
  assign w11253 = w4606 & ~w10887 ;
  assign w11254 = ( w10883 & ~w11252 ) | ( w10883 & w11253 ) | ( ~w11252 & w11253 ) ;
  assign w11255 = w10893 ^ w11139 ;
  assign w11256 = w10883 ^ w11255 ;
  assign w11257 = w4706 | w11139 ;
  assign w11258 = w11254 | w11256 ;
  assign w11259 = ( w4609 & w11254 ) | ( w4609 & w11258 ) | ( w11254 & w11258 ) ;
  assign w11260 = ( ~w11139 & w11257 ) | ( ~w11139 & w11259 ) | ( w11257 & w11259 ) ;
  assign w11261 = \pi23 ^ w11260 ;
  assign w11262 = w11155 ^ w11184 ;
  assign w11263 = w11165 ^ w11262 ;
  assign w11264 = ( w11251 & w11261 ) | ( w11251 & ~w11263 ) | ( w11261 & ~w11263 ) ;
  assign w11265 = w11231 ^ w11233 ;
  assign w11266 = w11241 ^ w11265 ;
  assign w11267 = w11220 ^ w11222 ;
  assign w11268 = w11230 ^ w11267 ;
  assign w11269 = w4143 | w10805 ;
  assign w11270 = w4052 & w10784 ;
  assign w11271 = ( ~w10805 & w11269 ) | ( ~w10805 & w11270 ) | ( w11269 & w11270 ) ;
  assign w11272 = ~w4147 & w11117 ;
  assign w11273 = w10807 & ~w11271 ;
  assign w11274 = ( w3964 & w11271 ) | ( w3964 & ~w11273 ) | ( w11271 & ~w11273 ) ;
  assign w11275 = ( w11117 & ~w11272 ) | ( w11117 & w11274 ) | ( ~w11272 & w11274 ) ;
  assign w11276 = \pi26 ^ w11275 ;
  assign w11277 = w9963 ^ w10043 ;
  assign w11278 = w9961 ^ w11277 ;
  assign w11279 = ( \pi29 & \pi31 ) | ( \pi29 & w9961 ) | ( \pi31 & w9961 ) ;
  assign w11280 = ( \pi29 & ~\pi30 ) | ( \pi29 & w11279 ) | ( ~\pi30 & w11279 ) ;
  assign w11281 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w11279 ) | ( \pi30 & w11279 ) ;
  assign w11282 = ( ~\pi29 & w9965 ) | ( ~\pi29 & w11281 ) | ( w9965 & w11281 ) ;
  assign w11283 = ( w9963 & ~w11281 ) | ( w9963 & w11282 ) | ( ~w11281 & w11282 ) ;
  assign w11284 = \pi31 | w11283 ;
  assign w11285 = ( w11280 & w11282 ) | ( w11280 & ~w11284 ) | ( w11282 & ~w11284 ) ;
  assign w11286 = ( w37 & ~w11278 ) | ( w37 & w11285 ) | ( ~w11278 & w11285 ) ;
  assign w11287 = w11285 | w11286 ;
  assign w11288 = ( w316 & w415 ) | ( w316 & ~w506 ) | ( w415 & ~w506 ) ;
  assign w11289 = w98 | w111 ;
  assign w11290 = ( ~w111 & w506 ) | ( ~w111 & w608 ) | ( w506 & w608 ) ;
  assign w11291 = w11289 | w11290 ;
  assign w11292 = w11288 | w11291 ;
  assign w11293 = ( w143 & ~w722 ) | ( w143 & w11292 ) | ( ~w722 & w11292 ) ;
  assign w11294 = w3630 | w5592 ;
  assign w11295 = ( w722 & w764 ) | ( w722 & ~w5592 ) | ( w764 & ~w5592 ) ;
  assign w11296 = w11294 | w11295 ;
  assign w11297 = w11293 | w11296 ;
  assign w11298 = w524 | w2092 ;
  assign w11299 = ( w147 & ~w2092 ) | ( w147 & w11297 ) | ( ~w2092 & w11297 ) ;
  assign w11300 = w11298 | w11299 ;
  assign w11301 = w886 | w888 ;
  assign w11302 = w343 | w11301 ;
  assign w11303 = ( ~w343 & w785 ) | ( ~w343 & w11300 ) | ( w785 & w11300 ) ;
  assign w11304 = w11302 | w11303 ;
  assign w11305 = w662 | w1340 ;
  assign w11306 = w131 | w11305 ;
  assign w11307 = ( ~w131 & w393 ) | ( ~w131 & w11304 ) | ( w393 & w11304 ) ;
  assign w11308 = w11306 | w11307 ;
  assign w11309 = w491 | w642 ;
  assign w11310 = w198 | w11309 ;
  assign w11311 = w3254 | w11310 ;
  assign w11312 = w1010 | w2501 ;
  assign w11313 = ( ~w1010 & w1836 ) | ( ~w1010 & w11311 ) | ( w1836 & w11311 ) ;
  assign w11314 = w11312 | w11313 ;
  assign w11315 = w860 | w1031 ;
  assign w11316 = w101 | w11315 ;
  assign w11317 = ( ~w101 & w315 ) | ( ~w101 & w11314 ) | ( w315 & w11314 ) ;
  assign w11318 = w11316 | w11317 ;
  assign w11319 = w2395 | w3782 ;
  assign w11320 = ( w527 & ~w3782 ) | ( w527 & w11318 ) | ( ~w3782 & w11318 ) ;
  assign w11321 = w11319 | w11320 ;
  assign w11322 = w956 | w1069 ;
  assign w11323 = w11321 | w11322 ;
  assign w11324 = ( w444 & w11308 ) | ( w444 & ~w11321 ) | ( w11308 & ~w11321 ) ;
  assign w11325 = w11323 | w11324 ;
  assign w11326 = w199 | w565 ;
  assign w11327 = w11325 | w11326 ;
  assign w11328 = ( w2167 & w4174 ) | ( w2167 & ~w11325 ) | ( w4174 & ~w11325 ) ;
  assign w11329 = w11327 | w11328 ;
  assign w11330 = ( w167 & w284 ) | ( w167 & ~w424 ) | ( w284 & ~w424 ) ;
  assign w11331 = w104 | w11329 ;
  assign w11332 = ( ~w104 & w424 ) | ( ~w104 & w1086 ) | ( w424 & w1086 ) ;
  assign w11333 = w11331 | w11332 ;
  assign w11334 = w11330 | w11333 ;
  assign w11335 = w128 | w664 ;
  assign w11336 = ( ~w128 & w176 ) | ( ~w128 & w11334 ) | ( w176 & w11334 ) ;
  assign w11337 = w11335 | w11336 ;
  assign w11338 = w9961 ^ w10042 ;
  assign w11339 = w9965 ^ w11338 ;
  assign w11340 = ( \pi29 & \pi31 ) | ( \pi29 & w9965 ) | ( \pi31 & w9965 ) ;
  assign w11341 = ( \pi29 & ~\pi30 ) | ( \pi29 & w11340 ) | ( ~\pi30 & w11340 ) ;
  assign w11342 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w11340 ) | ( \pi30 & w11340 ) ;
  assign w11343 = ( \pi29 & w9967 ) | ( \pi29 & ~w11342 ) | ( w9967 & ~w11342 ) ;
  assign w11344 = ( w9961 & w11342 ) | ( w9961 & w11343 ) | ( w11342 & w11343 ) ;
  assign w11345 = ~\pi31 & w11344 ;
  assign w11346 = ( w11341 & ~w11343 ) | ( w11341 & w11345 ) | ( ~w11343 & w11345 ) ;
  assign w11347 = ( w37 & w11339 ) | ( w37 & w11346 ) | ( w11339 & w11346 ) ;
  assign w11348 = w11346 | w11347 ;
  assign w11349 = ( ~w11058 & w11337 ) | ( ~w11058 & w11348 ) | ( w11337 & w11348 ) ;
  assign w11350 = w11058 ^ w11085 ;
  assign w11351 = w11081 ^ w11350 ;
  assign w11352 = ( w11287 & w11349 ) | ( w11287 & w11351 ) | ( w11349 & w11351 ) ;
  assign w11353 = w11086 ^ w11097 ;
  assign w11354 = w11040 ^ w11353 ;
  assign w11355 = ~w3717 & w9842 ;
  assign w11356 = w3649 & ~w9955 ;
  assign w11357 = ( w9842 & ~w11355 ) | ( w9842 & w11356 ) | ( ~w11355 & w11356 ) ;
  assign w11358 = ~w3549 & w9953 ;
  assign w11359 = w10965 | w11357 ;
  assign w11360 = ( w3448 & w11357 ) | ( w3448 & w11359 ) | ( w11357 & w11359 ) ;
  assign w11361 = ( w9953 & ~w11358 ) | ( w9953 & w11360 ) | ( ~w11358 & w11360 ) ;
  assign w11362 = \pi29 ^ w11361 ;
  assign w11363 = ( w11352 & w11354 ) | ( w11352 & w11362 ) | ( w11354 & w11362 ) ;
  assign w11364 = w11200 ^ w11219 ;
  assign w11365 = w11211 ^ w11364 ;
  assign w11366 = ~w4143 & w10784 ;
  assign w11367 = w4052 & w10211 ;
  assign w11368 = ( w10784 & ~w11366 ) | ( w10784 & w11367 ) | ( ~w11366 & w11367 ) ;
  assign w11369 = w4147 | w10855 ;
  assign w11370 = w10805 & ~w11368 ;
  assign w11371 = ( w3964 & w11368 ) | ( w3964 & ~w11370 ) | ( w11368 & ~w11370 ) ;
  assign w11372 = ( ~w10855 & w11369 ) | ( ~w10855 & w11371 ) | ( w11369 & w11371 ) ;
  assign w11373 = \pi26 ^ w11372 ;
  assign w11374 = ( w11363 & ~w11365 ) | ( w11363 & w11373 ) | ( ~w11365 & w11373 ) ;
  assign w11375 = ( w11268 & w11276 ) | ( w11268 & w11374 ) | ( w11276 & w11374 ) ;
  assign w11376 = w4651 | w10885 ;
  assign w11377 = w4606 & ~w10866 ;
  assign w11378 = ( ~w10885 & w11376 ) | ( ~w10885 & w11377 ) | ( w11376 & w11377 ) ;
  assign w11379 = w4706 | w10887 ;
  assign w11380 = w11131 & ~w11378 ;
  assign w11381 = ( w4609 & w11378 ) | ( w4609 & ~w11380 ) | ( w11378 & ~w11380 ) ;
  assign w11382 = ( ~w10887 & w11379 ) | ( ~w10887 & w11381 ) | ( w11379 & w11381 ) ;
  assign w11383 = \pi23 ^ w11382 ;
  assign w11384 = ( ~w11266 & w11375 ) | ( ~w11266 & w11383 ) | ( w11375 & w11383 ) ;
  assign w11385 = ( w4905 & w5343 ) | ( w4905 & ~w11138 ) | ( w5343 & ~w11138 ) ;
  assign w11386 = w5343 & ~w11385 ;
  assign w11387 = ( w5395 & ~w11385 ) | ( w5395 & w11386 ) | ( ~w11385 & w11386 ) ;
  assign w11388 = ( ~w10738 & w11385 ) | ( ~w10738 & w11387 ) | ( w11385 & w11387 ) ;
  assign w11389 = w11198 ^ w11242 ;
  assign w11390 = w11250 ^ w11389 ;
  assign w11391 = w11146 & ~w11388 ;
  assign w11392 = ( w4908 & w11388 ) | ( w4908 & ~w11391 ) | ( w11388 & ~w11391 ) ;
  assign w11393 = \pi20 ^ w11392 ;
  assign w11394 = ( w11384 & ~w11390 ) | ( w11384 & w11393 ) | ( ~w11390 & w11393 ) ;
  assign w11395 = w11251 ^ w11263 ;
  assign w11396 = w11261 ^ w11395 ;
  assign w11397 = w4908 & w11146 ;
  assign w11398 = ( w4908 & w11388 ) | ( w4908 & ~w11397 ) | ( w11388 & ~w11397 ) ;
  assign w11399 = w11390 ^ w11398 ;
  assign w11400 = \pi20 ^ w11384 ;
  assign w11401 = w11399 ^ w11400 ;
  assign w11402 = w11266 ^ w11375 ;
  assign w11403 = w11383 ^ w11402 ;
  assign w11404 = w11268 ^ w11374 ;
  assign w11405 = w11276 ^ w11404 ;
  assign w11406 = w4651 | w10866 ;
  assign w11407 = w4606 & w10801 ;
  assign w11408 = ( ~w10866 & w11406 ) | ( ~w10866 & w11407 ) | ( w11406 & w11407 ) ;
  assign w11409 = w4706 | w10885 ;
  assign w11410 = w11160 & ~w11408 ;
  assign w11411 = ( w4609 & w11408 ) | ( w4609 & ~w11410 ) | ( w11408 & ~w11410 ) ;
  assign w11412 = ( ~w10885 & w11409 ) | ( ~w10885 & w11411 ) | ( w11409 & w11411 ) ;
  assign w11413 = \pi23 ^ w11412 ;
  assign w11414 = w11363 ^ w11365 ;
  assign w11415 = w11373 ^ w11414 ;
  assign w11416 = w11287 ^ w11351 ;
  assign w11417 = w11349 ^ w11416 ;
  assign w11418 = w3717 | w9955 ;
  assign w11419 = w3649 & w9957 ;
  assign w11420 = ( ~w9955 & w11418 ) | ( ~w9955 & w11419 ) | ( w11418 & w11419 ) ;
  assign w11421 = ~w3549 & w9842 ;
  assign w11422 = w10976 & ~w11420 ;
  assign w11423 = ( w3448 & w11420 ) | ( w3448 & ~w11422 ) | ( w11420 & ~w11422 ) ;
  assign w11424 = ( w9842 & ~w11421 ) | ( w9842 & w11423 ) | ( ~w11421 & w11423 ) ;
  assign w11425 = \pi29 ^ w11424 ;
  assign w11426 = w11058 ^ w11348 ;
  assign w11427 = w11337 ^ w11426 ;
  assign w11428 = ( w313 & w415 ) | ( w313 & ~w524 ) | ( w415 & ~w524 ) ;
  assign w11429 = w1302 | w1646 ;
  assign w11430 = ( w524 & w899 ) | ( w524 & ~w1646 ) | ( w899 & ~w1646 ) ;
  assign w11431 = w11429 | w11430 ;
  assign w11432 = w11428 | w11431 ;
  assign w11433 = ( w490 & w512 ) | ( w490 & ~w560 ) | ( w512 & ~w560 ) ;
  assign w11434 = w90 | w11432 ;
  assign w11435 = ( ~w90 & w560 ) | ( ~w90 & w573 ) | ( w560 & w573 ) ;
  assign w11436 = w11434 | w11435 ;
  assign w11437 = w11433 | w11436 ;
  assign w11438 = ~w165 & w359 ;
  assign w11439 = ( ~w165 & w284 ) | ( ~w165 & w11437 ) | ( w284 & w11437 ) ;
  assign w11440 = w11438 & ~w11439 ;
  assign w11441 = ( w225 & w260 ) | ( w225 & ~w393 ) | ( w260 & ~w393 ) ;
  assign w11442 = w135 | w202 ;
  assign w11443 = ( ~w202 & w393 ) | ( ~w202 & w726 ) | ( w393 & w726 ) ;
  assign w11444 = w11442 | w11443 ;
  assign w11445 = w11441 | w11444 ;
  assign w11446 = w352 | w11445 ;
  assign w11447 = ( w265 & w388 ) | ( w265 & ~w593 ) | ( w388 & ~w593 ) ;
  assign w11448 = w139 | w226 ;
  assign w11449 = ( ~w226 & w593 ) | ( ~w226 & w1340 ) | ( w593 & w1340 ) ;
  assign w11450 = w11448 | w11449 ;
  assign w11451 = w11447 | w11450 ;
  assign w11452 = ( ~w2092 & w4207 ) | ( ~w2092 & w11446 ) | ( w4207 & w11446 ) ;
  assign w11453 = w2909 | w5854 ;
  assign w11454 = ( w2092 & ~w5854 ) | ( w2092 & w11451 ) | ( ~w5854 & w11451 ) ;
  assign w11455 = w11453 | w11454 ;
  assign w11456 = w11452 | w11455 ;
  assign w11457 = ( w1401 & w1421 ) | ( w1401 & ~w2705 ) | ( w1421 & ~w2705 ) ;
  assign w11458 = w11440 & ~w11456 ;
  assign w11459 = ( w413 & w2705 ) | ( w413 & w11440 ) | ( w2705 & w11440 ) ;
  assign w11460 = w11458 & ~w11459 ;
  assign w11461 = ~w11457 & w11460 ;
  assign w11462 = ( w263 & w324 ) | ( w263 & ~w361 ) | ( w324 & ~w361 ) ;
  assign w11463 = ~w254 & w11461 ;
  assign w11464 = ( ~w254 & w361 ) | ( ~w254 & w383 ) | ( w361 & w383 ) ;
  assign w11465 = w11463 & ~w11464 ;
  assign w11466 = ~w11462 & w11465 ;
  assign w11467 = ( w358 & ~w680 ) | ( w358 & w11466 ) | ( ~w680 & w11466 ) ;
  assign w11468 = ~w358 & w11467 ;
  assign w11469 = ( w92 & w127 ) | ( w92 & ~w568 ) | ( w127 & ~w568 ) ;
  assign w11470 = w1165 | w2295 ;
  assign w11471 = ( w568 & w625 ) | ( w568 & ~w2295 ) | ( w625 & ~w2295 ) ;
  assign w11472 = w11470 | w11471 ;
  assign w11473 = w11469 | w11472 ;
  assign w11474 = ( w310 & w496 ) | ( w310 & ~w515 ) | ( w496 & ~w515 ) ;
  assign w11475 = w56 | w111 ;
  assign w11476 = ( ~w111 & w515 ) | ( ~w111 & w640 ) | ( w515 & w640 ) ;
  assign w11477 = w11475 | w11476 ;
  assign w11478 = w11474 | w11477 ;
  assign w11479 = ( ~w389 & w596 ) | ( ~w389 & w11478 ) | ( w596 & w11478 ) ;
  assign w11480 = w389 | w11479 ;
  assign w11481 = ( ~w256 & w1145 ) | ( ~w256 & w11480 ) | ( w1145 & w11480 ) ;
  assign w11482 = w250 | w5562 ;
  assign w11483 = ( ~w250 & w256 ) | ( ~w250 & w530 ) | ( w256 & w530 ) ;
  assign w11484 = w11482 | w11483 ;
  assign w11485 = w11481 | w11484 ;
  assign w11486 = ( w952 & ~w3565 ) | ( w952 & w11473 ) | ( ~w3565 & w11473 ) ;
  assign w11487 = w3490 & ~w11485 ;
  assign w11488 = ( w3490 & w3565 ) | ( w3490 & w4381 ) | ( w3565 & w4381 ) ;
  assign w11489 = w11487 & ~w11488 ;
  assign w11490 = ~w11486 & w11489 ;
  assign w11491 = w180 | w390 ;
  assign w11492 = w114 | w11491 ;
  assign w11493 = ( w114 & ~w139 ) | ( w114 & w11490 ) | ( ~w139 & w11490 ) ;
  assign w11494 = ~w11492 & w11493 ;
  assign w11495 = ( \pi08 & \pi09 ) | ( \pi08 & ~\pi10 ) | ( \pi09 & ~\pi10 ) ;
  assign w11496 = ( \pi10 & ~\pi11 ) | ( \pi10 & w11495 ) | ( ~\pi11 & w11495 ) ;
  assign w11497 = w10738 ^ w11496 ;
  assign w11498 = ( \pi11 & w11496 ) | ( \pi11 & w11497 ) | ( w11496 & w11497 ) ;
  assign w11499 = ( w11468 & w11494 ) | ( w11468 & w11498 ) | ( w11494 & w11498 ) ;
  assign w11500 = w9965 ^ w10041 ;
  assign w11501 = w9967 ^ w11500 ;
  assign w11502 = w37 | w11501 ;
  assign w11503 = w3098 & w9971 ;
  assign w11504 = ( ~w11501 & w11502 ) | ( ~w11501 & w11503 ) | ( w11502 & w11503 ) ;
  assign w11505 = ( \pi29 & \pi30 ) | ( \pi29 & w9965 ) | ( \pi30 & w9965 ) ;
  assign w11506 = \pi31 | w11505 ;
  assign w11507 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w9967 ) | ( \pi30 & w9967 ) ;
  assign w11508 = ( \pi29 & \pi31 ) | ( \pi29 & w11507 ) | ( \pi31 & w11507 ) ;
  assign w11509 = ( w11504 & w11506 ) | ( w11504 & ~w11508 ) | ( w11506 & ~w11508 ) ;
  assign w11510 = ( w11058 & w11499 ) | ( w11058 & ~w11509 ) | ( w11499 & ~w11509 ) ;
  assign w11511 = w9967 ^ w10040 ;
  assign w11512 = w9971 ^ w11511 ;
  assign w11513 = ( \pi29 & \pi31 ) | ( \pi29 & w9971 ) | ( \pi31 & w9971 ) ;
  assign w11514 = ( \pi29 & ~\pi30 ) | ( \pi29 & w11513 ) | ( ~\pi30 & w11513 ) ;
  assign w11515 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w11513 ) | ( \pi30 & w11513 ) ;
  assign w11516 = ( \pi29 & w9973 ) | ( \pi29 & ~w11515 ) | ( w9973 & ~w11515 ) ;
  assign w11517 = ( ~w9967 & w11515 ) | ( ~w9967 & w11516 ) | ( w11515 & w11516 ) ;
  assign w11518 = ~\pi31 & w11517 ;
  assign w11519 = ( w11514 & ~w11516 ) | ( w11514 & w11518 ) | ( ~w11516 & w11518 ) ;
  assign w11520 = ( w37 & ~w11512 ) | ( w37 & w11519 ) | ( ~w11512 & w11519 ) ;
  assign w11521 = w11519 | w11520 ;
  assign w11522 = w11468 ^ w11498 ;
  assign w11523 = w11494 ^ w11522 ;
  assign w11524 = ( w571 & w623 ) | ( w571 & ~w1001 ) | ( w623 & ~w1001 ) ;
  assign w11525 = w84 | w672 ;
  assign w11526 = ( ~w84 & w1001 ) | ( ~w84 & w1094 ) | ( w1001 & w1094 ) ;
  assign w11527 = w11525 | w11526 ;
  assign w11528 = w11524 | w11527 ;
  assign w11529 = ( ~w141 & w674 ) | ( ~w141 & w11528 ) | ( w674 & w11528 ) ;
  assign w11530 = w141 | w11529 ;
  assign w11531 = w392 | w490 ;
  assign w11532 = w101 | w11531 ;
  assign w11533 = ( ~w101 & w361 ) | ( ~w101 & w11530 ) | ( w361 & w11530 ) ;
  assign w11534 = w11532 | w11533 ;
  assign w11535 = w252 | w1126 ;
  assign w11536 = ( w227 & ~w252 ) | ( w227 & w605 ) | ( ~w252 & w605 ) ;
  assign w11537 = w11535 | w11536 ;
  assign w11538 = w418 | w821 ;
  assign w11539 = ( ~w418 & w510 ) | ( ~w418 & w570 ) | ( w510 & w570 ) ;
  assign w11540 = w11538 | w11539 ;
  assign w11541 = ( w203 & w625 ) | ( w203 & ~w783 ) | ( w625 & ~w783 ) ;
  assign w11542 = w2784 | w11540 ;
  assign w11543 = ( w783 & w1153 ) | ( w783 & ~w11540 ) | ( w1153 & ~w11540 ) ;
  assign w11544 = w11542 | w11543 ;
  assign w11545 = w11541 | w11544 ;
  assign w11546 = ( w173 & ~w561 ) | ( w173 & w11537 ) | ( ~w561 & w11537 ) ;
  assign w11547 = w2003 & ~w11545 ;
  assign w11548 = ( w561 & w817 ) | ( w561 & ~w11545 ) | ( w817 & ~w11545 ) ;
  assign w11549 = w11547 & ~w11548 ;
  assign w11550 = ~w11546 & w11549 ;
  assign w11551 = ( w1302 & w1363 ) | ( w1302 & ~w1413 ) | ( w1363 & ~w1413 ) ;
  assign w11552 = ~w838 & w11550 ;
  assign w11553 = ( w388 & ~w838 ) | ( w388 & w1413 ) | ( ~w838 & w1413 ) ;
  assign w11554 = w11552 & ~w11553 ;
  assign w11555 = ~w11551 & w11554 ;
  assign w11556 = w260 | w1274 ;
  assign w11557 = w59 | w11556 ;
  assign w11558 = ( w59 & ~w92 ) | ( w59 & w11555 ) | ( ~w92 & w11555 ) ;
  assign w11559 = ~w11557 & w11558 ;
  assign w11560 = w681 | w899 ;
  assign w11561 = w272 | w11560 ;
  assign w11562 = ( ~w272 & w680 ) | ( ~w272 & w1689 ) | ( w680 & w1689 ) ;
  assign w11563 = w11561 | w11562 ;
  assign w11564 = w181 | w11563 ;
  assign w11565 = w4329 | w11564 ;
  assign w11566 = ( w4329 & ~w11534 ) | ( w4329 & w11559 ) | ( ~w11534 & w11559 ) ;
  assign w11567 = ~w11565 & w11566 ;
  assign w11568 = w524 | w663 ;
  assign w11569 = w147 | w11568 ;
  assign w11570 = ( w147 & ~w317 ) | ( w147 & w11567 ) | ( ~w317 & w11567 ) ;
  assign w11571 = ~w11569 & w11570 ;
  assign w11572 = w206 | w626 ;
  assign w11573 = w129 | w11572 ;
  assign w11574 = ( w129 & ~w343 ) | ( w129 & w11571 ) | ( ~w343 & w11571 ) ;
  assign w11575 = ~w11573 & w11574 ;
  assign w11576 = w225 | w408 ;
  assign w11577 = w86 | w11576 ;
  assign w11578 = ( w86 & ~w215 ) | ( w86 & w11575 ) | ( ~w215 & w11575 ) ;
  assign w11579 = ~w11577 & w11578 ;
  assign w11580 = ( w84 & w136 ) | ( w84 & ~w465 ) | ( w136 & ~w465 ) ;
  assign w11581 = w450 | w1617 ;
  assign w11582 = ( w465 & w980 ) | ( w465 & ~w1617 ) | ( w980 & ~w1617 ) ;
  assign w11583 = w11581 | w11582 ;
  assign w11584 = w11580 | w11583 ;
  assign w11585 = ( w252 & w573 ) | ( w252 & ~w596 ) | ( w573 & ~w596 ) ;
  assign w11586 = w101 | w11584 ;
  assign w11587 = ( ~w101 & w596 ) | ( ~w101 & w1030 ) | ( w596 & w1030 ) ;
  assign w11588 = w11586 | w11587 ;
  assign w11589 = w11585 | w11588 ;
  assign w11590 = ( w229 & w320 ) | ( w229 & ~w322 ) | ( w320 & ~w322 ) ;
  assign w11591 = w326 | w10938 ;
  assign w11592 = ( w322 & ~w326 ) | ( w322 & w509 ) | ( ~w326 & w509 ) ;
  assign w11593 = w11591 | w11592 ;
  assign w11594 = w11590 | w11593 ;
  assign w11595 = w821 | w1086 ;
  assign w11596 = w3494 | w11595 ;
  assign w11597 = ( w315 & ~w3494 ) | ( w315 & w11594 ) | ( ~w3494 & w11594 ) ;
  assign w11598 = w11596 | w11597 ;
  assign w11599 = w470 | w697 ;
  assign w11600 = ( ~w470 & w681 ) | ( ~w470 & w11598 ) | ( w681 & w11598 ) ;
  assign w11601 = w11599 | w11600 ;
  assign w11602 = ( w386 & w445 ) | ( w386 & ~w495 ) | ( w445 & ~w495 ) ;
  assign w11603 = w384 | w4210 ;
  assign w11604 = ( ~w384 & w495 ) | ( ~w384 & w496 ) | ( w495 & w496 ) ;
  assign w11605 = w11603 | w11604 ;
  assign w11606 = w11602 | w11605 ;
  assign w11607 = w204 | w4183 ;
  assign w11608 = ( ~w204 & w444 ) | ( ~w204 & w11606 ) | ( w444 & w11606 ) ;
  assign w11609 = w11607 | w11608 ;
  assign w11610 = ( w287 & w429 ) | ( w287 & ~w458 ) | ( w429 & ~w458 ) ;
  assign w11611 = w215 | w11609 ;
  assign w11612 = ( ~w215 & w458 ) | ( ~w215 & w817 ) | ( w458 & w817 ) ;
  assign w11613 = w11611 | w11612 ;
  assign w11614 = w11610 | w11613 ;
  assign w11615 = w3074 | w3618 ;
  assign w11616 = w3195 | w11615 ;
  assign w11617 = ( w2096 & w2420 ) | ( w2096 & ~w3195 ) | ( w2420 & ~w3195 ) ;
  assign w11618 = w11616 | w11617 ;
  assign w11619 = ( ~w2556 & w11589 ) | ( ~w2556 & w11614 ) | ( w11589 & w11614 ) ;
  assign w11620 = w11601 | w11618 ;
  assign w11621 = ( w2556 & w2760 ) | ( w2556 & ~w11601 ) | ( w2760 & ~w11601 ) ;
  assign w11622 = w11620 | w11621 ;
  assign w11623 = w11619 | w11622 ;
  assign w11624 = w169 | w1206 ;
  assign w11625 = w343 | w11624 ;
  assign w11626 = ( ~w343 & w731 ) | ( ~w343 & w11623 ) | ( w731 & w11623 ) ;
  assign w11627 = w11625 | w11626 ;
  assign w11628 = ( ~w92 & w317 ) | ( ~w92 & w11627 ) | ( w317 & w11627 ) ;
  assign w11629 = w92 | w11628 ;
  assign w11630 = ( w525 & w596 ) | ( w525 & ~w726 ) | ( w596 & ~w726 ) ;
  assign w11631 = w271 | w315 ;
  assign w11632 = ( ~w315 & w726 ) | ( ~w315 & w1274 ) | ( w726 & w1274 ) ;
  assign w11633 = w11631 | w11632 ;
  assign w11634 = w11630 | w11633 ;
  assign w11635 = w176 | w11634 ;
  assign w11636 = ( w1646 & ~w1744 ) | ( w1646 & w2082 ) | ( ~w1744 & w2082 ) ;
  assign w11637 = ~w1646 & w11636 ;
  assign w11638 = ( w120 & w254 ) | ( w120 & ~w268 ) | ( w254 & ~w268 ) ;
  assign w11639 = ~w822 & w11637 ;
  assign w11640 = ( w268 & w496 ) | ( w268 & ~w822 ) | ( w496 & ~w822 ) ;
  assign w11641 = w11639 & ~w11640 ;
  assign w11642 = ~w11638 & w11641 ;
  assign w11643 = ( w353 & w413 ) | ( w353 & ~w465 ) | ( w413 & ~w465 ) ;
  assign w11644 = w221 | w1957 ;
  assign w11645 = ( ~w221 & w465 ) | ( ~w221 & w533 ) | ( w465 & w533 ) ;
  assign w11646 = w11644 | w11645 ;
  assign w11647 = w11643 | w11646 ;
  assign w11648 = w285 | w512 ;
  assign w11649 = w1741 | w11648 ;
  assign w11650 = ( w227 & ~w1741 ) | ( w227 & w11647 ) | ( ~w1741 & w11647 ) ;
  assign w11651 = w11649 | w11650 ;
  assign w11652 = ( w11635 & w11642 ) | ( w11635 & ~w11651 ) | ( w11642 & ~w11651 ) ;
  assign w11653 = w1125 | w10623 ;
  assign w11654 = ( w87 & ~w10623 ) | ( w87 & w11635 ) | ( ~w10623 & w11635 ) ;
  assign w11655 = w11653 | w11654 ;
  assign w11656 = w11652 & ~w11655 ;
  assign w11657 = ( w344 & w345 ) | ( w344 & ~w388 ) | ( w345 & ~w388 ) ;
  assign w11658 = ~w180 & w11656 ;
  assign w11659 = ( ~w180 & w388 ) | ( ~w180 & w421 ) | ( w388 & w421 ) ;
  assign w11660 = w11658 & ~w11659 ;
  assign w11661 = ~w11657 & w11660 ;
  assign w11662 = w142 | w505 ;
  assign w11663 = ( w142 & ~w492 ) | ( w142 & w11661 ) | ( ~w492 & w11661 ) ;
  assign w11664 = ~w11662 & w11663 ;
  assign w11665 = ( \pi05 & \pi06 ) | ( \pi05 & ~\pi07 ) | ( \pi06 & ~\pi07 ) ;
  assign w11666 = ( \pi07 & ~\pi08 ) | ( \pi07 & w11665 ) | ( ~\pi08 & w11665 ) ;
  assign w11667 = w10738 ^ w11666 ;
  assign w11668 = ( \pi08 & w11666 ) | ( \pi08 & w11667 ) | ( w11666 & w11667 ) ;
  assign w11669 = ( ~w11629 & w11664 ) | ( ~w11629 & w11668 ) | ( w11664 & w11668 ) ;
  assign w11670 = w9973 ^ w10038 ;
  assign w11671 = w9975 ^ w11670 ;
  assign w11672 = w37 | w11671 ;
  assign w11673 = w3098 & w9977 ;
  assign w11674 = ( ~w11671 & w11672 ) | ( ~w11671 & w11673 ) | ( w11672 & w11673 ) ;
  assign w11675 = ( \pi29 & \pi30 ) | ( \pi29 & ~w9973 ) | ( \pi30 & ~w9973 ) ;
  assign w11676 = \pi31 | w11675 ;
  assign w11677 = ( \pi29 & ~\pi30 ) | ( \pi29 & w9975 ) | ( ~\pi30 & w9975 ) ;
  assign w11678 = ( \pi29 & \pi31 ) | ( \pi29 & ~w11677 ) | ( \pi31 & ~w11677 ) ;
  assign w11679 = ( w11674 & w11676 ) | ( w11674 & ~w11678 ) | ( w11676 & ~w11678 ) ;
  assign w11680 = ( w11468 & ~w11669 ) | ( w11468 & w11679 ) | ( ~w11669 & w11679 ) ;
  assign w11681 = ( w11468 & ~w11579 ) | ( w11468 & w11680 ) | ( ~w11579 & w11680 ) ;
  assign w11682 = ( w11521 & ~w11523 ) | ( w11521 & w11681 ) | ( ~w11523 & w11681 ) ;
  assign w11683 = w11499 ^ w11509 ;
  assign w11684 = w11058 ^ w11683 ;
  assign w11685 = w3549 & w9957 ;
  assign w11686 = ( w3717 & ~w9963 ) | ( w3717 & w11685 ) | ( ~w9963 & w11685 ) ;
  assign w11687 = w3649 | w11686 ;
  assign w11688 = ( w9961 & w11686 ) | ( w9961 & w11687 ) | ( w11686 & w11687 ) ;
  assign w11689 = w11685 | w11688 ;
  assign w11690 = w3448 | w11089 ;
  assign w11691 = ( ~w11089 & w11689 ) | ( ~w11089 & w11690 ) | ( w11689 & w11690 ) ;
  assign w11692 = \pi29 ^ w11691 ;
  assign w11693 = ( w11682 & w11684 ) | ( w11682 & w11692 ) | ( w11684 & w11692 ) ;
  assign w11694 = ( w11427 & w11510 ) | ( w11427 & ~w11693 ) | ( w11510 & ~w11693 ) ;
  assign w11695 = ( w11417 & w11425 ) | ( w11417 & ~w11694 ) | ( w11425 & ~w11694 ) ;
  assign w11696 = w11352 ^ w11354 ;
  assign w11697 = w11362 ^ w11696 ;
  assign w11698 = ~w4143 & w10211 ;
  assign w11699 = w4052 & w10114 ;
  assign w11700 = ( w10211 & ~w11698 ) | ( w10211 & w11699 ) | ( ~w11698 & w11699 ) ;
  assign w11701 = ~w4147 & w10789 ;
  assign w11702 = w10784 | w11700 ;
  assign w11703 = ( w3964 & w11700 ) | ( w3964 & w11702 ) | ( w11700 & w11702 ) ;
  assign w11704 = ( w10789 & ~w11701 ) | ( w10789 & w11703 ) | ( ~w11701 & w11703 ) ;
  assign w11705 = \pi26 ^ w11704 ;
  assign w11706 = ( w11695 & w11697 ) | ( w11695 & w11705 ) | ( w11697 & w11705 ) ;
  assign w11707 = ~w4651 & w10801 ;
  assign w11708 = w4606 & ~w10807 ;
  assign w11709 = ( w10801 & ~w11707 ) | ( w10801 & w11708 ) | ( ~w11707 & w11708 ) ;
  assign w11710 = w4706 | w10866 ;
  assign w11711 = w10874 | w11709 ;
  assign w11712 = ( w4609 & w11709 ) | ( w4609 & w11711 ) | ( w11709 & w11711 ) ;
  assign w11713 = ( ~w10866 & w11710 ) | ( ~w10866 & w11712 ) | ( w11710 & w11712 ) ;
  assign w11714 = \pi23 ^ w11713 ;
  assign w11715 = ( ~w11415 & w11706 ) | ( ~w11415 & w11714 ) | ( w11706 & w11714 ) ;
  assign w11716 = ( w11405 & w11413 ) | ( w11405 & w11715 ) | ( w11413 & w11715 ) ;
  assign w11717 = w5343 | w11139 ;
  assign w11718 = w4905 & w10883 ;
  assign w11719 = ( ~w11139 & w11717 ) | ( ~w11139 & w11718 ) | ( w11717 & w11718 ) ;
  assign w11720 = w5395 | w10738 ;
  assign w11721 = w11145 & ~w11719 ;
  assign w11722 = ( w4908 & w11719 ) | ( w4908 & ~w11721 ) | ( w11719 & ~w11721 ) ;
  assign w11723 = ( ~w10738 & w11720 ) | ( ~w10738 & w11722 ) | ( w11720 & w11722 ) ;
  assign w11724 = \pi20 ^ w11723 ;
  assign w11725 = ( ~w11403 & w11716 ) | ( ~w11403 & w11724 ) | ( w11716 & w11724 ) ;
  assign w11726 = w11403 ^ w11716 ;
  assign w11727 = w11724 ^ w11726 ;
  assign w11728 = w11415 ^ w11706 ;
  assign w11729 = w11714 ^ w11728 ;
  assign w11730 = w11695 ^ w11697 ;
  assign w11731 = w11705 ^ w11730 ;
  assign w11732 = w11417 ^ w11694 ;
  assign w11733 = w11425 ^ w11732 ;
  assign w11734 = ~w4143 & w10114 ;
  assign w11735 = w4052 & w9953 ;
  assign w11736 = ( w10114 & ~w11734 ) | ( w10114 & w11735 ) | ( ~w11734 & w11735 ) ;
  assign w11737 = ~w4147 & w10214 ;
  assign w11738 = w10211 | w11736 ;
  assign w11739 = ( w3964 & w11736 ) | ( w3964 & w11738 ) | ( w11736 & w11738 ) ;
  assign w11740 = ( w10214 & ~w11737 ) | ( w10214 & w11739 ) | ( ~w11737 & w11739 ) ;
  assign w11741 = \pi26 ^ w11740 ;
  assign w11742 = w11510 ^ w11693 ;
  assign w11743 = w11427 ^ w11742 ;
  assign w11744 = ~w3717 & w9957 ;
  assign w11745 = w3649 & ~w9963 ;
  assign w11746 = ( w9957 & ~w11744 ) | ( w9957 & w11745 ) | ( ~w11744 & w11745 ) ;
  assign w11747 = w3549 | w9955 ;
  assign w11748 = w11202 & ~w11746 ;
  assign w11749 = ( w3448 & w11746 ) | ( w3448 & ~w11748 ) | ( w11746 & ~w11748 ) ;
  assign w11750 = ( ~w9955 & w11747 ) | ( ~w9955 & w11749 ) | ( w11747 & w11749 ) ;
  assign w11751 = \pi29 ^ w11750 ;
  assign w11752 = ~w4143 & w9953 ;
  assign w11753 = w4052 & w9842 ;
  assign w11754 = ( w9953 & ~w11752 ) | ( w9953 & w11753 ) | ( ~w11752 & w11753 ) ;
  assign w11755 = ~w4147 & w10334 ;
  assign w11756 = w10114 | w11754 ;
  assign w11757 = ( w3964 & w11754 ) | ( w3964 & w11756 ) | ( w11754 & w11756 ) ;
  assign w11758 = ( w10334 & ~w11755 ) | ( w10334 & w11757 ) | ( ~w11755 & w11757 ) ;
  assign w11759 = \pi26 ^ w11758 ;
  assign w11760 = ( w11743 & w11751 ) | ( w11743 & w11759 ) | ( w11751 & w11759 ) ;
  assign w11761 = ( ~w11733 & w11741 ) | ( ~w11733 & w11760 ) | ( w11741 & w11760 ) ;
  assign w11762 = w4651 | w10807 ;
  assign w11763 = w4606 & ~w10805 ;
  assign w11764 = ( ~w10807 & w11762 ) | ( ~w10807 & w11763 ) | ( w11762 & w11763 ) ;
  assign w11765 = ~w4706 & w10801 ;
  assign w11766 = w10814 | w11764 ;
  assign w11767 = ( w4609 & w11764 ) | ( w4609 & w11766 ) | ( w11764 & w11766 ) ;
  assign w11768 = ( w10801 & ~w11765 ) | ( w10801 & w11767 ) | ( ~w11765 & w11767 ) ;
  assign w11769 = \pi23 ^ w11768 ;
  assign w11770 = ( w11731 & w11761 ) | ( w11731 & w11769 ) | ( w11761 & w11769 ) ;
  assign w11771 = w5343 | w10887 ;
  assign w11772 = w4905 & ~w10885 ;
  assign w11773 = ( ~w10887 & w11771 ) | ( ~w10887 & w11772 ) | ( w11771 & w11772 ) ;
  assign w11774 = ~w5395 & w10883 ;
  assign w11775 = w10895 | w11773 ;
  assign w11776 = ( w4908 & w11773 ) | ( w4908 & w11775 ) | ( w11773 & w11775 ) ;
  assign w11777 = ( w10883 & ~w11774 ) | ( w10883 & w11776 ) | ( ~w11774 & w11776 ) ;
  assign w11778 = \pi20 ^ w11777 ;
  assign w11779 = ( ~w11729 & w11770 ) | ( ~w11729 & w11778 ) | ( w11770 & w11778 ) ;
  assign w11780 = ~w5343 & w10883 ;
  assign w11781 = w4905 & ~w10887 ;
  assign w11782 = ( w10883 & ~w11780 ) | ( w10883 & w11781 ) | ( ~w11780 & w11781 ) ;
  assign w11783 = w5395 | w11139 ;
  assign w11784 = w11256 | w11782 ;
  assign w11785 = ( w4908 & w11782 ) | ( w4908 & w11784 ) | ( w11782 & w11784 ) ;
  assign w11786 = ( ~w11139 & w11783 ) | ( ~w11139 & w11785 ) | ( w11783 & w11785 ) ;
  assign w11787 = \pi20 ^ w11786 ;
  assign w11788 = w11405 ^ w11715 ;
  assign w11789 = w11413 ^ w11788 ;
  assign w11790 = ( w11779 & w11787 ) | ( w11779 & w11789 ) | ( w11787 & w11789 ) ;
  assign w11791 = w11731 ^ w11761 ;
  assign w11792 = w11769 ^ w11791 ;
  assign w11793 = w11733 ^ w11760 ;
  assign w11794 = w11741 ^ w11793 ;
  assign w11795 = w4651 | w10805 ;
  assign w11796 = w4606 & w10784 ;
  assign w11797 = ( ~w10805 & w11795 ) | ( ~w10805 & w11796 ) | ( w11795 & w11796 ) ;
  assign w11798 = w4706 | w10807 ;
  assign w11799 = w11117 | w11797 ;
  assign w11800 = ( w4609 & w11797 ) | ( w4609 & w11799 ) | ( w11797 & w11799 ) ;
  assign w11801 = ( ~w10807 & w11798 ) | ( ~w10807 & w11800 ) | ( w11798 & w11800 ) ;
  assign w11802 = \pi23 ^ w11801 ;
  assign w11803 = w11743 ^ w11759 ;
  assign w11804 = w11751 ^ w11803 ;
  assign w11805 = w11468 ^ w11680 ;
  assign w11806 = w11579 ^ w11805 ;
  assign w11807 = ( ~w9973 & w9975 ) | ( ~w9973 & w10038 ) | ( w9975 & w10038 ) ;
  assign w11808 = w9973 ^ w11807 ;
  assign w11809 = w9971 ^ w11808 ;
  assign w11810 = ( \pi29 & \pi31 ) | ( \pi29 & ~w9973 ) | ( \pi31 & ~w9973 ) ;
  assign w11811 = ( \pi29 & ~\pi30 ) | ( \pi29 & w11810 ) | ( ~\pi30 & w11810 ) ;
  assign w11812 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w11810 ) | ( \pi30 & w11810 ) ;
  assign w11813 = ( ~\pi29 & w9975 ) | ( ~\pi29 & w11812 ) | ( w9975 & w11812 ) ;
  assign w11814 = ( w9971 & w11812 ) | ( w9971 & ~w11813 ) | ( w11812 & ~w11813 ) ;
  assign w11815 = ~\pi31 & w11814 ;
  assign w11816 = ( w11811 & w11813 ) | ( w11811 & w11815 ) | ( w11813 & w11815 ) ;
  assign w11817 = ( w37 & ~w11809 ) | ( w37 & w11816 ) | ( ~w11809 & w11816 ) ;
  assign w11818 = w11816 | w11817 ;
  assign w11819 = w3549 & w9961 ;
  assign w11820 = ( w3717 & w9965 ) | ( w3717 & w11819 ) | ( w9965 & w11819 ) ;
  assign w11821 = w3649 | w11820 ;
  assign w11822 = ( ~w9967 & w11820 ) | ( ~w9967 & w11821 ) | ( w11820 & w11821 ) ;
  assign w11823 = w11819 | w11822 ;
  assign w11824 = ~w3448 & w11339 ;
  assign w11825 = ( w11339 & w11823 ) | ( w11339 & ~w11824 ) | ( w11823 & ~w11824 ) ;
  assign w11826 = \pi29 ^ w11825 ;
  assign w11827 = ( ~w11806 & w11818 ) | ( ~w11806 & w11826 ) | ( w11818 & w11826 ) ;
  assign w11828 = w11523 ^ w11681 ;
  assign w11829 = w11521 ^ w11828 ;
  assign w11830 = ~w3717 & w9961 ;
  assign w11831 = w3649 & w9965 ;
  assign w11832 = ( w9961 & ~w11830 ) | ( w9961 & w11831 ) | ( ~w11830 & w11831 ) ;
  assign w11833 = w3549 | w9963 ;
  assign w11834 = w11278 & ~w11832 ;
  assign w11835 = ( w3448 & w11832 ) | ( w3448 & ~w11834 ) | ( w11832 & ~w11834 ) ;
  assign w11836 = ( ~w9963 & w11833 ) | ( ~w9963 & w11835 ) | ( w11833 & w11835 ) ;
  assign w11837 = \pi29 ^ w11836 ;
  assign w11838 = ( w11827 & ~w11829 ) | ( w11827 & w11837 ) | ( ~w11829 & w11837 ) ;
  assign w11839 = w11682 ^ w11684 ;
  assign w11840 = w11692 ^ w11839 ;
  assign w11841 = ~w4143 & w9842 ;
  assign w11842 = w4052 & ~w9955 ;
  assign w11843 = ( w9842 & ~w11841 ) | ( w9842 & w11842 ) | ( ~w11841 & w11842 ) ;
  assign w11844 = ~w4147 & w10965 ;
  assign w11845 = w9953 | w11843 ;
  assign w11846 = ( w3964 & w11843 ) | ( w3964 & w11845 ) | ( w11843 & w11845 ) ;
  assign w11847 = ( w10965 & ~w11844 ) | ( w10965 & w11846 ) | ( ~w11844 & w11846 ) ;
  assign w11848 = \pi26 ^ w11847 ;
  assign w11849 = ( w11838 & w11840 ) | ( w11838 & w11848 ) | ( w11840 & w11848 ) ;
  assign w11850 = ~w4651 & w10784 ;
  assign w11851 = w4606 & w10211 ;
  assign w11852 = ( w10784 & ~w11850 ) | ( w10784 & w11851 ) | ( ~w11850 & w11851 ) ;
  assign w11853 = w4706 | w10805 ;
  assign w11854 = w10855 & ~w11852 ;
  assign w11855 = ( w4609 & w11852 ) | ( w4609 & ~w11854 ) | ( w11852 & ~w11854 ) ;
  assign w11856 = ( ~w10805 & w11853 ) | ( ~w10805 & w11855 ) | ( w11853 & w11855 ) ;
  assign w11857 = \pi23 ^ w11856 ;
  assign w11858 = ( w11804 & w11849 ) | ( w11804 & w11857 ) | ( w11849 & w11857 ) ;
  assign w11859 = ( ~w11794 & w11802 ) | ( ~w11794 & w11858 ) | ( w11802 & w11858 ) ;
  assign w11860 = w5343 | w10885 ;
  assign w11861 = w4905 & ~w10866 ;
  assign w11862 = ( ~w10885 & w11860 ) | ( ~w10885 & w11861 ) | ( w11860 & w11861 ) ;
  assign w11863 = w5395 | w10887 ;
  assign w11864 = w11131 & ~w11862 ;
  assign w11865 = ( w4908 & w11862 ) | ( w4908 & ~w11864 ) | ( w11862 & ~w11864 ) ;
  assign w11866 = ( ~w10887 & w11863 ) | ( ~w10887 & w11865 ) | ( w11863 & w11865 ) ;
  assign w11867 = \pi20 ^ w11866 ;
  assign w11868 = ( w11792 & w11859 ) | ( w11792 & w11867 ) | ( w11859 & w11867 ) ;
  assign w11869 = ( w5494 & w5710 ) | ( w5494 & ~w11138 ) | ( w5710 & ~w11138 ) ;
  assign w11870 = w5710 & ~w11869 ;
  assign w11871 = ( w5948 & ~w11869 ) | ( w5948 & w11870 ) | ( ~w11869 & w11870 ) ;
  assign w11872 = ( ~w10738 & w11869 ) | ( ~w10738 & w11871 ) | ( w11869 & w11871 ) ;
  assign w11873 = w11729 ^ w11770 ;
  assign w11874 = w11778 ^ w11873 ;
  assign w11875 = w11146 & ~w11872 ;
  assign w11876 = ( w5497 & w11872 ) | ( w5497 & ~w11875 ) | ( w11872 & ~w11875 ) ;
  assign w11877 = \pi17 ^ w11876 ;
  assign w11878 = ( w11868 & ~w11874 ) | ( w11868 & w11877 ) | ( ~w11874 & w11877 ) ;
  assign w11879 = w11779 ^ w11789 ;
  assign w11880 = w11787 ^ w11879 ;
  assign w11881 = w5497 & w11146 ;
  assign w11882 = ( w5497 & w11872 ) | ( w5497 & ~w11881 ) | ( w11872 & ~w11881 ) ;
  assign w11883 = w11868 ^ w11882 ;
  assign w11884 = \pi17 ^ w11874 ;
  assign w11885 = w11883 ^ w11884 ;
  assign w11886 = w11792 ^ w11859 ;
  assign w11887 = w11867 ^ w11886 ;
  assign w11888 = w11794 ^ w11858 ;
  assign w11889 = w11802 ^ w11888 ;
  assign w11890 = w5343 | w10866 ;
  assign w11891 = w4905 & w10801 ;
  assign w11892 = ( ~w10866 & w11890 ) | ( ~w10866 & w11891 ) | ( w11890 & w11891 ) ;
  assign w11893 = w5395 | w10885 ;
  assign w11894 = w11160 & ~w11892 ;
  assign w11895 = ( w4908 & w11892 ) | ( w4908 & ~w11894 ) | ( w11892 & ~w11894 ) ;
  assign w11896 = ( ~w10885 & w11893 ) | ( ~w10885 & w11895 ) | ( w11893 & w11895 ) ;
  assign w11897 = \pi20 ^ w11896 ;
  assign w11898 = w11804 ^ w11849 ;
  assign w11899 = w11857 ^ w11898 ;
  assign w11900 = w11838 ^ w11840 ;
  assign w11901 = w11848 ^ w11900 ;
  assign w11902 = w11827 ^ w11829 ;
  assign w11903 = w11837 ^ w11902 ;
  assign w11904 = w4143 | w9955 ;
  assign w11905 = w4052 & w9957 ;
  assign w11906 = ( ~w9955 & w11904 ) | ( ~w9955 & w11905 ) | ( w11904 & w11905 ) ;
  assign w11907 = w4147 | w10976 ;
  assign w11908 = w9842 | w11906 ;
  assign w11909 = ( w3964 & w11906 ) | ( w3964 & w11908 ) | ( w11906 & w11908 ) ;
  assign w11910 = ( ~w10976 & w11907 ) | ( ~w10976 & w11909 ) | ( w11907 & w11909 ) ;
  assign w11911 = \pi26 ^ w11910 ;
  assign w11912 = ( w9977 & w9979 ) | ( w9977 & w10036 ) | ( w9979 & w10036 ) ;
  assign w11913 = w9977 ^ w11912 ;
  assign w11914 = w9975 ^ w11913 ;
  assign w11915 = ( \pi29 & \pi31 ) | ( \pi29 & w9977 ) | ( \pi31 & w9977 ) ;
  assign w11916 = ( \pi29 & ~\pi30 ) | ( \pi29 & w11915 ) | ( ~\pi30 & w11915 ) ;
  assign w11917 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w11915 ) | ( \pi30 & w11915 ) ;
  assign w11918 = ( ~\pi29 & w9979 ) | ( ~\pi29 & w11917 ) | ( w9979 & w11917 ) ;
  assign w11919 = ( w9975 & w11917 ) | ( w9975 & ~w11918 ) | ( w11917 & ~w11918 ) ;
  assign w11920 = ~\pi31 & w11919 ;
  assign w11921 = ( w11916 & w11918 ) | ( w11916 & w11920 ) | ( w11918 & w11920 ) ;
  assign w11922 = ( w37 & w11914 ) | ( w37 & w11921 ) | ( w11914 & w11921 ) ;
  assign w11923 = w11921 | w11922 ;
  assign w11924 = w269 | w312 ;
  assign w11925 = w230 | w11924 ;
  assign w11926 = ( ~w230 & w232 ) | ( ~w230 & w1154 ) | ( w232 & w1154 ) ;
  assign w11927 = w11925 | w11926 ;
  assign w11928 = w901 | w1165 ;
  assign w11929 = ( w674 & ~w1165 ) | ( w674 & w11927 ) | ( ~w1165 & w11927 ) ;
  assign w11930 = w11928 | w11929 ;
  assign w11931 = ( ~w63 & w2872 ) | ( ~w63 & w11930 ) | ( w2872 & w11930 ) ;
  assign w11932 = w2022 & ~w3673 ;
  assign w11933 = ( w63 & w199 ) | ( w63 & ~w3673 ) | ( w199 & ~w3673 ) ;
  assign w11934 = w11932 & ~w11933 ;
  assign w11935 = ~w11931 & w11934 ;
  assign w11936 = ( w160 & w468 ) | ( w160 & ~w2253 ) | ( w468 & ~w2253 ) ;
  assign w11937 = ~w1917 & w11935 ;
  assign w11938 = ( w421 & w2253 ) | ( w421 & w11935 ) | ( w2253 & w11935 ) ;
  assign w11939 = w11937 & ~w11938 ;
  assign w11940 = ~w11936 & w11939 ;
  assign w11941 = ( w215 & w263 ) | ( w215 & ~w271 ) | ( w263 & ~w271 ) ;
  assign w11942 = ~w176 & w11940 ;
  assign w11943 = ( ~w176 & w271 ) | ( ~w176 & w560 ) | ( w271 & w560 ) ;
  assign w11944 = w11942 & ~w11943 ;
  assign w11945 = ~w11941 & w11944 ;
  assign w11946 = \pi02 ^ w10738 ;
  assign w11947 = \pi01 | w10738 ;
  assign w11948 = ( \pi00 & ~w11946 ) | ( \pi00 & w11947 ) | ( ~w11946 & w11947 ) ;
  assign w11949 = ~w11946 & w11948 ;
  assign w11950 = ( w221 & w229 ) | ( w221 & ~w509 ) | ( w229 & ~w509 ) ;
  assign w11951 = w101 | w133 ;
  assign w11952 = ( ~w133 & w509 ) | ( ~w133 & w640 ) | ( w509 & w640 ) ;
  assign w11953 = w11951 | w11952 ;
  assign w11954 = w11950 | w11953 ;
  assign w11955 = w257 | w317 ;
  assign w11956 = w3653 | w11955 ;
  assign w11957 = ( w432 & ~w3653 ) | ( w432 & w11954 ) | ( ~w3653 & w11954 ) ;
  assign w11958 = w11956 | w11957 ;
  assign w11959 = ( ~w139 & w392 ) | ( ~w139 & w11958 ) | ( w392 & w11958 ) ;
  assign w11960 = w139 | w11959 ;
  assign w11961 = ( w488 & w783 ) | ( w488 & ~w980 ) | ( w783 & ~w980 ) ;
  assign w11962 = w142 | w11960 ;
  assign w11963 = ( ~w142 & w980 ) | ( ~w142 & w1030 ) | ( w980 & w1030 ) ;
  assign w11964 = w11962 | w11963 ;
  assign w11965 = w11961 | w11964 ;
  assign w11966 = w283 | w11537 ;
  assign w11967 = ( w206 & w2782 ) | ( w206 & ~w11537 ) | ( w2782 & ~w11537 ) ;
  assign w11968 = w11966 | w11967 ;
  assign w11969 = w258 | w314 ;
  assign w11970 = w1565 | w11969 ;
  assign w11971 = ( w122 & w784 ) | ( w122 & ~w1565 ) | ( w784 & ~w1565 ) ;
  assign w11972 = w11970 | w11971 ;
  assign w11973 = w356 | w567 ;
  assign w11974 = ( w74 & ~w356 ) | ( w74 & w11972 ) | ( ~w356 & w11972 ) ;
  assign w11975 = w11973 | w11974 ;
  assign w11976 = ( w276 & ~w1835 ) | ( w276 & w11968 ) | ( ~w1835 & w11968 ) ;
  assign w11977 = w2713 | w11975 ;
  assign w11978 = ( w1835 & w10154 ) | ( w1835 & ~w11975 ) | ( w10154 & ~w11975 ) ;
  assign w11979 = w11977 | w11978 ;
  assign w11980 = w11976 | w11979 ;
  assign w11981 = w409 | w11980 ;
  assign w11982 = ( w1421 & w11965 ) | ( w1421 & ~w11980 ) | ( w11965 & ~w11980 ) ;
  assign w11983 = w11981 | w11982 ;
  assign w11984 = ( w103 & ~w104 ) | ( w103 & w507 ) | ( ~w104 & w507 ) ;
  assign w11985 = w5859 | w6309 ;
  assign w11986 = ( w104 & w1031 ) | ( w104 & ~w6309 ) | ( w1031 & ~w6309 ) ;
  assign w11987 = w11985 | w11986 ;
  assign w11988 = w11984 | w11987 ;
  assign w11989 = w1560 | w11988 ;
  assign w11990 = w11440 & ~w11989 ;
  assign w11991 = ( w9875 & w11440 ) | ( w9875 & w11983 ) | ( w11440 & w11983 ) ;
  assign w11992 = w11990 & ~w11991 ;
  assign w11993 = ( w203 & w223 ) | ( w203 & ~w224 ) | ( w223 & ~w224 ) ;
  assign w11994 = ~w144 & w11992 ;
  assign w11995 = ( ~w144 & w224 ) | ( ~w144 & w626 ) | ( w224 & w626 ) ;
  assign w11996 = w11994 & ~w11995 ;
  assign w11997 = ~w11993 & w11996 ;
  assign w11998 = w84 | w531 ;
  assign w11999 = ( w84 & ~w339 ) | ( w84 & w11997 ) | ( ~w339 & w11997 ) ;
  assign w12000 = ~w11998 & w11999 ;
  assign w12001 = w11949 ^ w12000 ;
  assign w12002 = ( ~\pi02 & \pi03 ) | ( ~\pi02 & \pi04 ) | ( \pi03 & \pi04 ) ;
  assign w12003 = ( \pi02 & ~\pi05 ) | ( \pi02 & w12002 ) | ( ~\pi05 & w12002 ) ;
  assign w12004 = w10738 ^ w12003 ;
  assign w12005 = ( \pi05 & w12003 ) | ( \pi05 & w12004 ) | ( w12003 & w12004 ) ;
  assign w12006 = w12001 & ~w12005 ;
  assign w12007 = ( w11949 & w12000 ) | ( w11949 & ~w12006 ) | ( w12000 & ~w12006 ) ;
  assign w12008 = ~w12006 & w12007 ;
  assign w12009 = w9979 ^ w10035 ;
  assign w12010 = w9981 ^ w12009 ;
  assign w12011 = ~w37 & w12010 ;
  assign w12012 = w3098 & w9983 ;
  assign w12013 = ( w12010 & ~w12011 ) | ( w12010 & w12012 ) | ( ~w12011 & w12012 ) ;
  assign w12014 = ( \pi29 & \pi30 ) | ( \pi29 & w9979 ) | ( \pi30 & w9979 ) ;
  assign w12015 = \pi31 | w12014 ;
  assign w12016 = ( \pi29 & ~\pi30 ) | ( \pi29 & w9981 ) | ( ~\pi30 & w9981 ) ;
  assign w12017 = ( \pi29 & \pi31 ) | ( \pi29 & ~w12016 ) | ( \pi31 & ~w12016 ) ;
  assign w12018 = ( w12013 & w12015 ) | ( w12013 & ~w12017 ) | ( w12015 & ~w12017 ) ;
  assign w12019 = ( w11629 & w12008 ) | ( w11629 & ~w12018 ) | ( w12008 & ~w12018 ) ;
  assign w12020 = ( w11629 & w11945 ) | ( w11629 & w12019 ) | ( w11945 & w12019 ) ;
  assign w12021 = w11629 ^ w11668 ;
  assign w12022 = w11664 ^ w12021 ;
  assign w12023 = ( w11923 & ~w12020 ) | ( w11923 & w12022 ) | ( ~w12020 & w12022 ) ;
  assign w12024 = w11669 ^ w11679 ;
  assign w12025 = w11468 ^ w12024 ;
  assign w12026 = w3549 & w9965 ;
  assign w12027 = ( w3717 & ~w9967 ) | ( w3717 & w12026 ) | ( ~w9967 & w12026 ) ;
  assign w12028 = w3649 | w12027 ;
  assign w12029 = ( w9971 & w12027 ) | ( w9971 & w12028 ) | ( w12027 & w12028 ) ;
  assign w12030 = w12026 | w12029 ;
  assign w12031 = w3448 | w11501 ;
  assign w12032 = ( ~w11501 & w12030 ) | ( ~w11501 & w12031 ) | ( w12030 & w12031 ) ;
  assign w12033 = \pi29 ^ w12032 ;
  assign w12034 = ( w12023 & ~w12025 ) | ( w12023 & w12033 ) | ( ~w12025 & w12033 ) ;
  assign w12035 = w11806 ^ w11826 ;
  assign w12036 = w11818 ^ w12035 ;
  assign w12037 = ~w4143 & w9957 ;
  assign w12038 = w4052 & ~w9963 ;
  assign w12039 = ( w9957 & ~w12037 ) | ( w9957 & w12038 ) | ( ~w12037 & w12038 ) ;
  assign w12040 = w4147 | w11202 ;
  assign w12041 = w9955 & ~w12039 ;
  assign w12042 = ( w3964 & w12039 ) | ( w3964 & ~w12041 ) | ( w12039 & ~w12041 ) ;
  assign w12043 = ( ~w11202 & w12040 ) | ( ~w11202 & w12042 ) | ( w12040 & w12042 ) ;
  assign w12044 = \pi26 ^ w12043 ;
  assign w12045 = ( w12034 & ~w12036 ) | ( w12034 & w12044 ) | ( ~w12036 & w12044 ) ;
  assign w12046 = ( ~w11903 & w11911 ) | ( ~w11903 & w12045 ) | ( w11911 & w12045 ) ;
  assign w12047 = ~w4651 & w10211 ;
  assign w12048 = w4606 & w10114 ;
  assign w12049 = ( w10211 & ~w12047 ) | ( w10211 & w12048 ) | ( ~w12047 & w12048 ) ;
  assign w12050 = ~w4706 & w10784 ;
  assign w12051 = w10789 | w12049 ;
  assign w12052 = ( w4609 & w12049 ) | ( w4609 & w12051 ) | ( w12049 & w12051 ) ;
  assign w12053 = ( w10784 & ~w12050 ) | ( w10784 & w12052 ) | ( ~w12050 & w12052 ) ;
  assign w12054 = \pi23 ^ w12053 ;
  assign w12055 = ( w11901 & w12046 ) | ( w11901 & w12054 ) | ( w12046 & w12054 ) ;
  assign w12056 = ~w5343 & w10801 ;
  assign w12057 = w4905 & ~w10807 ;
  assign w12058 = ( w10801 & ~w12056 ) | ( w10801 & w12057 ) | ( ~w12056 & w12057 ) ;
  assign w12059 = w5395 | w10866 ;
  assign w12060 = w10874 | w12058 ;
  assign w12061 = ( w4908 & w12058 ) | ( w4908 & w12060 ) | ( w12058 & w12060 ) ;
  assign w12062 = ( ~w10866 & w12059 ) | ( ~w10866 & w12061 ) | ( w12059 & w12061 ) ;
  assign w12063 = \pi20 ^ w12062 ;
  assign w12064 = ( w11899 & w12055 ) | ( w11899 & w12063 ) | ( w12055 & w12063 ) ;
  assign w12065 = ( ~w11889 & w11897 ) | ( ~w11889 & w12064 ) | ( w11897 & w12064 ) ;
  assign w12066 = w5710 | w11139 ;
  assign w12067 = w5494 & w10883 ;
  assign w12068 = ( ~w11139 & w12066 ) | ( ~w11139 & w12067 ) | ( w12066 & w12067 ) ;
  assign w12069 = w5948 | w10738 ;
  assign w12070 = w11145 & ~w12068 ;
  assign w12071 = ( w5497 & w12068 ) | ( w5497 & ~w12070 ) | ( w12068 & ~w12070 ) ;
  assign w12072 = ( ~w10738 & w12069 ) | ( ~w10738 & w12071 ) | ( w12069 & w12071 ) ;
  assign w12073 = \pi17 ^ w12072 ;
  assign w12074 = ( w11887 & w12065 ) | ( w11887 & w12073 ) | ( w12065 & w12073 ) ;
  assign w12075 = w11887 ^ w12065 ;
  assign w12076 = w12073 ^ w12075 ;
  assign w12077 = w11899 ^ w12055 ;
  assign w12078 = w12063 ^ w12077 ;
  assign w12079 = w11901 ^ w12046 ;
  assign w12080 = w12054 ^ w12079 ;
  assign w12081 = w11903 ^ w12045 ;
  assign w12082 = w11911 ^ w12081 ;
  assign w12083 = ~w4651 & w10114 ;
  assign w12084 = w4606 & w9953 ;
  assign w12085 = ( w10114 & ~w12083 ) | ( w10114 & w12084 ) | ( ~w12083 & w12084 ) ;
  assign w12086 = ~w4706 & w10211 ;
  assign w12087 = w10214 | w12085 ;
  assign w12088 = ( w4609 & w12085 ) | ( w4609 & w12087 ) | ( w12085 & w12087 ) ;
  assign w12089 = ( w10211 & ~w12086 ) | ( w10211 & w12088 ) | ( ~w12086 & w12088 ) ;
  assign w12090 = \pi23 ^ w12089 ;
  assign w12091 = w12034 ^ w12036 ;
  assign w12092 = w12044 ^ w12091 ;
  assign w12093 = w12020 ^ w12022 ;
  assign w12094 = w11923 ^ w12093 ;
  assign w12095 = ~w3717 & w9971 ;
  assign w12096 = w3649 & ~w9973 ;
  assign w12097 = ( w9971 & ~w12095 ) | ( w9971 & w12096 ) | ( ~w12095 & w12096 ) ;
  assign w12098 = w3549 | w9967 ;
  assign w12099 = w11512 & ~w12097 ;
  assign w12100 = ( w3448 & w12097 ) | ( w3448 & ~w12099 ) | ( w12097 & ~w12099 ) ;
  assign w12101 = ( ~w9967 & w12098 ) | ( ~w9967 & w12100 ) | ( w12098 & w12100 ) ;
  assign w12102 = \pi29 ^ w12101 ;
  assign w12103 = w11629 ^ w12019 ;
  assign w12104 = w11945 ^ w12103 ;
  assign w12105 = w9977 ^ w10036 ;
  assign w12106 = w9979 ^ w12105 ;
  assign w12107 = ( \pi29 & \pi31 ) | ( \pi29 & w9979 ) | ( \pi31 & w9979 ) ;
  assign w12108 = ( \pi29 & ~\pi30 ) | ( \pi29 & w12107 ) | ( ~\pi30 & w12107 ) ;
  assign w12109 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w12107 ) | ( \pi30 & w12107 ) ;
  assign w12110 = ( ~\pi29 & w9981 ) | ( ~\pi29 & w12109 ) | ( w9981 & w12109 ) ;
  assign w12111 = ( w9977 & w12109 ) | ( w9977 & ~w12110 ) | ( w12109 & ~w12110 ) ;
  assign w12112 = ~\pi31 & w12111 ;
  assign w12113 = ( w12108 & w12110 ) | ( w12108 & w12112 ) | ( w12110 & w12112 ) ;
  assign w12114 = ( w37 & w12106 ) | ( w37 & w12113 ) | ( w12106 & w12113 ) ;
  assign w12115 = w12113 | w12114 ;
  assign w12116 = ( w169 & ~w593 ) | ( w169 & w1955 ) | ( ~w593 & w1955 ) ;
  assign w12117 = w216 | w956 ;
  assign w12118 = ( w593 & ~w956 ) | ( w593 & w1274 ) | ( ~w956 & w1274 ) ;
  assign w12119 = w12117 | w12118 ;
  assign w12120 = w12116 | w12119 ;
  assign w12121 = ( w2915 & w5602 ) | ( w2915 & ~w12120 ) | ( w5602 & ~w12120 ) ;
  assign w12122 = w3776 | w3837 ;
  assign w12123 = ( w1206 & ~w3837 ) | ( w1206 & w12120 ) | ( ~w3837 & w12120 ) ;
  assign w12124 = w12122 | w12123 ;
  assign w12125 = w12121 | w12124 ;
  assign w12126 = ( w359 & ~w466 ) | ( w359 & w512 ) | ( ~w466 & w512 ) ;
  assign w12127 = w280 | w12125 ;
  assign w12128 = ( ~w280 & w512 ) | ( ~w280 & w1126 ) | ( w512 & w1126 ) ;
  assign w12129 = w12127 | w12128 ;
  assign w12130 = w12126 & ~w12129 ;
  assign w12131 = ( w277 & w524 ) | ( w277 & ~w595 ) | ( w524 & ~w595 ) ;
  assign w12132 = ~w127 & w12130 ;
  assign w12133 = ( ~w127 & w595 ) | ( ~w127 & w1130 ) | ( w595 & w1130 ) ;
  assign w12134 = w12132 & ~w12133 ;
  assign w12135 = ~w12131 & w12134 ;
  assign w12136 = w98 | w312 ;
  assign w12137 = ( ~w98 & w113 ) | ( ~w98 & w638 ) | ( w113 & w638 ) ;
  assign w12138 = w12136 | w12137 ;
  assign w12139 = ( w1759 & w10347 ) | ( w1759 & ~w12138 ) | ( w10347 & ~w12138 ) ;
  assign w12140 = w12138 | w12139 ;
  assign w12141 = ( ~w225 & w1977 ) | ( ~w225 & w12140 ) | ( w1977 & w12140 ) ;
  assign w12142 = w503 | w11983 ;
  assign w12143 = ( w225 & ~w503 ) | ( w225 & w511 ) | ( ~w503 & w511 ) ;
  assign w12144 = w12142 | w12143 ;
  assign w12145 = w12141 | w12144 ;
  assign w12146 = w1208 | w1837 ;
  assign w12147 = w741 | w12146 ;
  assign w12148 = ( w267 & ~w741 ) | ( w267 & w12145 ) | ( ~w741 & w12145 ) ;
  assign w12149 = w12147 | w12148 ;
  assign w12150 = w218 | w758 ;
  assign w12151 = w177 | w12150 ;
  assign w12152 = ( ~w177 & w4174 ) | ( ~w177 & w12149 ) | ( w4174 & w12149 ) ;
  assign w12153 = w12151 | w12152 ;
  assign w12154 = ( w320 & w449 ) | ( w320 & ~w897 ) | ( w449 & ~w897 ) ;
  assign w12155 = w167 | w12153 ;
  assign w12156 = ( ~w167 & w897 ) | ( ~w167 & w901 ) | ( w897 & w901 ) ;
  assign w12157 = w12155 | w12156 ;
  assign w12158 = w12154 | w12157 ;
  assign w12159 = ( w413 & w459 ) | ( w413 & ~w724 ) | ( w459 & ~w724 ) ;
  assign w12160 = w253 | w260 ;
  assign w12161 = ( ~w260 & w724 ) | ( ~w260 & w980 ) | ( w724 & w980 ) ;
  assign w12162 = w12160 | w12161 ;
  assign w12163 = w12159 | w12162 ;
  assign w12164 = w429 | w593 ;
  assign w12165 = ( ~w429 & w571 ) | ( ~w429 & w12163 ) | ( w571 & w12163 ) ;
  assign w12166 = w12164 | w12165 ;
  assign w12167 = ( w351 & w352 ) | ( w351 & ~w606 ) | ( w352 & ~w606 ) ;
  assign w12168 = w118 | w350 ;
  assign w12169 = ( ~w350 & w606 ) | ( ~w350 & w697 ) | ( w606 & w697 ) ;
  assign w12170 = w12168 | w12169 ;
  assign w12171 = w12167 | w12170 ;
  assign w12172 = ( w2452 & w5039 ) | ( w2452 & ~w9905 ) | ( w5039 & ~w9905 ) ;
  assign w12173 = w1778 | w12166 ;
  assign w12174 = ( w9905 & ~w12166 ) | ( w9905 & w12171 ) | ( ~w12166 & w12171 ) ;
  assign w12175 = w12173 | w12174 ;
  assign w12176 = w12172 | w12175 ;
  assign w12177 = ( w257 & w431 ) | ( w257 & ~w628 ) | ( w431 & ~w628 ) ;
  assign w12178 = w120 | w12176 ;
  assign w12179 = ( ~w120 & w628 ) | ( ~w120 & w1229 ) | ( w628 & w1229 ) ;
  assign w12180 = w12178 | w12179 ;
  assign w12181 = w12177 | w12180 ;
  assign w12182 = w278 | w341 ;
  assign w12183 = w1741 | w12182 ;
  assign w12184 = ( w139 & ~w1741 ) | ( w139 & w12181 ) | ( ~w1741 & w12181 ) ;
  assign w12185 = w12183 | w12184 ;
  assign w12186 = ( ~w531 & w1130 ) | ( ~w531 & w12185 ) | ( w1130 & w12185 ) ;
  assign w12187 = w531 | w12186 ;
  assign w12188 = ( w422 & w533 ) | ( w422 & ~w758 ) | ( w533 & ~w758 ) ;
  assign w12189 = w115 | w209 ;
  assign w12190 = ( ~w209 & w758 ) | ( ~w209 & w1340 ) | ( w758 & w1340 ) ;
  assign w12191 = w12189 | w12190 ;
  assign w12192 = w12188 | w12191 ;
  assign w12193 = w223 | w951 ;
  assign w12194 = w122 | w12193 ;
  assign w12195 = ( ~w122 & w178 ) | ( ~w122 & w12192 ) | ( w178 & w12192 ) ;
  assign w12196 = w12194 | w12195 ;
  assign w12197 = w443 | w470 ;
  assign w12198 = w161 | w12197 ;
  assign w12199 = ( ~w161 & w310 ) | ( ~w161 & w1565 ) | ( w310 & w1565 ) ;
  assign w12200 = w12198 | w12199 ;
  assign w12201 = ~w1813 & w2949 ;
  assign w12202 = ~w12196 & w12201 ;
  assign w12203 = ( w10306 & ~w12196 ) | ( w10306 & w12200 ) | ( ~w12196 & w12200 ) ;
  assign w12204 = w12202 & ~w12203 ;
  assign w12205 = ( ~w76 & w1265 ) | ( ~w76 & w11537 ) | ( w1265 & w11537 ) ;
  assign w12206 = ~w12187 & w12204 ;
  assign w12207 = ( w76 & w119 ) | ( w76 & w12204 ) | ( w119 & w12204 ) ;
  assign w12208 = w12206 & ~w12207 ;
  assign w12209 = ~w12205 & w12208 ;
  assign w12210 = ( w84 & w268 ) | ( w84 & ~w573 ) | ( w268 & ~w573 ) ;
  assign w12211 = ~w74 & w12209 ;
  assign w12212 = ( ~w74 & w573 ) | ( ~w74 & w595 ) | ( w573 & w595 ) ;
  assign w12213 = w12211 & ~w12212 ;
  assign w12214 = ~w12210 & w12213 ;
  assign w12215 = ( ~w9989 & w9991 ) | ( ~w9989 & w10030 ) | ( w9991 & w10030 ) ;
  assign w12216 = w9989 ^ w12215 ;
  assign w12217 = w9987 ^ w12216 ;
  assign w12218 = ( \pi29 & \pi31 ) | ( \pi29 & ~w9989 ) | ( \pi31 & ~w9989 ) ;
  assign w12219 = ( \pi29 & ~\pi30 ) | ( \pi29 & w12218 ) | ( ~\pi30 & w12218 ) ;
  assign w12220 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w12218 ) | ( \pi30 & w12218 ) ;
  assign w12221 = ( ~\pi29 & w9991 ) | ( ~\pi29 & w12220 ) | ( w9991 & w12220 ) ;
  assign w12222 = ( w9987 & w12220 ) | ( w9987 & ~w12221 ) | ( w12220 & ~w12221 ) ;
  assign w12223 = ~\pi31 & w12222 ;
  assign w12224 = ( w12219 & w12221 ) | ( w12219 & w12223 ) | ( w12221 & w12223 ) ;
  assign w12225 = ( w37 & ~w12217 ) | ( w37 & w12224 ) | ( ~w12217 & w12224 ) ;
  assign w12226 = w12224 | w12225 ;
  assign w12227 = ( w11949 & ~w12214 ) | ( w11949 & w12226 ) | ( ~w12214 & w12226 ) ;
  assign w12228 = ( w11949 & w12158 ) | ( w11949 & w12227 ) | ( w12158 & w12227 ) ;
  assign w12229 = ( w11949 & ~w12135 ) | ( w11949 & w12228 ) | ( ~w12135 & w12228 ) ;
  assign w12230 = ( \pi02 & ~\pi03 ) | ( \pi02 & \pi05 ) | ( ~\pi03 & \pi05 ) ;
  assign w12231 = ( \pi03 & ~\pi04 ) | ( \pi03 & w12230 ) | ( ~\pi04 & w12230 ) ;
  assign w12232 = \pi05 ^ w10738 ;
  assign w12233 = ( \pi04 & w12231 ) | ( \pi04 & ~w12232 ) | ( w12231 & ~w12232 ) ;
  assign w12234 = w12001 ^ w12233 ;
  assign w12235 = w9981 ^ w10034 ;
  assign w12236 = w9983 ^ w12235 ;
  assign w12237 = ( \pi29 & \pi31 ) | ( \pi29 & w9983 ) | ( \pi31 & w9983 ) ;
  assign w12238 = ( \pi29 & ~\pi30 ) | ( \pi29 & w12237 ) | ( ~\pi30 & w12237 ) ;
  assign w12239 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w12237 ) | ( \pi30 & w12237 ) ;
  assign w12240 = ( ~\pi29 & w9985 ) | ( ~\pi29 & w12239 ) | ( w9985 & w12239 ) ;
  assign w12241 = ( w9981 & w12239 ) | ( w9981 & ~w12240 ) | ( w12239 & ~w12240 ) ;
  assign w12242 = ~\pi31 & w12241 ;
  assign w12243 = ( w12238 & w12240 ) | ( w12238 & w12242 ) | ( w12240 & w12242 ) ;
  assign w12244 = ( w37 & w12236 ) | ( w37 & w12243 ) | ( w12236 & w12243 ) ;
  assign w12245 = w12243 | w12244 ;
  assign w12246 = ( w12229 & ~w12234 ) | ( w12229 & w12245 ) | ( ~w12234 & w12245 ) ;
  assign w12247 = w12008 ^ w12018 ;
  assign w12248 = w11629 ^ w12247 ;
  assign w12249 = w3549 & ~w9973 ;
  assign w12250 = ( w3717 & w9975 ) | ( w3717 & w12249 ) | ( w9975 & w12249 ) ;
  assign w12251 = w3649 | w12250 ;
  assign w12252 = ( w9977 & w12250 ) | ( w9977 & w12251 ) | ( w12250 & w12251 ) ;
  assign w12253 = w12249 | w12252 ;
  assign w12254 = w3448 | w11671 ;
  assign w12255 = ( ~w11671 & w12253 ) | ( ~w11671 & w12254 ) | ( w12253 & w12254 ) ;
  assign w12256 = \pi29 ^ w12255 ;
  assign w12257 = ( w12246 & w12248 ) | ( w12246 & w12256 ) | ( w12248 & w12256 ) ;
  assign w12258 = ( ~w12104 & w12115 ) | ( ~w12104 & w12257 ) | ( w12115 & w12257 ) ;
  assign w12259 = ( ~w12094 & w12102 ) | ( ~w12094 & w12258 ) | ( w12102 & w12258 ) ;
  assign w12260 = w12023 ^ w12025 ;
  assign w12261 = w12033 ^ w12260 ;
  assign w12262 = w4143 | w9963 ;
  assign w12263 = w4052 & w9961 ;
  assign w12264 = ( ~w9963 & w12262 ) | ( ~w9963 & w12263 ) | ( w12262 & w12263 ) ;
  assign w12265 = w4147 | w11089 ;
  assign w12266 = w9957 | w12264 ;
  assign w12267 = ( w3964 & w12264 ) | ( w3964 & w12266 ) | ( w12264 & w12266 ) ;
  assign w12268 = ( ~w11089 & w12265 ) | ( ~w11089 & w12267 ) | ( w12265 & w12267 ) ;
  assign w12269 = \pi26 ^ w12268 ;
  assign w12270 = ( w12259 & ~w12261 ) | ( w12259 & w12269 ) | ( ~w12261 & w12269 ) ;
  assign w12271 = ~w4651 & w9953 ;
  assign w12272 = w4606 & w9842 ;
  assign w12273 = ( w9953 & ~w12271 ) | ( w9953 & w12272 ) | ( ~w12271 & w12272 ) ;
  assign w12274 = ~w4706 & w10114 ;
  assign w12275 = w10334 | w12273 ;
  assign w12276 = ( w4609 & w12273 ) | ( w4609 & w12275 ) | ( w12273 & w12275 ) ;
  assign w12277 = ( w10114 & ~w12274 ) | ( w10114 & w12276 ) | ( ~w12274 & w12276 ) ;
  assign w12278 = \pi23 ^ w12277 ;
  assign w12279 = ( ~w12092 & w12270 ) | ( ~w12092 & w12278 ) | ( w12270 & w12278 ) ;
  assign w12280 = ( ~w12082 & w12090 ) | ( ~w12082 & w12279 ) | ( w12090 & w12279 ) ;
  assign w12281 = w5343 | w10807 ;
  assign w12282 = w4905 & ~w10805 ;
  assign w12283 = ( ~w10807 & w12281 ) | ( ~w10807 & w12282 ) | ( w12281 & w12282 ) ;
  assign w12284 = ~w5395 & w10801 ;
  assign w12285 = w10814 | w12283 ;
  assign w12286 = ( w4908 & w12283 ) | ( w4908 & w12285 ) | ( w12283 & w12285 ) ;
  assign w12287 = ( w10801 & ~w12284 ) | ( w10801 & w12286 ) | ( ~w12284 & w12286 ) ;
  assign w12288 = \pi20 ^ w12287 ;
  assign w12289 = ( w12080 & w12280 ) | ( w12080 & w12288 ) | ( w12280 & w12288 ) ;
  assign w12290 = w5710 | w10887 ;
  assign w12291 = w5494 & ~w10885 ;
  assign w12292 = ( ~w10887 & w12290 ) | ( ~w10887 & w12291 ) | ( w12290 & w12291 ) ;
  assign w12293 = ~w5948 & w10883 ;
  assign w12294 = w10895 | w12292 ;
  assign w12295 = ( w5497 & w12292 ) | ( w5497 & w12294 ) | ( w12292 & w12294 ) ;
  assign w12296 = ( w10883 & ~w12293 ) | ( w10883 & w12295 ) | ( ~w12293 & w12295 ) ;
  assign w12297 = \pi17 ^ w12296 ;
  assign w12298 = ( w12078 & w12289 ) | ( w12078 & w12297 ) | ( w12289 & w12297 ) ;
  assign w12299 = ~w5710 & w10883 ;
  assign w12300 = w5494 & ~w10887 ;
  assign w12301 = ( w10883 & ~w12299 ) | ( w10883 & w12300 ) | ( ~w12299 & w12300 ) ;
  assign w12302 = w5948 | w11139 ;
  assign w12303 = w11256 | w12301 ;
  assign w12304 = ( w5497 & w12301 ) | ( w5497 & w12303 ) | ( w12301 & w12303 ) ;
  assign w12305 = ( ~w11139 & w12302 ) | ( ~w11139 & w12304 ) | ( w12302 & w12304 ) ;
  assign w12306 = \pi17 ^ w12305 ;
  assign w12307 = w11889 ^ w12064 ;
  assign w12308 = w11897 ^ w12307 ;
  assign w12309 = ( w12298 & w12306 ) | ( w12298 & ~w12308 ) | ( w12306 & ~w12308 ) ;
  assign w12310 = w12080 ^ w12280 ;
  assign w12311 = w12288 ^ w12310 ;
  assign w12312 = w12082 ^ w12279 ;
  assign w12313 = w12090 ^ w12312 ;
  assign w12314 = w5343 | w10805 ;
  assign w12315 = w4905 & w10784 ;
  assign w12316 = ( ~w10805 & w12314 ) | ( ~w10805 & w12315 ) | ( w12314 & w12315 ) ;
  assign w12317 = w5395 | w10807 ;
  assign w12318 = w11117 | w12316 ;
  assign w12319 = ( w4908 & w12316 ) | ( w4908 & w12318 ) | ( w12316 & w12318 ) ;
  assign w12320 = ( ~w10807 & w12317 ) | ( ~w10807 & w12319 ) | ( w12317 & w12319 ) ;
  assign w12321 = \pi20 ^ w12320 ;
  assign w12322 = w12092 ^ w12270 ;
  assign w12323 = w12278 ^ w12322 ;
  assign w12324 = w12259 ^ w12261 ;
  assign w12325 = w12269 ^ w12324 ;
  assign w12326 = w12094 ^ w12258 ;
  assign w12327 = w12102 ^ w12326 ;
  assign w12328 = ~w4143 & w9961 ;
  assign w12329 = w4052 & w9965 ;
  assign w12330 = ( w9961 & ~w12328 ) | ( w9961 & w12329 ) | ( ~w12328 & w12329 ) ;
  assign w12331 = w4147 | w11278 ;
  assign w12332 = w9963 & ~w12330 ;
  assign w12333 = ( w3964 & w12330 ) | ( w3964 & ~w12332 ) | ( w12330 & ~w12332 ) ;
  assign w12334 = ( ~w11278 & w12331 ) | ( ~w11278 & w12333 ) | ( w12331 & w12333 ) ;
  assign w12335 = \pi26 ^ w12334 ;
  assign w12336 = w12104 ^ w12257 ;
  assign w12337 = w12115 ^ w12336 ;
  assign w12338 = w3717 | w9973 ;
  assign w12339 = w3649 & w9975 ;
  assign w12340 = ( ~w9973 & w12338 ) | ( ~w9973 & w12339 ) | ( w12338 & w12339 ) ;
  assign w12341 = ~w3549 & w9971 ;
  assign w12342 = w11809 & ~w12340 ;
  assign w12343 = ( w3448 & w12340 ) | ( w3448 & ~w12342 ) | ( w12340 & ~w12342 ) ;
  assign w12344 = ( w9971 & ~w12341 ) | ( w9971 & w12343 ) | ( ~w12341 & w12343 ) ;
  assign w12345 = \pi29 ^ w12344 ;
  assign w12346 = ~w4143 & w9965 ;
  assign w12347 = w4052 & ~w9967 ;
  assign w12348 = ( w9965 & ~w12346 ) | ( w9965 & w12347 ) | ( ~w12346 & w12347 ) ;
  assign w12349 = ~w4147 & w11339 ;
  assign w12350 = w9961 | w12348 ;
  assign w12351 = ( w3964 & w12348 ) | ( w3964 & w12350 ) | ( w12348 & w12350 ) ;
  assign w12352 = ( w11339 & ~w12349 ) | ( w11339 & w12351 ) | ( ~w12349 & w12351 ) ;
  assign w12353 = \pi26 ^ w12352 ;
  assign w12354 = ( ~w12337 & w12345 ) | ( ~w12337 & w12353 ) | ( w12345 & w12353 ) ;
  assign w12355 = ( ~w12327 & w12335 ) | ( ~w12327 & w12354 ) | ( w12335 & w12354 ) ;
  assign w12356 = ~w4651 & w9842 ;
  assign w12357 = w4606 & ~w9955 ;
  assign w12358 = ( w9842 & ~w12356 ) | ( w9842 & w12357 ) | ( ~w12356 & w12357 ) ;
  assign w12359 = ~w4706 & w9953 ;
  assign w12360 = w10965 | w12358 ;
  assign w12361 = ( w4609 & w12358 ) | ( w4609 & w12360 ) | ( w12358 & w12360 ) ;
  assign w12362 = ( w9953 & ~w12359 ) | ( w9953 & w12361 ) | ( ~w12359 & w12361 ) ;
  assign w12363 = \pi23 ^ w12362 ;
  assign w12364 = ( ~w12325 & w12355 ) | ( ~w12325 & w12363 ) | ( w12355 & w12363 ) ;
  assign w12365 = ~w5343 & w10784 ;
  assign w12366 = w4905 & w10211 ;
  assign w12367 = ( w10784 & ~w12365 ) | ( w10784 & w12366 ) | ( ~w12365 & w12366 ) ;
  assign w12368 = w5395 | w10805 ;
  assign w12369 = w10855 & ~w12367 ;
  assign w12370 = ( w4908 & w12367 ) | ( w4908 & ~w12369 ) | ( w12367 & ~w12369 ) ;
  assign w12371 = ( ~w10805 & w12368 ) | ( ~w10805 & w12370 ) | ( w12368 & w12370 ) ;
  assign w12372 = \pi20 ^ w12371 ;
  assign w12373 = ( ~w12323 & w12364 ) | ( ~w12323 & w12372 ) | ( w12364 & w12372 ) ;
  assign w12374 = ( ~w12313 & w12321 ) | ( ~w12313 & w12373 ) | ( w12321 & w12373 ) ;
  assign w12375 = w5710 | w10885 ;
  assign w12376 = w5494 & ~w10866 ;
  assign w12377 = ( ~w10885 & w12375 ) | ( ~w10885 & w12376 ) | ( w12375 & w12376 ) ;
  assign w12378 = w5948 | w10887 ;
  assign w12379 = w11131 & ~w12377 ;
  assign w12380 = ( w5497 & w12377 ) | ( w5497 & ~w12379 ) | ( w12377 & ~w12379 ) ;
  assign w12381 = ( ~w10887 & w12378 ) | ( ~w10887 & w12380 ) | ( w12378 & w12380 ) ;
  assign w12382 = \pi17 ^ w12381 ;
  assign w12383 = ( w12311 & w12374 ) | ( w12311 & w12382 ) | ( w12374 & w12382 ) ;
  assign w12384 = ( w6048 & w6549 ) | ( w6048 & ~w11138 ) | ( w6549 & ~w11138 ) ;
  assign w12385 = w6549 & ~w12384 ;
  assign w12386 = ( w6637 & ~w12384 ) | ( w6637 & w12385 ) | ( ~w12384 & w12385 ) ;
  assign w12387 = ( ~w10738 & w12384 ) | ( ~w10738 & w12386 ) | ( w12384 & w12386 ) ;
  assign w12388 = w12078 ^ w12289 ;
  assign w12389 = w12297 ^ w12388 ;
  assign w12390 = w11146 & ~w12387 ;
  assign w12391 = ( w6045 & w12387 ) | ( w6045 & ~w12390 ) | ( w12387 & ~w12390 ) ;
  assign w12392 = \pi14 ^ w12391 ;
  assign w12393 = ( w12383 & w12389 ) | ( w12383 & w12392 ) | ( w12389 & w12392 ) ;
  assign w12394 = w12298 ^ w12308 ;
  assign w12395 = w12306 ^ w12394 ;
  assign w12396 = w6045 & w11146 ;
  assign w12397 = ( w6045 & w12387 ) | ( w6045 & ~w12396 ) | ( w12387 & ~w12396 ) ;
  assign w12398 = w12383 ^ w12397 ;
  assign w12399 = \pi14 ^ w12389 ;
  assign w12400 = w12398 ^ w12399 ;
  assign w12401 = w12311 ^ w12374 ;
  assign w12402 = w12382 ^ w12401 ;
  assign w12403 = w12313 ^ w12373 ;
  assign w12404 = w12321 ^ w12403 ;
  assign w12405 = w5710 | w10866 ;
  assign w12406 = w5494 & w10801 ;
  assign w12407 = ( ~w10866 & w12405 ) | ( ~w10866 & w12406 ) | ( w12405 & w12406 ) ;
  assign w12408 = w5948 | w10885 ;
  assign w12409 = w11160 & ~w12407 ;
  assign w12410 = ( w5497 & w12407 ) | ( w5497 & ~w12409 ) | ( w12407 & ~w12409 ) ;
  assign w12411 = ( ~w10885 & w12408 ) | ( ~w10885 & w12410 ) | ( w12408 & w12410 ) ;
  assign w12412 = \pi17 ^ w12411 ;
  assign w12413 = w12323 ^ w12364 ;
  assign w12414 = w12372 ^ w12413 ;
  assign w12415 = w12325 ^ w12355 ;
  assign w12416 = w12363 ^ w12415 ;
  assign w12417 = w12327 ^ w12354 ;
  assign w12418 = w12335 ^ w12417 ;
  assign w12419 = w4651 | w9955 ;
  assign w12420 = w4606 & w9957 ;
  assign w12421 = ( ~w9955 & w12419 ) | ( ~w9955 & w12420 ) | ( w12419 & w12420 ) ;
  assign w12422 = ~w4706 & w9842 ;
  assign w12423 = w10976 & ~w12421 ;
  assign w12424 = ( w4609 & w12421 ) | ( w4609 & ~w12423 ) | ( w12421 & ~w12423 ) ;
  assign w12425 = ( w9842 & ~w12422 ) | ( w9842 & w12424 ) | ( ~w12422 & w12424 ) ;
  assign w12426 = \pi23 ^ w12425 ;
  assign w12427 = w12337 ^ w12353 ;
  assign w12428 = w12345 ^ w12427 ;
  assign w12429 = w11949 ^ w12228 ;
  assign w12430 = w12135 ^ w12429 ;
  assign w12431 = ( w9985 & w9987 ) | ( w9985 & w10032 ) | ( w9987 & w10032 ) ;
  assign w12432 = w9985 ^ w12431 ;
  assign w12433 = w9983 ^ w12432 ;
  assign w12434 = ( \pi29 & \pi31 ) | ( \pi29 & w9985 ) | ( \pi31 & w9985 ) ;
  assign w12435 = ( \pi29 & ~\pi30 ) | ( \pi29 & w12434 ) | ( ~\pi30 & w12434 ) ;
  assign w12436 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w12434 ) | ( \pi30 & w12434 ) ;
  assign w12437 = ( ~\pi29 & w9987 ) | ( ~\pi29 & w12436 ) | ( w9987 & w12436 ) ;
  assign w12438 = ( w9983 & w12436 ) | ( w9983 & ~w12437 ) | ( w12436 & ~w12437 ) ;
  assign w12439 = ~\pi31 & w12438 ;
  assign w12440 = ( w12435 & w12437 ) | ( w12435 & w12439 ) | ( w12437 & w12439 ) ;
  assign w12441 = ( w37 & w12433 ) | ( w37 & w12440 ) | ( w12433 & w12440 ) ;
  assign w12442 = w12440 | w12441 ;
  assign w12443 = w11949 ^ w12227 ;
  assign w12444 = w12158 ^ w12443 ;
  assign w12445 = w9985 ^ w10032 ;
  assign w12446 = w9987 ^ w12445 ;
  assign w12447 = ( \pi29 & \pi31 ) | ( \pi29 & w9987 ) | ( \pi31 & w9987 ) ;
  assign w12448 = ( \pi29 & ~\pi30 ) | ( \pi29 & w12447 ) | ( ~\pi30 & w12447 ) ;
  assign w12449 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w12447 ) | ( \pi30 & w12447 ) ;
  assign w12450 = ( \pi29 & w9989 ) | ( \pi29 & ~w12449 ) | ( w9989 & ~w12449 ) ;
  assign w12451 = ( w9985 & w12449 ) | ( w9985 & w12450 ) | ( w12449 & w12450 ) ;
  assign w12452 = ~\pi31 & w12451 ;
  assign w12453 = ( w12448 & ~w12450 ) | ( w12448 & w12452 ) | ( ~w12450 & w12452 ) ;
  assign w12454 = ( w37 & w12446 ) | ( w37 & w12453 ) | ( w12446 & w12453 ) ;
  assign w12455 = w12453 | w12454 ;
  assign w12456 = w11949 ^ w12226 ;
  assign w12457 = w12214 ^ w12456 ;
  assign w12458 = ( w252 & w271 ) | ( w252 & ~w287 ) | ( w271 & ~w287 ) ;
  assign w12459 = w144 | w10174 ;
  assign w12460 = ( ~w144 & w287 ) | ( ~w144 & w385 ) | ( w287 & w385 ) ;
  assign w12461 = w12459 | w12460 ;
  assign w12462 = w12458 | w12461 ;
  assign w12463 = ( w223 & w491 ) | ( w223 & ~w722 ) | ( w491 & ~w722 ) ;
  assign w12464 = w410 | w759 ;
  assign w12465 = ( w722 & ~w759 ) | ( w722 & w1030 ) | ( ~w759 & w1030 ) ;
  assign w12466 = w12464 | w12465 ;
  assign w12467 = w12463 | w12466 ;
  assign w12468 = w2957 | w12467 ;
  assign w12469 = ( w2169 & w2354 ) | ( w2169 & ~w12467 ) | ( w2354 & ~w12467 ) ;
  assign w12470 = w12468 | w12469 ;
  assign w12471 = w11446 | w12462 ;
  assign w12472 = w696 | w12471 ;
  assign w12473 = ( ~w696 & w4814 ) | ( ~w696 & w12470 ) | ( w4814 & w12470 ) ;
  assign w12474 = w12472 | w12473 ;
  assign w12475 = w118 | w343 ;
  assign w12476 = w82 | w12475 ;
  assign w12477 = ( ~w82 & w270 ) | ( ~w82 & w12474 ) | ( w270 & w12474 ) ;
  assign w12478 = w12476 | w12477 ;
  assign w12479 = w215 | w386 ;
  assign w12480 = w63 | w12479 ;
  assign w12481 = ( ~w63 & w138 ) | ( ~w63 & w12478 ) | ( w138 & w12478 ) ;
  assign w12482 = w12480 | w12481 ;
  assign w12483 = w9989 ^ w10030 ;
  assign w12484 = w9991 ^ w12483 ;
  assign w12485 = w37 | w12484 ;
  assign w12486 = w3098 & ~w9993 ;
  assign w12487 = ( ~w12484 & w12485 ) | ( ~w12484 & w12486 ) | ( w12485 & w12486 ) ;
  assign w12488 = ( \pi29 & \pi30 ) | ( \pi29 & ~w9989 ) | ( \pi30 & ~w9989 ) ;
  assign w12489 = \pi31 | w12488 ;
  assign w12490 = ( \pi29 & ~\pi30 ) | ( \pi29 & w9991 ) | ( ~\pi30 & w9991 ) ;
  assign w12491 = ( \pi29 & \pi31 ) | ( \pi29 & ~w12490 ) | ( \pi31 & ~w12490 ) ;
  assign w12492 = ( w12487 & w12489 ) | ( w12487 & ~w12491 ) | ( w12489 & ~w12491 ) ;
  assign w12493 = ( ~w161 & w663 ) | ( ~w161 & w1095 ) | ( w663 & w1095 ) ;
  assign w12494 = w161 | w12493 ;
  assign w12495 = ( w169 & w605 ) | ( w169 & ~w889 ) | ( w605 & ~w889 ) ;
  assign w12496 = w2535 | w12494 ;
  assign w12497 = ( w889 & w901 ) | ( w889 & ~w2535 ) | ( w901 & ~w2535 ) ;
  assign w12498 = w12496 | w12497 ;
  assign w12499 = w12495 | w12498 ;
  assign w12500 = w5773 | w12499 ;
  assign w12501 = w1063 | w12500 ;
  assign w12502 = ( w559 & ~w1063 ) | ( w559 & w10576 ) | ( ~w1063 & w10576 ) ;
  assign w12503 = w12501 | w12502 ;
  assign w12504 = w206 | w283 ;
  assign w12505 = w450 | w12504 ;
  assign w12506 = ( w205 & ~w450 ) | ( w205 & w12503 ) | ( ~w450 & w12503 ) ;
  assign w12507 = w12505 | w12506 ;
  assign w12508 = ( w63 & w423 ) | ( w63 & ~w726 ) | ( w423 & ~w726 ) ;
  assign w12509 = w51 | w12507 ;
  assign w12510 = ( ~w51 & w726 ) | ( ~w51 & w1126 ) | ( w726 & w1126 ) ;
  assign w12511 = w12509 | w12510 ;
  assign w12512 = w12508 | w12511 ;
  assign w12513 = w9991 ^ w10029 ;
  assign w12514 = w9993 ^ w12513 ;
  assign w12515 = w37 | w12514 ;
  assign w12516 = w3098 & w9995 ;
  assign w12517 = ( ~w12514 & w12515 ) | ( ~w12514 & w12516 ) | ( w12515 & w12516 ) ;
  assign w12518 = ( \pi29 & \pi30 ) | ( \pi29 & w9991 ) | ( \pi30 & w9991 ) ;
  assign w12519 = \pi31 | w12518 ;
  assign w12520 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w9993 ) | ( \pi30 & w9993 ) ;
  assign w12521 = ( \pi29 & \pi31 ) | ( \pi29 & w12520 ) | ( \pi31 & w12520 ) ;
  assign w12522 = ( w12517 & w12519 ) | ( w12517 & ~w12521 ) | ( w12519 & ~w12521 ) ;
  assign w12523 = ( ~w141 & w524 ) | ( ~w141 & w4076 ) | ( w524 & w4076 ) ;
  assign w12524 = w2734 | w12523 ;
  assign w12525 = ( ~w608 & w2676 ) | ( ~w608 & w12524 ) | ( w2676 & w12524 ) ;
  assign w12526 = w1808 | w12187 ;
  assign w12527 = ( w608 & w1031 ) | ( w608 & ~w1808 ) | ( w1031 & ~w1808 ) ;
  assign w12528 = w12526 | w12527 ;
  assign w12529 = w12525 | w12528 ;
  assign w12530 = w1512 | w4381 ;
  assign w12531 = w888 | w12530 ;
  assign w12532 = ( ~w888 & w1064 ) | ( ~w888 & w12529 ) | ( w1064 & w12529 ) ;
  assign w12533 = w12531 | w12532 ;
  assign w12534 = ( w263 & w642 ) | ( w263 & ~w664 ) | ( w642 & ~w664 ) ;
  assign w12535 = w142 | w12533 ;
  assign w12536 = ( ~w142 & w664 ) | ( ~w142 & w783 ) | ( w664 & w783 ) ;
  assign w12537 = w12535 | w12536 ;
  assign w12538 = w12534 | w12537 ;
  assign w12539 = ( w9995 & w9997 ) | ( w9995 & w10027 ) | ( w9997 & w10027 ) ;
  assign w12540 = w9995 ^ w12539 ;
  assign w12541 = w9993 ^ w12540 ;
  assign w12542 = w37 | w12541 ;
  assign w12543 = w3098 & w9997 ;
  assign w12544 = ( ~w12541 & w12542 ) | ( ~w12541 & w12543 ) | ( w12542 & w12543 ) ;
  assign w12545 = ( \pi29 & \pi30 ) | ( \pi29 & ~w9993 ) | ( \pi30 & ~w9993 ) ;
  assign w12546 = \pi31 | w12545 ;
  assign w12547 = ( \pi29 & ~\pi30 ) | ( \pi29 & w9995 ) | ( ~\pi30 & w9995 ) ;
  assign w12548 = ( \pi29 & \pi31 ) | ( \pi29 & ~w12547 ) | ( \pi31 & ~w12547 ) ;
  assign w12549 = ( w12544 & w12546 ) | ( w12544 & ~w12548 ) | ( w12546 & ~w12548 ) ;
  assign w12550 = ( w202 & w324 ) | ( w202 & ~w351 ) | ( w324 & ~w351 ) ;
  assign w12551 = w177 | w890 ;
  assign w12552 = ( w351 & w492 ) | ( w351 & ~w890 ) | ( w492 & ~w890 ) ;
  assign w12553 = w12551 | w12552 ;
  assign w12554 = w12550 | w12553 ;
  assign w12555 = w3313 | w4476 ;
  assign w12556 = ( w1629 & ~w3313 ) | ( w1629 & w9902 ) | ( ~w3313 & w9902 ) ;
  assign w12557 = w12555 | w12556 ;
  assign w12558 = ( w1512 & ~w1978 ) | ( w1512 & w3501 ) | ( ~w1978 & w3501 ) ;
  assign w12559 = w6429 | w12557 ;
  assign w12560 = ( w1978 & w6353 ) | ( w1978 & ~w6429 ) | ( w6353 & ~w6429 ) ;
  assign w12561 = w12559 | w12560 ;
  assign w12562 = w12558 | w12561 ;
  assign w12563 = ( w339 & ~w458 ) | ( w339 & w1566 ) | ( ~w458 & w1566 ) ;
  assign w12564 = w12554 | w12562 ;
  assign w12565 = ( w458 & w509 ) | ( w458 & ~w12554 ) | ( w509 & ~w12554 ) ;
  assign w12566 = w12564 | w12565 ;
  assign w12567 = w12563 | w12566 ;
  assign w12568 = w63 | w697 ;
  assign w12569 = ( ~w63 & w259 ) | ( ~w63 & w12567 ) | ( w259 & w12567 ) ;
  assign w12570 = w12568 | w12569 ;
  assign w12571 = w9995 ^ w10027 ;
  assign w12572 = w9997 ^ w12571 ;
  assign w12573 = ~w37 & w12572 ;
  assign w12574 = w3098 & w9999 ;
  assign w12575 = ( w12572 & ~w12573 ) | ( w12572 & w12574 ) | ( ~w12573 & w12574 ) ;
  assign w12576 = ( \pi29 & \pi30 ) | ( \pi29 & w9995 ) | ( \pi30 & w9995 ) ;
  assign w12577 = \pi31 | w12576 ;
  assign w12578 = ( \pi29 & ~\pi30 ) | ( \pi29 & w9997 ) | ( ~\pi30 & w9997 ) ;
  assign w12579 = ( \pi29 & \pi31 ) | ( \pi29 & ~w12578 ) | ( \pi31 & ~w12578 ) ;
  assign w12580 = ( w12575 & w12577 ) | ( w12575 & ~w12579 ) | ( w12577 & ~w12579 ) ;
  assign w12581 = ( w505 & w516 ) | ( w505 & ~w626 ) | ( w516 & ~w626 ) ;
  assign w12582 = w361 | w1421 ;
  assign w12583 = ( ~w361 & w626 ) | ( ~w361 & w1229 ) | ( w626 & w1229 ) ;
  assign w12584 = w12582 | w12583 ;
  assign w12585 = w12581 | w12584 ;
  assign w12586 = w164 | w697 ;
  assign w12587 = w12585 | w12586 ;
  assign w12588 = ( w3250 & w4174 ) | ( w3250 & ~w12585 ) | ( w4174 & ~w12585 ) ;
  assign w12589 = w12587 | w12588 ;
  assign w12590 = ( w199 & w218 ) | ( w199 & ~w565 ) | ( w218 & ~w565 ) ;
  assign w12591 = w6238 | w12589 ;
  assign w12592 = ( w565 & w606 ) | ( w565 & ~w12589 ) | ( w606 & ~w12589 ) ;
  assign w12593 = w12591 | w12592 ;
  assign w12594 = w12590 | w12593 ;
  assign w12595 = ( w226 & w277 ) | ( w226 & ~w322 ) | ( w277 & ~w322 ) ;
  assign w12596 = w138 | w12594 ;
  assign w12597 = ( ~w138 & w322 ) | ( ~w138 & w725 ) | ( w322 & w725 ) ;
  assign w12598 = w12596 | w12597 ;
  assign w12599 = w12595 | w12598 ;
  assign w12600 = ( w84 & w136 ) | ( w84 & ~w724 ) | ( w136 & ~w724 ) ;
  assign w12601 = w450 | w4104 ;
  assign w12602 = ( w724 & w980 ) | ( w724 & ~w4104 ) | ( w980 & ~w4104 ) ;
  assign w12603 = w12601 | w12602 ;
  assign w12604 = w12600 | w12603 ;
  assign w12605 = w268 | w459 ;
  assign w12606 = w6353 | w12605 ;
  assign w12607 = ( w141 & ~w6353 ) | ( w141 & w12604 ) | ( ~w6353 & w12604 ) ;
  assign w12608 = w12606 | w12607 ;
  assign w12609 = w956 | w2695 ;
  assign w12610 = w4080 | w12609 ;
  assign w12611 = ( w168 & ~w4080 ) | ( w168 & w12608 ) | ( ~w4080 & w12608 ) ;
  assign w12612 = w12610 | w12611 ;
  assign w12613 = ( w95 & w345 ) | ( w95 & ~w515 ) | ( w345 & ~w515 ) ;
  assign w12614 = w572 | w12612 ;
  assign w12615 = ( w515 & ~w572 ) | ( w515 & w681 ) | ( ~w572 & w681 ) ;
  assign w12616 = w12614 | w12615 ;
  assign w12617 = w12613 | w12616 ;
  assign w12618 = w209 | w787 ;
  assign w12619 = ( w44 & ~w209 ) | ( w44 & w383 ) | ( ~w209 & w383 ) ;
  assign w12620 = w12618 | w12619 ;
  assign w12621 = w389 | w623 ;
  assign w12622 = w2876 | w12621 ;
  assign w12623 = ( w532 & ~w2876 ) | ( w532 & w12620 ) | ( ~w2876 & w12620 ) ;
  assign w12624 = w12622 | w12623 ;
  assign w12625 = ( w1977 & ~w6139 ) | ( w1977 & w12624 ) | ( ~w6139 & w12624 ) ;
  assign w12626 = w11318 | w12617 ;
  assign w12627 = ( w2836 & w6139 ) | ( w2836 & ~w11318 ) | ( w6139 & ~w11318 ) ;
  assign w12628 = w12626 | w12627 ;
  assign w12629 = w12625 | w12628 ;
  assign w12630 = ( w177 & w1155 ) | ( w177 & ~w2705 ) | ( w1155 & ~w2705 ) ;
  assign w12631 = w12599 | w12629 ;
  assign w12632 = ( w340 & w2705 ) | ( w340 & ~w12629 ) | ( w2705 & ~w12629 ) ;
  assign w12633 = w12631 | w12632 ;
  assign w12634 = w12630 | w12633 ;
  assign w12635 = ( w358 & w362 ) | ( w358 & ~w495 ) | ( w362 & ~w495 ) ;
  assign w12636 = w120 | w12634 ;
  assign w12637 = ( ~w120 & w495 ) | ( ~w120 & w1130 ) | ( w495 & w1130 ) ;
  assign w12638 = w12636 | w12637 ;
  assign w12639 = w12635 | w12638 ;
  assign w12640 = w9997 ^ w10026 ;
  assign w12641 = w9999 ^ w12640 ;
  assign w12642 = ~w37 & w12641 ;
  assign w12643 = w3098 & w10001 ;
  assign w12644 = ( w12641 & ~w12642 ) | ( w12641 & w12643 ) | ( ~w12642 & w12643 ) ;
  assign w12645 = ( \pi29 & \pi30 ) | ( \pi29 & w9997 ) | ( \pi30 & w9997 ) ;
  assign w12646 = \pi31 | w12645 ;
  assign w12647 = ( \pi29 & ~\pi30 ) | ( \pi29 & w9999 ) | ( ~\pi30 & w9999 ) ;
  assign w12648 = ( \pi29 & \pi31 ) | ( \pi29 & ~w12647 ) | ( \pi31 & ~w12647 ) ;
  assign w12649 = ( w12644 & w12646 ) | ( w12644 & ~w12648 ) | ( w12646 & ~w12648 ) ;
  assign w12650 = ( w393 & w506 ) | ( w393 & ~w605 ) | ( w506 & ~w605 ) ;
  assign w12651 = w95 | w115 ;
  assign w12652 = ( ~w115 & w605 ) | ( ~w115 & w723 ) | ( w605 & w723 ) ;
  assign w12653 = w12651 | w12652 ;
  assign w12654 = w12650 | w12653 ;
  assign w12655 = ( w147 & w223 ) | ( w147 & ~w224 ) | ( w223 & ~w224 ) ;
  assign w12656 = w11642 & ~w12654 ;
  assign w12657 = ( w224 & w524 ) | ( w224 & ~w12654 ) | ( w524 & ~w12654 ) ;
  assign w12658 = w12656 & ~w12657 ;
  assign w12659 = ~w12655 & w12658 ;
  assign w12660 = w1208 | w1835 ;
  assign w12661 = w1297 | w12660 ;
  assign w12662 = ( ~w1087 & w1297 ) | ( ~w1087 & w12659 ) | ( w1297 & w12659 ) ;
  assign w12663 = ~w12661 & w12662 ;
  assign w12664 = ( w286 & ~w445 ) | ( w286 & w12663 ) | ( ~w445 & w12663 ) ;
  assign w12665 = ~w286 & w12664 ;
  assign w12666 = ( w342 & w384 ) | ( w342 & ~w697 ) | ( w384 & ~w697 ) ;
  assign w12667 = ~w638 & w12665 ;
  assign w12668 = ( ~w638 & w697 ) | ( ~w638 & w802 ) | ( w697 & w802 ) ;
  assign w12669 = w12667 & ~w12668 ;
  assign w12670 = ~w12666 & w12669 ;
  assign w12671 = ( ~w283 & w1853 ) | ( ~w283 & w2092 ) | ( w1853 & w2092 ) ;
  assign w12672 = w10149 | w10380 ;
  assign w12673 = ( w283 & w722 ) | ( w283 & ~w10149 ) | ( w722 & ~w10149 ) ;
  assign w12674 = w12672 | w12673 ;
  assign w12675 = w12671 | w12674 ;
  assign w12676 = ( ~w214 & w742 ) | ( ~w214 & w998 ) | ( w742 & w998 ) ;
  assign w12677 = w12670 & ~w12675 ;
  assign w12678 = ( w214 & w1274 ) | ( w214 & ~w12675 ) | ( w1274 & ~w12675 ) ;
  assign w12679 = w12677 & ~w12678 ;
  assign w12680 = ~w12676 & w12679 ;
  assign w12681 = ( w167 & w390 ) | ( w167 & ~w534 ) | ( w390 & ~w534 ) ;
  assign w12682 = ~w142 & w12680 ;
  assign w12683 = ( ~w142 & w534 ) | ( ~w142 & w606 ) | ( w534 & w606 ) ;
  assign w12684 = w12682 & ~w12683 ;
  assign w12685 = ~w12681 & w12684 ;
  assign w12686 = ( w10006 & ~w10016 ) | ( w10006 & w10021 ) | ( ~w10016 & w10021 ) ;
  assign w12687 = w10006 | w12686 ;
  assign w12688 = ( ~w10001 & w10016 ) | ( ~w10001 & w12687 ) | ( w10016 & w12687 ) ;
  assign w12689 = ( w10006 & ~w10011 ) | ( w10006 & w12688 ) | ( ~w10011 & w12688 ) ;
  assign w12690 = w9999 ^ w12689 ;
  assign w12691 = w10001 ^ w12690 ;
  assign w12692 = w37 | w12691 ;
  assign w12693 = w3098 & ~w10006 ;
  assign w12694 = ( ~w12691 & w12692 ) | ( ~w12691 & w12693 ) | ( w12692 & w12693 ) ;
  assign w12695 = ( \pi29 & \pi30 ) | ( \pi29 & w9999 ) | ( \pi30 & w9999 ) ;
  assign w12696 = \pi31 | w12695 ;
  assign w12697 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10001 ) | ( ~\pi30 & w10001 ) ;
  assign w12698 = ( \pi29 & \pi31 ) | ( \pi29 & ~w12697 ) | ( \pi31 & ~w12697 ) ;
  assign w12699 = ( w12694 & w12696 ) | ( w12694 & ~w12698 ) | ( w12696 & ~w12698 ) ;
  assign w12700 = ( w359 & ~w421 ) | ( w359 & w817 ) | ( ~w421 & w817 ) ;
  assign w12701 = w309 | w316 ;
  assign w12702 = ( ~w316 & w817 ) | ( ~w316 & w1031 ) | ( w817 & w1031 ) ;
  assign w12703 = w12701 | w12702 ;
  assign w12704 = w12700 & ~w12703 ;
  assign w12705 = ( w139 & ~w491 ) | ( w139 & w12704 ) | ( ~w491 & w12704 ) ;
  assign w12706 = ~w139 & w12705 ;
  assign w12707 = w339 | w837 ;
  assign w12708 = w144 | w12707 ;
  assign w12709 = ( w88 & ~w144 ) | ( w88 & w314 ) | ( ~w144 & w314 ) ;
  assign w12710 = w12708 | w12709 ;
  assign w12711 = ( ~w119 & w468 ) | ( ~w119 & w12710 ) | ( w468 & w12710 ) ;
  assign w12712 = ~w11534 & w12706 ;
  assign w12713 = ( w119 & w229 ) | ( w119 & w12706 ) | ( w229 & w12706 ) ;
  assign w12714 = w12712 & ~w12713 ;
  assign w12715 = ~w12711 & w12714 ;
  assign w12716 = ( w124 & ~w640 ) | ( w124 & w2556 ) | ( ~w640 & w2556 ) ;
  assign w12717 = ~w838 & w12715 ;
  assign w12718 = ( w640 & w758 ) | ( w640 & ~w838 ) | ( w758 & ~w838 ) ;
  assign w12719 = w12717 & ~w12718 ;
  assign w12720 = ~w12716 & w12719 ;
  assign w12721 = ( w284 & w350 ) | ( w284 & ~w463 ) | ( w350 & ~w463 ) ;
  assign w12722 = ~w256 & w12720 ;
  assign w12723 = ( ~w256 & w463 ) | ( ~w256 & w628 ) | ( w463 & w628 ) ;
  assign w12724 = w12722 & ~w12723 ;
  assign w12725 = ~w12721 & w12724 ;
  assign w12726 = ( w281 & w315 ) | ( w281 & ~w951 ) | ( w315 & ~w951 ) ;
  assign w12727 = w104 | w113 ;
  assign w12728 = ( ~w113 & w951 ) | ( ~w113 & w1126 ) | ( w951 & w1126 ) ;
  assign w12729 = w12727 | w12728 ;
  assign w12730 = w12726 | w12729 ;
  assign w12731 = ( w455 & w1157 ) | ( w455 & ~w4818 ) | ( w1157 & ~w4818 ) ;
  assign w12732 = w1589 | w2469 ;
  assign w12733 = ( ~w2469 & w4818 ) | ( ~w2469 & w12730 ) | ( w4818 & w12730 ) ;
  assign w12734 = w12732 | w12733 ;
  assign w12735 = w12731 | w12734 ;
  assign w12736 = w103 | w642 ;
  assign w12737 = w12725 & ~w12736 ;
  assign w12738 = ( w1282 & w12725 ) | ( w1282 & w12735 ) | ( w12725 & w12735 ) ;
  assign w12739 = w12737 & ~w12738 ;
  assign w12740 = w409 | w724 ;
  assign w12741 = ( w409 & ~w496 ) | ( w409 & w12739 ) | ( ~w496 & w12739 ) ;
  assign w12742 = ~w12740 & w12741 ;
  assign w12743 = ( w10006 & ~w10011 ) | ( w10006 & w10016 ) | ( ~w10011 & w10016 ) ;
  assign w12744 = ~w10011 & w10021 ;
  assign w12745 = w12743 | w12744 ;
  assign w12746 = w10001 ^ w10006 ;
  assign w12747 = w12745 ^ w12746 ;
  assign w12748 = ~w37 & w12747 ;
  assign w12749 = w3098 & w10011 ;
  assign w12750 = ( w12747 & ~w12748 ) | ( w12747 & w12749 ) | ( ~w12748 & w12749 ) ;
  assign w12751 = ( \pi29 & \pi30 ) | ( \pi29 & w10001 ) | ( \pi30 & w10001 ) ;
  assign w12752 = \pi31 | w12751 ;
  assign w12753 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10006 ) | ( \pi30 & w10006 ) ;
  assign w12754 = ( \pi29 & \pi31 ) | ( \pi29 & w12753 ) | ( \pi31 & w12753 ) ;
  assign w12755 = ( w12750 & w12752 ) | ( w12750 & ~w12754 ) | ( w12752 & ~w12754 ) ;
  assign w12756 = ( w317 & w459 ) | ( w317 & ~w511 ) | ( w459 & ~w511 ) ;
  assign w12757 = ( ~w98 & w511 ) | ( ~w98 & w530 ) | ( w511 & w530 ) ;
  assign w12758 = w2752 | w12757 ;
  assign w12759 = w12756 | w12758 ;
  assign w12760 = ( ~w179 & w6194 ) | ( ~w179 & w12759 ) | ( w6194 & w12759 ) ;
  assign w12761 = w3299 | w5274 ;
  assign w12762 = ( w179 & w596 ) | ( w179 & ~w5274 ) | ( w596 & ~w5274 ) ;
  assign w12763 = w12761 | w12762 ;
  assign w12764 = w12760 | w12763 ;
  assign w12765 = w1978 | w3993 ;
  assign w12766 = w10563 | w12765 ;
  assign w12767 = ( w10486 & ~w10563 ) | ( w10486 & w12764 ) | ( ~w10563 & w12764 ) ;
  assign w12768 = w12766 | w12767 ;
  assign w12769 = ( w119 & w465 ) | ( w119 & ~w567 ) | ( w465 & ~w567 ) ;
  assign w12770 = w2147 | w12768 ;
  assign w12771 = ( w567 & w726 ) | ( w567 & ~w2147 ) | ( w726 & ~w2147 ) ;
  assign w12772 = w12770 | w12771 ;
  assign w12773 = w12769 | w12772 ;
  assign w12774 = w10006 ^ w10016 ;
  assign w12775 = ~w10011 & w10016 ;
  assign w12776 = ( w10011 & w10021 ) | ( w10011 & ~w12775 ) | ( w10021 & ~w12775 ) ;
  assign w12777 = w12774 ^ w12776 ;
  assign w12778 = ~w37 & w12777 ;
  assign w12779 = w3098 & ~w10016 ;
  assign w12780 = ( w12777 & ~w12778 ) | ( w12777 & w12779 ) | ( ~w12778 & w12779 ) ;
  assign w12781 = ( \pi29 & \pi30 ) | ( \pi29 & ~w10006 ) | ( \pi30 & ~w10006 ) ;
  assign w12782 = \pi31 | w12781 ;
  assign w12783 = ( \pi29 & ~\pi30 ) | ( \pi29 & w10011 ) | ( ~\pi30 & w10011 ) ;
  assign w12784 = ( \pi29 & \pi31 ) | ( \pi29 & ~w12783 ) | ( \pi31 & ~w12783 ) ;
  assign w12785 = ( w12780 & w12782 ) | ( w12780 & ~w12784 ) | ( w12782 & ~w12784 ) ;
  assign w12786 = ( w593 & w637 ) | ( w593 & ~w723 ) | ( w637 & ~w723 ) ;
  assign w12787 = w119 | w1129 ;
  assign w12788 = ( ~w119 & w723 ) | ( ~w119 & w980 ) | ( w723 & w980 ) ;
  assign w12789 = w12787 | w12788 ;
  assign w12790 = w12786 | w12789 ;
  assign w12791 = w890 | w1514 ;
  assign w12792 = w742 | w12791 ;
  assign w12793 = ( ~w742 & w820 ) | ( ~w742 & w12790 ) | ( w820 & w12790 ) ;
  assign w12794 = w12792 | w12793 ;
  assign w12795 = ( w275 & w311 ) | ( w275 & ~w423 ) | ( w311 & ~w423 ) ;
  assign w12796 = w76 | w12794 ;
  assign w12797 = ( ~w76 & w423 ) | ( ~w76 & w424 ) | ( w423 & w424 ) ;
  assign w12798 = w12796 | w12797 ;
  assign w12799 = w12795 | w12798 ;
  assign w12800 = ( w286 & w322 ) | ( w286 & ~w339 ) | ( w322 & ~w339 ) ;
  assign w12801 = w201 | w414 ;
  assign w12802 = ( ~w201 & w339 ) | ( ~w201 & w724 ) | ( w339 & w724 ) ;
  assign w12803 = w12801 | w12802 ;
  assign w12804 = w12800 | w12803 ;
  assign w12805 = w664 | w3494 ;
  assign w12806 = ( w447 & ~w3494 ) | ( w447 & w12804 ) | ( ~w3494 & w12804 ) ;
  assign w12807 = w12805 | w12806 ;
  assign w12808 = ( ~w1275 & w12196 ) | ( ~w1275 & w12807 ) | ( w12196 & w12807 ) ;
  assign w12809 = w11559 & ~w12799 ;
  assign w12810 = ( w1275 & w5039 ) | ( w1275 & ~w12799 ) | ( w5039 & ~w12799 ) ;
  assign w12811 = w12809 & ~w12810 ;
  assign w12812 = ~w12808 & w12811 ;
  assign w12813 = ( w116 & w274 ) | ( w116 & ~w312 ) | ( w274 & ~w312 ) ;
  assign w12814 = ~w410 & w12812 ;
  assign w12815 = ( w312 & ~w410 ) | ( w312 & w511 ) | ( ~w410 & w511 ) ;
  assign w12816 = w12814 & ~w12815 ;
  assign w12817 = ~w12813 & w12816 ;
  assign w12818 = ( w385 & w430 ) | ( w385 & ~w512 ) | ( w430 & ~w512 ) ;
  assign w12819 = ~w198 & w12817 ;
  assign w12820 = ( ~w198 & w512 ) | ( ~w198 & w726 ) | ( w512 & w726 ) ;
  assign w12821 = w12819 & ~w12820 ;
  assign w12822 = ~w12818 & w12821 ;
  assign w12823 = w286 | w764 ;
  assign w12824 = w63 | w12823 ;
  assign w12825 = ( ~w63 & w275 ) | ( ~w63 & w2274 ) | ( w275 & w2274 ) ;
  assign w12826 = w12824 | w12825 ;
  assign w12827 = w218 | w447 ;
  assign w12828 = w115 | w12827 ;
  assign w12829 = ( ~w115 & w131 ) | ( ~w115 & w12826 ) | ( w131 & w12826 ) ;
  assign w12830 = w12828 | w12829 ;
  assign w12831 = ( w491 & ~w534 ) | ( w491 & w3985 ) | ( ~w534 & w3985 ) ;
  assign w12832 = w624 | w10626 ;
  assign w12833 = ( w534 & ~w624 ) | ( w534 & w860 ) | ( ~w624 & w860 ) ;
  assign w12834 = w12832 | w12833 ;
  assign w12835 = w12831 | w12834 ;
  assign w12836 = w264 | w800 ;
  assign w12837 = w12835 | w12836 ;
  assign w12838 = ( w12554 & w12830 ) | ( w12554 & ~w12835 ) | ( w12830 & ~w12835 ) ;
  assign w12839 = w12837 | w12838 ;
  assign w12840 = ( w44 & w74 ) | ( w44 & ~w208 ) | ( w74 & ~w208 ) ;
  assign w12841 = w838 | w12839 ;
  assign w12842 = ( w208 & w310 ) | ( w208 & ~w838 ) | ( w310 & ~w838 ) ;
  assign w12843 = w12841 | w12842 ;
  assign w12844 = w12840 | w12843 ;
  assign w12845 = w787 | w980 ;
  assign w12846 = w205 | w12845 ;
  assign w12847 = ( w205 & ~w637 ) | ( w205 & w2554 ) | ( ~w637 & w2554 ) ;
  assign w12848 = ~w12846 & w12847 ;
  assign w12849 = ( w2255 & ~w3869 ) | ( w2255 & w12848 ) | ( ~w3869 & w12848 ) ;
  assign w12850 = ~w2255 & w12849 ;
  assign w12851 = ( w2146 & ~w2190 ) | ( w2146 & w6304 ) | ( ~w2190 & w6304 ) ;
  assign w12852 = ~w12844 & w12850 ;
  assign w12853 = ( w2190 & w2452 ) | ( w2190 & ~w12844 ) | ( w2452 & ~w12844 ) ;
  assign w12854 = w12852 & ~w12853 ;
  assign w12855 = ~w12851 & w12854 ;
  assign w12856 = ( w167 & w274 ) | ( w167 & ~w430 ) | ( w274 & ~w430 ) ;
  assign w12857 = ~w144 & w12855 ;
  assign w12858 = ( ~w144 & w430 ) | ( ~w144 & w758 ) | ( w430 & w758 ) ;
  assign w12859 = w12857 & ~w12858 ;
  assign w12860 = ~w12856 & w12859 ;
  assign w12861 = ( \pi29 & \pi30 ) | ( \pi29 & ~w10016 ) | ( \pi30 & ~w10016 ) ;
  assign w12862 = \pi31 ^ w10021 ;
  assign w12863 = ( \pi31 & w6862 ) | ( \pi31 & w12862 ) | ( w6862 & w12862 ) ;
  assign w12864 = w12861 ^ w12863 ;
  assign w12865 = ~w12860 & w12864 ;
  assign w12866 = ~w10016 & w10021 ;
  assign w12867 = w10011 ^ w12866 ;
  assign w12868 = \pi31 & ~w10021 ;
  assign w12869 = w10011 ^ w12868 ;
  assign w12870 = ( \pi29 & \pi30 ) | ( \pi29 & w12869 ) | ( \pi30 & w12869 ) ;
  assign w12871 = \pi31 ^ w12870 ;
  assign w12872 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10021 ) | ( \pi30 & w10021 ) ;
  assign w12873 = w6462 & ~w12872 ;
  assign w12874 = ( ~w10016 & w12871 ) | ( ~w10016 & w12873 ) | ( w12871 & w12873 ) ;
  assign w12875 = w36 & w10011 ;
  assign w12876 = ( w10016 & w12873 ) | ( w10016 & w12875 ) | ( w12873 & w12875 ) ;
  assign w12877 = w12874 | w12876 ;
  assign w12878 = ( ~w12822 & w12865 ) | ( ~w12822 & w12877 ) | ( w12865 & w12877 ) ;
  assign w12879 = ( w12773 & w12785 ) | ( w12773 & w12878 ) | ( w12785 & w12878 ) ;
  assign w12880 = ( ~w12742 & w12755 ) | ( ~w12742 & w12879 ) | ( w12755 & w12879 ) ;
  assign w12881 = ( ~w12685 & w12699 ) | ( ~w12685 & w12880 ) | ( w12699 & w12880 ) ;
  assign w12882 = ( w12639 & w12649 ) | ( w12639 & w12881 ) | ( w12649 & w12881 ) ;
  assign w12883 = ( w12570 & w12580 ) | ( w12570 & w12882 ) | ( w12580 & w12882 ) ;
  assign w12884 = ( w12538 & w12549 ) | ( w12538 & w12883 ) | ( w12549 & w12883 ) ;
  assign w12885 = ( w12512 & w12522 ) | ( w12512 & w12884 ) | ( w12522 & w12884 ) ;
  assign w12886 = ( w12482 & w12492 ) | ( w12482 & w12885 ) | ( w12492 & w12885 ) ;
  assign w12887 = w3549 & w9981 ;
  assign w12888 = ( w3717 & w9983 ) | ( w3717 & w12887 ) | ( w9983 & w12887 ) ;
  assign w12889 = w3649 | w12888 ;
  assign w12890 = ( w9985 & w12888 ) | ( w9985 & w12889 ) | ( w12888 & w12889 ) ;
  assign w12891 = w12887 | w12890 ;
  assign w12892 = ~w3448 & w12236 ;
  assign w12893 = ( w12236 & w12891 ) | ( w12236 & ~w12892 ) | ( w12891 & ~w12892 ) ;
  assign w12894 = \pi29 ^ w12893 ;
  assign w12895 = ( ~w12457 & w12886 ) | ( ~w12457 & w12894 ) | ( w12886 & w12894 ) ;
  assign w12896 = ( w12444 & w12455 ) | ( w12444 & w12895 ) | ( w12455 & w12895 ) ;
  assign w12897 = ( ~w12430 & w12442 ) | ( ~w12430 & w12896 ) | ( w12442 & w12896 ) ;
  assign w12898 = w12229 ^ w12234 ;
  assign w12899 = w12245 ^ w12898 ;
  assign w12900 = ~w3717 & w9977 ;
  assign w12901 = w3649 & w9979 ;
  assign w12902 = ( w9977 & ~w12900 ) | ( w9977 & w12901 ) | ( ~w12900 & w12901 ) ;
  assign w12903 = ~w3549 & w9975 ;
  assign w12904 = w11914 | w12902 ;
  assign w12905 = ( w3448 & w12902 ) | ( w3448 & w12904 ) | ( w12902 & w12904 ) ;
  assign w12906 = ( w9975 & ~w12903 ) | ( w9975 & w12905 ) | ( ~w12903 & w12905 ) ;
  assign w12907 = \pi29 ^ w12906 ;
  assign w12908 = ( w12897 & ~w12899 ) | ( w12897 & w12907 ) | ( ~w12899 & w12907 ) ;
  assign w12909 = w12246 ^ w12248 ;
  assign w12910 = w12256 ^ w12909 ;
  assign w12911 = w4143 | w9967 ;
  assign w12912 = w4052 & w9971 ;
  assign w12913 = ( ~w9967 & w12911 ) | ( ~w9967 & w12912 ) | ( w12911 & w12912 ) ;
  assign w12914 = w4147 | w11501 ;
  assign w12915 = w9965 | w12913 ;
  assign w12916 = ( w3964 & w12913 ) | ( w3964 & w12915 ) | ( w12913 & w12915 ) ;
  assign w12917 = ( ~w11501 & w12914 ) | ( ~w11501 & w12916 ) | ( w12914 & w12916 ) ;
  assign w12918 = \pi26 ^ w12917 ;
  assign w12919 = ( w12908 & w12910 ) | ( w12908 & w12918 ) | ( w12910 & w12918 ) ;
  assign w12920 = ~w4651 & w9957 ;
  assign w12921 = w4606 & ~w9963 ;
  assign w12922 = ( w9957 & ~w12920 ) | ( w9957 & w12921 ) | ( ~w12920 & w12921 ) ;
  assign w12923 = w4706 | w9955 ;
  assign w12924 = w11202 & ~w12922 ;
  assign w12925 = ( w4609 & w12922 ) | ( w4609 & ~w12924 ) | ( w12922 & ~w12924 ) ;
  assign w12926 = ( ~w9955 & w12923 ) | ( ~w9955 & w12925 ) | ( w12923 & w12925 ) ;
  assign w12927 = \pi23 ^ w12926 ;
  assign w12928 = ( ~w12428 & w12919 ) | ( ~w12428 & w12927 ) | ( w12919 & w12927 ) ;
  assign w12929 = ( ~w12418 & w12426 ) | ( ~w12418 & w12928 ) | ( w12426 & w12928 ) ;
  assign w12930 = ~w5343 & w10211 ;
  assign w12931 = w4905 & w10114 ;
  assign w12932 = ( w10211 & ~w12930 ) | ( w10211 & w12931 ) | ( ~w12930 & w12931 ) ;
  assign w12933 = ~w5395 & w10784 ;
  assign w12934 = w10789 | w12932 ;
  assign w12935 = ( w4908 & w12932 ) | ( w4908 & w12934 ) | ( w12932 & w12934 ) ;
  assign w12936 = ( w10784 & ~w12933 ) | ( w10784 & w12935 ) | ( ~w12933 & w12935 ) ;
  assign w12937 = \pi20 ^ w12936 ;
  assign w12938 = ( ~w12416 & w12929 ) | ( ~w12416 & w12937 ) | ( w12929 & w12937 ) ;
  assign w12939 = ~w5710 & w10801 ;
  assign w12940 = w5494 & ~w10807 ;
  assign w12941 = ( w10801 & ~w12939 ) | ( w10801 & w12940 ) | ( ~w12939 & w12940 ) ;
  assign w12942 = w5948 | w10866 ;
  assign w12943 = w10874 | w12941 ;
  assign w12944 = ( w5497 & w12941 ) | ( w5497 & w12943 ) | ( w12941 & w12943 ) ;
  assign w12945 = ( ~w10866 & w12942 ) | ( ~w10866 & w12944 ) | ( w12942 & w12944 ) ;
  assign w12946 = \pi17 ^ w12945 ;
  assign w12947 = ( ~w12414 & w12938 ) | ( ~w12414 & w12946 ) | ( w12938 & w12946 ) ;
  assign w12948 = ( ~w12404 & w12412 ) | ( ~w12404 & w12947 ) | ( w12412 & w12947 ) ;
  assign w12949 = w6549 | w11139 ;
  assign w12950 = w6048 & w10883 ;
  assign w12951 = ( ~w11139 & w12949 ) | ( ~w11139 & w12950 ) | ( w12949 & w12950 ) ;
  assign w12952 = w6637 | w10738 ;
  assign w12953 = w11145 & ~w12951 ;
  assign w12954 = ( w6045 & w12951 ) | ( w6045 & ~w12953 ) | ( w12951 & ~w12953 ) ;
  assign w12955 = ( ~w10738 & w12952 ) | ( ~w10738 & w12954 ) | ( w12952 & w12954 ) ;
  assign w12956 = \pi14 ^ w12955 ;
  assign w12957 = ( w12402 & w12948 ) | ( w12402 & w12956 ) | ( w12948 & w12956 ) ;
  assign w12958 = w12402 ^ w12948 ;
  assign w12959 = w12956 ^ w12958 ;
  assign w12960 = w12414 ^ w12938 ;
  assign w12961 = w12946 ^ w12960 ;
  assign w12962 = w12416 ^ w12929 ;
  assign w12963 = w12937 ^ w12962 ;
  assign w12964 = w12418 ^ w12928 ;
  assign w12965 = w12426 ^ w12964 ;
  assign w12966 = ~w5343 & w10114 ;
  assign w12967 = w4905 & w9953 ;
  assign w12968 = ( w10114 & ~w12966 ) | ( w10114 & w12967 ) | ( ~w12966 & w12967 ) ;
  assign w12969 = ~w5395 & w10211 ;
  assign w12970 = w10214 | w12968 ;
  assign w12971 = ( w4908 & w12968 ) | ( w4908 & w12970 ) | ( w12968 & w12970 ) ;
  assign w12972 = ( w10211 & ~w12969 ) | ( w10211 & w12971 ) | ( ~w12969 & w12971 ) ;
  assign w12973 = \pi20 ^ w12972 ;
  assign w12974 = w12428 ^ w12919 ;
  assign w12975 = w12927 ^ w12974 ;
  assign w12976 = w12908 ^ w12910 ;
  assign w12977 = w12918 ^ w12976 ;
  assign w12978 = w12897 ^ w12899 ;
  assign w12979 = w12907 ^ w12978 ;
  assign w12980 = ~w4143 & w9971 ;
  assign w12981 = w4052 & ~w9973 ;
  assign w12982 = ( w9971 & ~w12980 ) | ( w9971 & w12981 ) | ( ~w12980 & w12981 ) ;
  assign w12983 = w4147 | w11512 ;
  assign w12984 = w9967 & ~w12982 ;
  assign w12985 = ( w3964 & w12982 ) | ( w3964 & ~w12984 ) | ( w12982 & ~w12984 ) ;
  assign w12986 = ( ~w11512 & w12983 ) | ( ~w11512 & w12985 ) | ( w12983 & w12985 ) ;
  assign w12987 = \pi26 ^ w12986 ;
  assign w12988 = w12430 ^ w12896 ;
  assign w12989 = w12442 ^ w12988 ;
  assign w12990 = ~w3717 & w9979 ;
  assign w12991 = w3649 & w9981 ;
  assign w12992 = ( w9979 & ~w12990 ) | ( w9979 & w12991 ) | ( ~w12990 & w12991 ) ;
  assign w12993 = ~w3549 & w9977 ;
  assign w12994 = w12106 | w12992 ;
  assign w12995 = ( w3448 & w12992 ) | ( w3448 & w12994 ) | ( w12992 & w12994 ) ;
  assign w12996 = ( w9977 & ~w12993 ) | ( w9977 & w12995 ) | ( ~w12993 & w12995 ) ;
  assign w12997 = \pi29 ^ w12996 ;
  assign w12998 = ~w3964 & w9971 ;
  assign w12999 = w4143 & ~w9973 ;
  assign w13000 = ( w9971 & ~w12998 ) | ( w9971 & w12999 ) | ( ~w12998 & w12999 ) ;
  assign w13001 = w4147 | w11809 ;
  assign w13002 = w9975 | w13000 ;
  assign w13003 = ( w4052 & w13000 ) | ( w4052 & w13002 ) | ( w13000 & w13002 ) ;
  assign w13004 = ( ~w11809 & w13001 ) | ( ~w11809 & w13003 ) | ( w13001 & w13003 ) ;
  assign w13005 = \pi26 ^ w13004 ;
  assign w13006 = ( ~w12989 & w12997 ) | ( ~w12989 & w13005 ) | ( w12997 & w13005 ) ;
  assign w13007 = ( ~w12979 & w12987 ) | ( ~w12979 & w13006 ) | ( w12987 & w13006 ) ;
  assign w13008 = w4651 | w9963 ;
  assign w13009 = w4606 & w9961 ;
  assign w13010 = ( ~w9963 & w13008 ) | ( ~w9963 & w13009 ) | ( w13008 & w13009 ) ;
  assign w13011 = ~w4706 & w9957 ;
  assign w13012 = w11089 & ~w13010 ;
  assign w13013 = ( w4609 & w13010 ) | ( w4609 & ~w13012 ) | ( w13010 & ~w13012 ) ;
  assign w13014 = ( w9957 & ~w13011 ) | ( w9957 & w13013 ) | ( ~w13011 & w13013 ) ;
  assign w13015 = \pi23 ^ w13014 ;
  assign w13016 = ( w12977 & w13007 ) | ( w12977 & w13015 ) | ( w13007 & w13015 ) ;
  assign w13017 = ~w5343 & w9953 ;
  assign w13018 = w4905 & w9842 ;
  assign w13019 = ( w9953 & ~w13017 ) | ( w9953 & w13018 ) | ( ~w13017 & w13018 ) ;
  assign w13020 = ~w5395 & w10114 ;
  assign w13021 = w10334 | w13019 ;
  assign w13022 = ( w4908 & w13019 ) | ( w4908 & w13021 ) | ( w13019 & w13021 ) ;
  assign w13023 = ( w10114 & ~w13020 ) | ( w10114 & w13022 ) | ( ~w13020 & w13022 ) ;
  assign w13024 = \pi20 ^ w13023 ;
  assign w13025 = ( ~w12975 & w13016 ) | ( ~w12975 & w13024 ) | ( w13016 & w13024 ) ;
  assign w13026 = ( ~w12965 & w12973 ) | ( ~w12965 & w13025 ) | ( w12973 & w13025 ) ;
  assign w13027 = w5710 | w10807 ;
  assign w13028 = w5494 & ~w10805 ;
  assign w13029 = ( ~w10807 & w13027 ) | ( ~w10807 & w13028 ) | ( w13027 & w13028 ) ;
  assign w13030 = ~w5948 & w10801 ;
  assign w13031 = w10814 | w13029 ;
  assign w13032 = ( w5497 & w13029 ) | ( w5497 & w13031 ) | ( w13029 & w13031 ) ;
  assign w13033 = ( w10801 & ~w13030 ) | ( w10801 & w13032 ) | ( ~w13030 & w13032 ) ;
  assign w13034 = \pi17 ^ w13033 ;
  assign w13035 = ( ~w12963 & w13026 ) | ( ~w12963 & w13034 ) | ( w13026 & w13034 ) ;
  assign w13036 = w6549 | w10887 ;
  assign w13037 = w6048 & ~w10885 ;
  assign w13038 = ( ~w10887 & w13036 ) | ( ~w10887 & w13037 ) | ( w13036 & w13037 ) ;
  assign w13039 = ~w6637 & w10883 ;
  assign w13040 = w10895 | w13038 ;
  assign w13041 = ( w6045 & w13038 ) | ( w6045 & w13040 ) | ( w13038 & w13040 ) ;
  assign w13042 = ( w10883 & ~w13039 ) | ( w10883 & w13041 ) | ( ~w13039 & w13041 ) ;
  assign w13043 = \pi14 ^ w13042 ;
  assign w13044 = ( ~w12961 & w13035 ) | ( ~w12961 & w13043 ) | ( w13035 & w13043 ) ;
  assign w13045 = ~w6549 & w10883 ;
  assign w13046 = w6048 & ~w10887 ;
  assign w13047 = ( w10883 & ~w13045 ) | ( w10883 & w13046 ) | ( ~w13045 & w13046 ) ;
  assign w13048 = w6637 | w11139 ;
  assign w13049 = w11256 | w13047 ;
  assign w13050 = ( w6045 & w13047 ) | ( w6045 & w13049 ) | ( w13047 & w13049 ) ;
  assign w13051 = ( ~w11139 & w13048 ) | ( ~w11139 & w13050 ) | ( w13048 & w13050 ) ;
  assign w13052 = \pi14 ^ w13051 ;
  assign w13053 = w12404 ^ w12947 ;
  assign w13054 = w12412 ^ w13053 ;
  assign w13055 = ( w13044 & w13052 ) | ( w13044 & ~w13054 ) | ( w13052 & ~w13054 ) ;
  assign w13056 = w12963 ^ w13026 ;
  assign w13057 = w13034 ^ w13056 ;
  assign w13058 = w12965 ^ w13025 ;
  assign w13059 = w12973 ^ w13058 ;
  assign w13060 = w5710 | w10805 ;
  assign w13061 = w5494 & w10784 ;
  assign w13062 = ( ~w10805 & w13060 ) | ( ~w10805 & w13061 ) | ( w13060 & w13061 ) ;
  assign w13063 = w5948 | w10807 ;
  assign w13064 = w11117 | w13062 ;
  assign w13065 = ( w5497 & w13062 ) | ( w5497 & w13064 ) | ( w13062 & w13064 ) ;
  assign w13066 = ( ~w10807 & w13063 ) | ( ~w10807 & w13065 ) | ( w13063 & w13065 ) ;
  assign w13067 = \pi17 ^ w13066 ;
  assign w13068 = w12975 ^ w13016 ;
  assign w13069 = w13024 ^ w13068 ;
  assign w13070 = w12977 ^ w13007 ;
  assign w13071 = w13015 ^ w13070 ;
  assign w13072 = w12979 ^ w13006 ;
  assign w13073 = w12987 ^ w13072 ;
  assign w13074 = ~w4651 & w9961 ;
  assign w13075 = w4606 & w9965 ;
  assign w13076 = ( w9961 & ~w13074 ) | ( w9961 & w13075 ) | ( ~w13074 & w13075 ) ;
  assign w13077 = w4706 | w9963 ;
  assign w13078 = w11278 & ~w13076 ;
  assign w13079 = ( w4609 & w13076 ) | ( w4609 & ~w13078 ) | ( w13076 & ~w13078 ) ;
  assign w13080 = ( ~w9963 & w13077 ) | ( ~w9963 & w13079 ) | ( w13077 & w13079 ) ;
  assign w13081 = \pi23 ^ w13080 ;
  assign w13082 = w12989 ^ w13005 ;
  assign w13083 = w12997 ^ w13082 ;
  assign w13084 = w12444 ^ w12895 ;
  assign w13085 = w12455 ^ w13084 ;
  assign w13086 = ~w3717 & w9981 ;
  assign w13087 = w3649 & w9983 ;
  assign w13088 = ( w9981 & ~w13086 ) | ( w9981 & w13087 ) | ( ~w13086 & w13087 ) ;
  assign w13089 = ~w3549 & w9979 ;
  assign w13090 = w12010 | w13088 ;
  assign w13091 = ( w3448 & w13088 ) | ( w3448 & w13090 ) | ( w13088 & w13090 ) ;
  assign w13092 = ( w9979 & ~w13089 ) | ( w9979 & w13091 ) | ( ~w13089 & w13091 ) ;
  assign w13093 = \pi29 ^ w13092 ;
  assign w13094 = w3964 | w9973 ;
  assign w13095 = w4052 & w9977 ;
  assign w13096 = ( ~w9973 & w13094 ) | ( ~w9973 & w13095 ) | ( w13094 & w13095 ) ;
  assign w13097 = w4147 | w11671 ;
  assign w13098 = w9975 | w13096 ;
  assign w13099 = ( w4143 & w13096 ) | ( w4143 & w13098 ) | ( w13096 & w13098 ) ;
  assign w13100 = ( ~w11671 & w13097 ) | ( ~w11671 & w13099 ) | ( w13097 & w13099 ) ;
  assign w13101 = \pi26 ^ w13100 ;
  assign w13102 = ( w13085 & w13093 ) | ( w13085 & w13101 ) | ( w13093 & w13101 ) ;
  assign w13103 = ~w4651 & w9965 ;
  assign w13104 = w4606 & ~w9967 ;
  assign w13105 = ( w9965 & ~w13103 ) | ( w9965 & w13104 ) | ( ~w13103 & w13104 ) ;
  assign w13106 = ~w4706 & w9961 ;
  assign w13107 = w11339 | w13105 ;
  assign w13108 = ( w4609 & w13105 ) | ( w4609 & w13107 ) | ( w13105 & w13107 ) ;
  assign w13109 = ( w9961 & ~w13106 ) | ( w9961 & w13108 ) | ( ~w13106 & w13108 ) ;
  assign w13110 = \pi23 ^ w13109 ;
  assign w13111 = ( ~w13083 & w13102 ) | ( ~w13083 & w13110 ) | ( w13102 & w13110 ) ;
  assign w13112 = ( ~w13073 & w13081 ) | ( ~w13073 & w13111 ) | ( w13081 & w13111 ) ;
  assign w13113 = ~w5343 & w9842 ;
  assign w13114 = w4905 & ~w9955 ;
  assign w13115 = ( w9842 & ~w13113 ) | ( w9842 & w13114 ) | ( ~w13113 & w13114 ) ;
  assign w13116 = ~w5395 & w9953 ;
  assign w13117 = w10965 | w13115 ;
  assign w13118 = ( w4908 & w13115 ) | ( w4908 & w13117 ) | ( w13115 & w13117 ) ;
  assign w13119 = ( w9953 & ~w13116 ) | ( w9953 & w13118 ) | ( ~w13116 & w13118 ) ;
  assign w13120 = \pi20 ^ w13119 ;
  assign w13121 = ( w13071 & w13112 ) | ( w13071 & w13120 ) | ( w13112 & w13120 ) ;
  assign w13122 = ~w5710 & w10784 ;
  assign w13123 = w5494 & w10211 ;
  assign w13124 = ( w10784 & ~w13122 ) | ( w10784 & w13123 ) | ( ~w13122 & w13123 ) ;
  assign w13125 = w5948 | w10805 ;
  assign w13126 = w10855 & ~w13124 ;
  assign w13127 = ( w5497 & w13124 ) | ( w5497 & ~w13126 ) | ( w13124 & ~w13126 ) ;
  assign w13128 = ( ~w10805 & w13125 ) | ( ~w10805 & w13127 ) | ( w13125 & w13127 ) ;
  assign w13129 = \pi17 ^ w13128 ;
  assign w13130 = ( ~w13069 & w13121 ) | ( ~w13069 & w13129 ) | ( w13121 & w13129 ) ;
  assign w13131 = ( ~w13059 & w13067 ) | ( ~w13059 & w13130 ) | ( w13067 & w13130 ) ;
  assign w13132 = w6549 | w10885 ;
  assign w13133 = w6048 & ~w10866 ;
  assign w13134 = ( ~w10885 & w13132 ) | ( ~w10885 & w13133 ) | ( w13132 & w13133 ) ;
  assign w13135 = w6637 | w10887 ;
  assign w13136 = w11131 & ~w13134 ;
  assign w13137 = ( w6045 & w13134 ) | ( w6045 & ~w13136 ) | ( w13134 & ~w13136 ) ;
  assign w13138 = ( ~w10887 & w13135 ) | ( ~w10887 & w13137 ) | ( w13135 & w13137 ) ;
  assign w13139 = \pi14 ^ w13138 ;
  assign w13140 = ( ~w13057 & w13131 ) | ( ~w13057 & w13139 ) | ( w13131 & w13139 ) ;
  assign w13141 = ( w6748 & w6949 ) | ( w6748 & ~w11138 ) | ( w6949 & ~w11138 ) ;
  assign w13142 = w6949 & ~w13141 ;
  assign w13143 = ( w7154 & ~w13141 ) | ( w7154 & w13142 ) | ( ~w13141 & w13142 ) ;
  assign w13144 = ( ~w10738 & w13141 ) | ( ~w10738 & w13143 ) | ( w13141 & w13143 ) ;
  assign w13145 = w12961 ^ w13035 ;
  assign w13146 = w13043 ^ w13145 ;
  assign w13147 = w11146 & ~w13144 ;
  assign w13148 = ( w6751 & w13144 ) | ( w6751 & ~w13147 ) | ( w13144 & ~w13147 ) ;
  assign w13149 = \pi11 ^ w13148 ;
  assign w13150 = ( w13140 & ~w13146 ) | ( w13140 & w13149 ) | ( ~w13146 & w13149 ) ;
  assign w13151 = w13044 ^ w13054 ;
  assign w13152 = w13052 ^ w13151 ;
  assign w13153 = w6751 & w11146 ;
  assign w13154 = ( w6751 & w13144 ) | ( w6751 & ~w13153 ) | ( w13144 & ~w13153 ) ;
  assign w13155 = w13140 ^ w13154 ;
  assign w13156 = \pi11 ^ w13146 ;
  assign w13157 = w13155 ^ w13156 ;
  assign w13158 = w13057 ^ w13131 ;
  assign w13159 = w13139 ^ w13158 ;
  assign w13160 = w13059 ^ w13130 ;
  assign w13161 = w13067 ^ w13160 ;
  assign w13162 = w6549 | w10866 ;
  assign w13163 = w6048 & w10801 ;
  assign w13164 = ( ~w10866 & w13162 ) | ( ~w10866 & w13163 ) | ( w13162 & w13163 ) ;
  assign w13165 = w6637 | w10885 ;
  assign w13166 = w11160 & ~w13164 ;
  assign w13167 = ( w6045 & w13164 ) | ( w6045 & ~w13166 ) | ( w13164 & ~w13166 ) ;
  assign w13168 = ( ~w10885 & w13165 ) | ( ~w10885 & w13167 ) | ( w13165 & w13167 ) ;
  assign w13169 = \pi14 ^ w13168 ;
  assign w13170 = w13069 ^ w13121 ;
  assign w13171 = w13129 ^ w13170 ;
  assign w13172 = w13071 ^ w13112 ;
  assign w13173 = w13120 ^ w13172 ;
  assign w13174 = w13073 ^ w13111 ;
  assign w13175 = w13081 ^ w13174 ;
  assign w13176 = w5343 | w9955 ;
  assign w13177 = w4905 & w9957 ;
  assign w13178 = ( ~w9955 & w13176 ) | ( ~w9955 & w13177 ) | ( w13176 & w13177 ) ;
  assign w13179 = ~w5395 & w9842 ;
  assign w13180 = w10976 & ~w13178 ;
  assign w13181 = ( w4908 & w13178 ) | ( w4908 & ~w13180 ) | ( w13178 & ~w13180 ) ;
  assign w13182 = ( w9842 & ~w13179 ) | ( w9842 & w13181 ) | ( ~w13179 & w13181 ) ;
  assign w13183 = \pi20 ^ w13182 ;
  assign w13184 = w13083 ^ w13102 ;
  assign w13185 = w13110 ^ w13184 ;
  assign w13186 = w13085 ^ w13101 ;
  assign w13187 = w13093 ^ w13186 ;
  assign w13188 = w12492 ^ w12885 ;
  assign w13189 = w12482 ^ w13188 ;
  assign w13190 = w3549 & w9983 ;
  assign w13191 = ( w3717 & w9985 ) | ( w3717 & w13190 ) | ( w9985 & w13190 ) ;
  assign w13192 = w3649 | w13191 ;
  assign w13193 = ( w9987 & w13191 ) | ( w9987 & w13192 ) | ( w13191 & w13192 ) ;
  assign w13194 = w13190 | w13193 ;
  assign w13195 = ~w3448 & w12433 ;
  assign w13196 = ( w12433 & w13194 ) | ( w12433 & ~w13195 ) | ( w13194 & ~w13195 ) ;
  assign w13197 = \pi29 ^ w13196 ;
  assign w13198 = w12522 ^ w12884 ;
  assign w13199 = w12512 ^ w13198 ;
  assign w13200 = w3549 & w9985 ;
  assign w13201 = ( w3717 & w9987 ) | ( w3717 & w13200 ) | ( w9987 & w13200 ) ;
  assign w13202 = w3649 | w13201 ;
  assign w13203 = ( ~w9989 & w13201 ) | ( ~w9989 & w13202 ) | ( w13201 & w13202 ) ;
  assign w13204 = w13200 | w13203 ;
  assign w13205 = ~w3448 & w12446 ;
  assign w13206 = ( w12446 & w13204 ) | ( w12446 & ~w13205 ) | ( w13204 & ~w13205 ) ;
  assign w13207 = \pi29 ^ w13206 ;
  assign w13208 = w12549 ^ w12883 ;
  assign w13209 = w12538 ^ w13208 ;
  assign w13210 = w3549 & w9987 ;
  assign w13211 = ( w3717 & ~w9989 ) | ( w3717 & w13210 ) | ( ~w9989 & w13210 ) ;
  assign w13212 = w3649 | w13211 ;
  assign w13213 = ( w9991 & w13211 ) | ( w9991 & w13212 ) | ( w13211 & w13212 ) ;
  assign w13214 = w13210 | w13213 ;
  assign w13215 = w3448 | w12217 ;
  assign w13216 = ( ~w12217 & w13214 ) | ( ~w12217 & w13215 ) | ( w13214 & w13215 ) ;
  assign w13217 = \pi29 ^ w13216 ;
  assign w13218 = w12580 ^ w12882 ;
  assign w13219 = w12570 ^ w13218 ;
  assign w13220 = w3549 & ~w9989 ;
  assign w13221 = ( w3717 & w9991 ) | ( w3717 & w13220 ) | ( w9991 & w13220 ) ;
  assign w13222 = w3649 | w13221 ;
  assign w13223 = ( ~w9993 & w13221 ) | ( ~w9993 & w13222 ) | ( w13221 & w13222 ) ;
  assign w13224 = w13220 | w13223 ;
  assign w13225 = w3448 | w12484 ;
  assign w13226 = ( ~w12484 & w13224 ) | ( ~w12484 & w13225 ) | ( w13224 & w13225 ) ;
  assign w13227 = \pi29 ^ w13226 ;
  assign w13228 = w12649 ^ w12881 ;
  assign w13229 = w12639 ^ w13228 ;
  assign w13230 = w3549 & w9991 ;
  assign w13231 = ( w3717 & ~w9993 ) | ( w3717 & w13230 ) | ( ~w9993 & w13230 ) ;
  assign w13232 = w3649 | w13231 ;
  assign w13233 = ( w9995 & w13231 ) | ( w9995 & w13232 ) | ( w13231 & w13232 ) ;
  assign w13234 = w13230 | w13233 ;
  assign w13235 = w3448 | w12514 ;
  assign w13236 = ( ~w12514 & w13234 ) | ( ~w12514 & w13235 ) | ( w13234 & w13235 ) ;
  assign w13237 = \pi29 ^ w13236 ;
  assign w13238 = ~w3717 & w9995 ;
  assign w13239 = w3649 & w9997 ;
  assign w13240 = ( w9995 & ~w13238 ) | ( w9995 & w13239 ) | ( ~w13238 & w13239 ) ;
  assign w13241 = w3549 | w9993 ;
  assign w13242 = w12541 & ~w13240 ;
  assign w13243 = ( w3448 & w13240 ) | ( w3448 & ~w13242 ) | ( w13240 & ~w13242 ) ;
  assign w13244 = ( ~w9993 & w13241 ) | ( ~w9993 & w13243 ) | ( w13241 & w13243 ) ;
  assign w13245 = \pi29 ^ w13244 ;
  assign w13246 = w12699 ^ w12880 ;
  assign w13247 = w12685 ^ w13246 ;
  assign w13248 = ~w3717 & w9997 ;
  assign w13249 = w3649 & w9999 ;
  assign w13250 = ( w9997 & ~w13248 ) | ( w9997 & w13249 ) | ( ~w13248 & w13249 ) ;
  assign w13251 = ~w3549 & w9995 ;
  assign w13252 = w12572 | w13250 ;
  assign w13253 = ( w3448 & w13250 ) | ( w3448 & w13252 ) | ( w13250 & w13252 ) ;
  assign w13254 = ( w9995 & ~w13251 ) | ( w9995 & w13253 ) | ( ~w13251 & w13253 ) ;
  assign w13255 = \pi29 ^ w13254 ;
  assign w13256 = w12755 ^ w12879 ;
  assign w13257 = w12742 ^ w13256 ;
  assign w13258 = ~w3717 & w9999 ;
  assign w13259 = w3649 & w10001 ;
  assign w13260 = ( w9999 & ~w13258 ) | ( w9999 & w13259 ) | ( ~w13258 & w13259 ) ;
  assign w13261 = ~w3549 & w9997 ;
  assign w13262 = w12641 | w13260 ;
  assign w13263 = ( w3448 & w13260 ) | ( w3448 & w13262 ) | ( w13260 & w13262 ) ;
  assign w13264 = ( w9997 & ~w13261 ) | ( w9997 & w13263 ) | ( ~w13261 & w13263 ) ;
  assign w13265 = \pi29 ^ w13264 ;
  assign w13266 = w12785 ^ w12878 ;
  assign w13267 = w12773 ^ w13266 ;
  assign w13268 = ~w3717 & w10001 ;
  assign w13269 = w3649 & ~w10006 ;
  assign w13270 = ( w10001 & ~w13268 ) | ( w10001 & w13269 ) | ( ~w13268 & w13269 ) ;
  assign w13271 = ~w3549 & w9999 ;
  assign w13272 = w12691 & ~w13270 ;
  assign w13273 = ( w3448 & w13270 ) | ( w3448 & ~w13272 ) | ( w13270 & ~w13272 ) ;
  assign w13274 = ( w9999 & ~w13271 ) | ( w9999 & w13273 ) | ( ~w13271 & w13273 ) ;
  assign w13275 = \pi29 ^ w13274 ;
  assign w13276 = w12865 ^ w12877 ;
  assign w13277 = w12822 ^ w13276 ;
  assign w13278 = w3717 | w10006 ;
  assign w13279 = w3649 & w10011 ;
  assign w13280 = ( ~w10006 & w13278 ) | ( ~w10006 & w13279 ) | ( w13278 & w13279 ) ;
  assign w13281 = ~w3549 & w10001 ;
  assign w13282 = w12747 | w13280 ;
  assign w13283 = ( w3448 & w13280 ) | ( w3448 & w13282 ) | ( w13280 & w13282 ) ;
  assign w13284 = ( w10001 & ~w13281 ) | ( w10001 & w13283 ) | ( ~w13281 & w13283 ) ;
  assign w13285 = \pi29 ^ w13284 ;
  assign w13286 = w12860 ^ w12864 ;
  assign w13287 = \pi29 & w10021 ;
  assign w13288 = w10016 & w13287 ;
  assign w13289 = ( \pi26 & \pi27 ) | ( \pi26 & ~w13288 ) | ( \pi27 & ~w13288 ) ;
  assign w13290 = ( \pi28 & \pi29 ) | ( \pi28 & ~w13289 ) | ( \pi29 & ~w13289 ) ;
  assign w13291 = ( \pi28 & ~w13287 ) | ( \pi28 & w13289 ) | ( ~w13287 & w13289 ) ;
  assign w13292 = ( w6866 & w13290 ) | ( w6866 & ~w13291 ) | ( w13290 & ~w13291 ) ;
  assign w13293 = w3549 & w10011 ;
  assign w13294 = ( w3717 & ~w10016 ) | ( w3717 & w13293 ) | ( ~w10016 & w13293 ) ;
  assign w13295 = w3649 | w13294 ;
  assign w13296 = ( ~w10021 & w13294 ) | ( ~w10021 & w13295 ) | ( w13294 & w13295 ) ;
  assign w13297 = w13293 | w13296 ;
  assign w13298 = ~w3448 & w12867 ;
  assign w13299 = ( w12867 & w13297 ) | ( w12867 & ~w13298 ) | ( w13297 & ~w13298 ) ;
  assign w13300 = \pi29 ^ w13299 ;
  assign w13301 = w13292 & w13300 ;
  assign w13302 = ~w3717 & w10011 ;
  assign w13303 = w3649 & ~w10016 ;
  assign w13304 = ( w10011 & ~w13302 ) | ( w10011 & w13303 ) | ( ~w13302 & w13303 ) ;
  assign w13305 = w3549 | w10006 ;
  assign w13306 = w12777 | w13304 ;
  assign w13307 = ( w3448 & w13304 ) | ( w3448 & w13306 ) | ( w13304 & w13306 ) ;
  assign w13308 = ( ~w10006 & w13305 ) | ( ~w10006 & w13307 ) | ( w13305 & w13307 ) ;
  assign w13309 = \pi29 ^ w13308 ;
  assign w13310 = w36 & ~w10021 ;
  assign w13311 = ( w13301 & w13309 ) | ( w13301 & w13310 ) | ( w13309 & w13310 ) ;
  assign w13312 = ( w13285 & ~w13286 ) | ( w13285 & w13311 ) | ( ~w13286 & w13311 ) ;
  assign w13313 = ( w13275 & ~w13277 ) | ( w13275 & w13312 ) | ( ~w13277 & w13312 ) ;
  assign w13314 = ( w13265 & w13267 ) | ( w13265 & w13313 ) | ( w13267 & w13313 ) ;
  assign w13315 = ( w13255 & ~w13257 ) | ( w13255 & w13314 ) | ( ~w13257 & w13314 ) ;
  assign w13316 = ( w13245 & ~w13247 ) | ( w13245 & w13315 ) | ( ~w13247 & w13315 ) ;
  assign w13317 = ( w13229 & w13237 ) | ( w13229 & w13316 ) | ( w13237 & w13316 ) ;
  assign w13318 = ( w13219 & w13227 ) | ( w13219 & w13317 ) | ( w13227 & w13317 ) ;
  assign w13319 = ( w13209 & w13217 ) | ( w13209 & w13318 ) | ( w13217 & w13318 ) ;
  assign w13320 = ( w13199 & w13207 ) | ( w13199 & w13319 ) | ( w13207 & w13319 ) ;
  assign w13321 = ( w13189 & w13197 ) | ( w13189 & w13320 ) | ( w13197 & w13320 ) ;
  assign w13322 = w12457 ^ w12894 ;
  assign w13323 = w12886 ^ w13322 ;
  assign w13324 = ~w4143 & w9977 ;
  assign w13325 = w4052 & w9979 ;
  assign w13326 = ( w9977 & ~w13324 ) | ( w9977 & w13325 ) | ( ~w13324 & w13325 ) ;
  assign w13327 = ~w4147 & w11914 ;
  assign w13328 = w9975 | w13326 ;
  assign w13329 = ( w3964 & w13326 ) | ( w3964 & w13328 ) | ( w13326 & w13328 ) ;
  assign w13330 = ( w11914 & ~w13327 ) | ( w11914 & w13329 ) | ( ~w13327 & w13329 ) ;
  assign w13331 = \pi26 ^ w13330 ;
  assign w13332 = ( w13321 & ~w13323 ) | ( w13321 & w13331 ) | ( ~w13323 & w13331 ) ;
  assign w13333 = w4651 | w9967 ;
  assign w13334 = w4606 & w9971 ;
  assign w13335 = ( ~w9967 & w13333 ) | ( ~w9967 & w13334 ) | ( w13333 & w13334 ) ;
  assign w13336 = ~w4706 & w9965 ;
  assign w13337 = w11501 & ~w13335 ;
  assign w13338 = ( w4609 & w13335 ) | ( w4609 & ~w13337 ) | ( w13335 & ~w13337 ) ;
  assign w13339 = ( w9965 & ~w13336 ) | ( w9965 & w13338 ) | ( ~w13336 & w13338 ) ;
  assign w13340 = \pi23 ^ w13339 ;
  assign w13341 = ( w13187 & w13332 ) | ( w13187 & w13340 ) | ( w13332 & w13340 ) ;
  assign w13342 = ~w5343 & w9957 ;
  assign w13343 = w4905 & ~w9963 ;
  assign w13344 = ( w9957 & ~w13342 ) | ( w9957 & w13343 ) | ( ~w13342 & w13343 ) ;
  assign w13345 = w5395 | w9955 ;
  assign w13346 = w11202 & ~w13344 ;
  assign w13347 = ( w4908 & w13344 ) | ( w4908 & ~w13346 ) | ( w13344 & ~w13346 ) ;
  assign w13348 = ( ~w9955 & w13345 ) | ( ~w9955 & w13347 ) | ( w13345 & w13347 ) ;
  assign w13349 = \pi20 ^ w13348 ;
  assign w13350 = ( ~w13185 & w13341 ) | ( ~w13185 & w13349 ) | ( w13341 & w13349 ) ;
  assign w13351 = ( ~w13175 & w13183 ) | ( ~w13175 & w13350 ) | ( w13183 & w13350 ) ;
  assign w13352 = ~w5710 & w10211 ;
  assign w13353 = w5494 & w10114 ;
  assign w13354 = ( w10211 & ~w13352 ) | ( w10211 & w13353 ) | ( ~w13352 & w13353 ) ;
  assign w13355 = ~w5948 & w10784 ;
  assign w13356 = w10789 | w13354 ;
  assign w13357 = ( w5497 & w13354 ) | ( w5497 & w13356 ) | ( w13354 & w13356 ) ;
  assign w13358 = ( w10784 & ~w13355 ) | ( w10784 & w13357 ) | ( ~w13355 & w13357 ) ;
  assign w13359 = \pi17 ^ w13358 ;
  assign w13360 = ( w13173 & w13351 ) | ( w13173 & w13359 ) | ( w13351 & w13359 ) ;
  assign w13361 = ~w6549 & w10801 ;
  assign w13362 = w6048 & ~w10807 ;
  assign w13363 = ( w10801 & ~w13361 ) | ( w10801 & w13362 ) | ( ~w13361 & w13362 ) ;
  assign w13364 = w6637 | w10866 ;
  assign w13365 = w10874 | w13363 ;
  assign w13366 = ( w6045 & w13363 ) | ( w6045 & w13365 ) | ( w13363 & w13365 ) ;
  assign w13367 = ( ~w10866 & w13364 ) | ( ~w10866 & w13366 ) | ( w13364 & w13366 ) ;
  assign w13368 = \pi14 ^ w13367 ;
  assign w13369 = ( ~w13171 & w13360 ) | ( ~w13171 & w13368 ) | ( w13360 & w13368 ) ;
  assign w13370 = ( ~w13161 & w13169 ) | ( ~w13161 & w13369 ) | ( w13169 & w13369 ) ;
  assign w13371 = w6949 | w11139 ;
  assign w13372 = w6748 & w10883 ;
  assign w13373 = ( ~w11139 & w13371 ) | ( ~w11139 & w13372 ) | ( w13371 & w13372 ) ;
  assign w13374 = w7154 | w10738 ;
  assign w13375 = w11145 & ~w13373 ;
  assign w13376 = ( w6751 & w13373 ) | ( w6751 & ~w13375 ) | ( w13373 & ~w13375 ) ;
  assign w13377 = ( ~w10738 & w13374 ) | ( ~w10738 & w13376 ) | ( w13374 & w13376 ) ;
  assign w13378 = \pi11 ^ w13377 ;
  assign w13379 = ( ~w13159 & w13370 ) | ( ~w13159 & w13378 ) | ( w13370 & w13378 ) ;
  assign w13380 = w13159 ^ w13370 ;
  assign w13381 = w13378 ^ w13380 ;
  assign w13382 = w13171 ^ w13360 ;
  assign w13383 = w13368 ^ w13382 ;
  assign w13384 = w13173 ^ w13351 ;
  assign w13385 = w13359 ^ w13384 ;
  assign w13386 = w13175 ^ w13350 ;
  assign w13387 = w13183 ^ w13386 ;
  assign w13388 = ~w5710 & w10114 ;
  assign w13389 = w5494 & w9953 ;
  assign w13390 = ( w10114 & ~w13388 ) | ( w10114 & w13389 ) | ( ~w13388 & w13389 ) ;
  assign w13391 = ~w5948 & w10211 ;
  assign w13392 = w10214 | w13390 ;
  assign w13393 = ( w5497 & w13390 ) | ( w5497 & w13392 ) | ( w13390 & w13392 ) ;
  assign w13394 = ( w10211 & ~w13391 ) | ( w10211 & w13393 ) | ( ~w13391 & w13393 ) ;
  assign w13395 = \pi17 ^ w13394 ;
  assign w13396 = w13185 ^ w13341 ;
  assign w13397 = w13349 ^ w13396 ;
  assign w13398 = w13187 ^ w13332 ;
  assign w13399 = w13340 ^ w13398 ;
  assign w13400 = w13323 ^ w13331 ;
  assign w13401 = w13321 ^ w13400 ;
  assign w13402 = w13197 ^ w13320 ;
  assign w13403 = w13189 ^ w13402 ;
  assign w13404 = w3964 & w9977 ;
  assign w13405 = ( w4143 & w9979 ) | ( w4143 & w13404 ) | ( w9979 & w13404 ) ;
  assign w13406 = w4052 | w13405 ;
  assign w13407 = ( w9981 & w13405 ) | ( w9981 & w13406 ) | ( w13405 & w13406 ) ;
  assign w13408 = w13404 | w13407 ;
  assign w13409 = ~w4147 & w12106 ;
  assign w13410 = ( w12106 & w13408 ) | ( w12106 & ~w13409 ) | ( w13408 & ~w13409 ) ;
  assign w13411 = \pi26 ^ w13410 ;
  assign w13412 = w13207 ^ w13319 ;
  assign w13413 = w13199 ^ w13412 ;
  assign w13414 = w3964 & w9979 ;
  assign w13415 = ( w4143 & w9981 ) | ( w4143 & w13414 ) | ( w9981 & w13414 ) ;
  assign w13416 = w4052 | w13415 ;
  assign w13417 = ( w9983 & w13415 ) | ( w9983 & w13416 ) | ( w13415 & w13416 ) ;
  assign w13418 = w13414 | w13417 ;
  assign w13419 = ~w4147 & w12010 ;
  assign w13420 = ( w12010 & w13418 ) | ( w12010 & ~w13419 ) | ( w13418 & ~w13419 ) ;
  assign w13421 = \pi26 ^ w13420 ;
  assign w13422 = w13217 ^ w13318 ;
  assign w13423 = w13209 ^ w13422 ;
  assign w13424 = w3964 & w9981 ;
  assign w13425 = ( w4143 & w9983 ) | ( w4143 & w13424 ) | ( w9983 & w13424 ) ;
  assign w13426 = w4052 | w13425 ;
  assign w13427 = ( w9985 & w13425 ) | ( w9985 & w13426 ) | ( w13425 & w13426 ) ;
  assign w13428 = w13424 | w13427 ;
  assign w13429 = ~w4147 & w12236 ;
  assign w13430 = ( w12236 & w13428 ) | ( w12236 & ~w13429 ) | ( w13428 & ~w13429 ) ;
  assign w13431 = \pi26 ^ w13430 ;
  assign w13432 = w13227 ^ w13317 ;
  assign w13433 = w13219 ^ w13432 ;
  assign w13434 = w3964 & w9983 ;
  assign w13435 = ( w4143 & w9985 ) | ( w4143 & w13434 ) | ( w9985 & w13434 ) ;
  assign w13436 = w4052 | w13435 ;
  assign w13437 = ( w9987 & w13435 ) | ( w9987 & w13436 ) | ( w13435 & w13436 ) ;
  assign w13438 = w13434 | w13437 ;
  assign w13439 = ~w4147 & w12433 ;
  assign w13440 = ( w12433 & w13438 ) | ( w12433 & ~w13439 ) | ( w13438 & ~w13439 ) ;
  assign w13441 = \pi26 ^ w13440 ;
  assign w13442 = w13237 ^ w13316 ;
  assign w13443 = w13229 ^ w13442 ;
  assign w13444 = w3964 & w9985 ;
  assign w13445 = ( w4143 & w9987 ) | ( w4143 & w13444 ) | ( w9987 & w13444 ) ;
  assign w13446 = w4052 | w13445 ;
  assign w13447 = ( ~w9989 & w13445 ) | ( ~w9989 & w13446 ) | ( w13445 & w13446 ) ;
  assign w13448 = w13444 | w13447 ;
  assign w13449 = ~w4147 & w12446 ;
  assign w13450 = ( w12446 & w13448 ) | ( w12446 & ~w13449 ) | ( w13448 & ~w13449 ) ;
  assign w13451 = \pi26 ^ w13450 ;
  assign w13452 = w13245 ^ w13315 ;
  assign w13453 = w13247 ^ w13452 ;
  assign w13454 = w3964 & w9987 ;
  assign w13455 = ( w4143 & ~w9989 ) | ( w4143 & w13454 ) | ( ~w9989 & w13454 ) ;
  assign w13456 = w4052 | w13455 ;
  assign w13457 = ( w9991 & w13455 ) | ( w9991 & w13456 ) | ( w13455 & w13456 ) ;
  assign w13458 = w13454 | w13457 ;
  assign w13459 = w4147 | w12217 ;
  assign w13460 = ( ~w12217 & w13458 ) | ( ~w12217 & w13459 ) | ( w13458 & w13459 ) ;
  assign w13461 = \pi26 ^ w13460 ;
  assign w13462 = w13255 ^ w13314 ;
  assign w13463 = w13257 ^ w13462 ;
  assign w13464 = w3964 & ~w9989 ;
  assign w13465 = ( w4143 & w9991 ) | ( w4143 & w13464 ) | ( w9991 & w13464 ) ;
  assign w13466 = w4052 | w13465 ;
  assign w13467 = ( ~w9993 & w13465 ) | ( ~w9993 & w13466 ) | ( w13465 & w13466 ) ;
  assign w13468 = w13464 | w13467 ;
  assign w13469 = w4147 | w12484 ;
  assign w13470 = ( ~w12484 & w13468 ) | ( ~w12484 & w13469 ) | ( w13468 & w13469 ) ;
  assign w13471 = \pi26 ^ w13470 ;
  assign w13472 = w13265 ^ w13313 ;
  assign w13473 = w13267 ^ w13472 ;
  assign w13474 = w3964 & w9991 ;
  assign w13475 = ( w4143 & ~w9993 ) | ( w4143 & w13474 ) | ( ~w9993 & w13474 ) ;
  assign w13476 = w4052 | w13475 ;
  assign w13477 = ( w9995 & w13475 ) | ( w9995 & w13476 ) | ( w13475 & w13476 ) ;
  assign w13478 = w13474 | w13477 ;
  assign w13479 = w4147 | w12514 ;
  assign w13480 = ( ~w12514 & w13478 ) | ( ~w12514 & w13479 ) | ( w13478 & w13479 ) ;
  assign w13481 = \pi26 ^ w13480 ;
  assign w13482 = w13275 ^ w13312 ;
  assign w13483 = w13277 ^ w13482 ;
  assign w13484 = w3964 & ~w9993 ;
  assign w13485 = ( w4143 & w9995 ) | ( w4143 & w13484 ) | ( w9995 & w13484 ) ;
  assign w13486 = w4052 | w13485 ;
  assign w13487 = ( w9997 & w13485 ) | ( w9997 & w13486 ) | ( w13485 & w13486 ) ;
  assign w13488 = w13484 | w13487 ;
  assign w13489 = w4147 | w12541 ;
  assign w13490 = ( ~w12541 & w13488 ) | ( ~w12541 & w13489 ) | ( w13488 & w13489 ) ;
  assign w13491 = \pi26 ^ w13490 ;
  assign w13492 = w13285 ^ w13311 ;
  assign w13493 = w13286 ^ w13492 ;
  assign w13494 = w3964 & w9995 ;
  assign w13495 = ( w4143 & w9997 ) | ( w4143 & w13494 ) | ( w9997 & w13494 ) ;
  assign w13496 = w4052 | w13495 ;
  assign w13497 = ( w9999 & w13495 ) | ( w9999 & w13496 ) | ( w13495 & w13496 ) ;
  assign w13498 = w13494 | w13497 ;
  assign w13499 = ~w4147 & w12572 ;
  assign w13500 = ( w12572 & w13498 ) | ( w12572 & ~w13499 ) | ( w13498 & ~w13499 ) ;
  assign w13501 = \pi26 ^ w13500 ;
  assign w13502 = ~w3964 & w9997 ;
  assign w13503 = w4052 & w10001 ;
  assign w13504 = ( w9997 & ~w13502 ) | ( w9997 & w13503 ) | ( ~w13502 & w13503 ) ;
  assign w13505 = ~w4147 & w12641 ;
  assign w13506 = w9999 | w13504 ;
  assign w13507 = ( w4143 & w13504 ) | ( w4143 & w13506 ) | ( w13504 & w13506 ) ;
  assign w13508 = ( w12641 & ~w13505 ) | ( w12641 & w13507 ) | ( ~w13505 & w13507 ) ;
  assign w13509 = \pi26 ^ w13508 ;
  assign w13510 = w13301 ^ w13309 ;
  assign w13511 = w13310 ^ w13510 ;
  assign w13512 = ~w3964 & w9999 ;
  assign w13513 = w4143 & w10001 ;
  assign w13514 = ( w9999 & ~w13512 ) | ( w9999 & w13513 ) | ( ~w13512 & w13513 ) ;
  assign w13515 = w4147 | w12691 ;
  assign w13516 = w10006 & ~w13514 ;
  assign w13517 = ( w4052 & w13514 ) | ( w4052 & ~w13516 ) | ( w13514 & ~w13516 ) ;
  assign w13518 = ( ~w12691 & w13515 ) | ( ~w12691 & w13517 ) | ( w13515 & w13517 ) ;
  assign w13519 = \pi26 ^ w13518 ;
  assign w13520 = w13292 ^ w13300 ;
  assign w13521 = ( \pi26 & \pi27 ) | ( \pi26 & ~w10016 ) | ( \pi27 & ~w10016 ) ;
  assign w13522 = ( \pi26 & \pi27 ) | ( \pi26 & ~w10021 ) | ( \pi27 & ~w10021 ) ;
  assign w13523 = \pi28 ^ w10021 ;
  assign w13524 = ( \pi28 & w13522 ) | ( \pi28 & w13523 ) | ( w13522 & w13523 ) ;
  assign w13525 = w13521 ^ w13524 ;
  assign w13526 = w3964 & w10001 ;
  assign w13527 = ( w4143 & ~w10006 ) | ( w4143 & w13526 ) | ( ~w10006 & w13526 ) ;
  assign w13528 = w4052 | w13527 ;
  assign w13529 = ( w10011 & w13527 ) | ( w10011 & w13528 ) | ( w13527 & w13528 ) ;
  assign w13530 = w13526 | w13529 ;
  assign w13531 = ~w4147 & w12747 ;
  assign w13532 = ( w12747 & w13530 ) | ( w12747 & ~w13531 ) | ( w13530 & ~w13531 ) ;
  assign w13533 = \pi26 ^ w13532 ;
  assign w13534 = \pi26 & w10021 ;
  assign w13535 = w10016 & w13534 ;
  assign w13536 = ( \pi23 & \pi24 ) | ( \pi23 & ~w13535 ) | ( \pi24 & ~w13535 ) ;
  assign w13537 = ( \pi25 & \pi26 ) | ( \pi25 & ~w13536 ) | ( \pi26 & ~w13536 ) ;
  assign w13538 = ( \pi25 & ~w13534 ) | ( \pi25 & w13536 ) | ( ~w13534 & w13536 ) ;
  assign w13539 = ( w7079 & w13537 ) | ( w7079 & ~w13538 ) | ( w13537 & ~w13538 ) ;
  assign w13540 = w3964 & w10011 ;
  assign w13541 = ( w4143 & ~w10016 ) | ( w4143 & w13540 ) | ( ~w10016 & w13540 ) ;
  assign w13542 = w4052 | w13541 ;
  assign w13543 = ( ~w10021 & w13541 ) | ( ~w10021 & w13542 ) | ( w13541 & w13542 ) ;
  assign w13544 = w13540 | w13543 ;
  assign w13545 = ~w4147 & w12867 ;
  assign w13546 = ( w12867 & w13544 ) | ( w12867 & ~w13545 ) | ( w13544 & ~w13545 ) ;
  assign w13547 = \pi26 ^ w13546 ;
  assign w13548 = w13539 & w13547 ;
  assign w13549 = w3964 | w10006 ;
  assign w13550 = w4143 & w10011 ;
  assign w13551 = ( ~w10006 & w13549 ) | ( ~w10006 & w13550 ) | ( w13549 & w13550 ) ;
  assign w13552 = ~w4147 & w12777 ;
  assign w13553 = w10016 & ~w13551 ;
  assign w13554 = ( w4052 & w13551 ) | ( w4052 & ~w13553 ) | ( w13551 & ~w13553 ) ;
  assign w13555 = ( w12777 & ~w13552 ) | ( w12777 & w13554 ) | ( ~w13552 & w13554 ) ;
  assign w13556 = \pi26 ^ w13555 ;
  assign w13557 = w3447 & ~w10021 ;
  assign w13558 = ( w13548 & w13556 ) | ( w13548 & w13557 ) | ( w13556 & w13557 ) ;
  assign w13559 = ( w13525 & w13533 ) | ( w13525 & w13558 ) | ( w13533 & w13558 ) ;
  assign w13560 = ( w13519 & w13520 ) | ( w13519 & w13559 ) | ( w13520 & w13559 ) ;
  assign w13561 = ( w13509 & w13511 ) | ( w13509 & w13560 ) | ( w13511 & w13560 ) ;
  assign w13562 = ( ~w13493 & w13501 ) | ( ~w13493 & w13561 ) | ( w13501 & w13561 ) ;
  assign w13563 = ( ~w13483 & w13491 ) | ( ~w13483 & w13562 ) | ( w13491 & w13562 ) ;
  assign w13564 = ( w13473 & w13481 ) | ( w13473 & w13563 ) | ( w13481 & w13563 ) ;
  assign w13565 = ( ~w13463 & w13471 ) | ( ~w13463 & w13564 ) | ( w13471 & w13564 ) ;
  assign w13566 = ( ~w13453 & w13461 ) | ( ~w13453 & w13565 ) | ( w13461 & w13565 ) ;
  assign w13567 = ( w13443 & w13451 ) | ( w13443 & w13566 ) | ( w13451 & w13566 ) ;
  assign w13568 = ( w13433 & w13441 ) | ( w13433 & w13567 ) | ( w13441 & w13567 ) ;
  assign w13569 = ( w13423 & w13431 ) | ( w13423 & w13568 ) | ( w13431 & w13568 ) ;
  assign w13570 = ( w13413 & w13421 ) | ( w13413 & w13569 ) | ( w13421 & w13569 ) ;
  assign w13571 = ( w13403 & w13411 ) | ( w13403 & w13570 ) | ( w13411 & w13570 ) ;
  assign w13572 = ~w4651 & w9971 ;
  assign w13573 = w4606 & ~w9973 ;
  assign w13574 = ( w9971 & ~w13572 ) | ( w9971 & w13573 ) | ( ~w13572 & w13573 ) ;
  assign w13575 = w4706 | w9967 ;
  assign w13576 = w11512 & ~w13574 ;
  assign w13577 = ( w4609 & w13574 ) | ( w4609 & ~w13576 ) | ( w13574 & ~w13576 ) ;
  assign w13578 = ( ~w9967 & w13575 ) | ( ~w9967 & w13577 ) | ( w13575 & w13577 ) ;
  assign w13579 = \pi23 ^ w13578 ;
  assign w13580 = ( ~w13401 & w13571 ) | ( ~w13401 & w13579 ) | ( w13571 & w13579 ) ;
  assign w13581 = w5343 | w9963 ;
  assign w13582 = w4905 & w9961 ;
  assign w13583 = ( ~w9963 & w13581 ) | ( ~w9963 & w13582 ) | ( w13581 & w13582 ) ;
  assign w13584 = ~w5395 & w9957 ;
  assign w13585 = w11089 & ~w13583 ;
  assign w13586 = ( w4908 & w13583 ) | ( w4908 & ~w13585 ) | ( w13583 & ~w13585 ) ;
  assign w13587 = ( w9957 & ~w13584 ) | ( w9957 & w13586 ) | ( ~w13584 & w13586 ) ;
  assign w13588 = \pi20 ^ w13587 ;
  assign w13589 = ( w13399 & w13580 ) | ( w13399 & w13588 ) | ( w13580 & w13588 ) ;
  assign w13590 = ~w5710 & w9953 ;
  assign w13591 = w5494 & w9842 ;
  assign w13592 = ( w9953 & ~w13590 ) | ( w9953 & w13591 ) | ( ~w13590 & w13591 ) ;
  assign w13593 = ~w5948 & w10114 ;
  assign w13594 = w10334 | w13592 ;
  assign w13595 = ( w5497 & w13592 ) | ( w5497 & w13594 ) | ( w13592 & w13594 ) ;
  assign w13596 = ( w10114 & ~w13593 ) | ( w10114 & w13595 ) | ( ~w13593 & w13595 ) ;
  assign w13597 = \pi17 ^ w13596 ;
  assign w13598 = ( ~w13397 & w13589 ) | ( ~w13397 & w13597 ) | ( w13589 & w13597 ) ;
  assign w13599 = ( ~w13387 & w13395 ) | ( ~w13387 & w13598 ) | ( w13395 & w13598 ) ;
  assign w13600 = w6549 | w10807 ;
  assign w13601 = w6048 & ~w10805 ;
  assign w13602 = ( ~w10807 & w13600 ) | ( ~w10807 & w13601 ) | ( w13600 & w13601 ) ;
  assign w13603 = ~w6637 & w10801 ;
  assign w13604 = w10814 | w13602 ;
  assign w13605 = ( w6045 & w13602 ) | ( w6045 & w13604 ) | ( w13602 & w13604 ) ;
  assign w13606 = ( w10801 & ~w13603 ) | ( w10801 & w13605 ) | ( ~w13603 & w13605 ) ;
  assign w13607 = \pi14 ^ w13606 ;
  assign w13608 = ( w13385 & w13599 ) | ( w13385 & w13607 ) | ( w13599 & w13607 ) ;
  assign w13609 = w6949 | w10887 ;
  assign w13610 = w6748 & ~w10885 ;
  assign w13611 = ( ~w10887 & w13609 ) | ( ~w10887 & w13610 ) | ( w13609 & w13610 ) ;
  assign w13612 = ~w7154 & w10883 ;
  assign w13613 = w10895 | w13611 ;
  assign w13614 = ( w6751 & w13611 ) | ( w6751 & w13613 ) | ( w13611 & w13613 ) ;
  assign w13615 = ( w10883 & ~w13612 ) | ( w10883 & w13614 ) | ( ~w13612 & w13614 ) ;
  assign w13616 = \pi11 ^ w13615 ;
  assign w13617 = ( ~w13383 & w13608 ) | ( ~w13383 & w13616 ) | ( w13608 & w13616 ) ;
  assign w13618 = ~w6949 & w10883 ;
  assign w13619 = w6748 & ~w10887 ;
  assign w13620 = ( w10883 & ~w13618 ) | ( w10883 & w13619 ) | ( ~w13618 & w13619 ) ;
  assign w13621 = w7154 | w11139 ;
  assign w13622 = w11256 | w13620 ;
  assign w13623 = ( w6751 & w13620 ) | ( w6751 & w13622 ) | ( w13620 & w13622 ) ;
  assign w13624 = ( ~w11139 & w13621 ) | ( ~w11139 & w13623 ) | ( w13621 & w13623 ) ;
  assign w13625 = \pi11 ^ w13624 ;
  assign w13626 = w13161 ^ w13369 ;
  assign w13627 = w13169 ^ w13626 ;
  assign w13628 = ( w13617 & w13625 ) | ( w13617 & ~w13627 ) | ( w13625 & ~w13627 ) ;
  assign w13629 = w13385 ^ w13599 ;
  assign w13630 = w13607 ^ w13629 ;
  assign w13631 = w13387 ^ w13598 ;
  assign w13632 = w13395 ^ w13631 ;
  assign w13633 = w6549 | w10805 ;
  assign w13634 = w6048 & w10784 ;
  assign w13635 = ( ~w10805 & w13633 ) | ( ~w10805 & w13634 ) | ( w13633 & w13634 ) ;
  assign w13636 = w6637 | w10807 ;
  assign w13637 = w11117 | w13635 ;
  assign w13638 = ( w6045 & w13635 ) | ( w6045 & w13637 ) | ( w13635 & w13637 ) ;
  assign w13639 = ( ~w10807 & w13636 ) | ( ~w10807 & w13638 ) | ( w13636 & w13638 ) ;
  assign w13640 = \pi14 ^ w13639 ;
  assign w13641 = w13397 ^ w13589 ;
  assign w13642 = w13597 ^ w13641 ;
  assign w13643 = w13399 ^ w13580 ;
  assign w13644 = w13588 ^ w13643 ;
  assign w13645 = w13401 ^ w13579 ;
  assign w13646 = w13571 ^ w13645 ;
  assign w13647 = w4651 | w9973 ;
  assign w13648 = w4606 & w9975 ;
  assign w13649 = ( ~w9973 & w13647 ) | ( ~w9973 & w13648 ) | ( w13647 & w13648 ) ;
  assign w13650 = ~w4706 & w9971 ;
  assign w13651 = w11809 & ~w13649 ;
  assign w13652 = ( w4609 & w13649 ) | ( w4609 & ~w13651 ) | ( w13649 & ~w13651 ) ;
  assign w13653 = ( w9971 & ~w13650 ) | ( w9971 & w13652 ) | ( ~w13650 & w13652 ) ;
  assign w13654 = \pi23 ^ w13653 ;
  assign w13655 = w13411 ^ w13570 ;
  assign w13656 = w13403 ^ w13655 ;
  assign w13657 = ~w4651 & w9975 ;
  assign w13658 = w4606 & w9977 ;
  assign w13659 = ( w9975 & ~w13657 ) | ( w9975 & w13658 ) | ( ~w13657 & w13658 ) ;
  assign w13660 = w4706 | w9973 ;
  assign w13661 = w11671 & ~w13659 ;
  assign w13662 = ( w4609 & w13659 ) | ( w4609 & ~w13661 ) | ( w13659 & ~w13661 ) ;
  assign w13663 = ( ~w9973 & w13660 ) | ( ~w9973 & w13662 ) | ( w13660 & w13662 ) ;
  assign w13664 = \pi23 ^ w13663 ;
  assign w13665 = w13421 ^ w13569 ;
  assign w13666 = w13413 ^ w13665 ;
  assign w13667 = ~w4651 & w9977 ;
  assign w13668 = w4606 & w9979 ;
  assign w13669 = ( w9977 & ~w13667 ) | ( w9977 & w13668 ) | ( ~w13667 & w13668 ) ;
  assign w13670 = ~w4706 & w9975 ;
  assign w13671 = w11914 | w13669 ;
  assign w13672 = ( w4609 & w13669 ) | ( w4609 & w13671 ) | ( w13669 & w13671 ) ;
  assign w13673 = ( w9975 & ~w13670 ) | ( w9975 & w13672 ) | ( ~w13670 & w13672 ) ;
  assign w13674 = \pi23 ^ w13673 ;
  assign w13675 = w13431 ^ w13568 ;
  assign w13676 = w13423 ^ w13675 ;
  assign w13677 = ~w4651 & w9979 ;
  assign w13678 = w4606 & w9981 ;
  assign w13679 = ( w9979 & ~w13677 ) | ( w9979 & w13678 ) | ( ~w13677 & w13678 ) ;
  assign w13680 = ~w4706 & w9977 ;
  assign w13681 = w12106 | w13679 ;
  assign w13682 = ( w4609 & w13679 ) | ( w4609 & w13681 ) | ( w13679 & w13681 ) ;
  assign w13683 = ( w9977 & ~w13680 ) | ( w9977 & w13682 ) | ( ~w13680 & w13682 ) ;
  assign w13684 = \pi23 ^ w13683 ;
  assign w13685 = w13441 ^ w13567 ;
  assign w13686 = w13433 ^ w13685 ;
  assign w13687 = ~w4651 & w9981 ;
  assign w13688 = w4606 & w9983 ;
  assign w13689 = ( w9981 & ~w13687 ) | ( w9981 & w13688 ) | ( ~w13687 & w13688 ) ;
  assign w13690 = ~w4706 & w9979 ;
  assign w13691 = w12010 | w13689 ;
  assign w13692 = ( w4609 & w13689 ) | ( w4609 & w13691 ) | ( w13689 & w13691 ) ;
  assign w13693 = ( w9979 & ~w13690 ) | ( w9979 & w13692 ) | ( ~w13690 & w13692 ) ;
  assign w13694 = \pi23 ^ w13693 ;
  assign w13695 = w13451 ^ w13566 ;
  assign w13696 = w13443 ^ w13695 ;
  assign w13697 = ~w4651 & w9983 ;
  assign w13698 = w4606 & w9985 ;
  assign w13699 = ( w9983 & ~w13697 ) | ( w9983 & w13698 ) | ( ~w13697 & w13698 ) ;
  assign w13700 = ~w4706 & w9981 ;
  assign w13701 = w12236 | w13699 ;
  assign w13702 = ( w4609 & w13699 ) | ( w4609 & w13701 ) | ( w13699 & w13701 ) ;
  assign w13703 = ( w9981 & ~w13700 ) | ( w9981 & w13702 ) | ( ~w13700 & w13702 ) ;
  assign w13704 = \pi23 ^ w13703 ;
  assign w13705 = w13461 ^ w13565 ;
  assign w13706 = w13453 ^ w13705 ;
  assign w13707 = ~w4651 & w9985 ;
  assign w13708 = w4606 & w9987 ;
  assign w13709 = ( w9985 & ~w13707 ) | ( w9985 & w13708 ) | ( ~w13707 & w13708 ) ;
  assign w13710 = ~w4706 & w9983 ;
  assign w13711 = w12433 | w13709 ;
  assign w13712 = ( w4609 & w13709 ) | ( w4609 & w13711 ) | ( w13709 & w13711 ) ;
  assign w13713 = ( w9983 & ~w13710 ) | ( w9983 & w13712 ) | ( ~w13710 & w13712 ) ;
  assign w13714 = \pi23 ^ w13713 ;
  assign w13715 = w13471 ^ w13564 ;
  assign w13716 = w13463 ^ w13715 ;
  assign w13717 = ~w4651 & w9987 ;
  assign w13718 = w4606 & ~w9989 ;
  assign w13719 = ( w9987 & ~w13717 ) | ( w9987 & w13718 ) | ( ~w13717 & w13718 ) ;
  assign w13720 = ~w4706 & w9985 ;
  assign w13721 = w12446 | w13719 ;
  assign w13722 = ( w4609 & w13719 ) | ( w4609 & w13721 ) | ( w13719 & w13721 ) ;
  assign w13723 = ( w9985 & ~w13720 ) | ( w9985 & w13722 ) | ( ~w13720 & w13722 ) ;
  assign w13724 = \pi23 ^ w13723 ;
  assign w13725 = w13481 ^ w13563 ;
  assign w13726 = w13473 ^ w13725 ;
  assign w13727 = w4651 | w9989 ;
  assign w13728 = w4606 & w9991 ;
  assign w13729 = ( ~w9989 & w13727 ) | ( ~w9989 & w13728 ) | ( w13727 & w13728 ) ;
  assign w13730 = ~w4706 & w9987 ;
  assign w13731 = w12217 & ~w13729 ;
  assign w13732 = ( w4609 & w13729 ) | ( w4609 & ~w13731 ) | ( w13729 & ~w13731 ) ;
  assign w13733 = ( w9987 & ~w13730 ) | ( w9987 & w13732 ) | ( ~w13730 & w13732 ) ;
  assign w13734 = \pi23 ^ w13733 ;
  assign w13735 = w13491 ^ w13562 ;
  assign w13736 = w13483 ^ w13735 ;
  assign w13737 = ~w4651 & w9991 ;
  assign w13738 = w4606 & ~w9993 ;
  assign w13739 = ( w9991 & ~w13737 ) | ( w9991 & w13738 ) | ( ~w13737 & w13738 ) ;
  assign w13740 = w4706 | w9989 ;
  assign w13741 = w12484 & ~w13739 ;
  assign w13742 = ( w4609 & w13739 ) | ( w4609 & ~w13741 ) | ( w13739 & ~w13741 ) ;
  assign w13743 = ( ~w9989 & w13740 ) | ( ~w9989 & w13742 ) | ( w13740 & w13742 ) ;
  assign w13744 = \pi23 ^ w13743 ;
  assign w13745 = w13501 ^ w13561 ;
  assign w13746 = w13493 ^ w13745 ;
  assign w13747 = w13509 ^ w13560 ;
  assign w13748 = w13511 ^ w13747 ;
  assign w13749 = w4606 & w9995 ;
  assign w13750 = ( w4706 & w9991 ) | ( w4706 & w13749 ) | ( w9991 & w13749 ) ;
  assign w13751 = w4651 | w13750 ;
  assign w13752 = ( ~w9993 & w13750 ) | ( ~w9993 & w13751 ) | ( w13750 & w13751 ) ;
  assign w13753 = w13749 | w13752 ;
  assign w13754 = w4609 | w12514 ;
  assign w13755 = ( ~w12514 & w13753 ) | ( ~w12514 & w13754 ) | ( w13753 & w13754 ) ;
  assign w13756 = \pi23 ^ w13755 ;
  assign w13757 = w13519 ^ w13559 ;
  assign w13758 = w13520 ^ w13757 ;
  assign w13759 = w4606 & w9997 ;
  assign w13760 = ( w4706 & ~w9993 ) | ( w4706 & w13759 ) | ( ~w9993 & w13759 ) ;
  assign w13761 = w4651 | w13760 ;
  assign w13762 = ( w9995 & w13760 ) | ( w9995 & w13761 ) | ( w13760 & w13761 ) ;
  assign w13763 = w13759 | w13762 ;
  assign w13764 = w4609 | w12541 ;
  assign w13765 = ( ~w12541 & w13763 ) | ( ~w12541 & w13764 ) | ( w13763 & w13764 ) ;
  assign w13766 = \pi23 ^ w13765 ;
  assign w13767 = ~w4651 & w9997 ;
  assign w13768 = w4606 & w9999 ;
  assign w13769 = ( w9997 & ~w13767 ) | ( w9997 & w13768 ) | ( ~w13767 & w13768 ) ;
  assign w13770 = ~w4706 & w9995 ;
  assign w13771 = w12572 | w13769 ;
  assign w13772 = ( w4609 & w13769 ) | ( w4609 & w13771 ) | ( w13769 & w13771 ) ;
  assign w13773 = ( w9995 & ~w13770 ) | ( w9995 & w13772 ) | ( ~w13770 & w13772 ) ;
  assign w13774 = \pi23 ^ w13773 ;
  assign w13775 = w13533 ^ w13558 ;
  assign w13776 = w13525 ^ w13775 ;
  assign w13777 = w13548 ^ w13556 ;
  assign w13778 = w13557 ^ w13777 ;
  assign w13779 = w4606 & w10001 ;
  assign w13780 = ( w4706 & w9997 ) | ( w4706 & w13779 ) | ( w9997 & w13779 ) ;
  assign w13781 = w4651 | w13780 ;
  assign w13782 = ( w9999 & w13780 ) | ( w9999 & w13781 ) | ( w13780 & w13781 ) ;
  assign w13783 = w13779 | w13782 ;
  assign w13784 = ~w4609 & w12641 ;
  assign w13785 = ( w12641 & w13783 ) | ( w12641 & ~w13784 ) | ( w13783 & ~w13784 ) ;
  assign w13786 = \pi23 ^ w13785 ;
  assign w13787 = ~w4651 & w10001 ;
  assign w13788 = w4606 & ~w10006 ;
  assign w13789 = ( w10001 & ~w13787 ) | ( w10001 & w13788 ) | ( ~w13787 & w13788 ) ;
  assign w13790 = ~w4706 & w9999 ;
  assign w13791 = w12691 & ~w13789 ;
  assign w13792 = ( w4609 & w13789 ) | ( w4609 & ~w13791 ) | ( w13789 & ~w13791 ) ;
  assign w13793 = ( w9999 & ~w13790 ) | ( w9999 & w13792 ) | ( ~w13790 & w13792 ) ;
  assign w13794 = \pi23 ^ w13793 ;
  assign w13795 = w13539 ^ w13547 ;
  assign w13796 = ( \pi23 & \pi24 ) | ( \pi23 & ~w10016 ) | ( \pi24 & ~w10016 ) ;
  assign w13797 = ( \pi23 & \pi24 ) | ( \pi23 & ~w10021 ) | ( \pi24 & ~w10021 ) ;
  assign w13798 = \pi25 ^ w10021 ;
  assign w13799 = ( \pi25 & w13797 ) | ( \pi25 & w13798 ) | ( w13797 & w13798 ) ;
  assign w13800 = w13796 ^ w13799 ;
  assign w13801 = w4606 & w10011 ;
  assign w13802 = ( w4706 & w10001 ) | ( w4706 & w13801 ) | ( w10001 & w13801 ) ;
  assign w13803 = w4651 | w13802 ;
  assign w13804 = ( ~w10006 & w13802 ) | ( ~w10006 & w13803 ) | ( w13802 & w13803 ) ;
  assign w13805 = w13801 | w13804 ;
  assign w13806 = ~w4609 & w12747 ;
  assign w13807 = ( w12747 & w13805 ) | ( w12747 & ~w13806 ) | ( w13805 & ~w13806 ) ;
  assign w13808 = \pi23 ^ w13807 ;
  assign w13809 = \pi23 & w10021 ;
  assign w13810 = w10016 & w13809 ;
  assign w13811 = ( \pi20 & \pi21 ) | ( \pi20 & ~w13810 ) | ( \pi21 & ~w13810 ) ;
  assign w13812 = ( \pi22 & \pi23 ) | ( \pi22 & ~w13811 ) | ( \pi23 & ~w13811 ) ;
  assign w13813 = ( \pi22 & ~w13809 ) | ( \pi22 & w13811 ) | ( ~w13809 & w13811 ) ;
  assign w13814 = ( w7331 & w13812 ) | ( w7331 & ~w13813 ) | ( w13812 & ~w13813 ) ;
  assign w13815 = w4606 & ~w10021 ;
  assign w13816 = ( w4706 & w10011 ) | ( w4706 & w13815 ) | ( w10011 & w13815 ) ;
  assign w13817 = w4651 | w13816 ;
  assign w13818 = ( ~w10016 & w13816 ) | ( ~w10016 & w13817 ) | ( w13816 & w13817 ) ;
  assign w13819 = w13815 | w13818 ;
  assign w13820 = ~w4609 & w12867 ;
  assign w13821 = ( w12867 & w13819 ) | ( w12867 & ~w13820 ) | ( w13819 & ~w13820 ) ;
  assign w13822 = \pi23 ^ w13821 ;
  assign w13823 = w13814 & w13822 ;
  assign w13824 = ~w4651 & w10011 ;
  assign w13825 = w4606 & ~w10016 ;
  assign w13826 = ( w10011 & ~w13824 ) | ( w10011 & w13825 ) | ( ~w13824 & w13825 ) ;
  assign w13827 = w4706 | w10006 ;
  assign w13828 = w12777 | w13826 ;
  assign w13829 = ( w4609 & w13826 ) | ( w4609 & w13828 ) | ( w13826 & w13828 ) ;
  assign w13830 = ( ~w10006 & w13827 ) | ( ~w10006 & w13829 ) | ( w13827 & w13829 ) ;
  assign w13831 = \pi23 ^ w13830 ;
  assign w13832 = w2832 & ~w10021 ;
  assign w13833 = ( w13823 & w13831 ) | ( w13823 & w13832 ) | ( w13831 & w13832 ) ;
  assign w13834 = ( w13800 & w13808 ) | ( w13800 & w13833 ) | ( w13808 & w13833 ) ;
  assign w13835 = ( w13794 & w13795 ) | ( w13794 & w13834 ) | ( w13795 & w13834 ) ;
  assign w13836 = ( w13778 & w13786 ) | ( w13778 & w13835 ) | ( w13786 & w13835 ) ;
  assign w13837 = ( w13774 & w13776 ) | ( w13774 & w13836 ) | ( w13776 & w13836 ) ;
  assign w13838 = ( w13758 & w13766 ) | ( w13758 & w13837 ) | ( w13766 & w13837 ) ;
  assign w13839 = ( w13748 & w13756 ) | ( w13748 & w13838 ) | ( w13756 & w13838 ) ;
  assign w13840 = ( w13744 & ~w13746 ) | ( w13744 & w13839 ) | ( ~w13746 & w13839 ) ;
  assign w13841 = ( w13734 & ~w13736 ) | ( w13734 & w13840 ) | ( ~w13736 & w13840 ) ;
  assign w13842 = ( w13724 & w13726 ) | ( w13724 & w13841 ) | ( w13726 & w13841 ) ;
  assign w13843 = ( w13714 & ~w13716 ) | ( w13714 & w13842 ) | ( ~w13716 & w13842 ) ;
  assign w13844 = ( w13704 & ~w13706 ) | ( w13704 & w13843 ) | ( ~w13706 & w13843 ) ;
  assign w13845 = ( w13694 & w13696 ) | ( w13694 & w13844 ) | ( w13696 & w13844 ) ;
  assign w13846 = ( w13684 & w13686 ) | ( w13684 & w13845 ) | ( w13686 & w13845 ) ;
  assign w13847 = ( w13674 & w13676 ) | ( w13674 & w13846 ) | ( w13676 & w13846 ) ;
  assign w13848 = ( w13664 & w13666 ) | ( w13664 & w13847 ) | ( w13666 & w13847 ) ;
  assign w13849 = ( w13654 & w13656 ) | ( w13654 & w13848 ) | ( w13656 & w13848 ) ;
  assign w13850 = ~w5343 & w9961 ;
  assign w13851 = w4905 & w9965 ;
  assign w13852 = ( w9961 & ~w13850 ) | ( w9961 & w13851 ) | ( ~w13850 & w13851 ) ;
  assign w13853 = w5395 | w9963 ;
  assign w13854 = w11278 & ~w13852 ;
  assign w13855 = ( w4908 & w13852 ) | ( w4908 & ~w13854 ) | ( w13852 & ~w13854 ) ;
  assign w13856 = ( ~w9963 & w13853 ) | ( ~w9963 & w13855 ) | ( w13853 & w13855 ) ;
  assign w13857 = \pi20 ^ w13856 ;
  assign w13858 = ( ~w13646 & w13849 ) | ( ~w13646 & w13857 ) | ( w13849 & w13857 ) ;
  assign w13859 = ~w5710 & w9842 ;
  assign w13860 = w5494 & ~w9955 ;
  assign w13861 = ( w9842 & ~w13859 ) | ( w9842 & w13860 ) | ( ~w13859 & w13860 ) ;
  assign w13862 = ~w5948 & w9953 ;
  assign w13863 = w10965 | w13861 ;
  assign w13864 = ( w5497 & w13861 ) | ( w5497 & w13863 ) | ( w13861 & w13863 ) ;
  assign w13865 = ( w9953 & ~w13862 ) | ( w9953 & w13864 ) | ( ~w13862 & w13864 ) ;
  assign w13866 = \pi17 ^ w13865 ;
  assign w13867 = ( w13644 & w13858 ) | ( w13644 & w13866 ) | ( w13858 & w13866 ) ;
  assign w13868 = ~w6549 & w10784 ;
  assign w13869 = w6048 & w10211 ;
  assign w13870 = ( w10784 & ~w13868 ) | ( w10784 & w13869 ) | ( ~w13868 & w13869 ) ;
  assign w13871 = w6637 | w10805 ;
  assign w13872 = w10855 & ~w13870 ;
  assign w13873 = ( w6045 & w13870 ) | ( w6045 & ~w13872 ) | ( w13870 & ~w13872 ) ;
  assign w13874 = ( ~w10805 & w13871 ) | ( ~w10805 & w13873 ) | ( w13871 & w13873 ) ;
  assign w13875 = \pi14 ^ w13874 ;
  assign w13876 = ( ~w13642 & w13867 ) | ( ~w13642 & w13875 ) | ( w13867 & w13875 ) ;
  assign w13877 = ( ~w13632 & w13640 ) | ( ~w13632 & w13876 ) | ( w13640 & w13876 ) ;
  assign w13878 = w6949 | w10885 ;
  assign w13879 = w6748 & ~w10866 ;
  assign w13880 = ( ~w10885 & w13878 ) | ( ~w10885 & w13879 ) | ( w13878 & w13879 ) ;
  assign w13881 = w7154 | w10887 ;
  assign w13882 = w11131 & ~w13880 ;
  assign w13883 = ( w6751 & w13880 ) | ( w6751 & ~w13882 ) | ( w13880 & ~w13882 ) ;
  assign w13884 = ( ~w10887 & w13881 ) | ( ~w10887 & w13883 ) | ( w13881 & w13883 ) ;
  assign w13885 = \pi11 ^ w13884 ;
  assign w13886 = ( w13630 & w13877 ) | ( w13630 & w13885 ) | ( w13877 & w13885 ) ;
  assign w13887 = ( w7411 & w7673 ) | ( w7411 & ~w11138 ) | ( w7673 & ~w11138 ) ;
  assign w13888 = w7673 & ~w13887 ;
  assign w13889 = ( w7944 & ~w13887 ) | ( w7944 & w13888 ) | ( ~w13887 & w13888 ) ;
  assign w13890 = ( ~w10738 & w13887 ) | ( ~w10738 & w13889 ) | ( w13887 & w13889 ) ;
  assign w13891 = w13383 ^ w13608 ;
  assign w13892 = w13616 ^ w13891 ;
  assign w13893 = w11146 & ~w13890 ;
  assign w13894 = ( w7414 & w13890 ) | ( w7414 & ~w13893 ) | ( w13890 & ~w13893 ) ;
  assign w13895 = \pi08 ^ w13894 ;
  assign w13896 = ( w13886 & ~w13892 ) | ( w13886 & w13895 ) | ( ~w13892 & w13895 ) ;
  assign w13897 = w13617 ^ w13627 ;
  assign w13898 = w13625 ^ w13897 ;
  assign w13899 = w7414 & w11146 ;
  assign w13900 = ( w7414 & w13890 ) | ( w7414 & ~w13899 ) | ( w13890 & ~w13899 ) ;
  assign w13901 = w13892 ^ w13900 ;
  assign w13902 = \pi08 ^ w13886 ;
  assign w13903 = w13901 ^ w13902 ;
  assign w13904 = w13630 ^ w13877 ;
  assign w13905 = w13885 ^ w13904 ;
  assign w13906 = w13632 ^ w13876 ;
  assign w13907 = w13640 ^ w13906 ;
  assign w13908 = w6949 | w10866 ;
  assign w13909 = w6748 & w10801 ;
  assign w13910 = ( ~w10866 & w13908 ) | ( ~w10866 & w13909 ) | ( w13908 & w13909 ) ;
  assign w13911 = w7154 | w10885 ;
  assign w13912 = w11160 & ~w13910 ;
  assign w13913 = ( w6751 & w13910 ) | ( w6751 & ~w13912 ) | ( w13910 & ~w13912 ) ;
  assign w13914 = ( ~w10885 & w13911 ) | ( ~w10885 & w13913 ) | ( w13911 & w13913 ) ;
  assign w13915 = \pi11 ^ w13914 ;
  assign w13916 = w13642 ^ w13867 ;
  assign w13917 = w13875 ^ w13916 ;
  assign w13918 = w13644 ^ w13858 ;
  assign w13919 = w13866 ^ w13918 ;
  assign w13920 = w13646 ^ w13857 ;
  assign w13921 = w13849 ^ w13920 ;
  assign w13922 = w13654 ^ w13848 ;
  assign w13923 = w13656 ^ w13922 ;
  assign w13924 = w4905 & ~w9967 ;
  assign w13925 = ( w5395 & w9961 ) | ( w5395 & w13924 ) | ( w9961 & w13924 ) ;
  assign w13926 = w5343 | w13925 ;
  assign w13927 = ( w9965 & w13925 ) | ( w9965 & w13926 ) | ( w13925 & w13926 ) ;
  assign w13928 = w13924 | w13927 ;
  assign w13929 = ~w4908 & w11339 ;
  assign w13930 = ( w11339 & w13928 ) | ( w11339 & ~w13929 ) | ( w13928 & ~w13929 ) ;
  assign w13931 = \pi20 ^ w13930 ;
  assign w13932 = w13664 ^ w13847 ;
  assign w13933 = w13666 ^ w13932 ;
  assign w13934 = w4905 & w9971 ;
  assign w13935 = ( w5395 & w9965 ) | ( w5395 & w13934 ) | ( w9965 & w13934 ) ;
  assign w13936 = w5343 | w13935 ;
  assign w13937 = ( ~w9967 & w13935 ) | ( ~w9967 & w13936 ) | ( w13935 & w13936 ) ;
  assign w13938 = w13934 | w13937 ;
  assign w13939 = w4908 | w11501 ;
  assign w13940 = ( ~w11501 & w13938 ) | ( ~w11501 & w13939 ) | ( w13938 & w13939 ) ;
  assign w13941 = \pi20 ^ w13940 ;
  assign w13942 = w13674 ^ w13846 ;
  assign w13943 = w13676 ^ w13942 ;
  assign w13944 = w4905 & ~w9973 ;
  assign w13945 = ( w5395 & ~w9967 ) | ( w5395 & w13944 ) | ( ~w9967 & w13944 ) ;
  assign w13946 = w5343 | w13945 ;
  assign w13947 = ( w9971 & w13945 ) | ( w9971 & w13946 ) | ( w13945 & w13946 ) ;
  assign w13948 = w13944 | w13947 ;
  assign w13949 = w4908 | w11512 ;
  assign w13950 = ( ~w11512 & w13948 ) | ( ~w11512 & w13949 ) | ( w13948 & w13949 ) ;
  assign w13951 = \pi20 ^ w13950 ;
  assign w13952 = w13684 ^ w13845 ;
  assign w13953 = w13686 ^ w13952 ;
  assign w13954 = w4905 & w9975 ;
  assign w13955 = ( w5395 & w9971 ) | ( w5395 & w13954 ) | ( w9971 & w13954 ) ;
  assign w13956 = w5343 | w13955 ;
  assign w13957 = ( ~w9973 & w13955 ) | ( ~w9973 & w13956 ) | ( w13955 & w13956 ) ;
  assign w13958 = w13954 | w13957 ;
  assign w13959 = w4908 | w11809 ;
  assign w13960 = ( ~w11809 & w13958 ) | ( ~w11809 & w13959 ) | ( w13958 & w13959 ) ;
  assign w13961 = \pi20 ^ w13960 ;
  assign w13962 = w13694 ^ w13844 ;
  assign w13963 = w13696 ^ w13962 ;
  assign w13964 = w4905 & w9977 ;
  assign w13965 = ( w5395 & ~w9973 ) | ( w5395 & w13964 ) | ( ~w9973 & w13964 ) ;
  assign w13966 = w5343 | w13965 ;
  assign w13967 = ( w9975 & w13965 ) | ( w9975 & w13966 ) | ( w13965 & w13966 ) ;
  assign w13968 = w13964 | w13967 ;
  assign w13969 = w4908 | w11671 ;
  assign w13970 = ( ~w11671 & w13968 ) | ( ~w11671 & w13969 ) | ( w13968 & w13969 ) ;
  assign w13971 = \pi20 ^ w13970 ;
  assign w13972 = w13704 ^ w13843 ;
  assign w13973 = w13706 ^ w13972 ;
  assign w13974 = w4905 & w9979 ;
  assign w13975 = ( w5395 & w9975 ) | ( w5395 & w13974 ) | ( w9975 & w13974 ) ;
  assign w13976 = w5343 | w13975 ;
  assign w13977 = ( w9977 & w13975 ) | ( w9977 & w13976 ) | ( w13975 & w13976 ) ;
  assign w13978 = w13974 | w13977 ;
  assign w13979 = ~w4908 & w11914 ;
  assign w13980 = ( w11914 & w13978 ) | ( w11914 & ~w13979 ) | ( w13978 & ~w13979 ) ;
  assign w13981 = \pi20 ^ w13980 ;
  assign w13982 = w13714 ^ w13842 ;
  assign w13983 = w13716 ^ w13982 ;
  assign w13984 = w4905 & w9981 ;
  assign w13985 = ( w5395 & w9977 ) | ( w5395 & w13984 ) | ( w9977 & w13984 ) ;
  assign w13986 = w5343 | w13985 ;
  assign w13987 = ( w9979 & w13985 ) | ( w9979 & w13986 ) | ( w13985 & w13986 ) ;
  assign w13988 = w13984 | w13987 ;
  assign w13989 = ~w4908 & w12106 ;
  assign w13990 = ( w12106 & w13988 ) | ( w12106 & ~w13989 ) | ( w13988 & ~w13989 ) ;
  assign w13991 = \pi20 ^ w13990 ;
  assign w13992 = w13724 ^ w13841 ;
  assign w13993 = w13726 ^ w13992 ;
  assign w13994 = w4905 & w9983 ;
  assign w13995 = ( w5395 & w9979 ) | ( w5395 & w13994 ) | ( w9979 & w13994 ) ;
  assign w13996 = w5343 | w13995 ;
  assign w13997 = ( w9981 & w13995 ) | ( w9981 & w13996 ) | ( w13995 & w13996 ) ;
  assign w13998 = w13994 | w13997 ;
  assign w13999 = ~w4908 & w12010 ;
  assign w14000 = ( w12010 & w13998 ) | ( w12010 & ~w13999 ) | ( w13998 & ~w13999 ) ;
  assign w14001 = \pi20 ^ w14000 ;
  assign w14002 = w13734 ^ w13840 ;
  assign w14003 = w13736 ^ w14002 ;
  assign w14004 = w4905 & w9985 ;
  assign w14005 = ( w5395 & w9981 ) | ( w5395 & w14004 ) | ( w9981 & w14004 ) ;
  assign w14006 = w5343 | w14005 ;
  assign w14007 = ( w9983 & w14005 ) | ( w9983 & w14006 ) | ( w14005 & w14006 ) ;
  assign w14008 = w14004 | w14007 ;
  assign w14009 = ~w4908 & w12236 ;
  assign w14010 = ( w12236 & w14008 ) | ( w12236 & ~w14009 ) | ( w14008 & ~w14009 ) ;
  assign w14011 = \pi20 ^ w14010 ;
  assign w14012 = w13744 ^ w13839 ;
  assign w14013 = w13746 ^ w14012 ;
  assign w14014 = w4905 & w9987 ;
  assign w14015 = ( w5395 & w9983 ) | ( w5395 & w14014 ) | ( w9983 & w14014 ) ;
  assign w14016 = w5343 | w14015 ;
  assign w14017 = ( w9985 & w14015 ) | ( w9985 & w14016 ) | ( w14015 & w14016 ) ;
  assign w14018 = w14014 | w14017 ;
  assign w14019 = ~w4908 & w12433 ;
  assign w14020 = ( w12433 & w14018 ) | ( w12433 & ~w14019 ) | ( w14018 & ~w14019 ) ;
  assign w14021 = \pi20 ^ w14020 ;
  assign w14022 = ~w5343 & w9987 ;
  assign w14023 = w4905 & ~w9989 ;
  assign w14024 = ( w9987 & ~w14022 ) | ( w9987 & w14023 ) | ( ~w14022 & w14023 ) ;
  assign w14025 = ~w5395 & w9985 ;
  assign w14026 = w12446 | w14024 ;
  assign w14027 = ( w4908 & w14024 ) | ( w4908 & w14026 ) | ( w14024 & w14026 ) ;
  assign w14028 = ( w9985 & ~w14025 ) | ( w9985 & w14027 ) | ( ~w14025 & w14027 ) ;
  assign w14029 = \pi20 ^ w14028 ;
  assign w14030 = w13756 ^ w13838 ;
  assign w14031 = w13748 ^ w14030 ;
  assign w14032 = w5343 | w9989 ;
  assign w14033 = w4905 & w9991 ;
  assign w14034 = ( ~w9989 & w14032 ) | ( ~w9989 & w14033 ) | ( w14032 & w14033 ) ;
  assign w14035 = ~w5395 & w9987 ;
  assign w14036 = w12217 & ~w14034 ;
  assign w14037 = ( w4908 & w14034 ) | ( w4908 & ~w14036 ) | ( w14034 & ~w14036 ) ;
  assign w14038 = ( w9987 & ~w14035 ) | ( w9987 & w14037 ) | ( ~w14035 & w14037 ) ;
  assign w14039 = \pi20 ^ w14038 ;
  assign w14040 = w13766 ^ w13837 ;
  assign w14041 = w13758 ^ w14040 ;
  assign w14042 = w13774 ^ w13836 ;
  assign w14043 = w13776 ^ w14042 ;
  assign w14044 = w4905 & ~w9993 ;
  assign w14045 = ( w5395 & ~w9989 ) | ( w5395 & w14044 ) | ( ~w9989 & w14044 ) ;
  assign w14046 = w5343 | w14045 ;
  assign w14047 = ( w9991 & w14045 ) | ( w9991 & w14046 ) | ( w14045 & w14046 ) ;
  assign w14048 = w14044 | w14047 ;
  assign w14049 = w4908 | w12484 ;
  assign w14050 = ( ~w12484 & w14048 ) | ( ~w12484 & w14049 ) | ( w14048 & w14049 ) ;
  assign w14051 = \pi20 ^ w14050 ;
  assign w14052 = w13786 ^ w13835 ;
  assign w14053 = w13778 ^ w14052 ;
  assign w14054 = w4905 & w9995 ;
  assign w14055 = ( w5395 & w9991 ) | ( w5395 & w14054 ) | ( w9991 & w14054 ) ;
  assign w14056 = w5343 | w14055 ;
  assign w14057 = ( ~w9993 & w14055 ) | ( ~w9993 & w14056 ) | ( w14055 & w14056 ) ;
  assign w14058 = w14054 | w14057 ;
  assign w14059 = w4908 | w12514 ;
  assign w14060 = ( ~w12514 & w14058 ) | ( ~w12514 & w14059 ) | ( w14058 & w14059 ) ;
  assign w14061 = \pi20 ^ w14060 ;
  assign w14062 = w13794 ^ w13834 ;
  assign w14063 = w13795 ^ w14062 ;
  assign w14064 = w4905 & w9997 ;
  assign w14065 = ( w5395 & ~w9993 ) | ( w5395 & w14064 ) | ( ~w9993 & w14064 ) ;
  assign w14066 = w5343 | w14065 ;
  assign w14067 = ( w9995 & w14065 ) | ( w9995 & w14066 ) | ( w14065 & w14066 ) ;
  assign w14068 = w14064 | w14067 ;
  assign w14069 = w4908 | w12541 ;
  assign w14070 = ( ~w12541 & w14068 ) | ( ~w12541 & w14069 ) | ( w14068 & w14069 ) ;
  assign w14071 = \pi20 ^ w14070 ;
  assign w14072 = ~w5343 & w9997 ;
  assign w14073 = w4905 & w9999 ;
  assign w14074 = ( w9997 & ~w14072 ) | ( w9997 & w14073 ) | ( ~w14072 & w14073 ) ;
  assign w14075 = ~w5395 & w9995 ;
  assign w14076 = w12572 | w14074 ;
  assign w14077 = ( w4908 & w14074 ) | ( w4908 & w14076 ) | ( w14074 & w14076 ) ;
  assign w14078 = ( w9995 & ~w14075 ) | ( w9995 & w14077 ) | ( ~w14075 & w14077 ) ;
  assign w14079 = \pi20 ^ w14078 ;
  assign w14080 = w13808 ^ w13833 ;
  assign w14081 = w13800 ^ w14080 ;
  assign w14082 = w13823 ^ w13831 ;
  assign w14083 = w13832 ^ w14082 ;
  assign w14084 = w4905 & w10001 ;
  assign w14085 = ( w5395 & w9997 ) | ( w5395 & w14084 ) | ( w9997 & w14084 ) ;
  assign w14086 = w5343 | w14085 ;
  assign w14087 = ( w9999 & w14085 ) | ( w9999 & w14086 ) | ( w14085 & w14086 ) ;
  assign w14088 = w14084 | w14087 ;
  assign w14089 = ~w4908 & w12641 ;
  assign w14090 = ( w12641 & w14088 ) | ( w12641 & ~w14089 ) | ( w14088 & ~w14089 ) ;
  assign w14091 = \pi20 ^ w14090 ;
  assign w14092 = ~w5343 & w10001 ;
  assign w14093 = w4905 & ~w10006 ;
  assign w14094 = ( w10001 & ~w14092 ) | ( w10001 & w14093 ) | ( ~w14092 & w14093 ) ;
  assign w14095 = ~w5395 & w9999 ;
  assign w14096 = w12691 & ~w14094 ;
  assign w14097 = ( w4908 & w14094 ) | ( w4908 & ~w14096 ) | ( w14094 & ~w14096 ) ;
  assign w14098 = ( w9999 & ~w14095 ) | ( w9999 & w14097 ) | ( ~w14095 & w14097 ) ;
  assign w14099 = \pi20 ^ w14098 ;
  assign w14100 = w13814 ^ w13822 ;
  assign w14101 = ( \pi20 & \pi21 ) | ( \pi20 & ~w10016 ) | ( \pi21 & ~w10016 ) ;
  assign w14102 = ( \pi20 & \pi21 ) | ( \pi20 & ~w10021 ) | ( \pi21 & ~w10021 ) ;
  assign w14103 = \pi22 ^ w10021 ;
  assign w14104 = ( \pi22 & w14102 ) | ( \pi22 & w14103 ) | ( w14102 & w14103 ) ;
  assign w14105 = w14101 ^ w14104 ;
  assign w14106 = w4905 & w10011 ;
  assign w14107 = ( w5395 & w10001 ) | ( w5395 & w14106 ) | ( w10001 & w14106 ) ;
  assign w14108 = w5343 | w14107 ;
  assign w14109 = ( ~w10006 & w14107 ) | ( ~w10006 & w14108 ) | ( w14107 & w14108 ) ;
  assign w14110 = w14106 | w14109 ;
  assign w14111 = ~w4908 & w12747 ;
  assign w14112 = ( w12747 & w14110 ) | ( w12747 & ~w14111 ) | ( w14110 & ~w14111 ) ;
  assign w14113 = \pi20 ^ w14112 ;
  assign w14114 = \pi20 & w10021 ;
  assign w14115 = w10016 & w14114 ;
  assign w14116 = ( \pi17 & \pi18 ) | ( \pi17 & ~w14115 ) | ( \pi18 & ~w14115 ) ;
  assign w14117 = ( \pi19 & \pi20 ) | ( \pi19 & ~w14116 ) | ( \pi20 & ~w14116 ) ;
  assign w14118 = ( \pi19 & ~w14114 ) | ( \pi19 & w14116 ) | ( ~w14114 & w14116 ) ;
  assign w14119 = ( w7590 & w14117 ) | ( w7590 & ~w14118 ) | ( w14117 & ~w14118 ) ;
  assign w14120 = w4905 & ~w10021 ;
  assign w14121 = ( w5395 & w10011 ) | ( w5395 & w14120 ) | ( w10011 & w14120 ) ;
  assign w14122 = w5343 | w14121 ;
  assign w14123 = ( ~w10016 & w14121 ) | ( ~w10016 & w14122 ) | ( w14121 & w14122 ) ;
  assign w14124 = w14120 | w14123 ;
  assign w14125 = ~w4908 & w12867 ;
  assign w14126 = ( w12867 & w14124 ) | ( w12867 & ~w14125 ) | ( w14124 & ~w14125 ) ;
  assign w14127 = \pi20 ^ w14126 ;
  assign w14128 = w14119 & w14127 ;
  assign w14129 = ~w5343 & w10011 ;
  assign w14130 = w4905 & ~w10016 ;
  assign w14131 = ( w10011 & ~w14129 ) | ( w10011 & w14130 ) | ( ~w14129 & w14130 ) ;
  assign w14132 = w5395 | w10006 ;
  assign w14133 = w12777 | w14131 ;
  assign w14134 = ( w4908 & w14131 ) | ( w4908 & w14133 ) | ( w14131 & w14133 ) ;
  assign w14135 = ( ~w10006 & w14132 ) | ( ~w10006 & w14134 ) | ( w14132 & w14134 ) ;
  assign w14136 = \pi20 ^ w14135 ;
  assign w14137 = w4608 & ~w10021 ;
  assign w14138 = ( w14128 & w14136 ) | ( w14128 & w14137 ) | ( w14136 & w14137 ) ;
  assign w14139 = ( w14105 & w14113 ) | ( w14105 & w14138 ) | ( w14113 & w14138 ) ;
  assign w14140 = ( w14099 & w14100 ) | ( w14099 & w14139 ) | ( w14100 & w14139 ) ;
  assign w14141 = ( w14083 & w14091 ) | ( w14083 & w14140 ) | ( w14091 & w14140 ) ;
  assign w14142 = ( w14079 & w14081 ) | ( w14079 & w14141 ) | ( w14081 & w14141 ) ;
  assign w14143 = ( w14063 & w14071 ) | ( w14063 & w14142 ) | ( w14071 & w14142 ) ;
  assign w14144 = ( w14053 & w14061 ) | ( w14053 & w14143 ) | ( w14061 & w14143 ) ;
  assign w14145 = ( w14043 & w14051 ) | ( w14043 & w14144 ) | ( w14051 & w14144 ) ;
  assign w14146 = ( w14039 & w14041 ) | ( w14039 & w14145 ) | ( w14041 & w14145 ) ;
  assign w14147 = ( w14029 & w14031 ) | ( w14029 & w14146 ) | ( w14031 & w14146 ) ;
  assign w14148 = ( ~w14013 & w14021 ) | ( ~w14013 & w14147 ) | ( w14021 & w14147 ) ;
  assign w14149 = ( ~w14003 & w14011 ) | ( ~w14003 & w14148 ) | ( w14011 & w14148 ) ;
  assign w14150 = ( w13993 & w14001 ) | ( w13993 & w14149 ) | ( w14001 & w14149 ) ;
  assign w14151 = ( ~w13983 & w13991 ) | ( ~w13983 & w14150 ) | ( w13991 & w14150 ) ;
  assign w14152 = ( ~w13973 & w13981 ) | ( ~w13973 & w14151 ) | ( w13981 & w14151 ) ;
  assign w14153 = ( w13963 & w13971 ) | ( w13963 & w14152 ) | ( w13971 & w14152 ) ;
  assign w14154 = ( w13953 & w13961 ) | ( w13953 & w14153 ) | ( w13961 & w14153 ) ;
  assign w14155 = ( w13943 & w13951 ) | ( w13943 & w14154 ) | ( w13951 & w14154 ) ;
  assign w14156 = ( w13933 & w13941 ) | ( w13933 & w14155 ) | ( w13941 & w14155 ) ;
  assign w14157 = ( w13923 & w13931 ) | ( w13923 & w14156 ) | ( w13931 & w14156 ) ;
  assign w14158 = w5710 | w9955 ;
  assign w14159 = w5494 & w9957 ;
  assign w14160 = ( ~w9955 & w14158 ) | ( ~w9955 & w14159 ) | ( w14158 & w14159 ) ;
  assign w14161 = ~w5948 & w9842 ;
  assign w14162 = w10976 & ~w14160 ;
  assign w14163 = ( w5497 & w14160 ) | ( w5497 & ~w14162 ) | ( w14160 & ~w14162 ) ;
  assign w14164 = ( w9842 & ~w14161 ) | ( w9842 & w14163 ) | ( ~w14161 & w14163 ) ;
  assign w14165 = \pi17 ^ w14164 ;
  assign w14166 = ( ~w13921 & w14157 ) | ( ~w13921 & w14165 ) | ( w14157 & w14165 ) ;
  assign w14167 = ~w6549 & w10211 ;
  assign w14168 = w6048 & w10114 ;
  assign w14169 = ( w10211 & ~w14167 ) | ( w10211 & w14168 ) | ( ~w14167 & w14168 ) ;
  assign w14170 = ~w6637 & w10784 ;
  assign w14171 = w10789 | w14169 ;
  assign w14172 = ( w6045 & w14169 ) | ( w6045 & w14171 ) | ( w14169 & w14171 ) ;
  assign w14173 = ( w10784 & ~w14170 ) | ( w10784 & w14172 ) | ( ~w14170 & w14172 ) ;
  assign w14174 = \pi14 ^ w14173 ;
  assign w14175 = ( w13919 & w14166 ) | ( w13919 & w14174 ) | ( w14166 & w14174 ) ;
  assign w14176 = ~w6949 & w10801 ;
  assign w14177 = w6748 & ~w10807 ;
  assign w14178 = ( w10801 & ~w14176 ) | ( w10801 & w14177 ) | ( ~w14176 & w14177 ) ;
  assign w14179 = w7154 | w10866 ;
  assign w14180 = w10874 | w14178 ;
  assign w14181 = ( w6751 & w14178 ) | ( w6751 & w14180 ) | ( w14178 & w14180 ) ;
  assign w14182 = ( ~w10866 & w14179 ) | ( ~w10866 & w14181 ) | ( w14179 & w14181 ) ;
  assign w14183 = \pi11 ^ w14182 ;
  assign w14184 = ( ~w13917 & w14175 ) | ( ~w13917 & w14183 ) | ( w14175 & w14183 ) ;
  assign w14185 = ( ~w13907 & w13915 ) | ( ~w13907 & w14184 ) | ( w13915 & w14184 ) ;
  assign w14186 = w7673 | w11139 ;
  assign w14187 = w7411 & w10883 ;
  assign w14188 = ( ~w11139 & w14186 ) | ( ~w11139 & w14187 ) | ( w14186 & w14187 ) ;
  assign w14189 = w7944 | w10738 ;
  assign w14190 = w11145 & ~w14188 ;
  assign w14191 = ( w7414 & w14188 ) | ( w7414 & ~w14190 ) | ( w14188 & ~w14190 ) ;
  assign w14192 = ( ~w10738 & w14189 ) | ( ~w10738 & w14191 ) | ( w14189 & w14191 ) ;
  assign w14193 = \pi08 ^ w14192 ;
  assign w14194 = ( w13905 & w14185 ) | ( w13905 & w14193 ) | ( w14185 & w14193 ) ;
  assign w14195 = w13905 ^ w14185 ;
  assign w14196 = w14193 ^ w14195 ;
  assign w14197 = w13917 ^ w14175 ;
  assign w14198 = w14183 ^ w14197 ;
  assign w14199 = w13919 ^ w14166 ;
  assign w14200 = w14174 ^ w14199 ;
  assign w14201 = w13921 ^ w14165 ;
  assign w14202 = w14157 ^ w14201 ;
  assign w14203 = ~w5710 & w9957 ;
  assign w14204 = w5494 & ~w9963 ;
  assign w14205 = ( w9957 & ~w14203 ) | ( w9957 & w14204 ) | ( ~w14203 & w14204 ) ;
  assign w14206 = w5948 | w9955 ;
  assign w14207 = w11202 & ~w14205 ;
  assign w14208 = ( w5497 & w14205 ) | ( w5497 & ~w14207 ) | ( w14205 & ~w14207 ) ;
  assign w14209 = ( ~w9955 & w14206 ) | ( ~w9955 & w14208 ) | ( w14206 & w14208 ) ;
  assign w14210 = \pi17 ^ w14209 ;
  assign w14211 = w13931 ^ w14156 ;
  assign w14212 = w13923 ^ w14211 ;
  assign w14213 = w5710 | w9963 ;
  assign w14214 = w5494 & w9961 ;
  assign w14215 = ( ~w9963 & w14213 ) | ( ~w9963 & w14214 ) | ( w14213 & w14214 ) ;
  assign w14216 = ~w5948 & w9957 ;
  assign w14217 = w11089 & ~w14215 ;
  assign w14218 = ( w5497 & w14215 ) | ( w5497 & ~w14217 ) | ( w14215 & ~w14217 ) ;
  assign w14219 = ( w9957 & ~w14216 ) | ( w9957 & w14218 ) | ( ~w14216 & w14218 ) ;
  assign w14220 = \pi17 ^ w14219 ;
  assign w14221 = w13941 ^ w14155 ;
  assign w14222 = w13933 ^ w14221 ;
  assign w14223 = ~w5710 & w9961 ;
  assign w14224 = w5494 & w9965 ;
  assign w14225 = ( w9961 & ~w14223 ) | ( w9961 & w14224 ) | ( ~w14223 & w14224 ) ;
  assign w14226 = w5948 | w9963 ;
  assign w14227 = w11278 & ~w14225 ;
  assign w14228 = ( w5497 & w14225 ) | ( w5497 & ~w14227 ) | ( w14225 & ~w14227 ) ;
  assign w14229 = ( ~w9963 & w14226 ) | ( ~w9963 & w14228 ) | ( w14226 & w14228 ) ;
  assign w14230 = \pi17 ^ w14229 ;
  assign w14231 = w13951 ^ w14154 ;
  assign w14232 = w13943 ^ w14231 ;
  assign w14233 = ~w5710 & w9965 ;
  assign w14234 = w5494 & ~w9967 ;
  assign w14235 = ( w9965 & ~w14233 ) | ( w9965 & w14234 ) | ( ~w14233 & w14234 ) ;
  assign w14236 = ~w5948 & w9961 ;
  assign w14237 = w11339 | w14235 ;
  assign w14238 = ( w5497 & w14235 ) | ( w5497 & w14237 ) | ( w14235 & w14237 ) ;
  assign w14239 = ( w9961 & ~w14236 ) | ( w9961 & w14238 ) | ( ~w14236 & w14238 ) ;
  assign w14240 = \pi17 ^ w14239 ;
  assign w14241 = w13961 ^ w14153 ;
  assign w14242 = w13953 ^ w14241 ;
  assign w14243 = w5710 | w9967 ;
  assign w14244 = w5494 & w9971 ;
  assign w14245 = ( ~w9967 & w14243 ) | ( ~w9967 & w14244 ) | ( w14243 & w14244 ) ;
  assign w14246 = ~w5948 & w9965 ;
  assign w14247 = w11501 & ~w14245 ;
  assign w14248 = ( w5497 & w14245 ) | ( w5497 & ~w14247 ) | ( w14245 & ~w14247 ) ;
  assign w14249 = ( w9965 & ~w14246 ) | ( w9965 & w14248 ) | ( ~w14246 & w14248 ) ;
  assign w14250 = \pi17 ^ w14249 ;
  assign w14251 = w13971 ^ w14152 ;
  assign w14252 = w13963 ^ w14251 ;
  assign w14253 = ~w5710 & w9971 ;
  assign w14254 = w5494 & ~w9973 ;
  assign w14255 = ( w9971 & ~w14253 ) | ( w9971 & w14254 ) | ( ~w14253 & w14254 ) ;
  assign w14256 = w5948 | w9967 ;
  assign w14257 = w11512 & ~w14255 ;
  assign w14258 = ( w5497 & w14255 ) | ( w5497 & ~w14257 ) | ( w14255 & ~w14257 ) ;
  assign w14259 = ( ~w9967 & w14256 ) | ( ~w9967 & w14258 ) | ( w14256 & w14258 ) ;
  assign w14260 = \pi17 ^ w14259 ;
  assign w14261 = w13981 ^ w14151 ;
  assign w14262 = w13973 ^ w14261 ;
  assign w14263 = w5710 | w9973 ;
  assign w14264 = w5494 & w9975 ;
  assign w14265 = ( ~w9973 & w14263 ) | ( ~w9973 & w14264 ) | ( w14263 & w14264 ) ;
  assign w14266 = ~w5948 & w9971 ;
  assign w14267 = w11809 & ~w14265 ;
  assign w14268 = ( w5497 & w14265 ) | ( w5497 & ~w14267 ) | ( w14265 & ~w14267 ) ;
  assign w14269 = ( w9971 & ~w14266 ) | ( w9971 & w14268 ) | ( ~w14266 & w14268 ) ;
  assign w14270 = \pi17 ^ w14269 ;
  assign w14271 = w13991 ^ w14150 ;
  assign w14272 = w13983 ^ w14271 ;
  assign w14273 = ~w5710 & w9975 ;
  assign w14274 = w5494 & w9977 ;
  assign w14275 = ( w9975 & ~w14273 ) | ( w9975 & w14274 ) | ( ~w14273 & w14274 ) ;
  assign w14276 = w5948 | w9973 ;
  assign w14277 = w11671 & ~w14275 ;
  assign w14278 = ( w5497 & w14275 ) | ( w5497 & ~w14277 ) | ( w14275 & ~w14277 ) ;
  assign w14279 = ( ~w9973 & w14276 ) | ( ~w9973 & w14278 ) | ( w14276 & w14278 ) ;
  assign w14280 = \pi17 ^ w14279 ;
  assign w14281 = w14001 ^ w14149 ;
  assign w14282 = w13993 ^ w14281 ;
  assign w14283 = ~w5710 & w9977 ;
  assign w14284 = w5494 & w9979 ;
  assign w14285 = ( w9977 & ~w14283 ) | ( w9977 & w14284 ) | ( ~w14283 & w14284 ) ;
  assign w14286 = ~w5948 & w9975 ;
  assign w14287 = w11914 | w14285 ;
  assign w14288 = ( w5497 & w14285 ) | ( w5497 & w14287 ) | ( w14285 & w14287 ) ;
  assign w14289 = ( w9975 & ~w14286 ) | ( w9975 & w14288 ) | ( ~w14286 & w14288 ) ;
  assign w14290 = \pi17 ^ w14289 ;
  assign w14291 = w14011 ^ w14148 ;
  assign w14292 = w14003 ^ w14291 ;
  assign w14293 = ~w5710 & w9979 ;
  assign w14294 = w5494 & w9981 ;
  assign w14295 = ( w9979 & ~w14293 ) | ( w9979 & w14294 ) | ( ~w14293 & w14294 ) ;
  assign w14296 = ~w5948 & w9977 ;
  assign w14297 = w12106 | w14295 ;
  assign w14298 = ( w5497 & w14295 ) | ( w5497 & w14297 ) | ( w14295 & w14297 ) ;
  assign w14299 = ( w9977 & ~w14296 ) | ( w9977 & w14298 ) | ( ~w14296 & w14298 ) ;
  assign w14300 = \pi17 ^ w14299 ;
  assign w14301 = w14021 ^ w14147 ;
  assign w14302 = w14013 ^ w14301 ;
  assign w14303 = w14029 ^ w14146 ;
  assign w14304 = w14031 ^ w14303 ;
  assign w14305 = w5494 & w9983 ;
  assign w14306 = ( w5948 & w9979 ) | ( w5948 & w14305 ) | ( w9979 & w14305 ) ;
  assign w14307 = w5710 | w14306 ;
  assign w14308 = ( w9981 & w14306 ) | ( w9981 & w14307 ) | ( w14306 & w14307 ) ;
  assign w14309 = w14305 | w14308 ;
  assign w14310 = ~w5497 & w12010 ;
  assign w14311 = ( w12010 & w14309 ) | ( w12010 & ~w14310 ) | ( w14309 & ~w14310 ) ;
  assign w14312 = \pi17 ^ w14311 ;
  assign w14313 = w14039 ^ w14145 ;
  assign w14314 = w14041 ^ w14313 ;
  assign w14315 = w5494 & w9985 ;
  assign w14316 = ( w5948 & w9981 ) | ( w5948 & w14315 ) | ( w9981 & w14315 ) ;
  assign w14317 = w5710 | w14316 ;
  assign w14318 = ( w9983 & w14316 ) | ( w9983 & w14317 ) | ( w14316 & w14317 ) ;
  assign w14319 = w14315 | w14318 ;
  assign w14320 = ~w5497 & w12236 ;
  assign w14321 = ( w12236 & w14319 ) | ( w12236 & ~w14320 ) | ( w14319 & ~w14320 ) ;
  assign w14322 = \pi17 ^ w14321 ;
  assign w14323 = ~w5710 & w9985 ;
  assign w14324 = w5494 & w9987 ;
  assign w14325 = ( w9985 & ~w14323 ) | ( w9985 & w14324 ) | ( ~w14323 & w14324 ) ;
  assign w14326 = ~w5948 & w9983 ;
  assign w14327 = w12433 | w14325 ;
  assign w14328 = ( w5497 & w14325 ) | ( w5497 & w14327 ) | ( w14325 & w14327 ) ;
  assign w14329 = ( w9983 & ~w14326 ) | ( w9983 & w14328 ) | ( ~w14326 & w14328 ) ;
  assign w14330 = \pi17 ^ w14329 ;
  assign w14331 = w14051 ^ w14144 ;
  assign w14332 = w14043 ^ w14331 ;
  assign w14333 = ~w5710 & w9987 ;
  assign w14334 = w5494 & ~w9989 ;
  assign w14335 = ( w9987 & ~w14333 ) | ( w9987 & w14334 ) | ( ~w14333 & w14334 ) ;
  assign w14336 = ~w5948 & w9985 ;
  assign w14337 = w12446 | w14335 ;
  assign w14338 = ( w5497 & w14335 ) | ( w5497 & w14337 ) | ( w14335 & w14337 ) ;
  assign w14339 = ( w9985 & ~w14336 ) | ( w9985 & w14338 ) | ( ~w14336 & w14338 ) ;
  assign w14340 = \pi17 ^ w14339 ;
  assign w14341 = w14061 ^ w14143 ;
  assign w14342 = w14053 ^ w14341 ;
  assign w14343 = w5710 | w9989 ;
  assign w14344 = w5494 & w9991 ;
  assign w14345 = ( ~w9989 & w14343 ) | ( ~w9989 & w14344 ) | ( w14343 & w14344 ) ;
  assign w14346 = ~w5948 & w9987 ;
  assign w14347 = w12217 & ~w14345 ;
  assign w14348 = ( w5497 & w14345 ) | ( w5497 & ~w14347 ) | ( w14345 & ~w14347 ) ;
  assign w14349 = ( w9987 & ~w14346 ) | ( w9987 & w14348 ) | ( ~w14346 & w14348 ) ;
  assign w14350 = \pi17 ^ w14349 ;
  assign w14351 = w14071 ^ w14142 ;
  assign w14352 = w14063 ^ w14351 ;
  assign w14353 = w14079 ^ w14141 ;
  assign w14354 = w14081 ^ w14353 ;
  assign w14355 = w5494 & ~w9993 ;
  assign w14356 = ( w5948 & ~w9989 ) | ( w5948 & w14355 ) | ( ~w9989 & w14355 ) ;
  assign w14357 = w5710 | w14356 ;
  assign w14358 = ( w9991 & w14356 ) | ( w9991 & w14357 ) | ( w14356 & w14357 ) ;
  assign w14359 = w14355 | w14358 ;
  assign w14360 = w5497 | w12484 ;
  assign w14361 = ( ~w12484 & w14359 ) | ( ~w12484 & w14360 ) | ( w14359 & w14360 ) ;
  assign w14362 = \pi17 ^ w14361 ;
  assign w14363 = w14091 ^ w14140 ;
  assign w14364 = w14083 ^ w14363 ;
  assign w14365 = w5494 & w9995 ;
  assign w14366 = ( w5948 & w9991 ) | ( w5948 & w14365 ) | ( w9991 & w14365 ) ;
  assign w14367 = w5710 | w14366 ;
  assign w14368 = ( ~w9993 & w14366 ) | ( ~w9993 & w14367 ) | ( w14366 & w14367 ) ;
  assign w14369 = w14365 | w14368 ;
  assign w14370 = w5497 | w12514 ;
  assign w14371 = ( ~w12514 & w14369 ) | ( ~w12514 & w14370 ) | ( w14369 & w14370 ) ;
  assign w14372 = \pi17 ^ w14371 ;
  assign w14373 = w14099 ^ w14139 ;
  assign w14374 = w14100 ^ w14373 ;
  assign w14375 = w5494 & w9997 ;
  assign w14376 = ( w5948 & ~w9993 ) | ( w5948 & w14375 ) | ( ~w9993 & w14375 ) ;
  assign w14377 = w5710 | w14376 ;
  assign w14378 = ( w9995 & w14376 ) | ( w9995 & w14377 ) | ( w14376 & w14377 ) ;
  assign w14379 = w14375 | w14378 ;
  assign w14380 = w5497 | w12541 ;
  assign w14381 = ( ~w12541 & w14379 ) | ( ~w12541 & w14380 ) | ( w14379 & w14380 ) ;
  assign w14382 = \pi17 ^ w14381 ;
  assign w14383 = ~w5710 & w9997 ;
  assign w14384 = w5494 & w9999 ;
  assign w14385 = ( w9997 & ~w14383 ) | ( w9997 & w14384 ) | ( ~w14383 & w14384 ) ;
  assign w14386 = ~w5948 & w9995 ;
  assign w14387 = w12572 | w14385 ;
  assign w14388 = ( w5497 & w14385 ) | ( w5497 & w14387 ) | ( w14385 & w14387 ) ;
  assign w14389 = ( w9995 & ~w14386 ) | ( w9995 & w14388 ) | ( ~w14386 & w14388 ) ;
  assign w14390 = \pi17 ^ w14389 ;
  assign w14391 = w14113 ^ w14138 ;
  assign w14392 = w14105 ^ w14391 ;
  assign w14393 = w14128 ^ w14136 ;
  assign w14394 = w14137 ^ w14393 ;
  assign w14395 = w5494 & w10001 ;
  assign w14396 = ( w5948 & w9997 ) | ( w5948 & w14395 ) | ( w9997 & w14395 ) ;
  assign w14397 = w5710 | w14396 ;
  assign w14398 = ( w9999 & w14396 ) | ( w9999 & w14397 ) | ( w14396 & w14397 ) ;
  assign w14399 = w14395 | w14398 ;
  assign w14400 = ~w5497 & w12641 ;
  assign w14401 = ( w12641 & w14399 ) | ( w12641 & ~w14400 ) | ( w14399 & ~w14400 ) ;
  assign w14402 = \pi17 ^ w14401 ;
  assign w14403 = ~w5710 & w10001 ;
  assign w14404 = w5494 & ~w10006 ;
  assign w14405 = ( w10001 & ~w14403 ) | ( w10001 & w14404 ) | ( ~w14403 & w14404 ) ;
  assign w14406 = ~w5948 & w9999 ;
  assign w14407 = w12691 & ~w14405 ;
  assign w14408 = ( w5497 & w14405 ) | ( w5497 & ~w14407 ) | ( w14405 & ~w14407 ) ;
  assign w14409 = ( w9999 & ~w14406 ) | ( w9999 & w14408 ) | ( ~w14406 & w14408 ) ;
  assign w14410 = \pi17 ^ w14409 ;
  assign w14411 = w14119 ^ w14127 ;
  assign w14412 = ( \pi17 & \pi18 ) | ( \pi17 & ~w10016 ) | ( \pi18 & ~w10016 ) ;
  assign w14413 = ( \pi17 & \pi18 ) | ( \pi17 & ~w10021 ) | ( \pi18 & ~w10021 ) ;
  assign w14414 = \pi19 ^ w10021 ;
  assign w14415 = ( \pi19 & w14413 ) | ( \pi19 & w14414 ) | ( w14413 & w14414 ) ;
  assign w14416 = w14412 ^ w14415 ;
  assign w14417 = w5494 & w10011 ;
  assign w14418 = ( w5948 & w10001 ) | ( w5948 & w14417 ) | ( w10001 & w14417 ) ;
  assign w14419 = w5710 | w14418 ;
  assign w14420 = ( ~w10006 & w14418 ) | ( ~w10006 & w14419 ) | ( w14418 & w14419 ) ;
  assign w14421 = w14417 | w14420 ;
  assign w14422 = ~w5497 & w12747 ;
  assign w14423 = ( w12747 & w14421 ) | ( w12747 & ~w14422 ) | ( w14421 & ~w14422 ) ;
  assign w14424 = \pi17 ^ w14423 ;
  assign w14425 = \pi17 & w10021 ;
  assign w14426 = w10016 & w14425 ;
  assign w14427 = ( \pi14 & \pi15 ) | ( \pi14 & ~w14426 ) | ( \pi15 & ~w14426 ) ;
  assign w14428 = ( \pi16 & \pi17 ) | ( \pi16 & ~w14427 ) | ( \pi17 & ~w14427 ) ;
  assign w14429 = ( \pi16 & ~w14425 ) | ( \pi16 & w14427 ) | ( ~w14425 & w14427 ) ;
  assign w14430 = ( w7879 & w14428 ) | ( w7879 & ~w14429 ) | ( w14428 & ~w14429 ) ;
  assign w14431 = w5494 & ~w10021 ;
  assign w14432 = ( w5948 & w10011 ) | ( w5948 & w14431 ) | ( w10011 & w14431 ) ;
  assign w14433 = w5710 | w14432 ;
  assign w14434 = ( ~w10016 & w14432 ) | ( ~w10016 & w14433 ) | ( w14432 & w14433 ) ;
  assign w14435 = w14431 | w14434 ;
  assign w14436 = ~w5497 & w12867 ;
  assign w14437 = ( w12867 & w14435 ) | ( w12867 & ~w14436 ) | ( w14435 & ~w14436 ) ;
  assign w14438 = \pi17 ^ w14437 ;
  assign w14439 = w14430 & w14438 ;
  assign w14440 = ~w5710 & w10011 ;
  assign w14441 = w5494 & ~w10016 ;
  assign w14442 = ( w10011 & ~w14440 ) | ( w10011 & w14441 ) | ( ~w14440 & w14441 ) ;
  assign w14443 = w5948 | w10006 ;
  assign w14444 = w12777 | w14442 ;
  assign w14445 = ( w5497 & w14442 ) | ( w5497 & w14444 ) | ( w14442 & w14444 ) ;
  assign w14446 = ( ~w10006 & w14443 ) | ( ~w10006 & w14445 ) | ( w14443 & w14445 ) ;
  assign w14447 = \pi17 ^ w14446 ;
  assign w14448 = w4907 & ~w10021 ;
  assign w14449 = ( w14439 & w14447 ) | ( w14439 & w14448 ) | ( w14447 & w14448 ) ;
  assign w14450 = ( w14416 & w14424 ) | ( w14416 & w14449 ) | ( w14424 & w14449 ) ;
  assign w14451 = ( w14410 & w14411 ) | ( w14410 & w14450 ) | ( w14411 & w14450 ) ;
  assign w14452 = ( w14394 & w14402 ) | ( w14394 & w14451 ) | ( w14402 & w14451 ) ;
  assign w14453 = ( w14390 & w14392 ) | ( w14390 & w14452 ) | ( w14392 & w14452 ) ;
  assign w14454 = ( w14374 & w14382 ) | ( w14374 & w14453 ) | ( w14382 & w14453 ) ;
  assign w14455 = ( w14364 & w14372 ) | ( w14364 & w14454 ) | ( w14372 & w14454 ) ;
  assign w14456 = ( w14354 & w14362 ) | ( w14354 & w14455 ) | ( w14362 & w14455 ) ;
  assign w14457 = ( w14350 & w14352 ) | ( w14350 & w14456 ) | ( w14352 & w14456 ) ;
  assign w14458 = ( w14340 & w14342 ) | ( w14340 & w14457 ) | ( w14342 & w14457 ) ;
  assign w14459 = ( w14330 & w14332 ) | ( w14330 & w14458 ) | ( w14332 & w14458 ) ;
  assign w14460 = ( w14314 & w14322 ) | ( w14314 & w14459 ) | ( w14322 & w14459 ) ;
  assign w14461 = ( w14304 & w14312 ) | ( w14304 & w14460 ) | ( w14312 & w14460 ) ;
  assign w14462 = ( w14300 & ~w14302 ) | ( w14300 & w14461 ) | ( ~w14302 & w14461 ) ;
  assign w14463 = ( w14290 & ~w14292 ) | ( w14290 & w14462 ) | ( ~w14292 & w14462 ) ;
  assign w14464 = ( w14280 & w14282 ) | ( w14280 & w14463 ) | ( w14282 & w14463 ) ;
  assign w14465 = ( w14270 & ~w14272 ) | ( w14270 & w14464 ) | ( ~w14272 & w14464 ) ;
  assign w14466 = ( w14260 & ~w14262 ) | ( w14260 & w14465 ) | ( ~w14262 & w14465 ) ;
  assign w14467 = ( w14250 & w14252 ) | ( w14250 & w14466 ) | ( w14252 & w14466 ) ;
  assign w14468 = ( w14240 & w14242 ) | ( w14240 & w14467 ) | ( w14242 & w14467 ) ;
  assign w14469 = ( w14230 & w14232 ) | ( w14230 & w14468 ) | ( w14232 & w14468 ) ;
  assign w14470 = ( w14220 & w14222 ) | ( w14220 & w14469 ) | ( w14222 & w14469 ) ;
  assign w14471 = ( w14210 & w14212 ) | ( w14210 & w14470 ) | ( w14212 & w14470 ) ;
  assign w14472 = ~w6549 & w10114 ;
  assign w14473 = w6048 & w9953 ;
  assign w14474 = ( w10114 & ~w14472 ) | ( w10114 & w14473 ) | ( ~w14472 & w14473 ) ;
  assign w14475 = ~w6637 & w10211 ;
  assign w14476 = w10214 | w14474 ;
  assign w14477 = ( w6045 & w14474 ) | ( w6045 & w14476 ) | ( w14474 & w14476 ) ;
  assign w14478 = ( w10211 & ~w14475 ) | ( w10211 & w14477 ) | ( ~w14475 & w14477 ) ;
  assign w14479 = \pi14 ^ w14478 ;
  assign w14480 = ( ~w14202 & w14471 ) | ( ~w14202 & w14479 ) | ( w14471 & w14479 ) ;
  assign w14481 = w6949 | w10807 ;
  assign w14482 = w6748 & ~w10805 ;
  assign w14483 = ( ~w10807 & w14481 ) | ( ~w10807 & w14482 ) | ( w14481 & w14482 ) ;
  assign w14484 = ~w7154 & w10801 ;
  assign w14485 = w10814 | w14483 ;
  assign w14486 = ( w6751 & w14483 ) | ( w6751 & w14485 ) | ( w14483 & w14485 ) ;
  assign w14487 = ( w10801 & ~w14484 ) | ( w10801 & w14486 ) | ( ~w14484 & w14486 ) ;
  assign w14488 = \pi11 ^ w14487 ;
  assign w14489 = ( w14200 & w14480 ) | ( w14200 & w14488 ) | ( w14480 & w14488 ) ;
  assign w14490 = w7673 | w10887 ;
  assign w14491 = w7411 & ~w10885 ;
  assign w14492 = ( ~w10887 & w14490 ) | ( ~w10887 & w14491 ) | ( w14490 & w14491 ) ;
  assign w14493 = ~w7944 & w10883 ;
  assign w14494 = w10895 | w14492 ;
  assign w14495 = ( w7414 & w14492 ) | ( w7414 & w14494 ) | ( w14492 & w14494 ) ;
  assign w14496 = ( w10883 & ~w14493 ) | ( w10883 & w14495 ) | ( ~w14493 & w14495 ) ;
  assign w14497 = \pi08 ^ w14496 ;
  assign w14498 = ( ~w14198 & w14489 ) | ( ~w14198 & w14497 ) | ( w14489 & w14497 ) ;
  assign w14499 = ~w7673 & w10883 ;
  assign w14500 = w7411 & ~w10887 ;
  assign w14501 = ( w10883 & ~w14499 ) | ( w10883 & w14500 ) | ( ~w14499 & w14500 ) ;
  assign w14502 = w7944 | w11139 ;
  assign w14503 = w11256 | w14501 ;
  assign w14504 = ( w7414 & w14501 ) | ( w7414 & w14503 ) | ( w14501 & w14503 ) ;
  assign w14505 = ( ~w11139 & w14502 ) | ( ~w11139 & w14504 ) | ( w14502 & w14504 ) ;
  assign w14506 = \pi08 ^ w14505 ;
  assign w14507 = w13907 ^ w14184 ;
  assign w14508 = w13915 ^ w14507 ;
  assign w14509 = ( w14498 & w14506 ) | ( w14498 & ~w14508 ) | ( w14506 & ~w14508 ) ;
  assign w14510 = w14200 ^ w14480 ;
  assign w14511 = w14488 ^ w14510 ;
  assign w14512 = w14202 ^ w14479 ;
  assign w14513 = w14471 ^ w14512 ;
  assign w14514 = w14210 ^ w14470 ;
  assign w14515 = w14212 ^ w14514 ;
  assign w14516 = ~w6549 & w9953 ;
  assign w14517 = w6048 & w9842 ;
  assign w14518 = ( w9953 & ~w14516 ) | ( w9953 & w14517 ) | ( ~w14516 & w14517 ) ;
  assign w14519 = ~w6637 & w10114 ;
  assign w14520 = w10334 | w14518 ;
  assign w14521 = ( w6045 & w14518 ) | ( w6045 & w14520 ) | ( w14518 & w14520 ) ;
  assign w14522 = ( w10114 & ~w14519 ) | ( w10114 & w14521 ) | ( ~w14519 & w14521 ) ;
  assign w14523 = \pi14 ^ w14522 ;
  assign w14524 = w14220 ^ w14469 ;
  assign w14525 = w14222 ^ w14524 ;
  assign w14526 = ~w6549 & w9842 ;
  assign w14527 = w6048 & ~w9955 ;
  assign w14528 = ( w9842 & ~w14526 ) | ( w9842 & w14527 ) | ( ~w14526 & w14527 ) ;
  assign w14529 = ~w6637 & w9953 ;
  assign w14530 = w10965 | w14528 ;
  assign w14531 = ( w6045 & w14528 ) | ( w6045 & w14530 ) | ( w14528 & w14530 ) ;
  assign w14532 = ( w9953 & ~w14529 ) | ( w9953 & w14531 ) | ( ~w14529 & w14531 ) ;
  assign w14533 = \pi14 ^ w14532 ;
  assign w14534 = w14230 ^ w14468 ;
  assign w14535 = w14232 ^ w14534 ;
  assign w14536 = w6549 | w9955 ;
  assign w14537 = w6048 & w9957 ;
  assign w14538 = ( ~w9955 & w14536 ) | ( ~w9955 & w14537 ) | ( w14536 & w14537 ) ;
  assign w14539 = ~w6637 & w9842 ;
  assign w14540 = w10976 & ~w14538 ;
  assign w14541 = ( w6045 & w14538 ) | ( w6045 & ~w14540 ) | ( w14538 & ~w14540 ) ;
  assign w14542 = ( w9842 & ~w14539 ) | ( w9842 & w14541 ) | ( ~w14539 & w14541 ) ;
  assign w14543 = \pi14 ^ w14542 ;
  assign w14544 = w14240 ^ w14467 ;
  assign w14545 = w14242 ^ w14544 ;
  assign w14546 = w6048 & ~w9963 ;
  assign w14547 = ( w6637 & ~w9955 ) | ( w6637 & w14546 ) | ( ~w9955 & w14546 ) ;
  assign w14548 = w6549 | w14547 ;
  assign w14549 = ( w9957 & w14547 ) | ( w9957 & w14548 ) | ( w14547 & w14548 ) ;
  assign w14550 = w14546 | w14549 ;
  assign w14551 = w6045 | w11202 ;
  assign w14552 = ( ~w11202 & w14550 ) | ( ~w11202 & w14551 ) | ( w14550 & w14551 ) ;
  assign w14553 = \pi14 ^ w14552 ;
  assign w14554 = w14250 ^ w14466 ;
  assign w14555 = w14252 ^ w14554 ;
  assign w14556 = w6048 & w9961 ;
  assign w14557 = ( w6637 & w9957 ) | ( w6637 & w14556 ) | ( w9957 & w14556 ) ;
  assign w14558 = w6549 | w14557 ;
  assign w14559 = ( ~w9963 & w14557 ) | ( ~w9963 & w14558 ) | ( w14557 & w14558 ) ;
  assign w14560 = w14556 | w14559 ;
  assign w14561 = w6045 | w11089 ;
  assign w14562 = ( ~w11089 & w14560 ) | ( ~w11089 & w14561 ) | ( w14560 & w14561 ) ;
  assign w14563 = \pi14 ^ w14562 ;
  assign w14564 = w14260 ^ w14465 ;
  assign w14565 = w14262 ^ w14564 ;
  assign w14566 = w6048 & w9965 ;
  assign w14567 = ( w6637 & ~w9963 ) | ( w6637 & w14566 ) | ( ~w9963 & w14566 ) ;
  assign w14568 = w6549 | w14567 ;
  assign w14569 = ( w9961 & w14567 ) | ( w9961 & w14568 ) | ( w14567 & w14568 ) ;
  assign w14570 = w14566 | w14569 ;
  assign w14571 = w6045 | w11278 ;
  assign w14572 = ( ~w11278 & w14570 ) | ( ~w11278 & w14571 ) | ( w14570 & w14571 ) ;
  assign w14573 = \pi14 ^ w14572 ;
  assign w14574 = w14270 ^ w14464 ;
  assign w14575 = w14272 ^ w14574 ;
  assign w14576 = w6048 & ~w9967 ;
  assign w14577 = ( w6637 & w9961 ) | ( w6637 & w14576 ) | ( w9961 & w14576 ) ;
  assign w14578 = w6549 | w14577 ;
  assign w14579 = ( w9965 & w14577 ) | ( w9965 & w14578 ) | ( w14577 & w14578 ) ;
  assign w14580 = w14576 | w14579 ;
  assign w14581 = ~w6045 & w11339 ;
  assign w14582 = ( w11339 & w14580 ) | ( w11339 & ~w14581 ) | ( w14580 & ~w14581 ) ;
  assign w14583 = \pi14 ^ w14582 ;
  assign w14584 = w14280 ^ w14463 ;
  assign w14585 = w14282 ^ w14584 ;
  assign w14586 = w6048 & w9971 ;
  assign w14587 = ( w6637 & w9965 ) | ( w6637 & w14586 ) | ( w9965 & w14586 ) ;
  assign w14588 = w6549 | w14587 ;
  assign w14589 = ( ~w9967 & w14587 ) | ( ~w9967 & w14588 ) | ( w14587 & w14588 ) ;
  assign w14590 = w14586 | w14589 ;
  assign w14591 = w6045 | w11501 ;
  assign w14592 = ( ~w11501 & w14590 ) | ( ~w11501 & w14591 ) | ( w14590 & w14591 ) ;
  assign w14593 = \pi14 ^ w14592 ;
  assign w14594 = w14290 ^ w14462 ;
  assign w14595 = w14292 ^ w14594 ;
  assign w14596 = w6048 & ~w9973 ;
  assign w14597 = ( w6637 & ~w9967 ) | ( w6637 & w14596 ) | ( ~w9967 & w14596 ) ;
  assign w14598 = w6549 | w14597 ;
  assign w14599 = ( w9971 & w14597 ) | ( w9971 & w14598 ) | ( w14597 & w14598 ) ;
  assign w14600 = w14596 | w14599 ;
  assign w14601 = w6045 | w11512 ;
  assign w14602 = ( ~w11512 & w14600 ) | ( ~w11512 & w14601 ) | ( w14600 & w14601 ) ;
  assign w14603 = \pi14 ^ w14602 ;
  assign w14604 = w14300 ^ w14461 ;
  assign w14605 = w14302 ^ w14604 ;
  assign w14606 = w6048 & w9975 ;
  assign w14607 = ( w6637 & w9971 ) | ( w6637 & w14606 ) | ( w9971 & w14606 ) ;
  assign w14608 = w6549 | w14607 ;
  assign w14609 = ( ~w9973 & w14607 ) | ( ~w9973 & w14608 ) | ( w14607 & w14608 ) ;
  assign w14610 = w14606 | w14609 ;
  assign w14611 = w6045 | w11809 ;
  assign w14612 = ( ~w11809 & w14610 ) | ( ~w11809 & w14611 ) | ( w14610 & w14611 ) ;
  assign w14613 = \pi14 ^ w14612 ;
  assign w14614 = ~w6549 & w9975 ;
  assign w14615 = w6048 & w9977 ;
  assign w14616 = ( w9975 & ~w14614 ) | ( w9975 & w14615 ) | ( ~w14614 & w14615 ) ;
  assign w14617 = w6637 | w9973 ;
  assign w14618 = w11671 & ~w14616 ;
  assign w14619 = ( w6045 & w14616 ) | ( w6045 & ~w14618 ) | ( w14616 & ~w14618 ) ;
  assign w14620 = ( ~w9973 & w14617 ) | ( ~w9973 & w14619 ) | ( w14617 & w14619 ) ;
  assign w14621 = \pi14 ^ w14620 ;
  assign w14622 = w14312 ^ w14460 ;
  assign w14623 = w14304 ^ w14622 ;
  assign w14624 = ~w6549 & w9977 ;
  assign w14625 = w6048 & w9979 ;
  assign w14626 = ( w9977 & ~w14624 ) | ( w9977 & w14625 ) | ( ~w14624 & w14625 ) ;
  assign w14627 = ~w6637 & w9975 ;
  assign w14628 = w11914 | w14626 ;
  assign w14629 = ( w6045 & w14626 ) | ( w6045 & w14628 ) | ( w14626 & w14628 ) ;
  assign w14630 = ( w9975 & ~w14627 ) | ( w9975 & w14629 ) | ( ~w14627 & w14629 ) ;
  assign w14631 = \pi14 ^ w14630 ;
  assign w14632 = w14322 ^ w14459 ;
  assign w14633 = w14314 ^ w14632 ;
  assign w14634 = w14330 ^ w14458 ;
  assign w14635 = w14332 ^ w14634 ;
  assign w14636 = w6048 & w9981 ;
  assign w14637 = ( w6637 & w9977 ) | ( w6637 & w14636 ) | ( w9977 & w14636 ) ;
  assign w14638 = w6549 | w14637 ;
  assign w14639 = ( w9979 & w14637 ) | ( w9979 & w14638 ) | ( w14637 & w14638 ) ;
  assign w14640 = w14636 | w14639 ;
  assign w14641 = ~w6045 & w12106 ;
  assign w14642 = ( w12106 & w14640 ) | ( w12106 & ~w14641 ) | ( w14640 & ~w14641 ) ;
  assign w14643 = \pi14 ^ w14642 ;
  assign w14644 = w14340 ^ w14457 ;
  assign w14645 = w14342 ^ w14644 ;
  assign w14646 = w6048 & w9983 ;
  assign w14647 = ( w6637 & w9979 ) | ( w6637 & w14646 ) | ( w9979 & w14646 ) ;
  assign w14648 = w6549 | w14647 ;
  assign w14649 = ( w9981 & w14647 ) | ( w9981 & w14648 ) | ( w14647 & w14648 ) ;
  assign w14650 = w14646 | w14649 ;
  assign w14651 = ~w6045 & w12010 ;
  assign w14652 = ( w12010 & w14650 ) | ( w12010 & ~w14651 ) | ( w14650 & ~w14651 ) ;
  assign w14653 = \pi14 ^ w14652 ;
  assign w14654 = w14350 ^ w14456 ;
  assign w14655 = w14352 ^ w14654 ;
  assign w14656 = w6048 & w9985 ;
  assign w14657 = ( w6637 & w9981 ) | ( w6637 & w14656 ) | ( w9981 & w14656 ) ;
  assign w14658 = w6549 | w14657 ;
  assign w14659 = ( w9983 & w14657 ) | ( w9983 & w14658 ) | ( w14657 & w14658 ) ;
  assign w14660 = w14656 | w14659 ;
  assign w14661 = ~w6045 & w12236 ;
  assign w14662 = ( w12236 & w14660 ) | ( w12236 & ~w14661 ) | ( w14660 & ~w14661 ) ;
  assign w14663 = \pi14 ^ w14662 ;
  assign w14664 = ~w6549 & w9985 ;
  assign w14665 = w6048 & w9987 ;
  assign w14666 = ( w9985 & ~w14664 ) | ( w9985 & w14665 ) | ( ~w14664 & w14665 ) ;
  assign w14667 = ~w6637 & w9983 ;
  assign w14668 = w12433 | w14666 ;
  assign w14669 = ( w6045 & w14666 ) | ( w6045 & w14668 ) | ( w14666 & w14668 ) ;
  assign w14670 = ( w9983 & ~w14667 ) | ( w9983 & w14669 ) | ( ~w14667 & w14669 ) ;
  assign w14671 = \pi14 ^ w14670 ;
  assign w14672 = w14362 ^ w14455 ;
  assign w14673 = w14354 ^ w14672 ;
  assign w14674 = ~w6549 & w9987 ;
  assign w14675 = w6048 & ~w9989 ;
  assign w14676 = ( w9987 & ~w14674 ) | ( w9987 & w14675 ) | ( ~w14674 & w14675 ) ;
  assign w14677 = ~w6637 & w9985 ;
  assign w14678 = w12446 | w14676 ;
  assign w14679 = ( w6045 & w14676 ) | ( w6045 & w14678 ) | ( w14676 & w14678 ) ;
  assign w14680 = ( w9985 & ~w14677 ) | ( w9985 & w14679 ) | ( ~w14677 & w14679 ) ;
  assign w14681 = \pi14 ^ w14680 ;
  assign w14682 = w14372 ^ w14454 ;
  assign w14683 = w14364 ^ w14682 ;
  assign w14684 = w6549 | w9989 ;
  assign w14685 = w6048 & w9991 ;
  assign w14686 = ( ~w9989 & w14684 ) | ( ~w9989 & w14685 ) | ( w14684 & w14685 ) ;
  assign w14687 = ~w6637 & w9987 ;
  assign w14688 = w12217 & ~w14686 ;
  assign w14689 = ( w6045 & w14686 ) | ( w6045 & ~w14688 ) | ( w14686 & ~w14688 ) ;
  assign w14690 = ( w9987 & ~w14687 ) | ( w9987 & w14689 ) | ( ~w14687 & w14689 ) ;
  assign w14691 = \pi14 ^ w14690 ;
  assign w14692 = w14382 ^ w14453 ;
  assign w14693 = w14374 ^ w14692 ;
  assign w14694 = w14390 ^ w14452 ;
  assign w14695 = w14392 ^ w14694 ;
  assign w14696 = w6048 & ~w9993 ;
  assign w14697 = ( w6637 & ~w9989 ) | ( w6637 & w14696 ) | ( ~w9989 & w14696 ) ;
  assign w14698 = w6549 | w14697 ;
  assign w14699 = ( w9991 & w14697 ) | ( w9991 & w14698 ) | ( w14697 & w14698 ) ;
  assign w14700 = w14696 | w14699 ;
  assign w14701 = w6045 | w12484 ;
  assign w14702 = ( ~w12484 & w14700 ) | ( ~w12484 & w14701 ) | ( w14700 & w14701 ) ;
  assign w14703 = \pi14 ^ w14702 ;
  assign w14704 = w14402 ^ w14451 ;
  assign w14705 = w14394 ^ w14704 ;
  assign w14706 = w6048 & w9995 ;
  assign w14707 = ( w6637 & w9991 ) | ( w6637 & w14706 ) | ( w9991 & w14706 ) ;
  assign w14708 = w6549 | w14707 ;
  assign w14709 = ( ~w9993 & w14707 ) | ( ~w9993 & w14708 ) | ( w14707 & w14708 ) ;
  assign w14710 = w14706 | w14709 ;
  assign w14711 = w6045 | w12514 ;
  assign w14712 = ( ~w12514 & w14710 ) | ( ~w12514 & w14711 ) | ( w14710 & w14711 ) ;
  assign w14713 = \pi14 ^ w14712 ;
  assign w14714 = w14410 ^ w14450 ;
  assign w14715 = w14411 ^ w14714 ;
  assign w14716 = w6048 & w9997 ;
  assign w14717 = ( w6637 & ~w9993 ) | ( w6637 & w14716 ) | ( ~w9993 & w14716 ) ;
  assign w14718 = w6549 | w14717 ;
  assign w14719 = ( w9995 & w14717 ) | ( w9995 & w14718 ) | ( w14717 & w14718 ) ;
  assign w14720 = w14716 | w14719 ;
  assign w14721 = w6045 | w12541 ;
  assign w14722 = ( ~w12541 & w14720 ) | ( ~w12541 & w14721 ) | ( w14720 & w14721 ) ;
  assign w14723 = \pi14 ^ w14722 ;
  assign w14724 = ~w6549 & w9997 ;
  assign w14725 = w6048 & w9999 ;
  assign w14726 = ( w9997 & ~w14724 ) | ( w9997 & w14725 ) | ( ~w14724 & w14725 ) ;
  assign w14727 = ~w6637 & w9995 ;
  assign w14728 = w12572 | w14726 ;
  assign w14729 = ( w6045 & w14726 ) | ( w6045 & w14728 ) | ( w14726 & w14728 ) ;
  assign w14730 = ( w9995 & ~w14727 ) | ( w9995 & w14729 ) | ( ~w14727 & w14729 ) ;
  assign w14731 = \pi14 ^ w14730 ;
  assign w14732 = w14424 ^ w14449 ;
  assign w14733 = w14416 ^ w14732 ;
  assign w14734 = w14439 ^ w14447 ;
  assign w14735 = w14448 ^ w14734 ;
  assign w14736 = w6048 & w10001 ;
  assign w14737 = ( w6637 & w9997 ) | ( w6637 & w14736 ) | ( w9997 & w14736 ) ;
  assign w14738 = w6549 | w14737 ;
  assign w14739 = ( w9999 & w14737 ) | ( w9999 & w14738 ) | ( w14737 & w14738 ) ;
  assign w14740 = w14736 | w14739 ;
  assign w14741 = ~w6045 & w12641 ;
  assign w14742 = ( w12641 & w14740 ) | ( w12641 & ~w14741 ) | ( w14740 & ~w14741 ) ;
  assign w14743 = \pi14 ^ w14742 ;
  assign w14744 = ~w6549 & w10001 ;
  assign w14745 = w6048 & ~w10006 ;
  assign w14746 = ( w10001 & ~w14744 ) | ( w10001 & w14745 ) | ( ~w14744 & w14745 ) ;
  assign w14747 = ~w6637 & w9999 ;
  assign w14748 = w12691 & ~w14746 ;
  assign w14749 = ( w6045 & w14746 ) | ( w6045 & ~w14748 ) | ( w14746 & ~w14748 ) ;
  assign w14750 = ( w9999 & ~w14747 ) | ( w9999 & w14749 ) | ( ~w14747 & w14749 ) ;
  assign w14751 = \pi14 ^ w14750 ;
  assign w14752 = w14430 ^ w14438 ;
  assign w14753 = ( \pi14 & \pi15 ) | ( \pi14 & ~w10016 ) | ( \pi15 & ~w10016 ) ;
  assign w14754 = ( \pi14 & \pi15 ) | ( \pi14 & ~w10021 ) | ( \pi15 & ~w10021 ) ;
  assign w14755 = \pi16 ^ w10021 ;
  assign w14756 = ( \pi16 & w14754 ) | ( \pi16 & w14755 ) | ( w14754 & w14755 ) ;
  assign w14757 = w14753 ^ w14756 ;
  assign w14758 = w6048 & w10011 ;
  assign w14759 = ( w6637 & w10001 ) | ( w6637 & w14758 ) | ( w10001 & w14758 ) ;
  assign w14760 = w6549 | w14759 ;
  assign w14761 = ( ~w10006 & w14759 ) | ( ~w10006 & w14760 ) | ( w14759 & w14760 ) ;
  assign w14762 = w14758 | w14761 ;
  assign w14763 = ~w6045 & w12747 ;
  assign w14764 = ( w12747 & w14762 ) | ( w12747 & ~w14763 ) | ( w14762 & ~w14763 ) ;
  assign w14765 = \pi14 ^ w14764 ;
  assign w14766 = \pi14 & w10021 ;
  assign w14767 = w10016 & w14766 ;
  assign w14768 = ( \pi11 & \pi12 ) | ( \pi11 & ~w14767 ) | ( \pi12 & ~w14767 ) ;
  assign w14769 = ( \pi13 & \pi14 ) | ( \pi13 & ~w14768 ) | ( \pi14 & ~w14768 ) ;
  assign w14770 = ( \pi13 & ~w14766 ) | ( \pi13 & w14768 ) | ( ~w14766 & w14768 ) ;
  assign w14771 = ( w8192 & w14769 ) | ( w8192 & ~w14770 ) | ( w14769 & ~w14770 ) ;
  assign w14772 = w6048 & ~w10021 ;
  assign w14773 = ( w6637 & w10011 ) | ( w6637 & w14772 ) | ( w10011 & w14772 ) ;
  assign w14774 = w6549 | w14773 ;
  assign w14775 = ( ~w10016 & w14773 ) | ( ~w10016 & w14774 ) | ( w14773 & w14774 ) ;
  assign w14776 = w14772 | w14775 ;
  assign w14777 = ~w6045 & w12867 ;
  assign w14778 = ( w12867 & w14776 ) | ( w12867 & ~w14777 ) | ( w14776 & ~w14777 ) ;
  assign w14779 = \pi14 ^ w14778 ;
  assign w14780 = w14771 & w14779 ;
  assign w14781 = ~w6549 & w10011 ;
  assign w14782 = w6048 & ~w10016 ;
  assign w14783 = ( w10011 & ~w14781 ) | ( w10011 & w14782 ) | ( ~w14781 & w14782 ) ;
  assign w14784 = w6637 | w10006 ;
  assign w14785 = w12777 | w14783 ;
  assign w14786 = ( w6045 & w14783 ) | ( w6045 & w14785 ) | ( w14783 & w14785 ) ;
  assign w14787 = ( ~w10006 & w14784 ) | ( ~w10006 & w14786 ) | ( w14784 & w14786 ) ;
  assign w14788 = \pi14 ^ w14787 ;
  assign w14789 = w5496 & ~w10021 ;
  assign w14790 = ( w14780 & w14788 ) | ( w14780 & w14789 ) | ( w14788 & w14789 ) ;
  assign w14791 = ( w14757 & w14765 ) | ( w14757 & w14790 ) | ( w14765 & w14790 ) ;
  assign w14792 = ( w14751 & w14752 ) | ( w14751 & w14791 ) | ( w14752 & w14791 ) ;
  assign w14793 = ( w14735 & w14743 ) | ( w14735 & w14792 ) | ( w14743 & w14792 ) ;
  assign w14794 = ( w14731 & w14733 ) | ( w14731 & w14793 ) | ( w14733 & w14793 ) ;
  assign w14795 = ( w14715 & w14723 ) | ( w14715 & w14794 ) | ( w14723 & w14794 ) ;
  assign w14796 = ( w14705 & w14713 ) | ( w14705 & w14795 ) | ( w14713 & w14795 ) ;
  assign w14797 = ( w14695 & w14703 ) | ( w14695 & w14796 ) | ( w14703 & w14796 ) ;
  assign w14798 = ( w14691 & w14693 ) | ( w14691 & w14797 ) | ( w14693 & w14797 ) ;
  assign w14799 = ( w14681 & w14683 ) | ( w14681 & w14798 ) | ( w14683 & w14798 ) ;
  assign w14800 = ( w14671 & w14673 ) | ( w14671 & w14799 ) | ( w14673 & w14799 ) ;
  assign w14801 = ( w14655 & w14663 ) | ( w14655 & w14800 ) | ( w14663 & w14800 ) ;
  assign w14802 = ( w14645 & w14653 ) | ( w14645 & w14801 ) | ( w14653 & w14801 ) ;
  assign w14803 = ( w14635 & w14643 ) | ( w14635 & w14802 ) | ( w14643 & w14802 ) ;
  assign w14804 = ( w14631 & w14633 ) | ( w14631 & w14803 ) | ( w14633 & w14803 ) ;
  assign w14805 = ( w14621 & w14623 ) | ( w14621 & w14804 ) | ( w14623 & w14804 ) ;
  assign w14806 = ( ~w14605 & w14613 ) | ( ~w14605 & w14805 ) | ( w14613 & w14805 ) ;
  assign w14807 = ( ~w14595 & w14603 ) | ( ~w14595 & w14806 ) | ( w14603 & w14806 ) ;
  assign w14808 = ( w14585 & w14593 ) | ( w14585 & w14807 ) | ( w14593 & w14807 ) ;
  assign w14809 = ( ~w14575 & w14583 ) | ( ~w14575 & w14808 ) | ( w14583 & w14808 ) ;
  assign w14810 = ( ~w14565 & w14573 ) | ( ~w14565 & w14809 ) | ( w14573 & w14809 ) ;
  assign w14811 = ( w14555 & w14563 ) | ( w14555 & w14810 ) | ( w14563 & w14810 ) ;
  assign w14812 = ( w14545 & w14553 ) | ( w14545 & w14811 ) | ( w14553 & w14811 ) ;
  assign w14813 = ( w14535 & w14543 ) | ( w14535 & w14812 ) | ( w14543 & w14812 ) ;
  assign w14814 = ( w14525 & w14533 ) | ( w14525 & w14813 ) | ( w14533 & w14813 ) ;
  assign w14815 = ( w14515 & w14523 ) | ( w14515 & w14814 ) | ( w14523 & w14814 ) ;
  assign w14816 = w6949 | w10805 ;
  assign w14817 = w6748 & w10784 ;
  assign w14818 = ( ~w10805 & w14816 ) | ( ~w10805 & w14817 ) | ( w14816 & w14817 ) ;
  assign w14819 = w7154 | w10807 ;
  assign w14820 = w11117 | w14818 ;
  assign w14821 = ( w6751 & w14818 ) | ( w6751 & w14820 ) | ( w14818 & w14820 ) ;
  assign w14822 = ( ~w10807 & w14819 ) | ( ~w10807 & w14821 ) | ( w14819 & w14821 ) ;
  assign w14823 = \pi11 ^ w14822 ;
  assign w14824 = ( ~w14513 & w14815 ) | ( ~w14513 & w14823 ) | ( w14815 & w14823 ) ;
  assign w14825 = w7673 | w10885 ;
  assign w14826 = w7411 & ~w10866 ;
  assign w14827 = ( ~w10885 & w14825 ) | ( ~w10885 & w14826 ) | ( w14825 & w14826 ) ;
  assign w14828 = w7944 | w10887 ;
  assign w14829 = w11131 & ~w14827 ;
  assign w14830 = ( w7414 & w14827 ) | ( w7414 & ~w14829 ) | ( w14827 & ~w14829 ) ;
  assign w14831 = ( ~w10887 & w14828 ) | ( ~w10887 & w14830 ) | ( w14828 & w14830 ) ;
  assign w14832 = \pi08 ^ w14831 ;
  assign w14833 = ( w14511 & w14824 ) | ( w14511 & w14832 ) | ( w14824 & w14832 ) ;
  assign w14834 = ( w35 & w8262 ) | ( w35 & ~w11138 ) | ( w8262 & ~w11138 ) ;
  assign w14835 = w35 & ~w14834 ;
  assign w14836 = ( w8593 & ~w14834 ) | ( w8593 & w14835 ) | ( ~w14834 & w14835 ) ;
  assign w14837 = ( ~w10738 & w14834 ) | ( ~w10738 & w14836 ) | ( w14834 & w14836 ) ;
  assign w14838 = w14198 ^ w14489 ;
  assign w14839 = w14497 ^ w14838 ;
  assign w14840 = w11146 & ~w14837 ;
  assign w14841 = ( w8263 & w14837 ) | ( w8263 & ~w14840 ) | ( w14837 & ~w14840 ) ;
  assign w14842 = \pi05 ^ w14841 ;
  assign w14843 = ( w14833 & ~w14839 ) | ( w14833 & w14842 ) | ( ~w14839 & w14842 ) ;
  assign w14844 = w14498 ^ w14508 ;
  assign w14845 = w14506 ^ w14844 ;
  assign w14846 = w8263 & w11146 ;
  assign w14847 = ( w8263 & w14837 ) | ( w8263 & ~w14846 ) | ( w14837 & ~w14846 ) ;
  assign w14848 = w14839 ^ w14847 ;
  assign w14849 = \pi05 ^ w14833 ;
  assign w14850 = w14848 ^ w14849 ;
  assign w14851 = w14511 ^ w14824 ;
  assign w14852 = w14832 ^ w14851 ;
  assign w14853 = w14513 ^ w14823 ;
  assign w14854 = w14815 ^ w14853 ;
  assign w14855 = ~w6949 & w10784 ;
  assign w14856 = w6748 & w10211 ;
  assign w14857 = ( w10784 & ~w14855 ) | ( w10784 & w14856 ) | ( ~w14855 & w14856 ) ;
  assign w14858 = w7154 | w10805 ;
  assign w14859 = w10855 & ~w14857 ;
  assign w14860 = ( w6751 & w14857 ) | ( w6751 & ~w14859 ) | ( w14857 & ~w14859 ) ;
  assign w14861 = ( ~w10805 & w14858 ) | ( ~w10805 & w14860 ) | ( w14858 & w14860 ) ;
  assign w14862 = \pi11 ^ w14861 ;
  assign w14863 = w14523 ^ w14814 ;
  assign w14864 = w14515 ^ w14863 ;
  assign w14865 = ~w6949 & w10211 ;
  assign w14866 = w6748 & w10114 ;
  assign w14867 = ( w10211 & ~w14865 ) | ( w10211 & w14866 ) | ( ~w14865 & w14866 ) ;
  assign w14868 = ~w7154 & w10784 ;
  assign w14869 = w10789 | w14867 ;
  assign w14870 = ( w6751 & w14867 ) | ( w6751 & w14869 ) | ( w14867 & w14869 ) ;
  assign w14871 = ( w10784 & ~w14868 ) | ( w10784 & w14870 ) | ( ~w14868 & w14870 ) ;
  assign w14872 = \pi11 ^ w14871 ;
  assign w14873 = w14533 ^ w14813 ;
  assign w14874 = w14525 ^ w14873 ;
  assign w14875 = ~w6949 & w10114 ;
  assign w14876 = w6748 & w9953 ;
  assign w14877 = ( w10114 & ~w14875 ) | ( w10114 & w14876 ) | ( ~w14875 & w14876 ) ;
  assign w14878 = ~w7154 & w10211 ;
  assign w14879 = w10214 | w14877 ;
  assign w14880 = ( w6751 & w14877 ) | ( w6751 & w14879 ) | ( w14877 & w14879 ) ;
  assign w14881 = ( w10211 & ~w14878 ) | ( w10211 & w14880 ) | ( ~w14878 & w14880 ) ;
  assign w14882 = \pi11 ^ w14881 ;
  assign w14883 = w14543 ^ w14812 ;
  assign w14884 = w14535 ^ w14883 ;
  assign w14885 = ~w6949 & w9953 ;
  assign w14886 = w6748 & w9842 ;
  assign w14887 = ( w9953 & ~w14885 ) | ( w9953 & w14886 ) | ( ~w14885 & w14886 ) ;
  assign w14888 = ~w7154 & w10114 ;
  assign w14889 = w10334 | w14887 ;
  assign w14890 = ( w6751 & w14887 ) | ( w6751 & w14889 ) | ( w14887 & w14889 ) ;
  assign w14891 = ( w10114 & ~w14888 ) | ( w10114 & w14890 ) | ( ~w14888 & w14890 ) ;
  assign w14892 = \pi11 ^ w14891 ;
  assign w14893 = w14553 ^ w14811 ;
  assign w14894 = w14545 ^ w14893 ;
  assign w14895 = ~w6949 & w9842 ;
  assign w14896 = w6748 & ~w9955 ;
  assign w14897 = ( w9842 & ~w14895 ) | ( w9842 & w14896 ) | ( ~w14895 & w14896 ) ;
  assign w14898 = ~w7154 & w9953 ;
  assign w14899 = w10965 | w14897 ;
  assign w14900 = ( w6751 & w14897 ) | ( w6751 & w14899 ) | ( w14897 & w14899 ) ;
  assign w14901 = ( w9953 & ~w14898 ) | ( w9953 & w14900 ) | ( ~w14898 & w14900 ) ;
  assign w14902 = \pi11 ^ w14901 ;
  assign w14903 = w14563 ^ w14810 ;
  assign w14904 = w14555 ^ w14903 ;
  assign w14905 = w6949 | w9955 ;
  assign w14906 = w6748 & w9957 ;
  assign w14907 = ( ~w9955 & w14905 ) | ( ~w9955 & w14906 ) | ( w14905 & w14906 ) ;
  assign w14908 = ~w7154 & w9842 ;
  assign w14909 = w10976 & ~w14907 ;
  assign w14910 = ( w6751 & w14907 ) | ( w6751 & ~w14909 ) | ( w14907 & ~w14909 ) ;
  assign w14911 = ( w9842 & ~w14908 ) | ( w9842 & w14910 ) | ( ~w14908 & w14910 ) ;
  assign w14912 = \pi11 ^ w14911 ;
  assign w14913 = w14573 ^ w14809 ;
  assign w14914 = w14565 ^ w14913 ;
  assign w14915 = ~w6949 & w9957 ;
  assign w14916 = w6748 & ~w9963 ;
  assign w14917 = ( w9957 & ~w14915 ) | ( w9957 & w14916 ) | ( ~w14915 & w14916 ) ;
  assign w14918 = w7154 | w9955 ;
  assign w14919 = w11202 & ~w14917 ;
  assign w14920 = ( w6751 & w14917 ) | ( w6751 & ~w14919 ) | ( w14917 & ~w14919 ) ;
  assign w14921 = ( ~w9955 & w14918 ) | ( ~w9955 & w14920 ) | ( w14918 & w14920 ) ;
  assign w14922 = \pi11 ^ w14921 ;
  assign w14923 = w14583 ^ w14808 ;
  assign w14924 = w14575 ^ w14923 ;
  assign w14925 = w6949 | w9963 ;
  assign w14926 = w6748 & w9961 ;
  assign w14927 = ( ~w9963 & w14925 ) | ( ~w9963 & w14926 ) | ( w14925 & w14926 ) ;
  assign w14928 = ~w7154 & w9957 ;
  assign w14929 = w11089 & ~w14927 ;
  assign w14930 = ( w6751 & w14927 ) | ( w6751 & ~w14929 ) | ( w14927 & ~w14929 ) ;
  assign w14931 = ( w9957 & ~w14928 ) | ( w9957 & w14930 ) | ( ~w14928 & w14930 ) ;
  assign w14932 = \pi11 ^ w14931 ;
  assign w14933 = w14593 ^ w14807 ;
  assign w14934 = w14585 ^ w14933 ;
  assign w14935 = ~w6949 & w9961 ;
  assign w14936 = w6748 & w9965 ;
  assign w14937 = ( w9961 & ~w14935 ) | ( w9961 & w14936 ) | ( ~w14935 & w14936 ) ;
  assign w14938 = w7154 | w9963 ;
  assign w14939 = w11278 & ~w14937 ;
  assign w14940 = ( w6751 & w14937 ) | ( w6751 & ~w14939 ) | ( w14937 & ~w14939 ) ;
  assign w14941 = ( ~w9963 & w14938 ) | ( ~w9963 & w14940 ) | ( w14938 & w14940 ) ;
  assign w14942 = \pi11 ^ w14941 ;
  assign w14943 = w14603 ^ w14806 ;
  assign w14944 = w14595 ^ w14943 ;
  assign w14945 = ~w6949 & w9965 ;
  assign w14946 = w6748 & ~w9967 ;
  assign w14947 = ( w9965 & ~w14945 ) | ( w9965 & w14946 ) | ( ~w14945 & w14946 ) ;
  assign w14948 = ~w7154 & w9961 ;
  assign w14949 = w11339 | w14947 ;
  assign w14950 = ( w6751 & w14947 ) | ( w6751 & w14949 ) | ( w14947 & w14949 ) ;
  assign w14951 = ( w9961 & ~w14948 ) | ( w9961 & w14950 ) | ( ~w14948 & w14950 ) ;
  assign w14952 = \pi11 ^ w14951 ;
  assign w14953 = w14613 ^ w14805 ;
  assign w14954 = w14605 ^ w14953 ;
  assign w14955 = w14621 ^ w14804 ;
  assign w14956 = w14623 ^ w14955 ;
  assign w14957 = w6748 & w9971 ;
  assign w14958 = ( w7154 & w9965 ) | ( w7154 & w14957 ) | ( w9965 & w14957 ) ;
  assign w14959 = w6949 | w14958 ;
  assign w14960 = ( ~w9967 & w14958 ) | ( ~w9967 & w14959 ) | ( w14958 & w14959 ) ;
  assign w14961 = w14957 | w14960 ;
  assign w14962 = w6751 | w11501 ;
  assign w14963 = ( ~w11501 & w14961 ) | ( ~w11501 & w14962 ) | ( w14961 & w14962 ) ;
  assign w14964 = \pi11 ^ w14963 ;
  assign w14965 = w14631 ^ w14803 ;
  assign w14966 = w14633 ^ w14965 ;
  assign w14967 = w6748 & ~w9973 ;
  assign w14968 = ( w7154 & ~w9967 ) | ( w7154 & w14967 ) | ( ~w9967 & w14967 ) ;
  assign w14969 = w6949 | w14968 ;
  assign w14970 = ( w9971 & w14968 ) | ( w9971 & w14969 ) | ( w14968 & w14969 ) ;
  assign w14971 = w14967 | w14970 ;
  assign w14972 = w6751 | w11512 ;
  assign w14973 = ( ~w11512 & w14971 ) | ( ~w11512 & w14972 ) | ( w14971 & w14972 ) ;
  assign w14974 = \pi11 ^ w14973 ;
  assign w14975 = w6949 | w9973 ;
  assign w14976 = w6748 & w9975 ;
  assign w14977 = ( ~w9973 & w14975 ) | ( ~w9973 & w14976 ) | ( w14975 & w14976 ) ;
  assign w14978 = ~w7154 & w9971 ;
  assign w14979 = w11809 & ~w14977 ;
  assign w14980 = ( w6751 & w14977 ) | ( w6751 & ~w14979 ) | ( w14977 & ~w14979 ) ;
  assign w14981 = ( w9971 & ~w14978 ) | ( w9971 & w14980 ) | ( ~w14978 & w14980 ) ;
  assign w14982 = \pi11 ^ w14981 ;
  assign w14983 = w14643 ^ w14802 ;
  assign w14984 = w14635 ^ w14983 ;
  assign w14985 = ~w6949 & w9975 ;
  assign w14986 = w6748 & w9977 ;
  assign w14987 = ( w9975 & ~w14985 ) | ( w9975 & w14986 ) | ( ~w14985 & w14986 ) ;
  assign w14988 = w7154 | w9973 ;
  assign w14989 = w11671 & ~w14987 ;
  assign w14990 = ( w6751 & w14987 ) | ( w6751 & ~w14989 ) | ( w14987 & ~w14989 ) ;
  assign w14991 = ( ~w9973 & w14988 ) | ( ~w9973 & w14990 ) | ( w14988 & w14990 ) ;
  assign w14992 = \pi11 ^ w14991 ;
  assign w14993 = w14653 ^ w14801 ;
  assign w14994 = w14645 ^ w14993 ;
  assign w14995 = ~w6949 & w9977 ;
  assign w14996 = w6748 & w9979 ;
  assign w14997 = ( w9977 & ~w14995 ) | ( w9977 & w14996 ) | ( ~w14995 & w14996 ) ;
  assign w14998 = ~w7154 & w9975 ;
  assign w14999 = w11914 | w14997 ;
  assign w15000 = ( w6751 & w14997 ) | ( w6751 & w14999 ) | ( w14997 & w14999 ) ;
  assign w15001 = ( w9975 & ~w14998 ) | ( w9975 & w15000 ) | ( ~w14998 & w15000 ) ;
  assign w15002 = \pi11 ^ w15001 ;
  assign w15003 = w14663 ^ w14800 ;
  assign w15004 = w14655 ^ w15003 ;
  assign w15005 = w14671 ^ w14799 ;
  assign w15006 = w14673 ^ w15005 ;
  assign w15007 = w6748 & w9981 ;
  assign w15008 = ( w7154 & w9977 ) | ( w7154 & w15007 ) | ( w9977 & w15007 ) ;
  assign w15009 = w6949 | w15008 ;
  assign w15010 = ( w9979 & w15008 ) | ( w9979 & w15009 ) | ( w15008 & w15009 ) ;
  assign w15011 = w15007 | w15010 ;
  assign w15012 = ~w6751 & w12106 ;
  assign w15013 = ( w12106 & w15011 ) | ( w12106 & ~w15012 ) | ( w15011 & ~w15012 ) ;
  assign w15014 = \pi11 ^ w15013 ;
  assign w15015 = w14681 ^ w14798 ;
  assign w15016 = w14683 ^ w15015 ;
  assign w15017 = w6748 & w9983 ;
  assign w15018 = ( w7154 & w9979 ) | ( w7154 & w15017 ) | ( w9979 & w15017 ) ;
  assign w15019 = w6949 | w15018 ;
  assign w15020 = ( w9981 & w15018 ) | ( w9981 & w15019 ) | ( w15018 & w15019 ) ;
  assign w15021 = w15017 | w15020 ;
  assign w15022 = ~w6751 & w12010 ;
  assign w15023 = ( w12010 & w15021 ) | ( w12010 & ~w15022 ) | ( w15021 & ~w15022 ) ;
  assign w15024 = \pi11 ^ w15023 ;
  assign w15025 = w14691 ^ w14797 ;
  assign w15026 = w14693 ^ w15025 ;
  assign w15027 = w6748 & w9985 ;
  assign w15028 = ( w7154 & w9981 ) | ( w7154 & w15027 ) | ( w9981 & w15027 ) ;
  assign w15029 = w6949 | w15028 ;
  assign w15030 = ( w9983 & w15028 ) | ( w9983 & w15029 ) | ( w15028 & w15029 ) ;
  assign w15031 = w15027 | w15030 ;
  assign w15032 = ~w6751 & w12236 ;
  assign w15033 = ( w12236 & w15031 ) | ( w12236 & ~w15032 ) | ( w15031 & ~w15032 ) ;
  assign w15034 = \pi11 ^ w15033 ;
  assign w15035 = ~w6949 & w9985 ;
  assign w15036 = w6748 & w9987 ;
  assign w15037 = ( w9985 & ~w15035 ) | ( w9985 & w15036 ) | ( ~w15035 & w15036 ) ;
  assign w15038 = ~w7154 & w9983 ;
  assign w15039 = w12433 | w15037 ;
  assign w15040 = ( w6751 & w15037 ) | ( w6751 & w15039 ) | ( w15037 & w15039 ) ;
  assign w15041 = ( w9983 & ~w15038 ) | ( w9983 & w15040 ) | ( ~w15038 & w15040 ) ;
  assign w15042 = \pi11 ^ w15041 ;
  assign w15043 = w14703 ^ w14796 ;
  assign w15044 = w14695 ^ w15043 ;
  assign w15045 = ~w6949 & w9987 ;
  assign w15046 = w6748 & ~w9989 ;
  assign w15047 = ( w9987 & ~w15045 ) | ( w9987 & w15046 ) | ( ~w15045 & w15046 ) ;
  assign w15048 = ~w7154 & w9985 ;
  assign w15049 = w12446 | w15047 ;
  assign w15050 = ( w6751 & w15047 ) | ( w6751 & w15049 ) | ( w15047 & w15049 ) ;
  assign w15051 = ( w9985 & ~w15048 ) | ( w9985 & w15050 ) | ( ~w15048 & w15050 ) ;
  assign w15052 = \pi11 ^ w15051 ;
  assign w15053 = w14713 ^ w14795 ;
  assign w15054 = w14705 ^ w15053 ;
  assign w15055 = w6949 | w9989 ;
  assign w15056 = w6748 & w9991 ;
  assign w15057 = ( ~w9989 & w15055 ) | ( ~w9989 & w15056 ) | ( w15055 & w15056 ) ;
  assign w15058 = ~w7154 & w9987 ;
  assign w15059 = w12217 & ~w15057 ;
  assign w15060 = ( w6751 & w15057 ) | ( w6751 & ~w15059 ) | ( w15057 & ~w15059 ) ;
  assign w15061 = ( w9987 & ~w15058 ) | ( w9987 & w15060 ) | ( ~w15058 & w15060 ) ;
  assign w15062 = \pi11 ^ w15061 ;
  assign w15063 = w14723 ^ w14794 ;
  assign w15064 = w14715 ^ w15063 ;
  assign w15065 = w14731 ^ w14793 ;
  assign w15066 = w14733 ^ w15065 ;
  assign w15067 = w6748 & ~w9993 ;
  assign w15068 = ( w7154 & ~w9989 ) | ( w7154 & w15067 ) | ( ~w9989 & w15067 ) ;
  assign w15069 = w6949 | w15068 ;
  assign w15070 = ( w9991 & w15068 ) | ( w9991 & w15069 ) | ( w15068 & w15069 ) ;
  assign w15071 = w15067 | w15070 ;
  assign w15072 = w6751 | w12484 ;
  assign w15073 = ( ~w12484 & w15071 ) | ( ~w12484 & w15072 ) | ( w15071 & w15072 ) ;
  assign w15074 = \pi11 ^ w15073 ;
  assign w15075 = w14743 ^ w14792 ;
  assign w15076 = w14735 ^ w15075 ;
  assign w15077 = w6748 & w9995 ;
  assign w15078 = ( w7154 & w9991 ) | ( w7154 & w15077 ) | ( w9991 & w15077 ) ;
  assign w15079 = w6949 | w15078 ;
  assign w15080 = ( ~w9993 & w15078 ) | ( ~w9993 & w15079 ) | ( w15078 & w15079 ) ;
  assign w15081 = w15077 | w15080 ;
  assign w15082 = w6751 | w12514 ;
  assign w15083 = ( ~w12514 & w15081 ) | ( ~w12514 & w15082 ) | ( w15081 & w15082 ) ;
  assign w15084 = \pi11 ^ w15083 ;
  assign w15085 = w14751 ^ w14791 ;
  assign w15086 = w14752 ^ w15085 ;
  assign w15087 = w6748 & w9997 ;
  assign w15088 = ( w7154 & ~w9993 ) | ( w7154 & w15087 ) | ( ~w9993 & w15087 ) ;
  assign w15089 = w6949 | w15088 ;
  assign w15090 = ( w9995 & w15088 ) | ( w9995 & w15089 ) | ( w15088 & w15089 ) ;
  assign w15091 = w15087 | w15090 ;
  assign w15092 = w6751 | w12541 ;
  assign w15093 = ( ~w12541 & w15091 ) | ( ~w12541 & w15092 ) | ( w15091 & w15092 ) ;
  assign w15094 = \pi11 ^ w15093 ;
  assign w15095 = ~w6949 & w9997 ;
  assign w15096 = w6748 & w9999 ;
  assign w15097 = ( w9997 & ~w15095 ) | ( w9997 & w15096 ) | ( ~w15095 & w15096 ) ;
  assign w15098 = ~w7154 & w9995 ;
  assign w15099 = w12572 | w15097 ;
  assign w15100 = ( w6751 & w15097 ) | ( w6751 & w15099 ) | ( w15097 & w15099 ) ;
  assign w15101 = ( w9995 & ~w15098 ) | ( w9995 & w15100 ) | ( ~w15098 & w15100 ) ;
  assign w15102 = \pi11 ^ w15101 ;
  assign w15103 = w14765 ^ w14790 ;
  assign w15104 = w14757 ^ w15103 ;
  assign w15105 = w14780 ^ w14788 ;
  assign w15106 = w14789 ^ w15105 ;
  assign w15107 = w6748 & w10001 ;
  assign w15108 = ( w7154 & w9997 ) | ( w7154 & w15107 ) | ( w9997 & w15107 ) ;
  assign w15109 = w6949 | w15108 ;
  assign w15110 = ( w9999 & w15108 ) | ( w9999 & w15109 ) | ( w15108 & w15109 ) ;
  assign w15111 = w15107 | w15110 ;
  assign w15112 = ~w6751 & w12641 ;
  assign w15113 = ( w12641 & w15111 ) | ( w12641 & ~w15112 ) | ( w15111 & ~w15112 ) ;
  assign w15114 = \pi11 ^ w15113 ;
  assign w15115 = ~w6949 & w10001 ;
  assign w15116 = w6748 & ~w10006 ;
  assign w15117 = ( w10001 & ~w15115 ) | ( w10001 & w15116 ) | ( ~w15115 & w15116 ) ;
  assign w15118 = ~w7154 & w9999 ;
  assign w15119 = w12691 & ~w15117 ;
  assign w15120 = ( w6751 & w15117 ) | ( w6751 & ~w15119 ) | ( w15117 & ~w15119 ) ;
  assign w15121 = ( w9999 & ~w15118 ) | ( w9999 & w15120 ) | ( ~w15118 & w15120 ) ;
  assign w15122 = \pi11 ^ w15121 ;
  assign w15123 = w14771 ^ w14779 ;
  assign w15124 = ( \pi11 & \pi12 ) | ( \pi11 & ~w10016 ) | ( \pi12 & ~w10016 ) ;
  assign w15125 = ( \pi11 & \pi12 ) | ( \pi11 & ~w10021 ) | ( \pi12 & ~w10021 ) ;
  assign w15126 = \pi13 ^ w10021 ;
  assign w15127 = ( \pi13 & w15125 ) | ( \pi13 & w15126 ) | ( w15125 & w15126 ) ;
  assign w15128 = w15124 ^ w15127 ;
  assign w15129 = w6748 & w10011 ;
  assign w15130 = ( w7154 & w10001 ) | ( w7154 & w15129 ) | ( w10001 & w15129 ) ;
  assign w15131 = w6949 | w15130 ;
  assign w15132 = ( ~w10006 & w15130 ) | ( ~w10006 & w15131 ) | ( w15130 & w15131 ) ;
  assign w15133 = w15129 | w15132 ;
  assign w15134 = ~w6751 & w12747 ;
  assign w15135 = ( w12747 & w15133 ) | ( w12747 & ~w15134 ) | ( w15133 & ~w15134 ) ;
  assign w15136 = \pi11 ^ w15135 ;
  assign w15137 = \pi11 & w10021 ;
  assign w15138 = w10016 & w15137 ;
  assign w15139 = ( \pi08 & \pi09 ) | ( \pi08 & ~w15138 ) | ( \pi09 & ~w15138 ) ;
  assign w15140 = ( \pi10 & \pi11 ) | ( \pi10 & ~w15139 ) | ( \pi11 & ~w15139 ) ;
  assign w15141 = ( \pi10 & ~w15137 ) | ( \pi10 & w15139 ) | ( ~w15137 & w15139 ) ;
  assign w15142 = ( w8530 & w15140 ) | ( w8530 & ~w15141 ) | ( w15140 & ~w15141 ) ;
  assign w15143 = w6748 & ~w10021 ;
  assign w15144 = ( w7154 & w10011 ) | ( w7154 & w15143 ) | ( w10011 & w15143 ) ;
  assign w15145 = w6949 | w15144 ;
  assign w15146 = ( ~w10016 & w15144 ) | ( ~w10016 & w15145 ) | ( w15144 & w15145 ) ;
  assign w15147 = w15143 | w15146 ;
  assign w15148 = ~w6751 & w12867 ;
  assign w15149 = ( w12867 & w15147 ) | ( w12867 & ~w15148 ) | ( w15147 & ~w15148 ) ;
  assign w15150 = \pi11 ^ w15149 ;
  assign w15151 = w15142 & w15150 ;
  assign w15152 = ~w6949 & w10011 ;
  assign w15153 = w6748 & ~w10016 ;
  assign w15154 = ( w10011 & ~w15152 ) | ( w10011 & w15153 ) | ( ~w15152 & w15153 ) ;
  assign w15155 = w7154 | w10006 ;
  assign w15156 = w12777 | w15154 ;
  assign w15157 = ( w6751 & w15154 ) | ( w6751 & w15156 ) | ( w15154 & w15156 ) ;
  assign w15158 = ( ~w10006 & w15155 ) | ( ~w10006 & w15157 ) | ( w15155 & w15157 ) ;
  assign w15159 = \pi11 ^ w15158 ;
  assign w15160 = w6044 & ~w10021 ;
  assign w15161 = ( w15151 & w15159 ) | ( w15151 & w15160 ) | ( w15159 & w15160 ) ;
  assign w15162 = ( w15128 & w15136 ) | ( w15128 & w15161 ) | ( w15136 & w15161 ) ;
  assign w15163 = ( w15122 & w15123 ) | ( w15122 & w15162 ) | ( w15123 & w15162 ) ;
  assign w15164 = ( w15106 & w15114 ) | ( w15106 & w15163 ) | ( w15114 & w15163 ) ;
  assign w15165 = ( w15102 & w15104 ) | ( w15102 & w15164 ) | ( w15104 & w15164 ) ;
  assign w15166 = ( w15086 & w15094 ) | ( w15086 & w15165 ) | ( w15094 & w15165 ) ;
  assign w15167 = ( w15076 & w15084 ) | ( w15076 & w15166 ) | ( w15084 & w15166 ) ;
  assign w15168 = ( w15066 & w15074 ) | ( w15066 & w15167 ) | ( w15074 & w15167 ) ;
  assign w15169 = ( w15062 & w15064 ) | ( w15062 & w15168 ) | ( w15064 & w15168 ) ;
  assign w15170 = ( w15052 & w15054 ) | ( w15052 & w15169 ) | ( w15054 & w15169 ) ;
  assign w15171 = ( w15042 & w15044 ) | ( w15042 & w15170 ) | ( w15044 & w15170 ) ;
  assign w15172 = ( w15026 & w15034 ) | ( w15026 & w15171 ) | ( w15034 & w15171 ) ;
  assign w15173 = ( w15016 & w15024 ) | ( w15016 & w15172 ) | ( w15024 & w15172 ) ;
  assign w15174 = ( w15006 & w15014 ) | ( w15006 & w15173 ) | ( w15014 & w15173 ) ;
  assign w15175 = ( w15002 & w15004 ) | ( w15002 & w15174 ) | ( w15004 & w15174 ) ;
  assign w15176 = ( w14992 & w14994 ) | ( w14992 & w15175 ) | ( w14994 & w15175 ) ;
  assign w15177 = ( w14982 & w14984 ) | ( w14982 & w15176 ) | ( w14984 & w15176 ) ;
  assign w15178 = ( w14966 & w14974 ) | ( w14966 & w15177 ) | ( w14974 & w15177 ) ;
  assign w15179 = ( w14956 & w14964 ) | ( w14956 & w15178 ) | ( w14964 & w15178 ) ;
  assign w15180 = ( w14952 & ~w14954 ) | ( w14952 & w15179 ) | ( ~w14954 & w15179 ) ;
  assign w15181 = ( w14942 & ~w14944 ) | ( w14942 & w15180 ) | ( ~w14944 & w15180 ) ;
  assign w15182 = ( w14932 & w14934 ) | ( w14932 & w15181 ) | ( w14934 & w15181 ) ;
  assign w15183 = ( w14922 & ~w14924 ) | ( w14922 & w15182 ) | ( ~w14924 & w15182 ) ;
  assign w15184 = ( w14912 & ~w14914 ) | ( w14912 & w15183 ) | ( ~w14914 & w15183 ) ;
  assign w15185 = ( w14902 & w14904 ) | ( w14902 & w15184 ) | ( w14904 & w15184 ) ;
  assign w15186 = ( w14892 & w14894 ) | ( w14892 & w15185 ) | ( w14894 & w15185 ) ;
  assign w15187 = ( w14882 & w14884 ) | ( w14882 & w15186 ) | ( w14884 & w15186 ) ;
  assign w15188 = ( w14872 & w14874 ) | ( w14872 & w15187 ) | ( w14874 & w15187 ) ;
  assign w15189 = ( w14862 & w14864 ) | ( w14862 & w15188 ) | ( w14864 & w15188 ) ;
  assign w15190 = w7673 | w10866 ;
  assign w15191 = w7411 & w10801 ;
  assign w15192 = ( ~w10866 & w15190 ) | ( ~w10866 & w15191 ) | ( w15190 & w15191 ) ;
  assign w15193 = w7944 | w10885 ;
  assign w15194 = w11160 & ~w15192 ;
  assign w15195 = ( w7414 & w15192 ) | ( w7414 & ~w15194 ) | ( w15192 & ~w15194 ) ;
  assign w15196 = ( ~w10885 & w15193 ) | ( ~w10885 & w15195 ) | ( w15193 & w15195 ) ;
  assign w15197 = \pi08 ^ w15196 ;
  assign w15198 = ( ~w14854 & w15189 ) | ( ~w14854 & w15197 ) | ( w15189 & w15197 ) ;
  assign w15199 = w8593 | w11139 ;
  assign w15200 = w8262 & w10883 ;
  assign w15201 = ( ~w11139 & w15199 ) | ( ~w11139 & w15200 ) | ( w15199 & w15200 ) ;
  assign w15202 = w8263 | w11145 ;
  assign w15203 = w10738 & ~w15201 ;
  assign w15204 = ( w35 & w15201 ) | ( w35 & ~w15203 ) | ( w15201 & ~w15203 ) ;
  assign w15205 = ( ~w11145 & w15202 ) | ( ~w11145 & w15204 ) | ( w15202 & w15204 ) ;
  assign w15206 = \pi05 ^ w15205 ;
  assign w15207 = ( w14852 & w15198 ) | ( w14852 & w15206 ) | ( w15198 & w15206 ) ;
  assign w15208 = w14852 ^ w15198 ;
  assign w15209 = w15206 ^ w15208 ;
  assign w15210 = w14854 ^ w15197 ;
  assign w15211 = w15189 ^ w15210 ;
  assign w15212 = w14862 ^ w15188 ;
  assign w15213 = w14864 ^ w15212 ;
  assign w15214 = ~w7673 & w10801 ;
  assign w15215 = w7411 & ~w10807 ;
  assign w15216 = ( w10801 & ~w15214 ) | ( w10801 & w15215 ) | ( ~w15214 & w15215 ) ;
  assign w15217 = w7944 | w10866 ;
  assign w15218 = w10874 | w15216 ;
  assign w15219 = ( w7414 & w15216 ) | ( w7414 & w15218 ) | ( w15216 & w15218 ) ;
  assign w15220 = ( ~w10866 & w15217 ) | ( ~w10866 & w15219 ) | ( w15217 & w15219 ) ;
  assign w15221 = \pi08 ^ w15220 ;
  assign w15222 = w14872 ^ w15187 ;
  assign w15223 = w14874 ^ w15222 ;
  assign w15224 = w7673 | w10807 ;
  assign w15225 = w7411 & ~w10805 ;
  assign w15226 = ( ~w10807 & w15224 ) | ( ~w10807 & w15225 ) | ( w15224 & w15225 ) ;
  assign w15227 = ~w7944 & w10801 ;
  assign w15228 = w10814 | w15226 ;
  assign w15229 = ( w7414 & w15226 ) | ( w7414 & w15228 ) | ( w15226 & w15228 ) ;
  assign w15230 = ( w10801 & ~w15227 ) | ( w10801 & w15229 ) | ( ~w15227 & w15229 ) ;
  assign w15231 = \pi08 ^ w15230 ;
  assign w15232 = w14882 ^ w15186 ;
  assign w15233 = w14884 ^ w15232 ;
  assign w15234 = w7673 | w10805 ;
  assign w15235 = w7411 & w10784 ;
  assign w15236 = ( ~w10805 & w15234 ) | ( ~w10805 & w15235 ) | ( w15234 & w15235 ) ;
  assign w15237 = w7944 | w10807 ;
  assign w15238 = w11117 | w15236 ;
  assign w15239 = ( w7414 & w15236 ) | ( w7414 & w15238 ) | ( w15236 & w15238 ) ;
  assign w15240 = ( ~w10807 & w15237 ) | ( ~w10807 & w15239 ) | ( w15237 & w15239 ) ;
  assign w15241 = \pi08 ^ w15240 ;
  assign w15242 = w14892 ^ w15185 ;
  assign w15243 = w14894 ^ w15242 ;
  assign w15244 = ~w7673 & w10784 ;
  assign w15245 = w7411 & w10211 ;
  assign w15246 = ( w10784 & ~w15244 ) | ( w10784 & w15245 ) | ( ~w15244 & w15245 ) ;
  assign w15247 = w7944 | w10805 ;
  assign w15248 = w10855 & ~w15246 ;
  assign w15249 = ( w7414 & w15246 ) | ( w7414 & ~w15248 ) | ( w15246 & ~w15248 ) ;
  assign w15250 = ( ~w10805 & w15247 ) | ( ~w10805 & w15249 ) | ( w15247 & w15249 ) ;
  assign w15251 = \pi08 ^ w15250 ;
  assign w15252 = w14902 ^ w15184 ;
  assign w15253 = w14904 ^ w15252 ;
  assign w15254 = ~w7673 & w10211 ;
  assign w15255 = w7411 & w10114 ;
  assign w15256 = ( w10211 & ~w15254 ) | ( w10211 & w15255 ) | ( ~w15254 & w15255 ) ;
  assign w15257 = ~w7944 & w10784 ;
  assign w15258 = w10789 | w15256 ;
  assign w15259 = ( w7414 & w15256 ) | ( w7414 & w15258 ) | ( w15256 & w15258 ) ;
  assign w15260 = ( w10784 & ~w15257 ) | ( w10784 & w15259 ) | ( ~w15257 & w15259 ) ;
  assign w15261 = \pi08 ^ w15260 ;
  assign w15262 = w14912 ^ w15183 ;
  assign w15263 = w14914 ^ w15262 ;
  assign w15264 = ~w7673 & w10114 ;
  assign w15265 = w7411 & w9953 ;
  assign w15266 = ( w10114 & ~w15264 ) | ( w10114 & w15265 ) | ( ~w15264 & w15265 ) ;
  assign w15267 = ~w7944 & w10211 ;
  assign w15268 = w10214 | w15266 ;
  assign w15269 = ( w7414 & w15266 ) | ( w7414 & w15268 ) | ( w15266 & w15268 ) ;
  assign w15270 = ( w10211 & ~w15267 ) | ( w10211 & w15269 ) | ( ~w15267 & w15269 ) ;
  assign w15271 = \pi08 ^ w15270 ;
  assign w15272 = w14922 ^ w15182 ;
  assign w15273 = w14924 ^ w15272 ;
  assign w15274 = ~w7673 & w9953 ;
  assign w15275 = w7411 & w9842 ;
  assign w15276 = ( w9953 & ~w15274 ) | ( w9953 & w15275 ) | ( ~w15274 & w15275 ) ;
  assign w15277 = ~w7944 & w10114 ;
  assign w15278 = w10334 | w15276 ;
  assign w15279 = ( w7414 & w15276 ) | ( w7414 & w15278 ) | ( w15276 & w15278 ) ;
  assign w15280 = ( w10114 & ~w15277 ) | ( w10114 & w15279 ) | ( ~w15277 & w15279 ) ;
  assign w15281 = \pi08 ^ w15280 ;
  assign w15282 = w14932 ^ w15181 ;
  assign w15283 = w14934 ^ w15282 ;
  assign w15284 = ~w7673 & w9842 ;
  assign w15285 = w7411 & ~w9955 ;
  assign w15286 = ( w9842 & ~w15284 ) | ( w9842 & w15285 ) | ( ~w15284 & w15285 ) ;
  assign w15287 = ~w7944 & w9953 ;
  assign w15288 = w10965 | w15286 ;
  assign w15289 = ( w7414 & w15286 ) | ( w7414 & w15288 ) | ( w15286 & w15288 ) ;
  assign w15290 = ( w9953 & ~w15287 ) | ( w9953 & w15289 ) | ( ~w15287 & w15289 ) ;
  assign w15291 = \pi08 ^ w15290 ;
  assign w15292 = w14942 ^ w15180 ;
  assign w15293 = w14944 ^ w15292 ;
  assign w15294 = w7673 | w9955 ;
  assign w15295 = w7411 & w9957 ;
  assign w15296 = ( ~w9955 & w15294 ) | ( ~w9955 & w15295 ) | ( w15294 & w15295 ) ;
  assign w15297 = ~w7944 & w9842 ;
  assign w15298 = w10976 & ~w15296 ;
  assign w15299 = ( w7414 & w15296 ) | ( w7414 & ~w15298 ) | ( w15296 & ~w15298 ) ;
  assign w15300 = ( w9842 & ~w15297 ) | ( w9842 & w15299 ) | ( ~w15297 & w15299 ) ;
  assign w15301 = \pi08 ^ w15300 ;
  assign w15302 = w14952 ^ w15179 ;
  assign w15303 = w14954 ^ w15302 ;
  assign w15304 = w7411 & ~w9963 ;
  assign w15305 = ( w7944 & ~w9955 ) | ( w7944 & w15304 ) | ( ~w9955 & w15304 ) ;
  assign w15306 = w7673 | w15305 ;
  assign w15307 = ( w9957 & w15305 ) | ( w9957 & w15306 ) | ( w15305 & w15306 ) ;
  assign w15308 = w15304 | w15307 ;
  assign w15309 = w7414 | w11202 ;
  assign w15310 = ( ~w11202 & w15308 ) | ( ~w11202 & w15309 ) | ( w15308 & w15309 ) ;
  assign w15311 = \pi08 ^ w15310 ;
  assign w15312 = w7673 | w9963 ;
  assign w15313 = w7411 & w9961 ;
  assign w15314 = ( ~w9963 & w15312 ) | ( ~w9963 & w15313 ) | ( w15312 & w15313 ) ;
  assign w15315 = ~w7944 & w9957 ;
  assign w15316 = w11089 & ~w15314 ;
  assign w15317 = ( w7414 & w15314 ) | ( w7414 & ~w15316 ) | ( w15314 & ~w15316 ) ;
  assign w15318 = ( w9957 & ~w15315 ) | ( w9957 & w15317 ) | ( ~w15315 & w15317 ) ;
  assign w15319 = \pi08 ^ w15318 ;
  assign w15320 = w14964 ^ w15178 ;
  assign w15321 = w14956 ^ w15320 ;
  assign w15322 = ~w7673 & w9961 ;
  assign w15323 = w7411 & w9965 ;
  assign w15324 = ( w9961 & ~w15322 ) | ( w9961 & w15323 ) | ( ~w15322 & w15323 ) ;
  assign w15325 = w7944 | w9963 ;
  assign w15326 = w11278 & ~w15324 ;
  assign w15327 = ( w7414 & w15324 ) | ( w7414 & ~w15326 ) | ( w15324 & ~w15326 ) ;
  assign w15328 = ( ~w9963 & w15325 ) | ( ~w9963 & w15327 ) | ( w15325 & w15327 ) ;
  assign w15329 = \pi08 ^ w15328 ;
  assign w15330 = w14974 ^ w15177 ;
  assign w15331 = w14966 ^ w15330 ;
  assign w15332 = w14982 ^ w15176 ;
  assign w15333 = w14984 ^ w15332 ;
  assign w15334 = w7411 & ~w9967 ;
  assign w15335 = ( w7944 & w9961 ) | ( w7944 & w15334 ) | ( w9961 & w15334 ) ;
  assign w15336 = w7673 | w15335 ;
  assign w15337 = ( w9965 & w15335 ) | ( w9965 & w15336 ) | ( w15335 & w15336 ) ;
  assign w15338 = w15334 | w15337 ;
  assign w15339 = ~w7414 & w11339 ;
  assign w15340 = ( w11339 & w15338 ) | ( w11339 & ~w15339 ) | ( w15338 & ~w15339 ) ;
  assign w15341 = \pi08 ^ w15340 ;
  assign w15342 = w14992 ^ w15175 ;
  assign w15343 = w14994 ^ w15342 ;
  assign w15344 = w7411 & w9971 ;
  assign w15345 = ( w7944 & w9965 ) | ( w7944 & w15344 ) | ( w9965 & w15344 ) ;
  assign w15346 = w7673 | w15345 ;
  assign w15347 = ( ~w9967 & w15345 ) | ( ~w9967 & w15346 ) | ( w15345 & w15346 ) ;
  assign w15348 = w15344 | w15347 ;
  assign w15349 = w7414 | w11501 ;
  assign w15350 = ( ~w11501 & w15348 ) | ( ~w11501 & w15349 ) | ( w15348 & w15349 ) ;
  assign w15351 = \pi08 ^ w15350 ;
  assign w15352 = w15002 ^ w15174 ;
  assign w15353 = w15004 ^ w15352 ;
  assign w15354 = w7411 & ~w9973 ;
  assign w15355 = ( w7944 & ~w9967 ) | ( w7944 & w15354 ) | ( ~w9967 & w15354 ) ;
  assign w15356 = w7673 | w15355 ;
  assign w15357 = ( w9971 & w15355 ) | ( w9971 & w15356 ) | ( w15355 & w15356 ) ;
  assign w15358 = w15354 | w15357 ;
  assign w15359 = w7414 | w11512 ;
  assign w15360 = ( ~w11512 & w15358 ) | ( ~w11512 & w15359 ) | ( w15358 & w15359 ) ;
  assign w15361 = \pi08 ^ w15360 ;
  assign w15362 = w7673 | w9973 ;
  assign w15363 = w7411 & w9975 ;
  assign w15364 = ( ~w9973 & w15362 ) | ( ~w9973 & w15363 ) | ( w15362 & w15363 ) ;
  assign w15365 = ~w7944 & w9971 ;
  assign w15366 = w11809 & ~w15364 ;
  assign w15367 = ( w7414 & w15364 ) | ( w7414 & ~w15366 ) | ( w15364 & ~w15366 ) ;
  assign w15368 = ( w9971 & ~w15365 ) | ( w9971 & w15367 ) | ( ~w15365 & w15367 ) ;
  assign w15369 = \pi08 ^ w15368 ;
  assign w15370 = w15014 ^ w15173 ;
  assign w15371 = w15006 ^ w15370 ;
  assign w15372 = ~w7673 & w9975 ;
  assign w15373 = w7411 & w9977 ;
  assign w15374 = ( w9975 & ~w15372 ) | ( w9975 & w15373 ) | ( ~w15372 & w15373 ) ;
  assign w15375 = w7944 | w9973 ;
  assign w15376 = w11671 & ~w15374 ;
  assign w15377 = ( w7414 & w15374 ) | ( w7414 & ~w15376 ) | ( w15374 & ~w15376 ) ;
  assign w15378 = ( ~w9973 & w15375 ) | ( ~w9973 & w15377 ) | ( w15375 & w15377 ) ;
  assign w15379 = \pi08 ^ w15378 ;
  assign w15380 = w15024 ^ w15172 ;
  assign w15381 = w15016 ^ w15380 ;
  assign w15382 = ~w7673 & w9977 ;
  assign w15383 = w7411 & w9979 ;
  assign w15384 = ( w9977 & ~w15382 ) | ( w9977 & w15383 ) | ( ~w15382 & w15383 ) ;
  assign w15385 = ~w7944 & w9975 ;
  assign w15386 = w11914 | w15384 ;
  assign w15387 = ( w7414 & w15384 ) | ( w7414 & w15386 ) | ( w15384 & w15386 ) ;
  assign w15388 = ( w9975 & ~w15385 ) | ( w9975 & w15387 ) | ( ~w15385 & w15387 ) ;
  assign w15389 = \pi08 ^ w15388 ;
  assign w15390 = w15034 ^ w15171 ;
  assign w15391 = w15026 ^ w15390 ;
  assign w15392 = w15042 ^ w15170 ;
  assign w15393 = w15044 ^ w15392 ;
  assign w15394 = w7411 & w9981 ;
  assign w15395 = ( w7944 & w9977 ) | ( w7944 & w15394 ) | ( w9977 & w15394 ) ;
  assign w15396 = w7673 | w15395 ;
  assign w15397 = ( w9979 & w15395 ) | ( w9979 & w15396 ) | ( w15395 & w15396 ) ;
  assign w15398 = w15394 | w15397 ;
  assign w15399 = ~w7414 & w12106 ;
  assign w15400 = ( w12106 & w15398 ) | ( w12106 & ~w15399 ) | ( w15398 & ~w15399 ) ;
  assign w15401 = \pi08 ^ w15400 ;
  assign w15402 = w15052 ^ w15169 ;
  assign w15403 = w15054 ^ w15402 ;
  assign w15404 = w7411 & w9983 ;
  assign w15405 = ( w7944 & w9979 ) | ( w7944 & w15404 ) | ( w9979 & w15404 ) ;
  assign w15406 = w7673 | w15405 ;
  assign w15407 = ( w9981 & w15405 ) | ( w9981 & w15406 ) | ( w15405 & w15406 ) ;
  assign w15408 = w15404 | w15407 ;
  assign w15409 = ~w7414 & w12010 ;
  assign w15410 = ( w12010 & w15408 ) | ( w12010 & ~w15409 ) | ( w15408 & ~w15409 ) ;
  assign w15411 = \pi08 ^ w15410 ;
  assign w15412 = w15062 ^ w15168 ;
  assign w15413 = w15064 ^ w15412 ;
  assign w15414 = w7411 & w9985 ;
  assign w15415 = ( w7944 & w9981 ) | ( w7944 & w15414 ) | ( w9981 & w15414 ) ;
  assign w15416 = w7673 | w15415 ;
  assign w15417 = ( w9983 & w15415 ) | ( w9983 & w15416 ) | ( w15415 & w15416 ) ;
  assign w15418 = w15414 | w15417 ;
  assign w15419 = ~w7414 & w12236 ;
  assign w15420 = ( w12236 & w15418 ) | ( w12236 & ~w15419 ) | ( w15418 & ~w15419 ) ;
  assign w15421 = \pi08 ^ w15420 ;
  assign w15422 = ~w7673 & w9985 ;
  assign w15423 = w7411 & w9987 ;
  assign w15424 = ( w9985 & ~w15422 ) | ( w9985 & w15423 ) | ( ~w15422 & w15423 ) ;
  assign w15425 = ~w7944 & w9983 ;
  assign w15426 = w12433 | w15424 ;
  assign w15427 = ( w7414 & w15424 ) | ( w7414 & w15426 ) | ( w15424 & w15426 ) ;
  assign w15428 = ( w9983 & ~w15425 ) | ( w9983 & w15427 ) | ( ~w15425 & w15427 ) ;
  assign w15429 = \pi08 ^ w15428 ;
  assign w15430 = w15074 ^ w15167 ;
  assign w15431 = w15066 ^ w15430 ;
  assign w15432 = ~w7673 & w9987 ;
  assign w15433 = w7411 & ~w9989 ;
  assign w15434 = ( w9987 & ~w15432 ) | ( w9987 & w15433 ) | ( ~w15432 & w15433 ) ;
  assign w15435 = ~w7944 & w9985 ;
  assign w15436 = w12446 | w15434 ;
  assign w15437 = ( w7414 & w15434 ) | ( w7414 & w15436 ) | ( w15434 & w15436 ) ;
  assign w15438 = ( w9985 & ~w15435 ) | ( w9985 & w15437 ) | ( ~w15435 & w15437 ) ;
  assign w15439 = \pi08 ^ w15438 ;
  assign w15440 = w15084 ^ w15166 ;
  assign w15441 = w15076 ^ w15440 ;
  assign w15442 = w7673 | w9989 ;
  assign w15443 = w7411 & w9991 ;
  assign w15444 = ( ~w9989 & w15442 ) | ( ~w9989 & w15443 ) | ( w15442 & w15443 ) ;
  assign w15445 = ~w7944 & w9987 ;
  assign w15446 = w12217 & ~w15444 ;
  assign w15447 = ( w7414 & w15444 ) | ( w7414 & ~w15446 ) | ( w15444 & ~w15446 ) ;
  assign w15448 = ( w9987 & ~w15445 ) | ( w9987 & w15447 ) | ( ~w15445 & w15447 ) ;
  assign w15449 = \pi08 ^ w15448 ;
  assign w15450 = w15094 ^ w15165 ;
  assign w15451 = w15086 ^ w15450 ;
  assign w15452 = w15102 ^ w15164 ;
  assign w15453 = w15104 ^ w15452 ;
  assign w15454 = w7411 & ~w9993 ;
  assign w15455 = ( w7944 & ~w9989 ) | ( w7944 & w15454 ) | ( ~w9989 & w15454 ) ;
  assign w15456 = w7673 | w15455 ;
  assign w15457 = ( w9991 & w15455 ) | ( w9991 & w15456 ) | ( w15455 & w15456 ) ;
  assign w15458 = w15454 | w15457 ;
  assign w15459 = w7414 | w12484 ;
  assign w15460 = ( ~w12484 & w15458 ) | ( ~w12484 & w15459 ) | ( w15458 & w15459 ) ;
  assign w15461 = \pi08 ^ w15460 ;
  assign w15462 = w15114 ^ w15163 ;
  assign w15463 = w15106 ^ w15462 ;
  assign w15464 = w7411 & w9995 ;
  assign w15465 = ( w7944 & w9991 ) | ( w7944 & w15464 ) | ( w9991 & w15464 ) ;
  assign w15466 = w7673 | w15465 ;
  assign w15467 = ( ~w9993 & w15465 ) | ( ~w9993 & w15466 ) | ( w15465 & w15466 ) ;
  assign w15468 = w15464 | w15467 ;
  assign w15469 = w7414 | w12514 ;
  assign w15470 = ( ~w12514 & w15468 ) | ( ~w12514 & w15469 ) | ( w15468 & w15469 ) ;
  assign w15471 = \pi08 ^ w15470 ;
  assign w15472 = w15122 ^ w15162 ;
  assign w15473 = w15123 ^ w15472 ;
  assign w15474 = w7411 & w9997 ;
  assign w15475 = ( w7944 & ~w9993 ) | ( w7944 & w15474 ) | ( ~w9993 & w15474 ) ;
  assign w15476 = w7673 | w15475 ;
  assign w15477 = ( w9995 & w15475 ) | ( w9995 & w15476 ) | ( w15475 & w15476 ) ;
  assign w15478 = w15474 | w15477 ;
  assign w15479 = w7414 | w12541 ;
  assign w15480 = ( ~w12541 & w15478 ) | ( ~w12541 & w15479 ) | ( w15478 & w15479 ) ;
  assign w15481 = \pi08 ^ w15480 ;
  assign w15482 = ~w7673 & w9997 ;
  assign w15483 = w7411 & w9999 ;
  assign w15484 = ( w9997 & ~w15482 ) | ( w9997 & w15483 ) | ( ~w15482 & w15483 ) ;
  assign w15485 = ~w7944 & w9995 ;
  assign w15486 = w12572 | w15484 ;
  assign w15487 = ( w7414 & w15484 ) | ( w7414 & w15486 ) | ( w15484 & w15486 ) ;
  assign w15488 = ( w9995 & ~w15485 ) | ( w9995 & w15487 ) | ( ~w15485 & w15487 ) ;
  assign w15489 = \pi08 ^ w15488 ;
  assign w15490 = w15136 ^ w15161 ;
  assign w15491 = w15128 ^ w15490 ;
  assign w15492 = w15151 ^ w15159 ;
  assign w15493 = w15160 ^ w15492 ;
  assign w15494 = w7411 & w10001 ;
  assign w15495 = ( w7944 & w9997 ) | ( w7944 & w15494 ) | ( w9997 & w15494 ) ;
  assign w15496 = w7673 | w15495 ;
  assign w15497 = ( w9999 & w15495 ) | ( w9999 & w15496 ) | ( w15495 & w15496 ) ;
  assign w15498 = w15494 | w15497 ;
  assign w15499 = ~w7414 & w12641 ;
  assign w15500 = ( w12641 & w15498 ) | ( w12641 & ~w15499 ) | ( w15498 & ~w15499 ) ;
  assign w15501 = \pi08 ^ w15500 ;
  assign w15502 = ~w7673 & w10001 ;
  assign w15503 = w7411 & ~w10006 ;
  assign w15504 = ( w10001 & ~w15502 ) | ( w10001 & w15503 ) | ( ~w15502 & w15503 ) ;
  assign w15505 = ~w7944 & w9999 ;
  assign w15506 = w12691 & ~w15504 ;
  assign w15507 = ( w7414 & w15504 ) | ( w7414 & ~w15506 ) | ( w15504 & ~w15506 ) ;
  assign w15508 = ( w9999 & ~w15505 ) | ( w9999 & w15507 ) | ( ~w15505 & w15507 ) ;
  assign w15509 = \pi08 ^ w15508 ;
  assign w15510 = w15142 ^ w15150 ;
  assign w15511 = ( \pi08 & \pi09 ) | ( \pi08 & ~w10016 ) | ( \pi09 & ~w10016 ) ;
  assign w15512 = ( \pi08 & \pi09 ) | ( \pi08 & ~w10021 ) | ( \pi09 & ~w10021 ) ;
  assign w15513 = \pi10 ^ w10021 ;
  assign w15514 = ( \pi10 & w15512 ) | ( \pi10 & w15513 ) | ( w15512 & w15513 ) ;
  assign w15515 = w15511 ^ w15514 ;
  assign w15516 = w7411 & w10011 ;
  assign w15517 = ( w7944 & w10001 ) | ( w7944 & w15516 ) | ( w10001 & w15516 ) ;
  assign w15518 = w7673 | w15517 ;
  assign w15519 = ( ~w10006 & w15517 ) | ( ~w10006 & w15518 ) | ( w15517 & w15518 ) ;
  assign w15520 = w15516 | w15519 ;
  assign w15521 = ~w7414 & w12747 ;
  assign w15522 = ( w12747 & w15520 ) | ( w12747 & ~w15521 ) | ( w15520 & ~w15521 ) ;
  assign w15523 = \pi08 ^ w15522 ;
  assign w15524 = \pi08 & w10021 ;
  assign w15525 = w10016 & w15524 ;
  assign w15526 = ( \pi05 & \pi06 ) | ( \pi05 & ~w15525 ) | ( \pi06 & ~w15525 ) ;
  assign w15527 = ( \pi07 & \pi08 ) | ( \pi07 & ~w15526 ) | ( \pi08 & ~w15526 ) ;
  assign w15528 = ( \pi07 & ~w15524 ) | ( \pi07 & w15526 ) | ( ~w15524 & w15526 ) ;
  assign w15529 = ( w8885 & w15527 ) | ( w8885 & ~w15528 ) | ( w15527 & ~w15528 ) ;
  assign w15530 = w7411 & ~w10021 ;
  assign w15531 = ( w7944 & w10011 ) | ( w7944 & w15530 ) | ( w10011 & w15530 ) ;
  assign w15532 = w7673 | w15531 ;
  assign w15533 = ( ~w10016 & w15531 ) | ( ~w10016 & w15532 ) | ( w15531 & w15532 ) ;
  assign w15534 = w15530 | w15533 ;
  assign w15535 = ~w7414 & w12867 ;
  assign w15536 = ( w12867 & w15534 ) | ( w12867 & ~w15535 ) | ( w15534 & ~w15535 ) ;
  assign w15537 = \pi08 ^ w15536 ;
  assign w15538 = w15529 & w15537 ;
  assign w15539 = ~w7673 & w10011 ;
  assign w15540 = w7411 & ~w10016 ;
  assign w15541 = ( w10011 & ~w15539 ) | ( w10011 & w15540 ) | ( ~w15539 & w15540 ) ;
  assign w15542 = w7944 | w10006 ;
  assign w15543 = w12777 | w15541 ;
  assign w15544 = ( w7414 & w15541 ) | ( w7414 & w15543 ) | ( w15541 & w15543 ) ;
  assign w15545 = ( ~w10006 & w15542 ) | ( ~w10006 & w15544 ) | ( w15542 & w15544 ) ;
  assign w15546 = \pi08 ^ w15545 ;
  assign w15547 = w6750 & ~w10021 ;
  assign w15548 = ( w15538 & w15546 ) | ( w15538 & w15547 ) | ( w15546 & w15547 ) ;
  assign w15549 = ( w15515 & w15523 ) | ( w15515 & w15548 ) | ( w15523 & w15548 ) ;
  assign w15550 = ( w15509 & w15510 ) | ( w15509 & w15549 ) | ( w15510 & w15549 ) ;
  assign w15551 = ( w15493 & w15501 ) | ( w15493 & w15550 ) | ( w15501 & w15550 ) ;
  assign w15552 = ( w15489 & w15491 ) | ( w15489 & w15551 ) | ( w15491 & w15551 ) ;
  assign w15553 = ( w15473 & w15481 ) | ( w15473 & w15552 ) | ( w15481 & w15552 ) ;
  assign w15554 = ( w15463 & w15471 ) | ( w15463 & w15553 ) | ( w15471 & w15553 ) ;
  assign w15555 = ( w15453 & w15461 ) | ( w15453 & w15554 ) | ( w15461 & w15554 ) ;
  assign w15556 = ( w15449 & w15451 ) | ( w15449 & w15555 ) | ( w15451 & w15555 ) ;
  assign w15557 = ( w15439 & w15441 ) | ( w15439 & w15556 ) | ( w15441 & w15556 ) ;
  assign w15558 = ( w15429 & w15431 ) | ( w15429 & w15557 ) | ( w15431 & w15557 ) ;
  assign w15559 = ( w15413 & w15421 ) | ( w15413 & w15558 ) | ( w15421 & w15558 ) ;
  assign w15560 = ( w15403 & w15411 ) | ( w15403 & w15559 ) | ( w15411 & w15559 ) ;
  assign w15561 = ( w15393 & w15401 ) | ( w15393 & w15560 ) | ( w15401 & w15560 ) ;
  assign w15562 = ( w15389 & w15391 ) | ( w15389 & w15561 ) | ( w15391 & w15561 ) ;
  assign w15563 = ( w15379 & w15381 ) | ( w15379 & w15562 ) | ( w15381 & w15562 ) ;
  assign w15564 = ( w15369 & w15371 ) | ( w15369 & w15563 ) | ( w15371 & w15563 ) ;
  assign w15565 = ( w15353 & w15361 ) | ( w15353 & w15564 ) | ( w15361 & w15564 ) ;
  assign w15566 = ( w15343 & w15351 ) | ( w15343 & w15565 ) | ( w15351 & w15565 ) ;
  assign w15567 = ( w15333 & w15341 ) | ( w15333 & w15566 ) | ( w15341 & w15566 ) ;
  assign w15568 = ( w15329 & w15331 ) | ( w15329 & w15567 ) | ( w15331 & w15567 ) ;
  assign w15569 = ( w15319 & w15321 ) | ( w15319 & w15568 ) | ( w15321 & w15568 ) ;
  assign w15570 = ( ~w15303 & w15311 ) | ( ~w15303 & w15569 ) | ( w15311 & w15569 ) ;
  assign w15571 = ( ~w15293 & w15301 ) | ( ~w15293 & w15570 ) | ( w15301 & w15570 ) ;
  assign w15572 = ( w15283 & w15291 ) | ( w15283 & w15571 ) | ( w15291 & w15571 ) ;
  assign w15573 = ( ~w15273 & w15281 ) | ( ~w15273 & w15572 ) | ( w15281 & w15572 ) ;
  assign w15574 = ( ~w15263 & w15271 ) | ( ~w15263 & w15573 ) | ( w15271 & w15573 ) ;
  assign w15575 = ( w15253 & w15261 ) | ( w15253 & w15574 ) | ( w15261 & w15574 ) ;
  assign w15576 = ( w15243 & w15251 ) | ( w15243 & w15575 ) | ( w15251 & w15575 ) ;
  assign w15577 = ( w15233 & w15241 ) | ( w15233 & w15576 ) | ( w15241 & w15576 ) ;
  assign w15578 = ( w15223 & w15231 ) | ( w15223 & w15577 ) | ( w15231 & w15577 ) ;
  assign w15579 = ( w15213 & w15221 ) | ( w15213 & w15578 ) | ( w15221 & w15578 ) ;
  assign w15580 = ~w8593 & w10883 ;
  assign w15581 = w8262 & ~w10887 ;
  assign w15582 = ( w10883 & ~w15580 ) | ( w10883 & w15581 ) | ( ~w15580 & w15581 ) ;
  assign w15583 = ~w8263 & w11256 ;
  assign w15584 = w11139 & ~w15582 ;
  assign w15585 = ( w35 & w15582 ) | ( w35 & ~w15584 ) | ( w15582 & ~w15584 ) ;
  assign w15586 = ( w11256 & ~w15583 ) | ( w11256 & w15585 ) | ( ~w15583 & w15585 ) ;
  assign w15587 = \pi05 ^ w15586 ;
  assign w15588 = ( ~w15211 & w15579 ) | ( ~w15211 & w15587 ) | ( w15579 & w15587 ) ;
  assign w15589 = w15211 ^ w15587 ;
  assign w15590 = w15579 ^ w15589 ;
  assign w15591 = w8593 | w10887 ;
  assign w15592 = w8262 & ~w10885 ;
  assign w15593 = ( ~w10887 & w15591 ) | ( ~w10887 & w15592 ) | ( w15591 & w15592 ) ;
  assign w15594 = ~w8263 & w10895 ;
  assign w15595 = w10883 | w15593 ;
  assign w15596 = ( w35 & w15593 ) | ( w35 & w15595 ) | ( w15593 & w15595 ) ;
  assign w15597 = ( w10895 & ~w15594 ) | ( w10895 & w15596 ) | ( ~w15594 & w15596 ) ;
  assign w15598 = \pi05 ^ w15597 ;
  assign w15599 = w15221 ^ w15578 ;
  assign w15600 = w15213 ^ w15599 ;
  assign w15601 = w15598 ^ w15600 ;
  assign w15602 = \pi00 ^ w10738 ;
  assign w15603 = ( w10738 & w11146 ) | ( w10738 & w15602 ) | ( w11146 & w15602 ) ;
  assign w15604 = ( \pi02 & ~w10738 ) | ( \pi02 & w15603 ) | ( ~w10738 & w15603 ) ;
  assign w15605 = \pi01 & ~w11146 ;
  assign w15606 = ( \pi02 & w10738 ) | ( \pi02 & w11138 ) | ( w10738 & w11138 ) ;
  assign w15607 = ( \pi00 & w15604 ) | ( \pi00 & ~w15606 ) | ( w15604 & ~w15606 ) ;
  assign w15608 = ( ~w15603 & w15605 ) | ( ~w15603 & w15607 ) | ( w15605 & w15607 ) ;
  assign w15609 = ( \pi01 & ~w10738 ) | ( \pi01 & w15608 ) | ( ~w10738 & w15608 ) ;
  assign w15610 = w15604 ^ w15609 ;
  assign w15611 = ( w15598 & w15600 ) | ( w15598 & w15610 ) | ( w15600 & w15610 ) ;
  assign w15612 = w8593 | w10885 ;
  assign w15613 = w8262 & ~w10866 ;
  assign w15614 = ( ~w10885 & w15612 ) | ( ~w10885 & w15613 ) | ( w15612 & w15613 ) ;
  assign w15615 = w8263 | w11131 ;
  assign w15616 = w10887 & ~w15614 ;
  assign w15617 = ( w35 & w15614 ) | ( w35 & ~w15616 ) | ( w15614 & ~w15616 ) ;
  assign w15618 = ( ~w11131 & w15615 ) | ( ~w11131 & w15617 ) | ( w15615 & w15617 ) ;
  assign w15619 = \pi05 ^ w15618 ;
  assign w15620 = w15231 ^ w15577 ;
  assign w15621 = w15223 ^ w15620 ;
  assign w15622 = w8593 | w10866 ;
  assign w15623 = w8262 & w10801 ;
  assign w15624 = ( ~w10866 & w15622 ) | ( ~w10866 & w15623 ) | ( w15622 & w15623 ) ;
  assign w15625 = w8263 | w11160 ;
  assign w15626 = w10885 & ~w15624 ;
  assign w15627 = ( w35 & w15624 ) | ( w35 & ~w15626 ) | ( w15624 & ~w15626 ) ;
  assign w15628 = ( ~w11160 & w15625 ) | ( ~w11160 & w15627 ) | ( w15625 & w15627 ) ;
  assign w15629 = \pi05 ^ w15628 ;
  assign w15630 = w15241 ^ w15576 ;
  assign w15631 = w15233 ^ w15630 ;
  assign w15632 = ~w8593 & w10801 ;
  assign w15633 = w8262 & ~w10807 ;
  assign w15634 = ( w10801 & ~w15632 ) | ( w10801 & w15633 ) | ( ~w15632 & w15633 ) ;
  assign w15635 = ~w8263 & w10874 ;
  assign w15636 = w10866 & ~w15634 ;
  assign w15637 = ( w35 & w15634 ) | ( w35 & ~w15636 ) | ( w15634 & ~w15636 ) ;
  assign w15638 = ( w10874 & ~w15635 ) | ( w10874 & w15637 ) | ( ~w15635 & w15637 ) ;
  assign w15639 = \pi05 ^ w15638 ;
  assign w15640 = w15251 ^ w15575 ;
  assign w15641 = w15243 ^ w15640 ;
  assign w15642 = w8593 | w10807 ;
  assign w15643 = w8262 & ~w10805 ;
  assign w15644 = ( ~w10807 & w15642 ) | ( ~w10807 & w15643 ) | ( w15642 & w15643 ) ;
  assign w15645 = ~w8263 & w10814 ;
  assign w15646 = w10801 | w15644 ;
  assign w15647 = ( w35 & w15644 ) | ( w35 & w15646 ) | ( w15644 & w15646 ) ;
  assign w15648 = ( w10814 & ~w15645 ) | ( w10814 & w15647 ) | ( ~w15645 & w15647 ) ;
  assign w15649 = \pi05 ^ w15648 ;
  assign w15650 = w15261 ^ w15574 ;
  assign w15651 = w15253 ^ w15650 ;
  assign w15652 = w8593 | w10805 ;
  assign w15653 = w8262 & w10784 ;
  assign w15654 = ( ~w10805 & w15652 ) | ( ~w10805 & w15653 ) | ( w15652 & w15653 ) ;
  assign w15655 = ~w8263 & w11117 ;
  assign w15656 = w10807 & ~w15654 ;
  assign w15657 = ( w35 & w15654 ) | ( w35 & ~w15656 ) | ( w15654 & ~w15656 ) ;
  assign w15658 = ( w11117 & ~w15655 ) | ( w11117 & w15657 ) | ( ~w15655 & w15657 ) ;
  assign w15659 = \pi05 ^ w15658 ;
  assign w15660 = w15271 ^ w15573 ;
  assign w15661 = w15263 ^ w15660 ;
  assign w15662 = ~w8593 & w10784 ;
  assign w15663 = w8262 & w10211 ;
  assign w15664 = ( w10784 & ~w15662 ) | ( w10784 & w15663 ) | ( ~w15662 & w15663 ) ;
  assign w15665 = w8263 | w10855 ;
  assign w15666 = w10805 & ~w15664 ;
  assign w15667 = ( w35 & w15664 ) | ( w35 & ~w15666 ) | ( w15664 & ~w15666 ) ;
  assign w15668 = ( ~w10855 & w15665 ) | ( ~w10855 & w15667 ) | ( w15665 & w15667 ) ;
  assign w15669 = \pi05 ^ w15668 ;
  assign w15670 = w15281 ^ w15572 ;
  assign w15671 = w15273 ^ w15670 ;
  assign w15672 = ~w8593 & w10211 ;
  assign w15673 = w8262 & w10114 ;
  assign w15674 = ( w10211 & ~w15672 ) | ( w10211 & w15673 ) | ( ~w15672 & w15673 ) ;
  assign w15675 = ~w8263 & w10789 ;
  assign w15676 = w10784 | w15674 ;
  assign w15677 = ( w35 & w15674 ) | ( w35 & w15676 ) | ( w15674 & w15676 ) ;
  assign w15678 = ( w10789 & ~w15675 ) | ( w10789 & w15677 ) | ( ~w15675 & w15677 ) ;
  assign w15679 = \pi05 ^ w15678 ;
  assign w15680 = w15291 ^ w15571 ;
  assign w15681 = w15283 ^ w15680 ;
  assign w15682 = ~w8593 & w10114 ;
  assign w15683 = w8262 & w9953 ;
  assign w15684 = ( w10114 & ~w15682 ) | ( w10114 & w15683 ) | ( ~w15682 & w15683 ) ;
  assign w15685 = ~w8263 & w10214 ;
  assign w15686 = w10211 | w15684 ;
  assign w15687 = ( w35 & w15684 ) | ( w35 & w15686 ) | ( w15684 & w15686 ) ;
  assign w15688 = ( w10214 & ~w15685 ) | ( w10214 & w15687 ) | ( ~w15685 & w15687 ) ;
  assign w15689 = \pi05 ^ w15688 ;
  assign w15690 = w15301 ^ w15570 ;
  assign w15691 = w15293 ^ w15690 ;
  assign w15692 = ~w8593 & w9953 ;
  assign w15693 = w8262 & w9842 ;
  assign w15694 = ( w9953 & ~w15692 ) | ( w9953 & w15693 ) | ( ~w15692 & w15693 ) ;
  assign w15695 = ~w8263 & w10334 ;
  assign w15696 = w10114 | w15694 ;
  assign w15697 = ( w35 & w15694 ) | ( w35 & w15696 ) | ( w15694 & w15696 ) ;
  assign w15698 = ( w10334 & ~w15695 ) | ( w10334 & w15697 ) | ( ~w15695 & w15697 ) ;
  assign w15699 = \pi05 ^ w15698 ;
  assign w15700 = w15311 ^ w15569 ;
  assign w15701 = w15303 ^ w15700 ;
  assign w15702 = w15319 ^ w15568 ;
  assign w15703 = w15321 ^ w15702 ;
  assign w15704 = ~w8593 & w9842 ;
  assign w15705 = w8262 & ~w9955 ;
  assign w15706 = ( w9842 & ~w15704 ) | ( w9842 & w15705 ) | ( ~w15704 & w15705 ) ;
  assign w15707 = ~w8263 & w10965 ;
  assign w15708 = w9953 | w15706 ;
  assign w15709 = ( w35 & w15706 ) | ( w35 & w15708 ) | ( w15706 & w15708 ) ;
  assign w15710 = ( w10965 & ~w15707 ) | ( w10965 & w15709 ) | ( ~w15707 & w15709 ) ;
  assign w15711 = \pi05 ^ w15710 ;
  assign w15712 = w15329 ^ w15567 ;
  assign w15713 = w15331 ^ w15712 ;
  assign w15714 = w8593 | w9955 ;
  assign w15715 = w8262 & w9957 ;
  assign w15716 = ( ~w9955 & w15714 ) | ( ~w9955 & w15715 ) | ( w15714 & w15715 ) ;
  assign w15717 = w8263 | w10976 ;
  assign w15718 = w9842 | w15716 ;
  assign w15719 = ( w35 & w15716 ) | ( w35 & w15718 ) | ( w15716 & w15718 ) ;
  assign w15720 = ( ~w10976 & w15717 ) | ( ~w10976 & w15719 ) | ( w15717 & w15719 ) ;
  assign w15721 = \pi05 ^ w15720 ;
  assign w15722 = ~w8593 & w9957 ;
  assign w15723 = w8262 & ~w9963 ;
  assign w15724 = ( w9957 & ~w15722 ) | ( w9957 & w15723 ) | ( ~w15722 & w15723 ) ;
  assign w15725 = w8263 | w11202 ;
  assign w15726 = w9955 & ~w15724 ;
  assign w15727 = ( w35 & w15724 ) | ( w35 & ~w15726 ) | ( w15724 & ~w15726 ) ;
  assign w15728 = ( ~w11202 & w15725 ) | ( ~w11202 & w15727 ) | ( w15725 & w15727 ) ;
  assign w15729 = \pi05 ^ w15728 ;
  assign w15730 = w15341 ^ w15566 ;
  assign w15731 = w15333 ^ w15730 ;
  assign w15732 = w8593 | w9963 ;
  assign w15733 = w8262 & w9961 ;
  assign w15734 = ( ~w9963 & w15732 ) | ( ~w9963 & w15733 ) | ( w15732 & w15733 ) ;
  assign w15735 = w8263 | w11089 ;
  assign w15736 = w9957 | w15734 ;
  assign w15737 = ( w35 & w15734 ) | ( w35 & w15736 ) | ( w15734 & w15736 ) ;
  assign w15738 = ( ~w11089 & w15735 ) | ( ~w11089 & w15737 ) | ( w15735 & w15737 ) ;
  assign w15739 = \pi05 ^ w15738 ;
  assign w15740 = w15351 ^ w15565 ;
  assign w15741 = w15343 ^ w15740 ;
  assign w15742 = ~w8593 & w9961 ;
  assign w15743 = w8262 & w9965 ;
  assign w15744 = ( w9961 & ~w15742 ) | ( w9961 & w15743 ) | ( ~w15742 & w15743 ) ;
  assign w15745 = w8263 | w11278 ;
  assign w15746 = w9963 & ~w15744 ;
  assign w15747 = ( w35 & w15744 ) | ( w35 & ~w15746 ) | ( w15744 & ~w15746 ) ;
  assign w15748 = ( ~w11278 & w15745 ) | ( ~w11278 & w15747 ) | ( w15745 & w15747 ) ;
  assign w15749 = \pi05 ^ w15748 ;
  assign w15750 = w15361 ^ w15564 ;
  assign w15751 = w15353 ^ w15750 ;
  assign w15752 = w15369 ^ w15563 ;
  assign w15753 = w15371 ^ w15752 ;
  assign w15754 = w35 & w9961 ;
  assign w15755 = ( w8593 & w9965 ) | ( w8593 & w15754 ) | ( w9965 & w15754 ) ;
  assign w15756 = w8262 | w15755 ;
  assign w15757 = ( ~w9967 & w15755 ) | ( ~w9967 & w15756 ) | ( w15755 & w15756 ) ;
  assign w15758 = w15754 | w15757 ;
  assign w15759 = ~w8263 & w11339 ;
  assign w15760 = ( w11339 & w15758 ) | ( w11339 & ~w15759 ) | ( w15758 & ~w15759 ) ;
  assign w15761 = \pi05 ^ w15760 ;
  assign w15762 = w15379 ^ w15562 ;
  assign w15763 = w15381 ^ w15762 ;
  assign w15764 = w35 & w9965 ;
  assign w15765 = ( w8593 & ~w9967 ) | ( w8593 & w15764 ) | ( ~w9967 & w15764 ) ;
  assign w15766 = w8262 | w15765 ;
  assign w15767 = ( w9971 & w15765 ) | ( w9971 & w15766 ) | ( w15765 & w15766 ) ;
  assign w15768 = w15764 | w15767 ;
  assign w15769 = w8263 | w11501 ;
  assign w15770 = ( ~w11501 & w15768 ) | ( ~w11501 & w15769 ) | ( w15768 & w15769 ) ;
  assign w15771 = \pi05 ^ w15770 ;
  assign w15772 = w15389 ^ w15561 ;
  assign w15773 = w15391 ^ w15772 ;
  assign w15774 = w35 & ~w9967 ;
  assign w15775 = ( w8593 & w9971 ) | ( w8593 & w15774 ) | ( w9971 & w15774 ) ;
  assign w15776 = w8262 | w15775 ;
  assign w15777 = ( ~w9973 & w15775 ) | ( ~w9973 & w15776 ) | ( w15775 & w15776 ) ;
  assign w15778 = w15774 | w15777 ;
  assign w15779 = w8263 | w11512 ;
  assign w15780 = ( ~w11512 & w15778 ) | ( ~w11512 & w15779 ) | ( w15778 & w15779 ) ;
  assign w15781 = \pi05 ^ w15780 ;
  assign w15782 = w8593 | w9973 ;
  assign w15783 = w8262 & w9975 ;
  assign w15784 = ( ~w9973 & w15782 ) | ( ~w9973 & w15783 ) | ( w15782 & w15783 ) ;
  assign w15785 = w8263 | w11809 ;
  assign w15786 = w9971 | w15784 ;
  assign w15787 = ( w35 & w15784 ) | ( w35 & w15786 ) | ( w15784 & w15786 ) ;
  assign w15788 = ( ~w11809 & w15785 ) | ( ~w11809 & w15787 ) | ( w15785 & w15787 ) ;
  assign w15789 = \pi05 ^ w15788 ;
  assign w15790 = w15401 ^ w15560 ;
  assign w15791 = w15393 ^ w15790 ;
  assign w15792 = ~w8593 & w9975 ;
  assign w15793 = w8262 & w9977 ;
  assign w15794 = ( w9975 & ~w15792 ) | ( w9975 & w15793 ) | ( ~w15792 & w15793 ) ;
  assign w15795 = w8263 | w11671 ;
  assign w15796 = w9973 & ~w15794 ;
  assign w15797 = ( w35 & w15794 ) | ( w35 & ~w15796 ) | ( w15794 & ~w15796 ) ;
  assign w15798 = ( ~w11671 & w15795 ) | ( ~w11671 & w15797 ) | ( w15795 & w15797 ) ;
  assign w15799 = \pi05 ^ w15798 ;
  assign w15800 = w15411 ^ w15559 ;
  assign w15801 = w15403 ^ w15800 ;
  assign w15802 = ~w8593 & w9977 ;
  assign w15803 = w8262 & w9979 ;
  assign w15804 = ( w9977 & ~w15802 ) | ( w9977 & w15803 ) | ( ~w15802 & w15803 ) ;
  assign w15805 = ~w8263 & w11914 ;
  assign w15806 = w9975 | w15804 ;
  assign w15807 = ( w35 & w15804 ) | ( w35 & w15806 ) | ( w15804 & w15806 ) ;
  assign w15808 = ( w11914 & ~w15805 ) | ( w11914 & w15807 ) | ( ~w15805 & w15807 ) ;
  assign w15809 = \pi05 ^ w15808 ;
  assign w15810 = w15421 ^ w15558 ;
  assign w15811 = w15413 ^ w15810 ;
  assign w15812 = w15429 ^ w15557 ;
  assign w15813 = w15431 ^ w15812 ;
  assign w15814 = w35 & w9977 ;
  assign w15815 = ( w8593 & w9979 ) | ( w8593 & w15814 ) | ( w9979 & w15814 ) ;
  assign w15816 = w8262 | w15815 ;
  assign w15817 = ( w9981 & w15815 ) | ( w9981 & w15816 ) | ( w15815 & w15816 ) ;
  assign w15818 = w15814 | w15817 ;
  assign w15819 = ~w8263 & w12106 ;
  assign w15820 = ( w12106 & w15818 ) | ( w12106 & ~w15819 ) | ( w15818 & ~w15819 ) ;
  assign w15821 = \pi05 ^ w15820 ;
  assign w15822 = w15439 ^ w15556 ;
  assign w15823 = w15441 ^ w15822 ;
  assign w15824 = w35 & w9979 ;
  assign w15825 = ( w8593 & w9981 ) | ( w8593 & w15824 ) | ( w9981 & w15824 ) ;
  assign w15826 = w8262 | w15825 ;
  assign w15827 = ( w9983 & w15825 ) | ( w9983 & w15826 ) | ( w15825 & w15826 ) ;
  assign w15828 = w15824 | w15827 ;
  assign w15829 = ~w8263 & w12010 ;
  assign w15830 = ( w12010 & w15828 ) | ( w12010 & ~w15829 ) | ( w15828 & ~w15829 ) ;
  assign w15831 = \pi05 ^ w15830 ;
  assign w15832 = w15449 ^ w15555 ;
  assign w15833 = w15451 ^ w15832 ;
  assign w15834 = w35 & w9981 ;
  assign w15835 = ( w8593 & w9983 ) | ( w8593 & w15834 ) | ( w9983 & w15834 ) ;
  assign w15836 = w8262 | w15835 ;
  assign w15837 = ( w9985 & w15835 ) | ( w9985 & w15836 ) | ( w15835 & w15836 ) ;
  assign w15838 = w15834 | w15837 ;
  assign w15839 = ~w8263 & w12236 ;
  assign w15840 = ( w12236 & w15838 ) | ( w12236 & ~w15839 ) | ( w15838 & ~w15839 ) ;
  assign w15841 = \pi05 ^ w15840 ;
  assign w15842 = ~w8593 & w9985 ;
  assign w15843 = w8262 & w9987 ;
  assign w15844 = ( w9985 & ~w15842 ) | ( w9985 & w15843 ) | ( ~w15842 & w15843 ) ;
  assign w15845 = ~w8263 & w12433 ;
  assign w15846 = w9983 | w15844 ;
  assign w15847 = ( w35 & w15844 ) | ( w35 & w15846 ) | ( w15844 & w15846 ) ;
  assign w15848 = ( w12433 & ~w15845 ) | ( w12433 & w15847 ) | ( ~w15845 & w15847 ) ;
  assign w15849 = \pi05 ^ w15848 ;
  assign w15850 = w15461 ^ w15554 ;
  assign w15851 = w15453 ^ w15850 ;
  assign w15852 = ~w8593 & w9987 ;
  assign w15853 = w8262 & ~w9989 ;
  assign w15854 = ( w9987 & ~w15852 ) | ( w9987 & w15853 ) | ( ~w15852 & w15853 ) ;
  assign w15855 = ~w8263 & w12446 ;
  assign w15856 = w9985 | w15854 ;
  assign w15857 = ( w35 & w15854 ) | ( w35 & w15856 ) | ( w15854 & w15856 ) ;
  assign w15858 = ( w12446 & ~w15855 ) | ( w12446 & w15857 ) | ( ~w15855 & w15857 ) ;
  assign w15859 = \pi05 ^ w15858 ;
  assign w15860 = w15471 ^ w15553 ;
  assign w15861 = w15463 ^ w15860 ;
  assign w15862 = w8593 | w9989 ;
  assign w15863 = w8262 & w9991 ;
  assign w15864 = ( ~w9989 & w15862 ) | ( ~w9989 & w15863 ) | ( w15862 & w15863 ) ;
  assign w15865 = w8263 | w12217 ;
  assign w15866 = w9987 | w15864 ;
  assign w15867 = ( w35 & w15864 ) | ( w35 & w15866 ) | ( w15864 & w15866 ) ;
  assign w15868 = ( ~w12217 & w15865 ) | ( ~w12217 & w15867 ) | ( w15865 & w15867 ) ;
  assign w15869 = \pi05 ^ w15868 ;
  assign w15870 = w15481 ^ w15552 ;
  assign w15871 = w15473 ^ w15870 ;
  assign w15872 = w15489 ^ w15551 ;
  assign w15873 = w15491 ^ w15872 ;
  assign w15874 = w35 & ~w9989 ;
  assign w15875 = ( w8593 & w9991 ) | ( w8593 & w15874 ) | ( w9991 & w15874 ) ;
  assign w15876 = w8262 | w15875 ;
  assign w15877 = ( ~w9993 & w15875 ) | ( ~w9993 & w15876 ) | ( w15875 & w15876 ) ;
  assign w15878 = w15874 | w15877 ;
  assign w15879 = w8263 | w12484 ;
  assign w15880 = ( ~w12484 & w15878 ) | ( ~w12484 & w15879 ) | ( w15878 & w15879 ) ;
  assign w15881 = \pi05 ^ w15880 ;
  assign w15882 = w15501 ^ w15550 ;
  assign w15883 = w15493 ^ w15882 ;
  assign w15884 = w35 & w9991 ;
  assign w15885 = ( w8593 & ~w9993 ) | ( w8593 & w15884 ) | ( ~w9993 & w15884 ) ;
  assign w15886 = w8262 | w15885 ;
  assign w15887 = ( w9995 & w15885 ) | ( w9995 & w15886 ) | ( w15885 & w15886 ) ;
  assign w15888 = w15884 | w15887 ;
  assign w15889 = w8263 | w12514 ;
  assign w15890 = ( ~w12514 & w15888 ) | ( ~w12514 & w15889 ) | ( w15888 & w15889 ) ;
  assign w15891 = \pi05 ^ w15890 ;
  assign w15892 = w15509 ^ w15549 ;
  assign w15893 = w15510 ^ w15892 ;
  assign w15894 = w35 & ~w9993 ;
  assign w15895 = ( w8593 & w9995 ) | ( w8593 & w15894 ) | ( w9995 & w15894 ) ;
  assign w15896 = w8262 | w15895 ;
  assign w15897 = ( w9997 & w15895 ) | ( w9997 & w15896 ) | ( w15895 & w15896 ) ;
  assign w15898 = w15894 | w15897 ;
  assign w15899 = w8263 | w12541 ;
  assign w15900 = ( ~w12541 & w15898 ) | ( ~w12541 & w15899 ) | ( w15898 & w15899 ) ;
  assign w15901 = \pi05 ^ w15900 ;
  assign w15902 = ~w8593 & w9997 ;
  assign w15903 = w8262 & w9999 ;
  assign w15904 = ( w9997 & ~w15902 ) | ( w9997 & w15903 ) | ( ~w15902 & w15903 ) ;
  assign w15905 = ~w8263 & w12572 ;
  assign w15906 = w9995 | w15904 ;
  assign w15907 = ( w35 & w15904 ) | ( w35 & w15906 ) | ( w15904 & w15906 ) ;
  assign w15908 = ( w12572 & ~w15905 ) | ( w12572 & w15907 ) | ( ~w15905 & w15907 ) ;
  assign w15909 = \pi05 ^ w15908 ;
  assign w15910 = w15523 ^ w15548 ;
  assign w15911 = w15515 ^ w15910 ;
  assign w15912 = w15538 ^ w15546 ;
  assign w15913 = w15547 ^ w15912 ;
  assign w15914 = w35 & w9997 ;
  assign w15915 = ( w8593 & w9999 ) | ( w8593 & w15914 ) | ( w9999 & w15914 ) ;
  assign w15916 = w8262 | w15915 ;
  assign w15917 = ( w10001 & w15915 ) | ( w10001 & w15916 ) | ( w15915 & w15916 ) ;
  assign w15918 = w15914 | w15917 ;
  assign w15919 = ~w8263 & w12641 ;
  assign w15920 = ( w12641 & w15918 ) | ( w12641 & ~w15919 ) | ( w15918 & ~w15919 ) ;
  assign w15921 = \pi05 ^ w15920 ;
  assign w15922 = ~w8593 & w10001 ;
  assign w15923 = w8262 & ~w10006 ;
  assign w15924 = ( w10001 & ~w15922 ) | ( w10001 & w15923 ) | ( ~w15922 & w15923 ) ;
  assign w15925 = w8263 | w12691 ;
  assign w15926 = w9999 | w15924 ;
  assign w15927 = ( w35 & w15924 ) | ( w35 & w15926 ) | ( w15924 & w15926 ) ;
  assign w15928 = ( ~w12691 & w15925 ) | ( ~w12691 & w15927 ) | ( w15925 & w15927 ) ;
  assign w15929 = \pi05 ^ w15928 ;
  assign w15930 = w15529 ^ w15537 ;
  assign w15931 = ( \pi05 & \pi06 ) | ( \pi05 & ~w10016 ) | ( \pi06 & ~w10016 ) ;
  assign w15932 = ( \pi05 & \pi06 ) | ( \pi05 & ~w10021 ) | ( \pi06 & ~w10021 ) ;
  assign w15933 = \pi07 ^ w10021 ;
  assign w15934 = ( \pi07 & w15932 ) | ( \pi07 & w15933 ) | ( w15932 & w15933 ) ;
  assign w15935 = w15931 ^ w15934 ;
  assign w15936 = w35 & w10001 ;
  assign w15937 = ( w8593 & ~w10006 ) | ( w8593 & w15936 ) | ( ~w10006 & w15936 ) ;
  assign w15938 = w8262 | w15937 ;
  assign w15939 = ( w10011 & w15937 ) | ( w10011 & w15938 ) | ( w15937 & w15938 ) ;
  assign w15940 = w15936 | w15939 ;
  assign w15941 = ~w8263 & w12747 ;
  assign w15942 = ( w12747 & w15940 ) | ( w12747 & ~w15941 ) | ( w15940 & ~w15941 ) ;
  assign w15943 = \pi05 ^ w15942 ;
  assign w15944 = w10016 ^ w10021 ;
  assign w15945 = ( w8593 & ~w10016 ) | ( w8593 & w15944 ) | ( ~w10016 & w15944 ) ;
  assign w15946 = ( ~w8263 & w10016 ) | ( ~w8263 & w10021 ) | ( w10016 & w10021 ) ;
  assign w15947 = w35 | w10016 ;
  assign w15948 = ( w15945 & ~w15946 ) | ( w15945 & w15947 ) | ( ~w15946 & w15947 ) ;
  assign w15949 = w34 & ~w10021 ;
  assign w15950 = ( \pi05 & ~w15948 ) | ( \pi05 & w15949 ) | ( ~w15948 & w15949 ) ;
  assign w15951 = ~w15949 & w15950 ;
  assign w15952 = w35 & w10011 ;
  assign w15953 = ( w8593 & ~w10016 ) | ( w8593 & w15952 ) | ( ~w10016 & w15952 ) ;
  assign w15954 = w8262 | w15953 ;
  assign w15955 = ( ~w10021 & w15953 ) | ( ~w10021 & w15954 ) | ( w15953 & w15954 ) ;
  assign w15956 = w15952 | w15955 ;
  assign w15957 = ~w8263 & w12867 ;
  assign w15958 = ( w12867 & w15956 ) | ( w12867 & ~w15957 ) | ( w15956 & ~w15957 ) ;
  assign w15959 = \pi05 ^ w15958 ;
  assign w15960 = w15951 & w15959 ;
  assign w15961 = ~w8593 & w10011 ;
  assign w15962 = w8262 & ~w10016 ;
  assign w15963 = ( w10011 & ~w15961 ) | ( w10011 & w15962 ) | ( ~w15961 & w15962 ) ;
  assign w15964 = ~w8263 & w12777 ;
  assign w15965 = w10006 & ~w15963 ;
  assign w15966 = ( w35 & w15963 ) | ( w35 & ~w15965 ) | ( w15963 & ~w15965 ) ;
  assign w15967 = ( w12777 & ~w15964 ) | ( w12777 & w15966 ) | ( ~w15964 & w15966 ) ;
  assign w15968 = \pi05 ^ w15967 ;
  assign w15969 = w7413 & ~w10021 ;
  assign w15970 = ( w15960 & w15968 ) | ( w15960 & w15969 ) | ( w15968 & w15969 ) ;
  assign w15971 = ( w15935 & w15943 ) | ( w15935 & w15970 ) | ( w15943 & w15970 ) ;
  assign w15972 = ( w15929 & w15930 ) | ( w15929 & w15971 ) | ( w15930 & w15971 ) ;
  assign w15973 = ( w15913 & w15921 ) | ( w15913 & w15972 ) | ( w15921 & w15972 ) ;
  assign w15974 = ( w15909 & w15911 ) | ( w15909 & w15973 ) | ( w15911 & w15973 ) ;
  assign w15975 = ( w15893 & w15901 ) | ( w15893 & w15974 ) | ( w15901 & w15974 ) ;
  assign w15976 = ( w15883 & w15891 ) | ( w15883 & w15975 ) | ( w15891 & w15975 ) ;
  assign w15977 = ( w15873 & w15881 ) | ( w15873 & w15976 ) | ( w15881 & w15976 ) ;
  assign w15978 = ( w15869 & w15871 ) | ( w15869 & w15977 ) | ( w15871 & w15977 ) ;
  assign w15979 = ( w15859 & w15861 ) | ( w15859 & w15978 ) | ( w15861 & w15978 ) ;
  assign w15980 = ( w15849 & w15851 ) | ( w15849 & w15979 ) | ( w15851 & w15979 ) ;
  assign w15981 = ( w15833 & w15841 ) | ( w15833 & w15980 ) | ( w15841 & w15980 ) ;
  assign w15982 = ( w15823 & w15831 ) | ( w15823 & w15981 ) | ( w15831 & w15981 ) ;
  assign w15983 = ( w15813 & w15821 ) | ( w15813 & w15982 ) | ( w15821 & w15982 ) ;
  assign w15984 = ( w15809 & w15811 ) | ( w15809 & w15983 ) | ( w15811 & w15983 ) ;
  assign w15985 = ( w15799 & w15801 ) | ( w15799 & w15984 ) | ( w15801 & w15984 ) ;
  assign w15986 = ( w15789 & w15791 ) | ( w15789 & w15985 ) | ( w15791 & w15985 ) ;
  assign w15987 = ( w15773 & w15781 ) | ( w15773 & w15986 ) | ( w15781 & w15986 ) ;
  assign w15988 = ( w15763 & w15771 ) | ( w15763 & w15987 ) | ( w15771 & w15987 ) ;
  assign w15989 = ( w15753 & w15761 ) | ( w15753 & w15988 ) | ( w15761 & w15988 ) ;
  assign w15990 = ( w15749 & w15751 ) | ( w15749 & w15989 ) | ( w15751 & w15989 ) ;
  assign w15991 = ( w15739 & w15741 ) | ( w15739 & w15990 ) | ( w15741 & w15990 ) ;
  assign w15992 = ( w15729 & w15731 ) | ( w15729 & w15991 ) | ( w15731 & w15991 ) ;
  assign w15993 = ( w15713 & w15721 ) | ( w15713 & w15992 ) | ( w15721 & w15992 ) ;
  assign w15994 = ( w15703 & w15711 ) | ( w15703 & w15993 ) | ( w15711 & w15993 ) ;
  assign w15995 = ( w15699 & ~w15701 ) | ( w15699 & w15994 ) | ( ~w15701 & w15994 ) ;
  assign w15996 = ( w15689 & ~w15691 ) | ( w15689 & w15995 ) | ( ~w15691 & w15995 ) ;
  assign w15997 = ( w15679 & w15681 ) | ( w15679 & w15996 ) | ( w15681 & w15996 ) ;
  assign w15998 = ( w15669 & ~w15671 ) | ( w15669 & w15997 ) | ( ~w15671 & w15997 ) ;
  assign w15999 = ( w15659 & ~w15661 ) | ( w15659 & w15998 ) | ( ~w15661 & w15998 ) ;
  assign w16000 = ( w15649 & w15651 ) | ( w15649 & w15999 ) | ( w15651 & w15999 ) ;
  assign w16001 = ( w15639 & w15641 ) | ( w15639 & w16000 ) | ( w15641 & w16000 ) ;
  assign w16002 = ( w15629 & w15631 ) | ( w15629 & w16001 ) | ( w15631 & w16001 ) ;
  assign w16003 = ( w15619 & w15621 ) | ( w15619 & w16002 ) | ( w15621 & w16002 ) ;
  assign w16004 = w15619 ^ w16002 ;
  assign w16005 = w15621 ^ w16004 ;
  assign w16006 = \pi00 | \pi01 ;
  assign w16007 = w10431 & ~w16006 ;
  assign w16008 = w10736 ^ w16007 ;
  assign w16009 = ( ~w10402 & w10431 ) | ( ~w10402 & w10736 ) | ( w10431 & w10736 ) ;
  assign w16010 = w16008 & ~w16009 ;
  assign w16011 = ( \pi00 & \pi01 ) | ( \pi00 & ~\pi02 ) | ( \pi01 & ~\pi02 ) ;
  assign w16012 = ( \pi01 & w10431 ) | ( \pi01 & w10736 ) | ( w10431 & w10736 ) ;
  assign w16013 = ( \pi01 & w10736 ) | ( \pi01 & ~w16012 ) | ( w10736 & ~w16012 ) ;
  assign w16014 = ( w10402 & w10431 ) | ( w10402 & ~w16012 ) | ( w10431 & ~w16012 ) ;
  assign w16015 = w16013 | w16014 ;
  assign w16016 = ~\pi00 & w16015 ;
  assign w16017 = ( \pi02 & w16011 ) | ( \pi02 & w16016 ) | ( w16011 & w16016 ) ;
  assign w16018 = ~\pi01 & w16011 ;
  assign w16019 = ( ~w16010 & w16017 ) | ( ~w16010 & w16018 ) | ( w16017 & w16018 ) ;
  assign w16020 = w15629 ^ w16001 ;
  assign w16021 = w15631 ^ w16020 ;
  assign w16022 = ( \pi02 & ~w10883 ) | ( \pi02 & w11139 ) | ( ~w10883 & w11139 ) ;
  assign w16023 = \pi00 ^ w16022 ;
  assign w16024 = ( \pi02 & ~w11139 ) | ( \pi02 & w16023 ) | ( ~w11139 & w16023 ) ;
  assign w16025 = ( \pi02 & w10883 ) | ( \pi02 & ~w16023 ) | ( w10883 & ~w16023 ) ;
  assign w16026 = \pi01 & w16025 ;
  assign w16027 = ( \pi00 & w10887 ) | ( \pi00 & ~w16026 ) | ( w10887 & ~w16026 ) ;
  assign w16028 = ( \pi01 & \pi02 ) | ( \pi01 & w16027 ) | ( \pi02 & w16027 ) ;
  assign w16029 = ( w16024 & w16026 ) | ( w16024 & ~w16028 ) | ( w16026 & ~w16028 ) ;
  assign w16030 = w15639 ^ w16000 ;
  assign w16031 = w15641 ^ w16030 ;
  assign w16032 = ( \pi02 & ~w10883 ) | ( \pi02 & w10887 ) | ( ~w10883 & w10887 ) ;
  assign w16033 = \pi00 ^ w16032 ;
  assign w16034 = ( \pi02 & w10883 ) | ( \pi02 & w16033 ) | ( w10883 & w16033 ) ;
  assign w16035 = ( ~\pi02 & w10887 ) | ( ~\pi02 & w16033 ) | ( w10887 & w16033 ) ;
  assign w16036 = \pi01 & ~w16035 ;
  assign w16037 = ( \pi00 & w10885 ) | ( \pi00 & ~w16036 ) | ( w10885 & ~w16036 ) ;
  assign w16038 = ( \pi01 & \pi02 ) | ( \pi01 & w16037 ) | ( \pi02 & w16037 ) ;
  assign w16039 = ( w16034 & w16036 ) | ( w16034 & ~w16038 ) | ( w16036 & ~w16038 ) ;
  assign w16040 = w15649 ^ w15999 ;
  assign w16041 = w15651 ^ w16040 ;
  assign w16042 = ( \pi02 & w10885 ) | ( \pi02 & w10887 ) | ( w10885 & w10887 ) ;
  assign w16043 = \pi00 ^ w16042 ;
  assign w16044 = ( \pi02 & ~w10887 ) | ( \pi02 & w16043 ) | ( ~w10887 & w16043 ) ;
  assign w16045 = ( ~\pi02 & w10885 ) | ( ~\pi02 & w16043 ) | ( w10885 & w16043 ) ;
  assign w16046 = \pi01 & ~w16045 ;
  assign w16047 = ( \pi00 & w10866 ) | ( \pi00 & ~w16046 ) | ( w10866 & ~w16046 ) ;
  assign w16048 = ( \pi01 & \pi02 ) | ( \pi01 & w16047 ) | ( \pi02 & w16047 ) ;
  assign w16049 = ( w16044 & w16046 ) | ( w16044 & ~w16048 ) | ( w16046 & ~w16048 ) ;
  assign w16050 = w15659 ^ w15998 ;
  assign w16051 = w15661 ^ w16050 ;
  assign w16052 = ( \pi02 & w10866 ) | ( \pi02 & w10885 ) | ( w10866 & w10885 ) ;
  assign w16053 = \pi00 ^ w16052 ;
  assign w16054 = ( \pi02 & ~w10885 ) | ( \pi02 & w16053 ) | ( ~w10885 & w16053 ) ;
  assign w16055 = ( ~\pi02 & w10866 ) | ( ~\pi02 & w16053 ) | ( w10866 & w16053 ) ;
  assign w16056 = \pi01 & ~w16055 ;
  assign w16057 = ( ~\pi00 & w10801 ) | ( ~\pi00 & w16056 ) | ( w10801 & w16056 ) ;
  assign w16058 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16057 ) | ( \pi02 & ~w16057 ) ;
  assign w16059 = ( w16054 & w16056 ) | ( w16054 & ~w16058 ) | ( w16056 & ~w16058 ) ;
  assign w16060 = w15669 ^ w15997 ;
  assign w16061 = w15671 ^ w16060 ;
  assign w16062 = ( \pi02 & ~w10801 ) | ( \pi02 & w10866 ) | ( ~w10801 & w10866 ) ;
  assign w16063 = \pi00 ^ w16062 ;
  assign w16064 = ( \pi02 & ~w10866 ) | ( \pi02 & w16063 ) | ( ~w10866 & w16063 ) ;
  assign w16065 = ( \pi02 & w10801 ) | ( \pi02 & ~w16063 ) | ( w10801 & ~w16063 ) ;
  assign w16066 = \pi01 & w16065 ;
  assign w16067 = ( \pi00 & w10807 ) | ( \pi00 & ~w16066 ) | ( w10807 & ~w16066 ) ;
  assign w16068 = ( \pi01 & \pi02 ) | ( \pi01 & w16067 ) | ( \pi02 & w16067 ) ;
  assign w16069 = ( w16064 & w16066 ) | ( w16064 & ~w16068 ) | ( w16066 & ~w16068 ) ;
  assign w16070 = ~w8954 & w10874 ;
  assign w16071 = ( w10874 & w16069 ) | ( w10874 & ~w16070 ) | ( w16069 & ~w16070 ) ;
  assign w16072 = \pi02 ^ w16071 ;
  assign w16073 = w15679 ^ w15996 ;
  assign w16074 = w15681 ^ w16073 ;
  assign w16075 = ( \pi02 & ~w10801 ) | ( \pi02 & w10807 ) | ( ~w10801 & w10807 ) ;
  assign w16076 = \pi00 ^ w16075 ;
  assign w16077 = ( \pi02 & w10801 ) | ( \pi02 & w16076 ) | ( w10801 & w16076 ) ;
  assign w16078 = ( ~\pi02 & w10807 ) | ( ~\pi02 & w16076 ) | ( w10807 & w16076 ) ;
  assign w16079 = \pi01 & ~w16078 ;
  assign w16080 = ( \pi00 & w10805 ) | ( \pi00 & ~w16079 ) | ( w10805 & ~w16079 ) ;
  assign w16081 = ( \pi01 & \pi02 ) | ( \pi01 & w16080 ) | ( \pi02 & w16080 ) ;
  assign w16082 = ( w16077 & w16079 ) | ( w16077 & ~w16081 ) | ( w16079 & ~w16081 ) ;
  assign w16083 = ~w8954 & w10814 ;
  assign w16084 = ( w10814 & w16082 ) | ( w10814 & ~w16083 ) | ( w16082 & ~w16083 ) ;
  assign w16085 = \pi02 ^ w16084 ;
  assign w16086 = w15689 ^ w15995 ;
  assign w16087 = w15691 ^ w16086 ;
  assign w16088 = ( \pi02 & w10805 ) | ( \pi02 & w10807 ) | ( w10805 & w10807 ) ;
  assign w16089 = \pi00 ^ w16088 ;
  assign w16090 = ( \pi02 & ~w10807 ) | ( \pi02 & w16089 ) | ( ~w10807 & w16089 ) ;
  assign w16091 = ( ~\pi02 & w10805 ) | ( ~\pi02 & w16089 ) | ( w10805 & w16089 ) ;
  assign w16092 = \pi01 & ~w16091 ;
  assign w16093 = ( ~\pi00 & w10784 ) | ( ~\pi00 & w16092 ) | ( w10784 & w16092 ) ;
  assign w16094 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16093 ) | ( \pi02 & ~w16093 ) ;
  assign w16095 = ( w16090 & w16092 ) | ( w16090 & ~w16094 ) | ( w16092 & ~w16094 ) ;
  assign w16096 = ~w8954 & w11117 ;
  assign w16097 = ( w11117 & w16095 ) | ( w11117 & ~w16096 ) | ( w16095 & ~w16096 ) ;
  assign w16098 = \pi02 ^ w16097 ;
  assign w16099 = w15699 ^ w15994 ;
  assign w16100 = w15701 ^ w16099 ;
  assign w16101 = ( \pi02 & ~w10784 ) | ( \pi02 & w10805 ) | ( ~w10784 & w10805 ) ;
  assign w16102 = \pi00 ^ w16101 ;
  assign w16103 = ( \pi02 & ~w10805 ) | ( \pi02 & w16102 ) | ( ~w10805 & w16102 ) ;
  assign w16104 = ( \pi02 & w10784 ) | ( \pi02 & ~w16102 ) | ( w10784 & ~w16102 ) ;
  assign w16105 = \pi01 & w16104 ;
  assign w16106 = ( ~\pi00 & w10211 ) | ( ~\pi00 & w16105 ) | ( w10211 & w16105 ) ;
  assign w16107 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16106 ) | ( \pi02 & ~w16106 ) ;
  assign w16108 = ( w16103 & w16105 ) | ( w16103 & ~w16107 ) | ( w16105 & ~w16107 ) ;
  assign w16109 = w8954 | w10855 ;
  assign w16110 = ( ~w10855 & w16108 ) | ( ~w10855 & w16109 ) | ( w16108 & w16109 ) ;
  assign w16111 = \pi02 ^ w16110 ;
  assign w16112 = \pi00 ^ w10011 ;
  assign w16113 = ( \pi01 & w10011 ) | ( \pi01 & ~w16112 ) | ( w10011 & ~w16112 ) ;
  assign w16114 = ( \pi00 & ~w10016 ) | ( \pi00 & w16113 ) | ( ~w10016 & w16113 ) ;
  assign w16115 = ( \pi02 & ~w10021 ) | ( \pi02 & w16114 ) | ( ~w10021 & w16114 ) ;
  assign w16116 = \pi02 & ~w16115 ;
  assign w16117 = ( \pi02 & w10006 ) | ( \pi02 & ~w10011 ) | ( w10006 & ~w10011 ) ;
  assign w16118 = \pi00 ^ w16117 ;
  assign w16119 = ( \pi02 & ~w10006 ) | ( \pi02 & w16118 ) | ( ~w10006 & w16118 ) ;
  assign w16120 = ( \pi02 & w10011 ) | ( \pi02 & ~w16118 ) | ( w10011 & ~w16118 ) ;
  assign w16121 = \pi01 & w16120 ;
  assign w16122 = ( \pi00 & w10016 ) | ( \pi00 & ~w16121 ) | ( w10016 & ~w16121 ) ;
  assign w16123 = ( \pi01 & \pi02 ) | ( \pi01 & w16122 ) | ( \pi02 & w16122 ) ;
  assign w16124 = ( w16119 & w16121 ) | ( w16119 & ~w16123 ) | ( w16121 & ~w16123 ) ;
  assign w16125 = w12777 | w16124 ;
  assign w16126 = ( w8954 & w16124 ) | ( w8954 & w16125 ) | ( w16124 & w16125 ) ;
  assign w16127 = \pi02 ^ w16126 ;
  assign w16128 = ( w15949 & w16116 ) | ( w15949 & w16127 ) | ( w16116 & w16127 ) ;
  assign w16129 = ( \pi02 & ~w10001 ) | ( \pi02 & w10006 ) | ( ~w10001 & w10006 ) ;
  assign w16130 = \pi00 ^ w16129 ;
  assign w16131 = ( \pi02 & w10001 ) | ( \pi02 & w16130 ) | ( w10001 & w16130 ) ;
  assign w16132 = ( ~\pi02 & w10006 ) | ( ~\pi02 & w16130 ) | ( w10006 & w16130 ) ;
  assign w16133 = \pi01 & ~w16132 ;
  assign w16134 = ( ~\pi00 & w10011 ) | ( ~\pi00 & w16133 ) | ( w10011 & w16133 ) ;
  assign w16135 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16134 ) | ( \pi02 & ~w16134 ) ;
  assign w16136 = ( w16131 & w16133 ) | ( w16131 & ~w16135 ) | ( w16133 & ~w16135 ) ;
  assign w16137 = ~w8954 & w12747 ;
  assign w16138 = ( w12747 & w16136 ) | ( w12747 & ~w16137 ) | ( w16136 & ~w16137 ) ;
  assign w16139 = \pi02 ^ w16138 ;
  assign w16140 = \pi05 & w15949 ;
  assign w16141 = w15948 ^ w16140 ;
  assign w16142 = ( w16128 & w16139 ) | ( w16128 & w16141 ) | ( w16139 & w16141 ) ;
  assign w16143 = ( ~\pi02 & w9999 ) | ( ~\pi02 & w10001 ) | ( w9999 & w10001 ) ;
  assign w16144 = \pi00 ^ w16143 ;
  assign w16145 = ( \pi02 & w9999 ) | ( \pi02 & ~w16144 ) | ( w9999 & ~w16144 ) ;
  assign w16146 = ( \pi02 & w10001 ) | ( \pi02 & w16144 ) | ( w10001 & w16144 ) ;
  assign w16147 = \pi01 & w16146 ;
  assign w16148 = ( \pi00 & w10006 ) | ( \pi00 & ~w16147 ) | ( w10006 & ~w16147 ) ;
  assign w16149 = ( \pi01 & \pi02 ) | ( \pi01 & w16148 ) | ( \pi02 & w16148 ) ;
  assign w16150 = ( w16145 & w16147 ) | ( w16145 & ~w16149 ) | ( w16147 & ~w16149 ) ;
  assign w16151 = w8954 | w12691 ;
  assign w16152 = ( ~w12691 & w16150 ) | ( ~w12691 & w16151 ) | ( w16150 & w16151 ) ;
  assign w16153 = \pi02 ^ w16152 ;
  assign w16154 = w15951 ^ w15959 ;
  assign w16155 = ( w16142 & w16153 ) | ( w16142 & w16154 ) | ( w16153 & w16154 ) ;
  assign w16156 = ( ~\pi02 & w9997 ) | ( ~\pi02 & w9999 ) | ( w9997 & w9999 ) ;
  assign w16157 = \pi00 ^ w16156 ;
  assign w16158 = ( \pi02 & w9997 ) | ( \pi02 & ~w16157 ) | ( w9997 & ~w16157 ) ;
  assign w16159 = ( \pi02 & w9999 ) | ( \pi02 & w16157 ) | ( w9999 & w16157 ) ;
  assign w16160 = \pi01 & w16159 ;
  assign w16161 = ( ~\pi00 & w10001 ) | ( ~\pi00 & w16160 ) | ( w10001 & w16160 ) ;
  assign w16162 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16161 ) | ( \pi02 & ~w16161 ) ;
  assign w16163 = ( w16158 & w16160 ) | ( w16158 & ~w16162 ) | ( w16160 & ~w16162 ) ;
  assign w16164 = w15960 ^ w15968 ;
  assign w16165 = w15969 ^ w16164 ;
  assign w16166 = w12641 | w16163 ;
  assign w16167 = ( w8954 & w16163 ) | ( w8954 & w16166 ) | ( w16163 & w16166 ) ;
  assign w16168 = \pi02 ^ w16167 ;
  assign w16169 = ( w16155 & w16165 ) | ( w16155 & w16168 ) | ( w16165 & w16168 ) ;
  assign w16170 = ( ~\pi02 & w9995 ) | ( ~\pi02 & w9997 ) | ( w9995 & w9997 ) ;
  assign w16171 = \pi00 ^ w16170 ;
  assign w16172 = ( \pi02 & w9995 ) | ( \pi02 & ~w16171 ) | ( w9995 & ~w16171 ) ;
  assign w16173 = ( \pi02 & w9997 ) | ( \pi02 & w16171 ) | ( w9997 & w16171 ) ;
  assign w16174 = \pi01 & w16173 ;
  assign w16175 = ( ~\pi00 & w9999 ) | ( ~\pi00 & w16174 ) | ( w9999 & w16174 ) ;
  assign w16176 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16175 ) | ( \pi02 & ~w16175 ) ;
  assign w16177 = ( w16172 & w16174 ) | ( w16172 & ~w16176 ) | ( w16174 & ~w16176 ) ;
  assign w16178 = ~w8954 & w12572 ;
  assign w16179 = ( w12572 & w16177 ) | ( w12572 & ~w16178 ) | ( w16177 & ~w16178 ) ;
  assign w16180 = \pi02 ^ w16179 ;
  assign w16181 = w15943 ^ w15970 ;
  assign w16182 = w15935 ^ w16181 ;
  assign w16183 = ( w16169 & w16180 ) | ( w16169 & w16182 ) | ( w16180 & w16182 ) ;
  assign w16184 = ( \pi02 & w9993 ) | ( \pi02 & ~w9995 ) | ( w9993 & ~w9995 ) ;
  assign w16185 = \pi00 ^ w16184 ;
  assign w16186 = ( \pi02 & ~w9993 ) | ( \pi02 & w16185 ) | ( ~w9993 & w16185 ) ;
  assign w16187 = ( \pi02 & w9995 ) | ( \pi02 & ~w16185 ) | ( w9995 & ~w16185 ) ;
  assign w16188 = \pi01 & w16187 ;
  assign w16189 = ( ~\pi00 & w9997 ) | ( ~\pi00 & w16188 ) | ( w9997 & w16188 ) ;
  assign w16190 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16189 ) | ( \pi02 & ~w16189 ) ;
  assign w16191 = ( w16186 & w16188 ) | ( w16186 & ~w16190 ) | ( w16188 & ~w16190 ) ;
  assign w16192 = w8954 | w12541 ;
  assign w16193 = ( ~w12541 & w16191 ) | ( ~w12541 & w16192 ) | ( w16191 & w16192 ) ;
  assign w16194 = \pi02 ^ w16193 ;
  assign w16195 = w15929 ^ w15971 ;
  assign w16196 = w15930 ^ w16195 ;
  assign w16197 = ( w16183 & w16194 ) | ( w16183 & w16196 ) | ( w16194 & w16196 ) ;
  assign w16198 = ( \pi02 & ~w9991 ) | ( \pi02 & w9993 ) | ( ~w9991 & w9993 ) ;
  assign w16199 = \pi00 ^ w16198 ;
  assign w16200 = ( \pi02 & w9991 ) | ( \pi02 & w16199 ) | ( w9991 & w16199 ) ;
  assign w16201 = ( ~\pi02 & w9993 ) | ( ~\pi02 & w16199 ) | ( w9993 & w16199 ) ;
  assign w16202 = \pi01 & ~w16201 ;
  assign w16203 = ( ~\pi00 & w9995 ) | ( ~\pi00 & w16202 ) | ( w9995 & w16202 ) ;
  assign w16204 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16203 ) | ( \pi02 & ~w16203 ) ;
  assign w16205 = ( w16200 & w16202 ) | ( w16200 & ~w16204 ) | ( w16202 & ~w16204 ) ;
  assign w16206 = w8954 | w12514 ;
  assign w16207 = ( ~w12514 & w16205 ) | ( ~w12514 & w16206 ) | ( w16205 & w16206 ) ;
  assign w16208 = \pi02 ^ w16207 ;
  assign w16209 = w15921 ^ w15972 ;
  assign w16210 = w15913 ^ w16209 ;
  assign w16211 = ( w16197 & w16208 ) | ( w16197 & w16210 ) | ( w16208 & w16210 ) ;
  assign w16212 = ( \pi02 & w9989 ) | ( \pi02 & ~w9991 ) | ( w9989 & ~w9991 ) ;
  assign w16213 = \pi00 ^ w16212 ;
  assign w16214 = ( \pi02 & ~w9989 ) | ( \pi02 & w16213 ) | ( ~w9989 & w16213 ) ;
  assign w16215 = ( \pi02 & w9991 ) | ( \pi02 & ~w16213 ) | ( w9991 & ~w16213 ) ;
  assign w16216 = \pi01 & w16215 ;
  assign w16217 = ( \pi00 & w9993 ) | ( \pi00 & ~w16216 ) | ( w9993 & ~w16216 ) ;
  assign w16218 = ( \pi01 & \pi02 ) | ( \pi01 & w16217 ) | ( \pi02 & w16217 ) ;
  assign w16219 = ( w16214 & w16216 ) | ( w16214 & ~w16218 ) | ( w16216 & ~w16218 ) ;
  assign w16220 = w8954 | w12484 ;
  assign w16221 = ( ~w12484 & w16219 ) | ( ~w12484 & w16220 ) | ( w16219 & w16220 ) ;
  assign w16222 = \pi02 ^ w16221 ;
  assign w16223 = w15909 ^ w15973 ;
  assign w16224 = w15911 ^ w16223 ;
  assign w16225 = ( w16211 & w16222 ) | ( w16211 & w16224 ) | ( w16222 & w16224 ) ;
  assign w16226 = ( \pi02 & ~w9987 ) | ( \pi02 & w9989 ) | ( ~w9987 & w9989 ) ;
  assign w16227 = \pi00 ^ w16226 ;
  assign w16228 = ( \pi02 & w9987 ) | ( \pi02 & w16227 ) | ( w9987 & w16227 ) ;
  assign w16229 = ( ~\pi02 & w9989 ) | ( ~\pi02 & w16227 ) | ( w9989 & w16227 ) ;
  assign w16230 = \pi01 & ~w16229 ;
  assign w16231 = ( ~\pi00 & w9991 ) | ( ~\pi00 & w16230 ) | ( w9991 & w16230 ) ;
  assign w16232 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16231 ) | ( \pi02 & ~w16231 ) ;
  assign w16233 = ( w16228 & w16230 ) | ( w16228 & ~w16232 ) | ( w16230 & ~w16232 ) ;
  assign w16234 = w8954 | w12217 ;
  assign w16235 = ( ~w12217 & w16233 ) | ( ~w12217 & w16234 ) | ( w16233 & w16234 ) ;
  assign w16236 = \pi02 ^ w16235 ;
  assign w16237 = w15901 ^ w15974 ;
  assign w16238 = w15893 ^ w16237 ;
  assign w16239 = ( w16225 & w16236 ) | ( w16225 & w16238 ) | ( w16236 & w16238 ) ;
  assign w16240 = ( ~\pi02 & w9985 ) | ( ~\pi02 & w9987 ) | ( w9985 & w9987 ) ;
  assign w16241 = \pi00 ^ w16240 ;
  assign w16242 = ( \pi02 & w9985 ) | ( \pi02 & ~w16241 ) | ( w9985 & ~w16241 ) ;
  assign w16243 = ( \pi02 & w9987 ) | ( \pi02 & w16241 ) | ( w9987 & w16241 ) ;
  assign w16244 = \pi01 & w16243 ;
  assign w16245 = ( \pi00 & w9989 ) | ( \pi00 & ~w16244 ) | ( w9989 & ~w16244 ) ;
  assign w16246 = ( \pi01 & \pi02 ) | ( \pi01 & w16245 ) | ( \pi02 & w16245 ) ;
  assign w16247 = ( w16242 & w16244 ) | ( w16242 & ~w16246 ) | ( w16244 & ~w16246 ) ;
  assign w16248 = ~w8954 & w12446 ;
  assign w16249 = ( w12446 & w16247 ) | ( w12446 & ~w16248 ) | ( w16247 & ~w16248 ) ;
  assign w16250 = \pi02 ^ w16249 ;
  assign w16251 = w15891 ^ w15975 ;
  assign w16252 = w15883 ^ w16251 ;
  assign w16253 = ( w16239 & w16250 ) | ( w16239 & w16252 ) | ( w16250 & w16252 ) ;
  assign w16254 = ( ~\pi02 & w9983 ) | ( ~\pi02 & w9985 ) | ( w9983 & w9985 ) ;
  assign w16255 = \pi00 ^ w16254 ;
  assign w16256 = ( \pi02 & w9983 ) | ( \pi02 & ~w16255 ) | ( w9983 & ~w16255 ) ;
  assign w16257 = ( \pi02 & w9985 ) | ( \pi02 & w16255 ) | ( w9985 & w16255 ) ;
  assign w16258 = \pi01 & w16257 ;
  assign w16259 = ( ~\pi00 & w9987 ) | ( ~\pi00 & w16258 ) | ( w9987 & w16258 ) ;
  assign w16260 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16259 ) | ( \pi02 & ~w16259 ) ;
  assign w16261 = ( w16256 & w16258 ) | ( w16256 & ~w16260 ) | ( w16258 & ~w16260 ) ;
  assign w16262 = ~w8954 & w12433 ;
  assign w16263 = ( w12433 & w16261 ) | ( w12433 & ~w16262 ) | ( w16261 & ~w16262 ) ;
  assign w16264 = \pi02 ^ w16263 ;
  assign w16265 = w15881 ^ w15976 ;
  assign w16266 = w15873 ^ w16265 ;
  assign w16267 = ( w16253 & w16264 ) | ( w16253 & w16266 ) | ( w16264 & w16266 ) ;
  assign w16268 = ( ~\pi02 & w9981 ) | ( ~\pi02 & w9983 ) | ( w9981 & w9983 ) ;
  assign w16269 = \pi00 ^ w16268 ;
  assign w16270 = ( \pi02 & w9981 ) | ( \pi02 & ~w16269 ) | ( w9981 & ~w16269 ) ;
  assign w16271 = ( \pi02 & w9983 ) | ( \pi02 & w16269 ) | ( w9983 & w16269 ) ;
  assign w16272 = \pi01 & w16271 ;
  assign w16273 = ( ~\pi00 & w9985 ) | ( ~\pi00 & w16272 ) | ( w9985 & w16272 ) ;
  assign w16274 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16273 ) | ( \pi02 & ~w16273 ) ;
  assign w16275 = ( w16270 & w16272 ) | ( w16270 & ~w16274 ) | ( w16272 & ~w16274 ) ;
  assign w16276 = ~w8954 & w12236 ;
  assign w16277 = ( w12236 & w16275 ) | ( w12236 & ~w16276 ) | ( w16275 & ~w16276 ) ;
  assign w16278 = \pi02 ^ w16277 ;
  assign w16279 = w15869 ^ w15977 ;
  assign w16280 = w15871 ^ w16279 ;
  assign w16281 = ( w16267 & w16278 ) | ( w16267 & w16280 ) | ( w16278 & w16280 ) ;
  assign w16282 = ( ~\pi02 & w9979 ) | ( ~\pi02 & w9981 ) | ( w9979 & w9981 ) ;
  assign w16283 = \pi00 ^ w16282 ;
  assign w16284 = ( \pi02 & w9979 ) | ( \pi02 & ~w16283 ) | ( w9979 & ~w16283 ) ;
  assign w16285 = ( \pi02 & w9981 ) | ( \pi02 & w16283 ) | ( w9981 & w16283 ) ;
  assign w16286 = \pi01 & w16285 ;
  assign w16287 = ( ~\pi00 & w9983 ) | ( ~\pi00 & w16286 ) | ( w9983 & w16286 ) ;
  assign w16288 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16287 ) | ( \pi02 & ~w16287 ) ;
  assign w16289 = ( w16284 & w16286 ) | ( w16284 & ~w16288 ) | ( w16286 & ~w16288 ) ;
  assign w16290 = ~w8954 & w12010 ;
  assign w16291 = ( w12010 & w16289 ) | ( w12010 & ~w16290 ) | ( w16289 & ~w16290 ) ;
  assign w16292 = \pi02 ^ w16291 ;
  assign w16293 = w15859 ^ w15978 ;
  assign w16294 = w15861 ^ w16293 ;
  assign w16295 = ( w16281 & w16292 ) | ( w16281 & w16294 ) | ( w16292 & w16294 ) ;
  assign w16296 = ( ~\pi02 & w9977 ) | ( ~\pi02 & w9979 ) | ( w9977 & w9979 ) ;
  assign w16297 = \pi00 ^ w16296 ;
  assign w16298 = ( \pi02 & w9977 ) | ( \pi02 & ~w16297 ) | ( w9977 & ~w16297 ) ;
  assign w16299 = ( \pi02 & w9979 ) | ( \pi02 & w16297 ) | ( w9979 & w16297 ) ;
  assign w16300 = \pi01 & w16299 ;
  assign w16301 = ( ~\pi00 & w9981 ) | ( ~\pi00 & w16300 ) | ( w9981 & w16300 ) ;
  assign w16302 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16301 ) | ( \pi02 & ~w16301 ) ;
  assign w16303 = ( w16298 & w16300 ) | ( w16298 & ~w16302 ) | ( w16300 & ~w16302 ) ;
  assign w16304 = ~w8954 & w12106 ;
  assign w16305 = ( w12106 & w16303 ) | ( w12106 & ~w16304 ) | ( w16303 & ~w16304 ) ;
  assign w16306 = \pi02 ^ w16305 ;
  assign w16307 = w15849 ^ w15979 ;
  assign w16308 = w15851 ^ w16307 ;
  assign w16309 = ( w16295 & w16306 ) | ( w16295 & w16308 ) | ( w16306 & w16308 ) ;
  assign w16310 = ( ~\pi02 & w9975 ) | ( ~\pi02 & w9977 ) | ( w9975 & w9977 ) ;
  assign w16311 = \pi00 ^ w16310 ;
  assign w16312 = ( \pi02 & w9975 ) | ( \pi02 & ~w16311 ) | ( w9975 & ~w16311 ) ;
  assign w16313 = ( \pi02 & w9977 ) | ( \pi02 & w16311 ) | ( w9977 & w16311 ) ;
  assign w16314 = \pi01 & w16313 ;
  assign w16315 = ( ~\pi00 & w9979 ) | ( ~\pi00 & w16314 ) | ( w9979 & w16314 ) ;
  assign w16316 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16315 ) | ( \pi02 & ~w16315 ) ;
  assign w16317 = ( w16312 & w16314 ) | ( w16312 & ~w16316 ) | ( w16314 & ~w16316 ) ;
  assign w16318 = ~w8954 & w11914 ;
  assign w16319 = ( w11914 & w16317 ) | ( w11914 & ~w16318 ) | ( w16317 & ~w16318 ) ;
  assign w16320 = \pi02 ^ w16319 ;
  assign w16321 = w15841 ^ w15980 ;
  assign w16322 = w15833 ^ w16321 ;
  assign w16323 = ( w16309 & w16320 ) | ( w16309 & w16322 ) | ( w16320 & w16322 ) ;
  assign w16324 = ( \pi02 & w9973 ) | ( \pi02 & ~w9975 ) | ( w9973 & ~w9975 ) ;
  assign w16325 = \pi00 ^ w16324 ;
  assign w16326 = ( \pi02 & ~w9973 ) | ( \pi02 & w16325 ) | ( ~w9973 & w16325 ) ;
  assign w16327 = ( \pi02 & w9975 ) | ( \pi02 & ~w16325 ) | ( w9975 & ~w16325 ) ;
  assign w16328 = \pi01 & w16327 ;
  assign w16329 = ( ~\pi00 & w9977 ) | ( ~\pi00 & w16328 ) | ( w9977 & w16328 ) ;
  assign w16330 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16329 ) | ( \pi02 & ~w16329 ) ;
  assign w16331 = ( w16326 & w16328 ) | ( w16326 & ~w16330 ) | ( w16328 & ~w16330 ) ;
  assign w16332 = w8954 | w11671 ;
  assign w16333 = ( ~w11671 & w16331 ) | ( ~w11671 & w16332 ) | ( w16331 & w16332 ) ;
  assign w16334 = \pi02 ^ w16333 ;
  assign w16335 = w15831 ^ w15981 ;
  assign w16336 = w15823 ^ w16335 ;
  assign w16337 = ( w16323 & w16334 ) | ( w16323 & w16336 ) | ( w16334 & w16336 ) ;
  assign w16338 = ( \pi02 & ~w9971 ) | ( \pi02 & w9973 ) | ( ~w9971 & w9973 ) ;
  assign w16339 = \pi00 ^ w16338 ;
  assign w16340 = ( \pi02 & w9971 ) | ( \pi02 & w16339 ) | ( w9971 & w16339 ) ;
  assign w16341 = ( ~\pi02 & w9973 ) | ( ~\pi02 & w16339 ) | ( w9973 & w16339 ) ;
  assign w16342 = \pi01 & ~w16341 ;
  assign w16343 = ( ~\pi00 & w9975 ) | ( ~\pi00 & w16342 ) | ( w9975 & w16342 ) ;
  assign w16344 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16343 ) | ( \pi02 & ~w16343 ) ;
  assign w16345 = ( w16340 & w16342 ) | ( w16340 & ~w16344 ) | ( w16342 & ~w16344 ) ;
  assign w16346 = w8954 | w11809 ;
  assign w16347 = ( ~w11809 & w16345 ) | ( ~w11809 & w16346 ) | ( w16345 & w16346 ) ;
  assign w16348 = \pi02 ^ w16347 ;
  assign w16349 = w15821 ^ w15982 ;
  assign w16350 = w15813 ^ w16349 ;
  assign w16351 = ( w16337 & w16348 ) | ( w16337 & w16350 ) | ( w16348 & w16350 ) ;
  assign w16352 = ( \pi02 & w9967 ) | ( \pi02 & ~w9971 ) | ( w9967 & ~w9971 ) ;
  assign w16353 = \pi00 ^ w16352 ;
  assign w16354 = ( \pi02 & ~w9967 ) | ( \pi02 & w16353 ) | ( ~w9967 & w16353 ) ;
  assign w16355 = ( \pi02 & w9971 ) | ( \pi02 & ~w16353 ) | ( w9971 & ~w16353 ) ;
  assign w16356 = \pi01 & w16355 ;
  assign w16357 = ( \pi00 & w9973 ) | ( \pi00 & ~w16356 ) | ( w9973 & ~w16356 ) ;
  assign w16358 = ( \pi01 & \pi02 ) | ( \pi01 & w16357 ) | ( \pi02 & w16357 ) ;
  assign w16359 = ( w16354 & w16356 ) | ( w16354 & ~w16358 ) | ( w16356 & ~w16358 ) ;
  assign w16360 = w8954 | w11512 ;
  assign w16361 = ( ~w11512 & w16359 ) | ( ~w11512 & w16360 ) | ( w16359 & w16360 ) ;
  assign w16362 = \pi02 ^ w16361 ;
  assign w16363 = w15809 ^ w15983 ;
  assign w16364 = w15811 ^ w16363 ;
  assign w16365 = ( w16351 & w16362 ) | ( w16351 & w16364 ) | ( w16362 & w16364 ) ;
  assign w16366 = ( \pi02 & ~w9965 ) | ( \pi02 & w9967 ) | ( ~w9965 & w9967 ) ;
  assign w16367 = \pi00 ^ w16366 ;
  assign w16368 = ( \pi02 & w9965 ) | ( \pi02 & w16367 ) | ( w9965 & w16367 ) ;
  assign w16369 = ( ~\pi02 & w9967 ) | ( ~\pi02 & w16367 ) | ( w9967 & w16367 ) ;
  assign w16370 = \pi01 & ~w16369 ;
  assign w16371 = ( ~\pi00 & w9971 ) | ( ~\pi00 & w16370 ) | ( w9971 & w16370 ) ;
  assign w16372 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16371 ) | ( \pi02 & ~w16371 ) ;
  assign w16373 = ( w16368 & w16370 ) | ( w16368 & ~w16372 ) | ( w16370 & ~w16372 ) ;
  assign w16374 = w8954 | w11501 ;
  assign w16375 = ( ~w11501 & w16373 ) | ( ~w11501 & w16374 ) | ( w16373 & w16374 ) ;
  assign w16376 = \pi02 ^ w16375 ;
  assign w16377 = w15799 ^ w15984 ;
  assign w16378 = w15801 ^ w16377 ;
  assign w16379 = ( w16365 & w16376 ) | ( w16365 & w16378 ) | ( w16376 & w16378 ) ;
  assign w16380 = ( ~\pi02 & w9961 ) | ( ~\pi02 & w9965 ) | ( w9961 & w9965 ) ;
  assign w16381 = \pi00 ^ w16380 ;
  assign w16382 = ( \pi02 & w9961 ) | ( \pi02 & ~w16381 ) | ( w9961 & ~w16381 ) ;
  assign w16383 = ( \pi02 & w9965 ) | ( \pi02 & w16381 ) | ( w9965 & w16381 ) ;
  assign w16384 = \pi01 & w16383 ;
  assign w16385 = ( \pi00 & w9967 ) | ( \pi00 & ~w16384 ) | ( w9967 & ~w16384 ) ;
  assign w16386 = ( \pi01 & \pi02 ) | ( \pi01 & w16385 ) | ( \pi02 & w16385 ) ;
  assign w16387 = ( w16382 & w16384 ) | ( w16382 & ~w16386 ) | ( w16384 & ~w16386 ) ;
  assign w16388 = ~w8954 & w11339 ;
  assign w16389 = ( w11339 & w16387 ) | ( w11339 & ~w16388 ) | ( w16387 & ~w16388 ) ;
  assign w16390 = \pi02 ^ w16389 ;
  assign w16391 = w15789 ^ w15985 ;
  assign w16392 = w15791 ^ w16391 ;
  assign w16393 = ( w16379 & w16390 ) | ( w16379 & w16392 ) | ( w16390 & w16392 ) ;
  assign w16394 = ( \pi02 & ~w9961 ) | ( \pi02 & w9963 ) | ( ~w9961 & w9963 ) ;
  assign w16395 = \pi00 ^ w16394 ;
  assign w16396 = ( \pi02 & ~w9963 ) | ( \pi02 & w16395 ) | ( ~w9963 & w16395 ) ;
  assign w16397 = ( \pi02 & w9961 ) | ( \pi02 & ~w16395 ) | ( w9961 & ~w16395 ) ;
  assign w16398 = \pi01 & w16397 ;
  assign w16399 = ( ~\pi00 & w9965 ) | ( ~\pi00 & w16398 ) | ( w9965 & w16398 ) ;
  assign w16400 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16399 ) | ( \pi02 & ~w16399 ) ;
  assign w16401 = ( w16396 & w16398 ) | ( w16396 & ~w16400 ) | ( w16398 & ~w16400 ) ;
  assign w16402 = w8954 | w11278 ;
  assign w16403 = ( ~w11278 & w16401 ) | ( ~w11278 & w16402 ) | ( w16401 & w16402 ) ;
  assign w16404 = \pi02 ^ w16403 ;
  assign w16405 = w15781 ^ w15986 ;
  assign w16406 = w15773 ^ w16405 ;
  assign w16407 = ( w16393 & w16404 ) | ( w16393 & w16406 ) | ( w16404 & w16406 ) ;
  assign w16408 = ( \pi02 & ~w9957 ) | ( \pi02 & w9963 ) | ( ~w9957 & w9963 ) ;
  assign w16409 = \pi00 ^ w16408 ;
  assign w16410 = ( \pi02 & w9957 ) | ( \pi02 & w16409 ) | ( w9957 & w16409 ) ;
  assign w16411 = ( ~\pi02 & w9963 ) | ( ~\pi02 & w16409 ) | ( w9963 & w16409 ) ;
  assign w16412 = \pi01 & ~w16411 ;
  assign w16413 = ( ~\pi00 & w9961 ) | ( ~\pi00 & w16412 ) | ( w9961 & w16412 ) ;
  assign w16414 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16413 ) | ( \pi02 & ~w16413 ) ;
  assign w16415 = ( w16410 & w16412 ) | ( w16410 & ~w16414 ) | ( w16412 & ~w16414 ) ;
  assign w16416 = w8954 | w11089 ;
  assign w16417 = ( ~w11089 & w16415 ) | ( ~w11089 & w16416 ) | ( w16415 & w16416 ) ;
  assign w16418 = \pi02 ^ w16417 ;
  assign w16419 = w15771 ^ w15987 ;
  assign w16420 = w15763 ^ w16419 ;
  assign w16421 = ( w16407 & w16418 ) | ( w16407 & w16420 ) | ( w16418 & w16420 ) ;
  assign w16422 = ( \pi02 & w9955 ) | ( \pi02 & ~w9957 ) | ( w9955 & ~w9957 ) ;
  assign w16423 = \pi00 ^ w16422 ;
  assign w16424 = ( \pi02 & ~w9955 ) | ( \pi02 & w16423 ) | ( ~w9955 & w16423 ) ;
  assign w16425 = ( \pi02 & w9957 ) | ( \pi02 & ~w16423 ) | ( w9957 & ~w16423 ) ;
  assign w16426 = \pi01 & w16425 ;
  assign w16427 = ( \pi00 & w9963 ) | ( \pi00 & ~w16426 ) | ( w9963 & ~w16426 ) ;
  assign w16428 = ( \pi01 & \pi02 ) | ( \pi01 & w16427 ) | ( \pi02 & w16427 ) ;
  assign w16429 = ( w16424 & w16426 ) | ( w16424 & ~w16428 ) | ( w16426 & ~w16428 ) ;
  assign w16430 = w8954 | w11202 ;
  assign w16431 = ( ~w11202 & w16429 ) | ( ~w11202 & w16430 ) | ( w16429 & w16430 ) ;
  assign w16432 = \pi02 ^ w16431 ;
  assign w16433 = w15761 ^ w15988 ;
  assign w16434 = w15753 ^ w16433 ;
  assign w16435 = ( w16421 & w16432 ) | ( w16421 & w16434 ) | ( w16432 & w16434 ) ;
  assign w16436 = ( \pi02 & ~w9842 ) | ( \pi02 & w9955 ) | ( ~w9842 & w9955 ) ;
  assign w16437 = \pi00 ^ w16436 ;
  assign w16438 = ( \pi02 & w9842 ) | ( \pi02 & w16437 ) | ( w9842 & w16437 ) ;
  assign w16439 = ( ~\pi02 & w9955 ) | ( ~\pi02 & w16437 ) | ( w9955 & w16437 ) ;
  assign w16440 = \pi01 & ~w16439 ;
  assign w16441 = ( ~\pi00 & w9957 ) | ( ~\pi00 & w16440 ) | ( w9957 & w16440 ) ;
  assign w16442 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16441 ) | ( \pi02 & ~w16441 ) ;
  assign w16443 = ( w16438 & w16440 ) | ( w16438 & ~w16442 ) | ( w16440 & ~w16442 ) ;
  assign w16444 = w8954 | w10976 ;
  assign w16445 = ( ~w10976 & w16443 ) | ( ~w10976 & w16444 ) | ( w16443 & w16444 ) ;
  assign w16446 = \pi02 ^ w16445 ;
  assign w16447 = w15749 ^ w15989 ;
  assign w16448 = w15751 ^ w16447 ;
  assign w16449 = ( w16435 & w16446 ) | ( w16435 & w16448 ) | ( w16446 & w16448 ) ;
  assign w16450 = ( ~\pi02 & w9842 ) | ( ~\pi02 & w9953 ) | ( w9842 & w9953 ) ;
  assign w16451 = \pi00 ^ w16450 ;
  assign w16452 = ( \pi02 & w9953 ) | ( \pi02 & ~w16451 ) | ( w9953 & ~w16451 ) ;
  assign w16453 = ( \pi02 & w9842 ) | ( \pi02 & w16451 ) | ( w9842 & w16451 ) ;
  assign w16454 = \pi01 & w16453 ;
  assign w16455 = ( \pi00 & w9955 ) | ( \pi00 & ~w16454 ) | ( w9955 & ~w16454 ) ;
  assign w16456 = ( \pi01 & \pi02 ) | ( \pi01 & w16455 ) | ( \pi02 & w16455 ) ;
  assign w16457 = ( w16452 & w16454 ) | ( w16452 & ~w16456 ) | ( w16454 & ~w16456 ) ;
  assign w16458 = ~w8954 & w10965 ;
  assign w16459 = ( w10965 & w16457 ) | ( w10965 & ~w16458 ) | ( w16457 & ~w16458 ) ;
  assign w16460 = \pi02 ^ w16459 ;
  assign w16461 = w15739 ^ w15990 ;
  assign w16462 = w15741 ^ w16461 ;
  assign w16463 = ( w16449 & w16460 ) | ( w16449 & w16462 ) | ( w16460 & w16462 ) ;
  assign w16464 = ( ~\pi02 & w9953 ) | ( ~\pi02 & w10114 ) | ( w9953 & w10114 ) ;
  assign w16465 = \pi00 ^ w16464 ;
  assign w16466 = ( \pi02 & w10114 ) | ( \pi02 & ~w16465 ) | ( w10114 & ~w16465 ) ;
  assign w16467 = ( \pi02 & w9953 ) | ( \pi02 & w16465 ) | ( w9953 & w16465 ) ;
  assign w16468 = \pi01 & w16467 ;
  assign w16469 = ( ~\pi00 & w9842 ) | ( ~\pi00 & w16468 ) | ( w9842 & w16468 ) ;
  assign w16470 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16469 ) | ( \pi02 & ~w16469 ) ;
  assign w16471 = ( w16466 & w16468 ) | ( w16466 & ~w16470 ) | ( w16468 & ~w16470 ) ;
  assign w16472 = ~w8954 & w10334 ;
  assign w16473 = ( w10334 & w16471 ) | ( w10334 & ~w16472 ) | ( w16471 & ~w16472 ) ;
  assign w16474 = \pi02 ^ w16473 ;
  assign w16475 = w15729 ^ w15991 ;
  assign w16476 = w15731 ^ w16475 ;
  assign w16477 = ( w16463 & w16474 ) | ( w16463 & w16476 ) | ( w16474 & w16476 ) ;
  assign w16478 = ( ~\pi02 & w10114 ) | ( ~\pi02 & w10211 ) | ( w10114 & w10211 ) ;
  assign w16479 = \pi00 ^ w16478 ;
  assign w16480 = ( \pi02 & w10211 ) | ( \pi02 & ~w16479 ) | ( w10211 & ~w16479 ) ;
  assign w16481 = ( \pi02 & w10114 ) | ( \pi02 & w16479 ) | ( w10114 & w16479 ) ;
  assign w16482 = \pi01 & w16481 ;
  assign w16483 = ( ~\pi00 & w9953 ) | ( ~\pi00 & w16482 ) | ( w9953 & w16482 ) ;
  assign w16484 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16483 ) | ( \pi02 & ~w16483 ) ;
  assign w16485 = ( w16480 & w16482 ) | ( w16480 & ~w16484 ) | ( w16482 & ~w16484 ) ;
  assign w16486 = ~w8954 & w10214 ;
  assign w16487 = ( w10214 & w16485 ) | ( w10214 & ~w16486 ) | ( w16485 & ~w16486 ) ;
  assign w16488 = \pi02 ^ w16487 ;
  assign w16489 = w15721 ^ w15992 ;
  assign w16490 = w15713 ^ w16489 ;
  assign w16491 = ( w16477 & w16488 ) | ( w16477 & w16490 ) | ( w16488 & w16490 ) ;
  assign w16492 = ( ~\pi02 & w10211 ) | ( ~\pi02 & w10784 ) | ( w10211 & w10784 ) ;
  assign w16493 = \pi00 ^ w16492 ;
  assign w16494 = ( \pi02 & w10784 ) | ( \pi02 & ~w16493 ) | ( w10784 & ~w16493 ) ;
  assign w16495 = ( \pi02 & w10211 ) | ( \pi02 & w16493 ) | ( w10211 & w16493 ) ;
  assign w16496 = \pi01 & w16495 ;
  assign w16497 = ( ~\pi00 & w10114 ) | ( ~\pi00 & w16496 ) | ( w10114 & w16496 ) ;
  assign w16498 = ( \pi01 & \pi02 ) | ( \pi01 & ~w16497 ) | ( \pi02 & ~w16497 ) ;
  assign w16499 = ( w16494 & w16496 ) | ( w16494 & ~w16498 ) | ( w16496 & ~w16498 ) ;
  assign w16500 = ~w8954 & w10789 ;
  assign w16501 = ( w10789 & w16499 ) | ( w10789 & ~w16500 ) | ( w16499 & ~w16500 ) ;
  assign w16502 = \pi02 ^ w16501 ;
  assign w16503 = w15711 ^ w15993 ;
  assign w16504 = w15703 ^ w16503 ;
  assign w16505 = ( w16491 & w16502 ) | ( w16491 & w16504 ) | ( w16502 & w16504 ) ;
  assign w16506 = ( ~w16100 & w16111 ) | ( ~w16100 & w16505 ) | ( w16111 & w16505 ) ;
  assign w16507 = ( ~w16087 & w16098 ) | ( ~w16087 & w16506 ) | ( w16098 & w16506 ) ;
  assign w16508 = ( w16074 & w16085 ) | ( w16074 & w16507 ) | ( w16085 & w16507 ) ;
  assign w16509 = ( ~w16061 & w16072 ) | ( ~w16061 & w16508 ) | ( w16072 & w16508 ) ;
  assign w16510 = w11160 & ~w16059 ;
  assign w16511 = ( w8954 & w16059 ) | ( w8954 & ~w16510 ) | ( w16059 & ~w16510 ) ;
  assign w16512 = \pi02 ^ w16511 ;
  assign w16513 = ( ~w16051 & w16509 ) | ( ~w16051 & w16512 ) | ( w16509 & w16512 ) ;
  assign w16514 = w11131 & ~w16049 ;
  assign w16515 = ( w8954 & w16049 ) | ( w8954 & ~w16514 ) | ( w16049 & ~w16514 ) ;
  assign w16516 = \pi02 ^ w16515 ;
  assign w16517 = ( w16041 & w16513 ) | ( w16041 & w16516 ) | ( w16513 & w16516 ) ;
  assign w16518 = w10895 | w16039 ;
  assign w16519 = ( w8954 & w16039 ) | ( w8954 & w16518 ) | ( w16039 & w16518 ) ;
  assign w16520 = \pi02 ^ w16519 ;
  assign w16521 = ( w16031 & w16517 ) | ( w16031 & w16520 ) | ( w16517 & w16520 ) ;
  assign w16522 = w11256 | w16029 ;
  assign w16523 = ( w8954 & w16029 ) | ( w8954 & w16522 ) | ( w16029 & w16522 ) ;
  assign w16524 = \pi02 ^ w16523 ;
  assign w16525 = ( w16021 & w16521 ) | ( w16021 & w16524 ) | ( w16521 & w16524 ) ;
  assign w16526 = w11145 & ~w16019 ;
  assign w16527 = ( w8954 & w16019 ) | ( w8954 & ~w16526 ) | ( w16019 & ~w16526 ) ;
  assign w16528 = \pi02 ^ w16527 ;
  assign w16529 = ( w16005 & w16525 ) | ( w16005 & w16528 ) | ( w16525 & w16528 ) ;
  assign w16530 = w15601 ^ w15610 ;
  assign w16531 = ( w16003 & w16529 ) | ( w16003 & w16530 ) | ( w16529 & w16530 ) ;
  assign w16532 = ( ~w15590 & w15611 ) | ( ~w15590 & w16531 ) | ( w15611 & w16531 ) ;
  assign w16533 = ( w15209 & w15588 ) | ( w15209 & w16532 ) | ( w15588 & w16532 ) ;
  assign w16534 = ( ~w14850 & w15207 ) | ( ~w14850 & w16533 ) | ( w15207 & w16533 ) ;
  assign w16535 = ( w14843 & ~w14845 ) | ( w14843 & w16534 ) | ( ~w14845 & w16534 ) ;
  assign w16536 = ( w14196 & w14509 ) | ( w14196 & w16535 ) | ( w14509 & w16535 ) ;
  assign w16537 = ( ~w13903 & w14194 ) | ( ~w13903 & w16536 ) | ( w14194 & w16536 ) ;
  assign w16538 = ( w13896 & ~w13898 ) | ( w13896 & w16537 ) | ( ~w13898 & w16537 ) ;
  assign w16539 = ( ~w13381 & w13628 ) | ( ~w13381 & w16538 ) | ( w13628 & w16538 ) ;
  assign w16540 = ( ~w13157 & w13379 ) | ( ~w13157 & w16539 ) | ( w13379 & w16539 ) ;
  assign w16541 = ( w13150 & ~w13152 ) | ( w13150 & w16540 ) | ( ~w13152 & w16540 ) ;
  assign w16542 = ( w12959 & w13055 ) | ( w12959 & w16541 ) | ( w13055 & w16541 ) ;
  assign w16543 = ( w12400 & w12957 ) | ( w12400 & w16542 ) | ( w12957 & w16542 ) ;
  assign w16544 = ( w12393 & ~w12395 ) | ( w12393 & w16543 ) | ( ~w12395 & w16543 ) ;
  assign w16545 = ( w12076 & w12309 ) | ( w12076 & w16544 ) | ( w12309 & w16544 ) ;
  assign w16546 = ( ~w11885 & w12074 ) | ( ~w11885 & w16545 ) | ( w12074 & w16545 ) ;
  assign w16547 = ( w11878 & w11880 ) | ( w11878 & w16546 ) | ( w11880 & w16546 ) ;
  assign w16548 = ( ~w11727 & w11790 ) | ( ~w11727 & w16547 ) | ( w11790 & w16547 ) ;
  assign w16549 = ( ~w11401 & w11725 ) | ( ~w11401 & w16548 ) | ( w11725 & w16548 ) ;
  assign w16550 = ( w11394 & ~w11396 ) | ( w11394 & w16549 ) | ( ~w11396 & w16549 ) ;
  assign w16551 = ( w11196 & w11264 ) | ( w11196 & w16550 ) | ( w11264 & w16550 ) ;
  assign w16552 = ( w11151 & w11194 ) | ( w11151 & w16551 ) | ( w11194 & w16551 ) ;
  assign w16553 = ~w11143 & w11146 ;
  assign w16554 = ( w4609 & w11143 ) | ( w4609 & ~w16553 ) | ( w11143 & ~w16553 ) ;
  assign w16555 = \pi23 ^ w16554 ;
  assign w16556 = ( w10902 & w11137 ) | ( w10902 & w16555 ) | ( w11137 & w16555 ) ;
  assign w16557 = ( w10820 & w10881 ) | ( w10820 & w10900 ) | ( w10881 & w10900 ) ;
  assign w16558 = ~w4143 & w10883 ;
  assign w16559 = w4052 & ~w10887 ;
  assign w16560 = ( w10883 & ~w16558 ) | ( w10883 & w16559 ) | ( ~w16558 & w16559 ) ;
  assign w16561 = ~w4147 & w11256 ;
  assign w16562 = w11139 & ~w16560 ;
  assign w16563 = ( w3964 & w16560 ) | ( w3964 & ~w16562 ) | ( w16560 & ~w16562 ) ;
  assign w16564 = ( w11256 & ~w16561 ) | ( w11256 & w16563 ) | ( ~w16561 & w16563 ) ;
  assign w16565 = \pi26 ^ w16564 ;
  assign w16566 = ( \pi29 & \pi31 ) | ( \pi29 & ~w10805 ) | ( \pi31 & ~w10805 ) ;
  assign w16567 = ( \pi29 & ~\pi30 ) | ( \pi29 & w16566 ) | ( ~\pi30 & w16566 ) ;
  assign w16568 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w16566 ) | ( \pi30 & w16566 ) ;
  assign w16569 = ( ~\pi29 & w10784 ) | ( ~\pi29 & w16568 ) | ( w10784 & w16568 ) ;
  assign w16570 = ( w10807 & ~w16568 ) | ( w10807 & w16569 ) | ( ~w16568 & w16569 ) ;
  assign w16571 = \pi31 | w16570 ;
  assign w16572 = ( w16567 & w16569 ) | ( w16567 & ~w16571 ) | ( w16569 & ~w16571 ) ;
  assign w16573 = ( w37 & w11117 ) | ( w37 & w16572 ) | ( w11117 & w16572 ) ;
  assign w16574 = w16572 | w16573 ;
  assign w16575 = ( \pi20 & \pi21 ) | ( \pi20 & ~\pi22 ) | ( \pi21 & ~\pi22 ) ;
  assign w16576 = ( \pi22 & ~\pi23 ) | ( \pi22 & w16575 ) | ( ~\pi23 & w16575 ) ;
  assign w16577 = w10738 ^ w16576 ;
  assign w16578 = ( \pi23 & w16576 ) | ( \pi23 & w16577 ) | ( w16576 & w16577 ) ;
  assign w16579 = w283 | w663 ;
  assign w16580 = ( w161 & ~w283 ) | ( w161 & w284 ) | ( ~w283 & w284 ) ;
  assign w16581 = w16579 | w16580 ;
  assign w16582 = ( ~w266 & w1154 ) | ( ~w266 & w16581 ) | ( w1154 & w16581 ) ;
  assign w16583 = w4830 | w12799 ;
  assign w16584 = ( w266 & w456 ) | ( w266 & ~w12799 ) | ( w456 & ~w12799 ) ;
  assign w16585 = w16583 | w16584 ;
  assign w16586 = w16582 | w16585 ;
  assign w16587 = w785 | w11601 ;
  assign w16588 = ( w11018 & ~w11601 ) | ( w11018 & w16586 ) | ( ~w11601 & w16586 ) ;
  assign w16589 = w16587 | w16588 ;
  assign w16590 = w860 | w1302 ;
  assign w16591 = w3826 | w16590 ;
  assign w16592 = ( w468 & ~w3826 ) | ( w468 & w16589 ) | ( ~w3826 & w16589 ) ;
  assign w16593 = w16591 | w16592 ;
  assign w16594 = ( w203 & w252 ) | ( w203 & ~w287 ) | ( w252 & ~w287 ) ;
  assign w16595 = w128 | w16593 ;
  assign w16596 = ( ~w128 & w287 ) | ( ~w128 & w353 ) | ( w287 & w353 ) ;
  assign w16597 = w16595 | w16596 ;
  assign w16598 = w16594 | w16597 ;
  assign w16599 = w16578 ^ w16598 ;
  assign w16600 = w10850 ^ w16599 ;
  assign w16601 = w10851 ^ w16600 ;
  assign w16602 = w16574 ^ w16601 ;
  assign w16603 = ( w10853 & w10864 ) | ( w10853 & w10879 ) | ( w10864 & w10879 ) ;
  assign w16604 = w3717 | w10866 ;
  assign w16605 = w3649 & w10801 ;
  assign w16606 = ( ~w10866 & w16604 ) | ( ~w10866 & w16605 ) | ( w16604 & w16605 ) ;
  assign w16607 = w3549 | w10885 ;
  assign w16608 = w11160 & ~w16606 ;
  assign w16609 = ( w3448 & w16606 ) | ( w3448 & ~w16608 ) | ( w16606 & ~w16608 ) ;
  assign w16610 = ( ~w10885 & w16607 ) | ( ~w10885 & w16609 ) | ( w16607 & w16609 ) ;
  assign w16611 = \pi29 ^ w16610 ;
  assign w16612 = w16602 ^ w16603 ;
  assign w16613 = w16611 ^ w16612 ;
  assign w16614 = w16557 ^ w16613 ;
  assign w16615 = w16565 ^ w16614 ;
  assign w16616 = w16552 ^ w16556 ;
  assign w16617 = w16615 ^ w16616 ;
  assign w16618 = w11196 ^ w16550 ;
  assign w16619 = w11264 ^ w16618 ;
  assign w16620 = w11151 ^ w16551 ;
  assign w16621 = w11194 ^ w16620 ;
  assign w16622 = ~w8593 & w16621 ;
  assign w16623 = w8262 & w16619 ;
  assign w16624 = ( w16621 & ~w16622 ) | ( w16621 & w16623 ) | ( ~w16622 & w16623 ) ;
  assign w16625 = w11394 ^ w16549 ;
  assign w16626 = w11396 ^ w16625 ;
  assign w16627 = w11725 ^ w16548 ;
  assign w16628 = w11401 ^ w16627 ;
  assign w16629 = w11727 ^ w16547 ;
  assign w16630 = w11790 ^ w16629 ;
  assign w16631 = w11878 ^ w16546 ;
  assign w16632 = w11880 ^ w16631 ;
  assign w16633 = w12074 ^ w16545 ;
  assign w16634 = w11885 ^ w16633 ;
  assign w16635 = w12076 ^ w16544 ;
  assign w16636 = w12309 ^ w16635 ;
  assign w16637 = w12393 ^ w16543 ;
  assign w16638 = w12395 ^ w16637 ;
  assign w16639 = w12400 ^ w16542 ;
  assign w16640 = w12957 ^ w16639 ;
  assign w16641 = w12959 ^ w16541 ;
  assign w16642 = w13055 ^ w16641 ;
  assign w16643 = w13150 ^ w16540 ;
  assign w16644 = w13152 ^ w16643 ;
  assign w16645 = w13157 ^ w16539 ;
  assign w16646 = w13379 ^ w16645 ;
  assign w16647 = w13381 ^ w16538 ;
  assign w16648 = w13628 ^ w16647 ;
  assign w16649 = w13896 ^ w16537 ;
  assign w16650 = w13898 ^ w16649 ;
  assign w16651 = w13903 ^ w16536 ;
  assign w16652 = w14194 ^ w16651 ;
  assign w16653 = w14196 ^ w16535 ;
  assign w16654 = w14509 ^ w16653 ;
  assign w16655 = w14843 ^ w16534 ;
  assign w16656 = w14845 ^ w16655 ;
  assign w16657 = w14850 ^ w16533 ;
  assign w16658 = w15207 ^ w16657 ;
  assign w16659 = w15209 ^ w16532 ;
  assign w16660 = w15588 ^ w16659 ;
  assign w16661 = w15590 ^ w16531 ;
  assign w16662 = w15611 ^ w16661 ;
  assign w16663 = w15601 ^ w16003 ;
  assign w16664 = w16529 ^ w16663 ;
  assign w16665 = w15610 ^ w16664 ;
  assign w16666 = w8954 & w11145 ;
  assign w16667 = ( w8954 & w16019 ) | ( w8954 & ~w16666 ) | ( w16019 & ~w16666 ) ;
  assign w16668 = w16525 ^ w16667 ;
  assign w16669 = \pi02 ^ w16005 ;
  assign w16670 = w16668 ^ w16669 ;
  assign w16671 = w8954 & ~w11256 ;
  assign w16672 = ( w8954 & w16029 ) | ( w8954 & ~w16671 ) | ( w16029 & ~w16671 ) ;
  assign w16673 = w16521 ^ w16672 ;
  assign w16674 = \pi02 ^ w16021 ;
  assign w16675 = w16673 ^ w16674 ;
  assign w16676 = w8954 & ~w10895 ;
  assign w16677 = ( w8954 & w16039 ) | ( w8954 & ~w16676 ) | ( w16039 & ~w16676 ) ;
  assign w16678 = w16517 ^ w16677 ;
  assign w16679 = \pi02 ^ w16031 ;
  assign w16680 = w16678 ^ w16679 ;
  assign w16681 = w8954 & w11131 ;
  assign w16682 = ( w8954 & w16049 ) | ( w8954 & ~w16681 ) | ( w16049 & ~w16681 ) ;
  assign w16683 = w16513 ^ w16682 ;
  assign w16684 = \pi02 ^ w16041 ;
  assign w16685 = w16683 ^ w16684 ;
  assign w16686 = w8954 & w11160 ;
  assign w16687 = ( w8954 & w16059 ) | ( w8954 & ~w16686 ) | ( w16059 & ~w16686 ) ;
  assign w16688 = w16509 ^ w16687 ;
  assign w16689 = \pi02 ^ w16051 ;
  assign w16690 = w16688 ^ w16689 ;
  assign w16691 = w16072 ^ w16508 ;
  assign w16692 = w16061 ^ w16691 ;
  assign w16693 = w16085 ^ w16507 ;
  assign w16694 = w16074 ^ w16693 ;
  assign w16695 = w16098 ^ w16506 ;
  assign w16696 = w16087 ^ w16695 ;
  assign w16697 = w16111 ^ w16505 ;
  assign w16698 = w16100 ^ w16697 ;
  assign w16699 = ( ~w16685 & w16690 ) | ( ~w16685 & w16692 ) | ( w16690 & w16692 ) ;
  assign w16700 = w16690 | w16696 ;
  assign w16701 = ( w16696 & w16698 ) | ( w16696 & w16700 ) | ( w16698 & w16700 ) ;
  assign w16702 = ( w16690 & w16694 ) | ( w16690 & ~w16701 ) | ( w16694 & ~w16701 ) ;
  assign w16703 = ( w16690 & w16699 ) | ( w16690 & ~w16702 ) | ( w16699 & ~w16702 ) ;
  assign w16704 = ( w16680 & w16685 ) | ( w16680 & ~w16703 ) | ( w16685 & ~w16703 ) ;
  assign w16705 = ( w16675 & w16680 ) | ( w16675 & w16704 ) | ( w16680 & w16704 ) ;
  assign w16706 = ( w16670 & w16675 ) | ( w16670 & w16705 ) | ( w16675 & w16705 ) ;
  assign w16707 = ( w16665 & w16670 ) | ( w16665 & w16706 ) | ( w16670 & w16706 ) ;
  assign w16708 = ( w16660 & ~w16662 ) | ( w16660 & w16707 ) | ( ~w16662 & w16707 ) ;
  assign w16709 = ( ~w16662 & w16665 ) | ( ~w16662 & w16708 ) | ( w16665 & w16708 ) ;
  assign w16710 = ( ~w16658 & w16660 ) | ( ~w16658 & w16709 ) | ( w16660 & w16709 ) ;
  assign w16711 = ( w16656 & w16658 ) | ( w16656 & ~w16710 ) | ( w16658 & ~w16710 ) ;
  assign w16712 = ( ~w16654 & w16656 ) | ( ~w16654 & w16711 ) | ( w16656 & w16711 ) ;
  assign w16713 = ( w16650 & w16652 ) | ( w16650 & w16712 ) | ( w16652 & w16712 ) ;
  assign w16714 = ( w16652 & ~w16654 ) | ( w16652 & w16713 ) | ( ~w16654 & w16713 ) ;
  assign w16715 = ( w16648 & w16650 ) | ( w16648 & w16714 ) | ( w16650 & w16714 ) ;
  assign w16716 = ( w16644 & w16646 ) | ( w16644 & w16715 ) | ( w16646 & w16715 ) ;
  assign w16717 = ( w16646 & w16648 ) | ( w16646 & w16716 ) | ( w16648 & w16716 ) ;
  assign w16718 = ( ~w16642 & w16644 ) | ( ~w16642 & w16717 ) | ( w16644 & w16717 ) ;
  assign w16719 = ( w16638 & ~w16640 ) | ( w16638 & w16718 ) | ( ~w16640 & w16718 ) ;
  assign w16720 = ( w16640 & w16642 ) | ( w16640 & ~w16719 ) | ( w16642 & ~w16719 ) ;
  assign w16721 = ( w16636 & ~w16638 ) | ( w16636 & w16720 ) | ( ~w16638 & w16720 ) ;
  assign w16722 = ( w16632 & ~w16634 ) | ( w16632 & w16721 ) | ( ~w16634 & w16721 ) ;
  assign w16723 = ( ~w16634 & w16636 ) | ( ~w16634 & w16722 ) | ( w16636 & w16722 ) ;
  assign w16724 = ( ~w16630 & w16632 ) | ( ~w16630 & w16723 ) | ( w16632 & w16723 ) ;
  assign w16725 = ( w16626 & w16628 ) | ( w16626 & ~w16724 ) | ( w16628 & ~w16724 ) ;
  assign w16726 = ( w16628 & w16630 ) | ( w16628 & w16725 ) | ( w16630 & w16725 ) ;
  assign w16727 = ( ~w16619 & w16626 ) | ( ~w16619 & w16726 ) | ( w16626 & w16726 ) ;
  assign w16728 = ( w16617 & w16621 ) | ( w16617 & ~w16727 ) | ( w16621 & ~w16727 ) ;
  assign w16729 = ( w16619 & w16621 ) | ( w16619 & w16728 ) | ( w16621 & w16728 ) ;
  assign w16730 = ( w16619 & w16621 ) | ( w16619 & ~w16727 ) | ( w16621 & ~w16727 ) ;
  assign w16731 = w16621 ^ w16730 ;
  assign w16732 = w16617 ^ w16731 ;
  assign w16733 = ~w8263 & w16732 ;
  assign w16734 = w16617 | w16624 ;
  assign w16735 = ( w35 & w16624 ) | ( w35 & w16734 ) | ( w16624 & w16734 ) ;
  assign w16736 = ( w16732 & ~w16733 ) | ( w16732 & w16735 ) | ( ~w16733 & w16735 ) ;
  assign w16737 = \pi05 ^ w16736 ;
  assign w16738 = ~w6949 & w16636 ;
  assign w16739 = w6748 & ~w16638 ;
  assign w16740 = ( w16636 & ~w16738 ) | ( w16636 & w16739 ) | ( ~w16738 & w16739 ) ;
  assign w16741 = w16634 ^ w16721 ;
  assign w16742 = w16636 ^ w16741 ;
  assign w16743 = w7154 | w16634 ;
  assign w16744 = ~w16740 & w16742 ;
  assign w16745 = ( w6751 & w16740 ) | ( w6751 & ~w16744 ) | ( w16740 & ~w16744 ) ;
  assign w16746 = ( ~w16634 & w16743 ) | ( ~w16634 & w16745 ) | ( w16743 & w16745 ) ;
  assign w16747 = \pi11 ^ w16746 ;
  assign w16748 = w5710 | w16650 ;
  assign w16749 = w5494 & ~w16652 ;
  assign w16750 = ( ~w16650 & w16748 ) | ( ~w16650 & w16749 ) | ( w16748 & w16749 ) ;
  assign w16751 = w16648 ^ w16714 ;
  assign w16752 = w16650 ^ w16751 ;
  assign w16753 = w5948 | w16648 ;
  assign w16754 = ~w16750 & w16752 ;
  assign w16755 = ( w5497 & w16750 ) | ( w5497 & ~w16754 ) | ( w16750 & ~w16754 ) ;
  assign w16756 = ( ~w16648 & w16753 ) | ( ~w16648 & w16755 ) | ( w16753 & w16755 ) ;
  assign w16757 = \pi17 ^ w16756 ;
  assign w16758 = ~w4651 & w16665 ;
  assign w16759 = w4606 & w16670 ;
  assign w16760 = ( w16665 & ~w16758 ) | ( w16665 & w16759 ) | ( ~w16758 & w16759 ) ;
  assign w16761 = w16662 ^ w16707 ;
  assign w16762 = w16665 ^ w16761 ;
  assign w16763 = w4706 | w16662 ;
  assign w16764 = ~w16760 & w16762 ;
  assign w16765 = ( w4609 & w16760 ) | ( w4609 & ~w16764 ) | ( w16760 & ~w16764 ) ;
  assign w16766 = ( ~w16662 & w16763 ) | ( ~w16662 & w16765 ) | ( w16763 & w16765 ) ;
  assign w16767 = \pi23 ^ w16766 ;
  assign w16768 = ~w4143 & w16685 ;
  assign w16769 = w4052 & ~w16690 ;
  assign w16770 = ( w16685 & ~w16768 ) | ( w16685 & w16769 ) | ( ~w16768 & w16769 ) ;
  assign w16771 = w16680 ^ w16703 ;
  assign w16772 = w16685 ^ w16771 ;
  assign w16773 = w4147 | w16772 ;
  assign w16774 = w16680 | w16770 ;
  assign w16775 = ( w3964 & w16770 ) | ( w3964 & w16774 ) | ( w16770 & w16774 ) ;
  assign w16776 = ( ~w16772 & w16773 ) | ( ~w16772 & w16775 ) | ( w16773 & w16775 ) ;
  assign w16777 = \pi26 ^ w16776 ;
  assign w16778 = ~w3717 & w16694 ;
  assign w16779 = w3649 & ~w16696 ;
  assign w16780 = ( w16694 & ~w16778 ) | ( w16694 & w16779 ) | ( ~w16778 & w16779 ) ;
  assign w16781 = w16692 ^ w16696 ;
  assign w16782 = ~w16694 & w16696 ;
  assign w16783 = ( w16694 & w16698 ) | ( w16694 & ~w16782 ) | ( w16698 & ~w16782 ) ;
  assign w16784 = w16781 ^ w16783 ;
  assign w16785 = w3549 | w16692 ;
  assign w16786 = w16780 | w16784 ;
  assign w16787 = ( w3448 & w16780 ) | ( w3448 & w16786 ) | ( w16780 & w16786 ) ;
  assign w16788 = ( ~w16692 & w16785 ) | ( ~w16692 & w16787 ) | ( w16785 & w16787 ) ;
  assign w16789 = \pi29 ^ w16788 ;
  assign w16790 = \pi29 & w16698 ;
  assign w16791 = w16696 & w16790 ;
  assign w16792 = ( \pi26 & \pi27 ) | ( \pi26 & ~w16791 ) | ( \pi27 & ~w16791 ) ;
  assign w16793 = ( \pi28 & \pi29 ) | ( \pi28 & ~w16792 ) | ( \pi29 & ~w16792 ) ;
  assign w16794 = ( \pi28 & ~w16790 ) | ( \pi28 & w16792 ) | ( ~w16790 & w16792 ) ;
  assign w16795 = ( w6866 & w16793 ) | ( w6866 & ~w16794 ) | ( w16793 & ~w16794 ) ;
  assign w16796 = w3549 & w16694 ;
  assign w16797 = ( w3717 & ~w16696 ) | ( w3717 & w16796 ) | ( ~w16696 & w16796 ) ;
  assign w16798 = w3649 | w16797 ;
  assign w16799 = ( ~w16698 & w16797 ) | ( ~w16698 & w16798 ) | ( w16797 & w16798 ) ;
  assign w16800 = w16796 | w16799 ;
  assign w16801 = ~w16696 & w16698 ;
  assign w16802 = w16694 ^ w16801 ;
  assign w16803 = w3448 & ~w16802 ;
  assign w16804 = ( w3448 & w16800 ) | ( w3448 & ~w16803 ) | ( w16800 & ~w16803 ) ;
  assign w16805 = \pi29 ^ w16804 ;
  assign w16806 = w16795 & w16805 ;
  assign w16807 = w36 & ~w16698 ;
  assign w16808 = w16789 ^ w16806 ;
  assign w16809 = w16807 ^ w16808 ;
  assign w16810 = w4143 | w16690 ;
  assign w16811 = w4052 & ~w16692 ;
  assign w16812 = ( ~w16690 & w16810 ) | ( ~w16690 & w16811 ) | ( w16810 & w16811 ) ;
  assign w16813 = ( w16692 & ~w16696 ) | ( w16692 & w16698 ) | ( ~w16696 & w16698 ) ;
  assign w16814 = w16692 | w16813 ;
  assign w16815 = ( w16690 & w16696 ) | ( w16690 & w16814 ) | ( w16696 & w16814 ) ;
  assign w16816 = ( w16692 & ~w16694 ) | ( w16692 & w16815 ) | ( ~w16694 & w16815 ) ;
  assign w16817 = w16685 ^ w16816 ;
  assign w16818 = w16690 ^ w16817 ;
  assign w16819 = ~w4147 & w16818 ;
  assign w16820 = w16685 | w16812 ;
  assign w16821 = ( w3964 & w16812 ) | ( w3964 & w16820 ) | ( w16812 & w16820 ) ;
  assign w16822 = ( w16818 & ~w16819 ) | ( w16818 & w16821 ) | ( ~w16819 & w16821 ) ;
  assign w16823 = \pi26 ^ w16822 ;
  assign w16824 = w16795 ^ w16805 ;
  assign w16825 = ( \pi26 & \pi27 ) | ( \pi26 & ~w16696 ) | ( \pi27 & ~w16696 ) ;
  assign w16826 = ( \pi26 & \pi27 ) | ( \pi26 & ~w16698 ) | ( \pi27 & ~w16698 ) ;
  assign w16827 = \pi28 ^ w16698 ;
  assign w16828 = ( \pi28 & w16826 ) | ( \pi28 & w16827 ) | ( w16826 & w16827 ) ;
  assign w16829 = w16825 ^ w16828 ;
  assign w16830 = w3964 & ~w16690 ;
  assign w16831 = ( w4143 & ~w16692 ) | ( w4143 & w16830 ) | ( ~w16692 & w16830 ) ;
  assign w16832 = w4052 | w16831 ;
  assign w16833 = ( w16694 & w16831 ) | ( w16694 & w16832 ) | ( w16831 & w16832 ) ;
  assign w16834 = w16830 | w16833 ;
  assign w16835 = ( w16692 & ~w16694 ) | ( w16692 & w16696 ) | ( ~w16694 & w16696 ) ;
  assign w16836 = ~w16694 & w16698 ;
  assign w16837 = w16835 | w16836 ;
  assign w16838 = w16690 ^ w16692 ;
  assign w16839 = w16837 ^ w16838 ;
  assign w16840 = w4147 & w16839 ;
  assign w16841 = ( w4147 & w16834 ) | ( w4147 & ~w16840 ) | ( w16834 & ~w16840 ) ;
  assign w16842 = \pi26 ^ w16841 ;
  assign w16843 = \pi26 & w16698 ;
  assign w16844 = w16696 & w16843 ;
  assign w16845 = ( \pi23 & \pi24 ) | ( \pi23 & ~w16844 ) | ( \pi24 & ~w16844 ) ;
  assign w16846 = ( \pi25 & \pi26 ) | ( \pi25 & ~w16845 ) | ( \pi26 & ~w16845 ) ;
  assign w16847 = ( \pi25 & ~w16843 ) | ( \pi25 & w16845 ) | ( ~w16843 & w16845 ) ;
  assign w16848 = ( w7079 & w16846 ) | ( w7079 & ~w16847 ) | ( w16846 & ~w16847 ) ;
  assign w16849 = w3964 & w16694 ;
  assign w16850 = ( w4143 & ~w16696 ) | ( w4143 & w16849 ) | ( ~w16696 & w16849 ) ;
  assign w16851 = w4052 | w16850 ;
  assign w16852 = ( ~w16698 & w16850 ) | ( ~w16698 & w16851 ) | ( w16850 & w16851 ) ;
  assign w16853 = w16849 | w16852 ;
  assign w16854 = ~w4147 & w16802 ;
  assign w16855 = ( w16802 & w16853 ) | ( w16802 & ~w16854 ) | ( w16853 & ~w16854 ) ;
  assign w16856 = \pi26 ^ w16855 ;
  assign w16857 = w16848 & w16856 ;
  assign w16858 = ~w4143 & w16694 ;
  assign w16859 = w4052 & ~w16696 ;
  assign w16860 = ( w16694 & ~w16858 ) | ( w16694 & w16859 ) | ( ~w16858 & w16859 ) ;
  assign w16861 = ~w4147 & w16784 ;
  assign w16862 = w16692 & ~w16860 ;
  assign w16863 = ( w3964 & w16860 ) | ( w3964 & ~w16862 ) | ( w16860 & ~w16862 ) ;
  assign w16864 = ( w16784 & ~w16861 ) | ( w16784 & w16863 ) | ( ~w16861 & w16863 ) ;
  assign w16865 = \pi26 ^ w16864 ;
  assign w16866 = w3447 & ~w16698 ;
  assign w16867 = ( w16857 & w16865 ) | ( w16857 & w16866 ) | ( w16865 & w16866 ) ;
  assign w16868 = ( w16829 & w16842 ) | ( w16829 & w16867 ) | ( w16842 & w16867 ) ;
  assign w16869 = ( w16823 & w16824 ) | ( w16823 & w16868 ) | ( w16824 & w16868 ) ;
  assign w16870 = ( w16777 & w16809 ) | ( w16777 & w16869 ) | ( w16809 & w16869 ) ;
  assign w16871 = w3717 | w16692 ;
  assign w16872 = w3649 & w16694 ;
  assign w16873 = ( ~w16692 & w16871 ) | ( ~w16692 & w16872 ) | ( w16871 & w16872 ) ;
  assign w16874 = w3549 | w16690 ;
  assign w16875 = w16839 & ~w16873 ;
  assign w16876 = ( w3448 & w16873 ) | ( w3448 & ~w16875 ) | ( w16873 & ~w16875 ) ;
  assign w16877 = ( ~w16690 & w16874 ) | ( ~w16690 & w16876 ) | ( w16874 & w16876 ) ;
  assign w16878 = \pi29 ^ w16877 ;
  assign w16879 = w430 | w2169 ;
  assign w16880 = ( w429 & w900 ) | ( w429 & ~w2169 ) | ( w900 & ~w2169 ) ;
  assign w16881 = w16879 | w16880 ;
  assign w16882 = ( w68 & w74 ) | ( w68 & ~w118 ) | ( w74 & ~w118 ) ;
  assign w16883 = w1401 | w16881 ;
  assign w16884 = ( w118 & w459 ) | ( w118 & ~w1401 ) | ( w459 & ~w1401 ) ;
  assign w16885 = w16883 | w16884 ;
  assign w16886 = w16882 | w16885 ;
  assign w16887 = ( w408 & w722 ) | ( w408 & ~w802 ) | ( w722 & ~w802 ) ;
  assign w16888 = w205 | w16886 ;
  assign w16889 = ( ~w205 & w802 ) | ( ~w205 & w1001 ) | ( w802 & w1001 ) ;
  assign w16890 = w16888 | w16889 ;
  assign w16891 = w16887 | w16890 ;
  assign w16892 = w313 | w423 ;
  assign w16893 = w201 | w16892 ;
  assign w16894 = ( ~w201 & w208 ) | ( ~w201 & w594 ) | ( w208 & w594 ) ;
  assign w16895 = w16893 | w16894 ;
  assign w16896 = ( w2949 & w4177 ) | ( w2949 & w16895 ) | ( w4177 & w16895 ) ;
  assign w16897 = w2949 & ~w16896 ;
  assign w16898 = w310 | w511 ;
  assign w16899 = w3251 | w16898 ;
  assign w16900 = ( w3251 & ~w11292 ) | ( w3251 & w16897 ) | ( ~w11292 & w16897 ) ;
  assign w16901 = ~w16899 & w16900 ;
  assign w16902 = ( ~w354 & w638 ) | ( ~w354 & w2374 ) | ( w638 & w2374 ) ;
  assign w16903 = ~w410 & w16901 ;
  assign w16904 = ( w354 & ~w410 ) | ( w354 & w534 ) | ( ~w410 & w534 ) ;
  assign w16905 = w16903 & ~w16904 ;
  assign w16906 = ~w16902 & w16905 ;
  assign w16907 = w490 | w593 ;
  assign w16908 = w133 | w16907 ;
  assign w16909 = ( w133 & ~w445 ) | ( w133 & w16906 ) | ( ~w445 & w16906 ) ;
  assign w16910 = ~w16908 & w16909 ;
  assign w16911 = ( w225 & w533 ) | ( w225 & ~w663 ) | ( w533 & ~w663 ) ;
  assign w16912 = w1068 | w2147 ;
  assign w16913 = ( w663 & w1130 ) | ( w663 & ~w2147 ) | ( w1130 & ~w2147 ) ;
  assign w16914 = w16912 | w16913 ;
  assign w16915 = w16911 | w16914 ;
  assign w16916 = w12710 | w16915 ;
  assign w16917 = ( ~w1185 & w16891 ) | ( ~w1185 & w16916 ) | ( w16891 & w16916 ) ;
  assign w16918 = ~w12599 & w16910 ;
  assign w16919 = ( w1185 & w1302 ) | ( w1185 & w16910 ) | ( w1302 & w16910 ) ;
  assign w16920 = w16918 & ~w16919 ;
  assign w16921 = ~w16917 & w16920 ;
  assign w16922 = w1154 | w1206 ;
  assign w16923 = w326 | w16922 ;
  assign w16924 = ( w326 & ~w822 ) | ( w326 & w16921 ) | ( ~w822 & w16921 ) ;
  assign w16925 = ~w16923 & w16924 ;
  assign w16926 = ( w163 & w315 ) | ( w163 & ~w352 ) | ( w315 & ~w352 ) ;
  assign w16927 = ~w113 & w16925 ;
  assign w16928 = ( ~w113 & w352 ) | ( ~w113 & w388 ) | ( w352 & w388 ) ;
  assign w16929 = w16927 & ~w16928 ;
  assign w16930 = ~w16926 & w16929 ;
  assign w16931 = ( \pi29 & \pi30 ) | ( \pi29 & ~w16696 ) | ( \pi30 & ~w16696 ) ;
  assign w16932 = \pi31 ^ w16698 ;
  assign w16933 = ( \pi31 & w6862 ) | ( \pi31 & w16932 ) | ( w6862 & w16932 ) ;
  assign w16934 = w16931 ^ w16933 ;
  assign w16935 = ~w16930 & w16934 ;
  assign w16936 = w16930 ^ w16934 ;
  assign w16937 = ( w16789 & w16806 ) | ( w16789 & w16807 ) | ( w16806 & w16807 ) ;
  assign w16938 = w16878 ^ w16937 ;
  assign w16939 = w16936 ^ w16938 ;
  assign w16940 = w3964 & w16675 ;
  assign w16941 = ( w4143 & w16680 ) | ( w4143 & w16940 ) | ( w16680 & w16940 ) ;
  assign w16942 = w4052 | w16941 ;
  assign w16943 = ( w16685 & w16941 ) | ( w16685 & w16942 ) | ( w16941 & w16942 ) ;
  assign w16944 = w16940 | w16943 ;
  assign w16945 = w16675 ^ w16704 ;
  assign w16946 = w16680 ^ w16945 ;
  assign w16947 = w4147 & ~w16946 ;
  assign w16948 = ( w4147 & w16944 ) | ( w4147 & ~w16947 ) | ( w16944 & ~w16947 ) ;
  assign w16949 = \pi26 ^ w16948 ;
  assign w16950 = w16870 ^ w16949 ;
  assign w16951 = w16939 ^ w16950 ;
  assign w16952 = w16777 ^ w16869 ;
  assign w16953 = w16809 ^ w16952 ;
  assign w16954 = w4606 & w16675 ;
  assign w16955 = ( w4706 & w16665 ) | ( w4706 & w16954 ) | ( w16665 & w16954 ) ;
  assign w16956 = w4651 | w16955 ;
  assign w16957 = ( w16670 & w16955 ) | ( w16670 & w16956 ) | ( w16955 & w16956 ) ;
  assign w16958 = w16954 | w16957 ;
  assign w16959 = w16665 ^ w16706 ;
  assign w16960 = w16670 ^ w16959 ;
  assign w16961 = w4609 & ~w16960 ;
  assign w16962 = ( w4609 & w16958 ) | ( w4609 & ~w16961 ) | ( w16958 & ~w16961 ) ;
  assign w16963 = \pi23 ^ w16962 ;
  assign w16964 = w16823 ^ w16868 ;
  assign w16965 = w16824 ^ w16964 ;
  assign w16966 = w4606 & w16680 ;
  assign w16967 = ( w4706 & w16670 ) | ( w4706 & w16966 ) | ( w16670 & w16966 ) ;
  assign w16968 = w4651 | w16967 ;
  assign w16969 = ( w16675 & w16967 ) | ( w16675 & w16968 ) | ( w16967 & w16968 ) ;
  assign w16970 = w16966 | w16969 ;
  assign w16971 = w16670 ^ w16705 ;
  assign w16972 = w16675 ^ w16971 ;
  assign w16973 = w4609 & ~w16972 ;
  assign w16974 = ( w4609 & w16970 ) | ( w4609 & ~w16973 ) | ( w16970 & ~w16973 ) ;
  assign w16975 = \pi23 ^ w16974 ;
  assign w16976 = ~w4651 & w16680 ;
  assign w16977 = w4606 & w16685 ;
  assign w16978 = ( w16680 & ~w16976 ) | ( w16680 & w16977 ) | ( ~w16976 & w16977 ) ;
  assign w16979 = ~w4706 & w16675 ;
  assign w16980 = w16946 | w16978 ;
  assign w16981 = ( w4609 & w16978 ) | ( w4609 & w16980 ) | ( w16978 & w16980 ) ;
  assign w16982 = ( w16675 & ~w16979 ) | ( w16675 & w16981 ) | ( ~w16979 & w16981 ) ;
  assign w16983 = \pi23 ^ w16982 ;
  assign w16984 = w16842 ^ w16867 ;
  assign w16985 = w16829 ^ w16984 ;
  assign w16986 = w16857 ^ w16865 ;
  assign w16987 = w16866 ^ w16986 ;
  assign w16988 = w4606 & ~w16690 ;
  assign w16989 = ( w4706 & w16680 ) | ( w4706 & w16988 ) | ( w16680 & w16988 ) ;
  assign w16990 = w4651 | w16989 ;
  assign w16991 = ( w16685 & w16989 ) | ( w16685 & w16990 ) | ( w16989 & w16990 ) ;
  assign w16992 = w16988 | w16991 ;
  assign w16993 = w4609 | w16772 ;
  assign w16994 = ( ~w16772 & w16992 ) | ( ~w16772 & w16993 ) | ( w16992 & w16993 ) ;
  assign w16995 = \pi23 ^ w16994 ;
  assign w16996 = w4651 | w16690 ;
  assign w16997 = w4606 & ~w16692 ;
  assign w16998 = ( ~w16690 & w16996 ) | ( ~w16690 & w16997 ) | ( w16996 & w16997 ) ;
  assign w16999 = ~w4706 & w16685 ;
  assign w17000 = w16818 | w16998 ;
  assign w17001 = ( w4609 & w16998 ) | ( w4609 & w17000 ) | ( w16998 & w17000 ) ;
  assign w17002 = ( w16685 & ~w16999 ) | ( w16685 & w17001 ) | ( ~w16999 & w17001 ) ;
  assign w17003 = \pi23 ^ w17002 ;
  assign w17004 = w16848 ^ w16856 ;
  assign w17005 = ( \pi23 & \pi24 ) | ( \pi23 & ~w16696 ) | ( \pi24 & ~w16696 ) ;
  assign w17006 = ( \pi23 & \pi24 ) | ( \pi23 & ~w16698 ) | ( \pi24 & ~w16698 ) ;
  assign w17007 = \pi25 ^ w16698 ;
  assign w17008 = ( \pi25 & w17006 ) | ( \pi25 & w17007 ) | ( w17006 & w17007 ) ;
  assign w17009 = w17005 ^ w17008 ;
  assign w17010 = w4606 & w16694 ;
  assign w17011 = ( w4706 & ~w16690 ) | ( w4706 & w17010 ) | ( ~w16690 & w17010 ) ;
  assign w17012 = w4651 | w17011 ;
  assign w17013 = ( ~w16692 & w17011 ) | ( ~w16692 & w17012 ) | ( w17011 & w17012 ) ;
  assign w17014 = w17010 | w17013 ;
  assign w17015 = w4609 | w16839 ;
  assign w17016 = ( ~w16839 & w17014 ) | ( ~w16839 & w17015 ) | ( w17014 & w17015 ) ;
  assign w17017 = \pi23 ^ w17016 ;
  assign w17018 = \pi23 & w16698 ;
  assign w17019 = w16696 & w17018 ;
  assign w17020 = ( \pi20 & \pi21 ) | ( \pi20 & ~w17019 ) | ( \pi21 & ~w17019 ) ;
  assign w17021 = ( \pi22 & \pi23 ) | ( \pi22 & ~w17020 ) | ( \pi23 & ~w17020 ) ;
  assign w17022 = ( \pi22 & ~w17018 ) | ( \pi22 & w17020 ) | ( ~w17018 & w17020 ) ;
  assign w17023 = ( w7331 & w17021 ) | ( w7331 & ~w17022 ) | ( w17021 & ~w17022 ) ;
  assign w17024 = w4606 & ~w16698 ;
  assign w17025 = ( w4706 & w16694 ) | ( w4706 & w17024 ) | ( w16694 & w17024 ) ;
  assign w17026 = w4651 | w17025 ;
  assign w17027 = ( ~w16696 & w17025 ) | ( ~w16696 & w17026 ) | ( w17025 & w17026 ) ;
  assign w17028 = w17024 | w17027 ;
  assign w17029 = ~w4609 & w16802 ;
  assign w17030 = ( w16802 & w17028 ) | ( w16802 & ~w17029 ) | ( w17028 & ~w17029 ) ;
  assign w17031 = \pi23 ^ w17030 ;
  assign w17032 = w17023 & w17031 ;
  assign w17033 = ~w4651 & w16694 ;
  assign w17034 = w4606 & ~w16696 ;
  assign w17035 = ( w16694 & ~w17033 ) | ( w16694 & w17034 ) | ( ~w17033 & w17034 ) ;
  assign w17036 = w4706 | w16692 ;
  assign w17037 = w16784 | w17035 ;
  assign w17038 = ( w4609 & w17035 ) | ( w4609 & w17037 ) | ( w17035 & w17037 ) ;
  assign w17039 = ( ~w16692 & w17036 ) | ( ~w16692 & w17038 ) | ( w17036 & w17038 ) ;
  assign w17040 = \pi23 ^ w17039 ;
  assign w17041 = w2832 & ~w16698 ;
  assign w17042 = ( w17032 & w17040 ) | ( w17032 & w17041 ) | ( w17040 & w17041 ) ;
  assign w17043 = ( w17009 & w17017 ) | ( w17009 & w17042 ) | ( w17017 & w17042 ) ;
  assign w17044 = ( w17003 & w17004 ) | ( w17003 & w17043 ) | ( w17004 & w17043 ) ;
  assign w17045 = ( w16987 & w16995 ) | ( w16987 & w17044 ) | ( w16995 & w17044 ) ;
  assign w17046 = ( w16983 & w16985 ) | ( w16983 & w17045 ) | ( w16985 & w17045 ) ;
  assign w17047 = ( w16965 & w16975 ) | ( w16965 & w17046 ) | ( w16975 & w17046 ) ;
  assign w17048 = ( w16953 & w16963 ) | ( w16953 & w17047 ) | ( w16963 & w17047 ) ;
  assign w17049 = w16767 ^ w17048 ;
  assign w17050 = w16951 ^ w17049 ;
  assign w17051 = w4905 & w16660 ;
  assign w17052 = ( w5395 & ~w16656 ) | ( w5395 & w17051 ) | ( ~w16656 & w17051 ) ;
  assign w17053 = w5343 | w17052 ;
  assign w17054 = ( ~w16658 & w17052 ) | ( ~w16658 & w17053 ) | ( w17052 & w17053 ) ;
  assign w17055 = w17051 | w17054 ;
  assign w17056 = w16656 ^ w16710 ;
  assign w17057 = w16658 ^ w17056 ;
  assign w17058 = w4908 & ~w17057 ;
  assign w17059 = ( w4908 & w17055 ) | ( w4908 & ~w17058 ) | ( w17055 & ~w17058 ) ;
  assign w17060 = \pi20 ^ w17059 ;
  assign w17061 = ~w5343 & w16660 ;
  assign w17062 = w4905 & ~w16662 ;
  assign w17063 = ( w16660 & ~w17061 ) | ( w16660 & w17062 ) | ( ~w17061 & w17062 ) ;
  assign w17064 = w16658 ^ w16709 ;
  assign w17065 = w16660 ^ w17064 ;
  assign w17066 = w5395 | w16658 ;
  assign w17067 = ~w17063 & w17065 ;
  assign w17068 = ( w4908 & w17063 ) | ( w4908 & ~w17067 ) | ( w17063 & ~w17067 ) ;
  assign w17069 = ( ~w16658 & w17066 ) | ( ~w16658 & w17068 ) | ( w17066 & w17068 ) ;
  assign w17070 = \pi20 ^ w17069 ;
  assign w17071 = w16963 ^ w17047 ;
  assign w17072 = w16953 ^ w17071 ;
  assign w17073 = w5343 | w16662 ;
  assign w17074 = w4905 & w16665 ;
  assign w17075 = ( ~w16662 & w17073 ) | ( ~w16662 & w17074 ) | ( w17073 & w17074 ) ;
  assign w17076 = ( ~w16662 & w16665 ) | ( ~w16662 & w16707 ) | ( w16665 & w16707 ) ;
  assign w17077 = w16662 ^ w17076 ;
  assign w17078 = w16660 ^ w17077 ;
  assign w17079 = ~w5395 & w16660 ;
  assign w17080 = ~w17075 & w17078 ;
  assign w17081 = ( w4908 & w17075 ) | ( w4908 & ~w17080 ) | ( w17075 & ~w17080 ) ;
  assign w17082 = ( w16660 & ~w17079 ) | ( w16660 & w17081 ) | ( ~w17079 & w17081 ) ;
  assign w17083 = \pi20 ^ w17082 ;
  assign w17084 = w16975 ^ w17046 ;
  assign w17085 = w16965 ^ w17084 ;
  assign w17086 = w16983 ^ w17045 ;
  assign w17087 = w16985 ^ w17086 ;
  assign w17088 = w4905 & w16670 ;
  assign w17089 = ( w5395 & ~w16662 ) | ( w5395 & w17088 ) | ( ~w16662 & w17088 ) ;
  assign w17090 = w5343 | w17089 ;
  assign w17091 = ( w16665 & w17089 ) | ( w16665 & w17090 ) | ( w17089 & w17090 ) ;
  assign w17092 = w17088 | w17091 ;
  assign w17093 = w4908 | w16762 ;
  assign w17094 = ( ~w16762 & w17092 ) | ( ~w16762 & w17093 ) | ( w17092 & w17093 ) ;
  assign w17095 = \pi20 ^ w17094 ;
  assign w17096 = w16995 ^ w17044 ;
  assign w17097 = w16987 ^ w17096 ;
  assign w17098 = w4905 & w16675 ;
  assign w17099 = ( w5395 & w16665 ) | ( w5395 & w17098 ) | ( w16665 & w17098 ) ;
  assign w17100 = w5343 | w17099 ;
  assign w17101 = ( w16670 & w17099 ) | ( w16670 & w17100 ) | ( w17099 & w17100 ) ;
  assign w17102 = w17098 | w17101 ;
  assign w17103 = ~w4908 & w16960 ;
  assign w17104 = ( w16960 & w17102 ) | ( w16960 & ~w17103 ) | ( w17102 & ~w17103 ) ;
  assign w17105 = \pi20 ^ w17104 ;
  assign w17106 = w17003 ^ w17043 ;
  assign w17107 = w17004 ^ w17106 ;
  assign w17108 = w4905 & w16680 ;
  assign w17109 = ( w5395 & w16670 ) | ( w5395 & w17108 ) | ( w16670 & w17108 ) ;
  assign w17110 = w5343 | w17109 ;
  assign w17111 = ( w16675 & w17109 ) | ( w16675 & w17110 ) | ( w17109 & w17110 ) ;
  assign w17112 = w17108 | w17111 ;
  assign w17113 = ~w4908 & w16972 ;
  assign w17114 = ( w16972 & w17112 ) | ( w16972 & ~w17113 ) | ( w17112 & ~w17113 ) ;
  assign w17115 = \pi20 ^ w17114 ;
  assign w17116 = ~w5343 & w16680 ;
  assign w17117 = w4905 & w16685 ;
  assign w17118 = ( w16680 & ~w17116 ) | ( w16680 & w17117 ) | ( ~w17116 & w17117 ) ;
  assign w17119 = ~w5395 & w16675 ;
  assign w17120 = w16946 | w17118 ;
  assign w17121 = ( w4908 & w17118 ) | ( w4908 & w17120 ) | ( w17118 & w17120 ) ;
  assign w17122 = ( w16675 & ~w17119 ) | ( w16675 & w17121 ) | ( ~w17119 & w17121 ) ;
  assign w17123 = \pi20 ^ w17122 ;
  assign w17124 = w17017 ^ w17042 ;
  assign w17125 = w17009 ^ w17124 ;
  assign w17126 = w17032 ^ w17040 ;
  assign w17127 = w17041 ^ w17126 ;
  assign w17128 = w4905 & ~w16690 ;
  assign w17129 = ( w5395 & w16680 ) | ( w5395 & w17128 ) | ( w16680 & w17128 ) ;
  assign w17130 = w5343 | w17129 ;
  assign w17131 = ( w16685 & w17129 ) | ( w16685 & w17130 ) | ( w17129 & w17130 ) ;
  assign w17132 = w17128 | w17131 ;
  assign w17133 = w4908 | w16772 ;
  assign w17134 = ( ~w16772 & w17132 ) | ( ~w16772 & w17133 ) | ( w17132 & w17133 ) ;
  assign w17135 = \pi20 ^ w17134 ;
  assign w17136 = w5343 | w16690 ;
  assign w17137 = w4905 & ~w16692 ;
  assign w17138 = ( ~w16690 & w17136 ) | ( ~w16690 & w17137 ) | ( w17136 & w17137 ) ;
  assign w17139 = ~w5395 & w16685 ;
  assign w17140 = w16818 | w17138 ;
  assign w17141 = ( w4908 & w17138 ) | ( w4908 & w17140 ) | ( w17138 & w17140 ) ;
  assign w17142 = ( w16685 & ~w17139 ) | ( w16685 & w17141 ) | ( ~w17139 & w17141 ) ;
  assign w17143 = \pi20 ^ w17142 ;
  assign w17144 = w17023 ^ w17031 ;
  assign w17145 = ( \pi20 & \pi21 ) | ( \pi20 & ~w16696 ) | ( \pi21 & ~w16696 ) ;
  assign w17146 = ( \pi20 & \pi21 ) | ( \pi20 & ~w16698 ) | ( \pi21 & ~w16698 ) ;
  assign w17147 = \pi22 ^ w16698 ;
  assign w17148 = ( \pi22 & w17146 ) | ( \pi22 & w17147 ) | ( w17146 & w17147 ) ;
  assign w17149 = w17145 ^ w17148 ;
  assign w17150 = w4905 & w16694 ;
  assign w17151 = ( w5395 & ~w16690 ) | ( w5395 & w17150 ) | ( ~w16690 & w17150 ) ;
  assign w17152 = w5343 | w17151 ;
  assign w17153 = ( ~w16692 & w17151 ) | ( ~w16692 & w17152 ) | ( w17151 & w17152 ) ;
  assign w17154 = w17150 | w17153 ;
  assign w17155 = w4908 | w16839 ;
  assign w17156 = ( ~w16839 & w17154 ) | ( ~w16839 & w17155 ) | ( w17154 & w17155 ) ;
  assign w17157 = \pi20 ^ w17156 ;
  assign w17158 = \pi20 & w16698 ;
  assign w17159 = w16696 & w17158 ;
  assign w17160 = ( \pi17 & \pi18 ) | ( \pi17 & ~w17159 ) | ( \pi18 & ~w17159 ) ;
  assign w17161 = ( \pi19 & \pi20 ) | ( \pi19 & ~w17160 ) | ( \pi20 & ~w17160 ) ;
  assign w17162 = ( \pi19 & ~w17158 ) | ( \pi19 & w17160 ) | ( ~w17158 & w17160 ) ;
  assign w17163 = ( w7590 & w17161 ) | ( w7590 & ~w17162 ) | ( w17161 & ~w17162 ) ;
  assign w17164 = w4905 & ~w16698 ;
  assign w17165 = ( w5395 & w16694 ) | ( w5395 & w17164 ) | ( w16694 & w17164 ) ;
  assign w17166 = w5343 | w17165 ;
  assign w17167 = ( ~w16696 & w17165 ) | ( ~w16696 & w17166 ) | ( w17165 & w17166 ) ;
  assign w17168 = w17164 | w17167 ;
  assign w17169 = ~w4908 & w16802 ;
  assign w17170 = ( w16802 & w17168 ) | ( w16802 & ~w17169 ) | ( w17168 & ~w17169 ) ;
  assign w17171 = \pi20 ^ w17170 ;
  assign w17172 = w17163 & w17171 ;
  assign w17173 = ~w5343 & w16694 ;
  assign w17174 = w4905 & ~w16696 ;
  assign w17175 = ( w16694 & ~w17173 ) | ( w16694 & w17174 ) | ( ~w17173 & w17174 ) ;
  assign w17176 = w5395 | w16692 ;
  assign w17177 = w16784 | w17175 ;
  assign w17178 = ( w4908 & w17175 ) | ( w4908 & w17177 ) | ( w17175 & w17177 ) ;
  assign w17179 = ( ~w16692 & w17176 ) | ( ~w16692 & w17178 ) | ( w17176 & w17178 ) ;
  assign w17180 = \pi20 ^ w17179 ;
  assign w17181 = w4608 & ~w16698 ;
  assign w17182 = ( w17172 & w17180 ) | ( w17172 & w17181 ) | ( w17180 & w17181 ) ;
  assign w17183 = ( w17149 & w17157 ) | ( w17149 & w17182 ) | ( w17157 & w17182 ) ;
  assign w17184 = ( w17143 & w17144 ) | ( w17143 & w17183 ) | ( w17144 & w17183 ) ;
  assign w17185 = ( w17127 & w17135 ) | ( w17127 & w17184 ) | ( w17135 & w17184 ) ;
  assign w17186 = ( w17123 & w17125 ) | ( w17123 & w17185 ) | ( w17125 & w17185 ) ;
  assign w17187 = ( w17107 & w17115 ) | ( w17107 & w17186 ) | ( w17115 & w17186 ) ;
  assign w17188 = ( w17097 & w17105 ) | ( w17097 & w17187 ) | ( w17105 & w17187 ) ;
  assign w17189 = ( w17087 & w17095 ) | ( w17087 & w17188 ) | ( w17095 & w17188 ) ;
  assign w17190 = ( w17083 & w17085 ) | ( w17083 & w17189 ) | ( w17085 & w17189 ) ;
  assign w17191 = ( w17070 & w17072 ) | ( w17070 & w17190 ) | ( w17072 & w17190 ) ;
  assign w17192 = ( ~w17050 & w17060 ) | ( ~w17050 & w17191 ) | ( w17060 & w17191 ) ;
  assign w17193 = w4651 | w16662 ;
  assign w17194 = w4606 & w16665 ;
  assign w17195 = ( ~w16662 & w17193 ) | ( ~w16662 & w17194 ) | ( w17193 & w17194 ) ;
  assign w17196 = ~w4706 & w16660 ;
  assign w17197 = w17078 & ~w17195 ;
  assign w17198 = ( w4609 & w17195 ) | ( w4609 & ~w17197 ) | ( w17195 & ~w17197 ) ;
  assign w17199 = ( w16660 & ~w17196 ) | ( w16660 & w17198 ) | ( ~w17196 & w17198 ) ;
  assign w17200 = \pi23 ^ w17199 ;
  assign w17201 = ( w16870 & ~w16939 ) | ( w16870 & w16949 ) | ( ~w16939 & w16949 ) ;
  assign w17202 = w3717 | w16690 ;
  assign w17203 = w3649 & ~w16692 ;
  assign w17204 = ( ~w16690 & w17202 ) | ( ~w16690 & w17203 ) | ( w17202 & w17203 ) ;
  assign w17205 = ~w3549 & w16685 ;
  assign w17206 = w16818 | w17204 ;
  assign w17207 = ( w3448 & w17204 ) | ( w3448 & w17206 ) | ( w17204 & w17206 ) ;
  assign w17208 = ( w16685 & ~w17205 ) | ( w16685 & w17207 ) | ( ~w17205 & w17207 ) ;
  assign w17209 = \pi29 ^ w17208 ;
  assign w17210 = \pi31 & ~w16698 ;
  assign w17211 = w16694 ^ w17210 ;
  assign w17212 = ( \pi29 & \pi30 ) | ( \pi29 & w17211 ) | ( \pi30 & w17211 ) ;
  assign w17213 = \pi31 ^ w17212 ;
  assign w17214 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w16698 ) | ( \pi30 & w16698 ) ;
  assign w17215 = w6462 & ~w17214 ;
  assign w17216 = ( ~w16696 & w17213 ) | ( ~w16696 & w17215 ) | ( w17213 & w17215 ) ;
  assign w17217 = w36 & w16694 ;
  assign w17218 = ( w16696 & w17215 ) | ( w16696 & w17217 ) | ( w17215 & w17217 ) ;
  assign w17219 = w17216 | w17218 ;
  assign w17220 = w210 | w316 ;
  assign w17221 = w98 | w17220 ;
  assign w17222 = ( w51 & ~w98 ) | ( w51 & w113 ) | ( ~w98 & w113 ) ;
  assign w17223 = w17221 | w17222 ;
  assign w17224 = w358 | w470 ;
  assign w17225 = w3115 | w17224 ;
  assign w17226 = ( ~w3115 & w9856 ) | ( ~w3115 & w17223 ) | ( w9856 & w17223 ) ;
  assign w17227 = w17225 | w17226 ;
  assign w17228 = ( w276 & ~w987 ) | ( w276 & w5161 ) | ( ~w987 & w5161 ) ;
  assign w17229 = w6262 | w17227 ;
  assign w17230 = ( w276 & w3350 ) | ( w276 & ~w17227 ) | ( w3350 & ~w17227 ) ;
  assign w17231 = w17229 | w17230 ;
  assign w17232 = w17228 & ~w17231 ;
  assign w17233 = w413 | w1155 ;
  assign w17234 = w12599 | w17233 ;
  assign w17235 = ( ~w742 & w12599 ) | ( ~w742 & w17232 ) | ( w12599 & w17232 ) ;
  assign w17236 = ~w17234 & w17235 ;
  assign w17237 = ( w262 & w569 ) | ( w262 & ~w681 ) | ( w569 & ~w681 ) ;
  assign w17238 = ~w205 & w17236 ;
  assign w17239 = ( ~w205 & w681 ) | ( ~w205 & w1001 ) | ( w681 & w1001 ) ;
  assign w17240 = w17238 & ~w17239 ;
  assign w17241 = ~w17237 & w17240 ;
  assign w17242 = w16935 ^ w17219 ;
  assign w17243 = w17241 ^ w17242 ;
  assign w17244 = ( w16878 & ~w16936 ) | ( w16878 & w16937 ) | ( ~w16936 & w16937 ) ;
  assign w17245 = w17209 ^ w17244 ;
  assign w17246 = w17243 ^ w17245 ;
  assign w17247 = w3964 & w16670 ;
  assign w17248 = ( w4143 & w16675 ) | ( w4143 & w17247 ) | ( w16675 & w17247 ) ;
  assign w17249 = w4052 | w17248 ;
  assign w17250 = ( w16680 & w17248 ) | ( w16680 & w17249 ) | ( w17248 & w17249 ) ;
  assign w17251 = w17247 | w17250 ;
  assign w17252 = ~w4147 & w16972 ;
  assign w17253 = ( w16972 & w17251 ) | ( w16972 & ~w17252 ) | ( w17251 & ~w17252 ) ;
  assign w17254 = \pi26 ^ w17253 ;
  assign w17255 = w17201 ^ w17254 ;
  assign w17256 = w17246 ^ w17255 ;
  assign w17257 = ( w16767 & ~w16951 ) | ( w16767 & w17048 ) | ( ~w16951 & w17048 ) ;
  assign w17258 = w17200 ^ w17257 ;
  assign w17259 = w17256 ^ w17258 ;
  assign w17260 = w4905 & ~w16658 ;
  assign w17261 = ( w5395 & w16654 ) | ( w5395 & w17260 ) | ( w16654 & w17260 ) ;
  assign w17262 = w5343 | w17261 ;
  assign w17263 = ( ~w16656 & w17261 ) | ( ~w16656 & w17262 ) | ( w17261 & w17262 ) ;
  assign w17264 = w17260 | w17263 ;
  assign w17265 = w16654 ^ w16711 ;
  assign w17266 = w16656 ^ w17265 ;
  assign w17267 = w4908 & ~w17266 ;
  assign w17268 = ( w4908 & w17264 ) | ( w4908 & ~w17267 ) | ( w17264 & ~w17267 ) ;
  assign w17269 = \pi20 ^ w17268 ;
  assign w17270 = w17192 ^ w17269 ;
  assign w17271 = w17259 ^ w17270 ;
  assign w17272 = w5710 | w16652 ;
  assign w17273 = w5494 & w16654 ;
  assign w17274 = ( ~w16652 & w17272 ) | ( ~w16652 & w17273 ) | ( w17272 & w17273 ) ;
  assign w17275 = ( w16652 & ~w16654 ) | ( w16652 & w16712 ) | ( ~w16654 & w16712 ) ;
  assign w17276 = w16652 ^ w17275 ;
  assign w17277 = w16650 ^ w17276 ;
  assign w17278 = w5948 | w16650 ;
  assign w17279 = ~w17274 & w17277 ;
  assign w17280 = ( w5497 & w17274 ) | ( w5497 & ~w17279 ) | ( w17274 & ~w17279 ) ;
  assign w17281 = ( ~w16650 & w17278 ) | ( ~w16650 & w17280 ) | ( w17278 & w17280 ) ;
  assign w17282 = \pi17 ^ w17281 ;
  assign w17283 = w17060 ^ w17191 ;
  assign w17284 = w17050 ^ w17283 ;
  assign w17285 = w17070 ^ w17190 ;
  assign w17286 = w17072 ^ w17285 ;
  assign w17287 = w5494 & ~w16656 ;
  assign w17288 = ( w5948 & ~w16652 ) | ( w5948 & w17287 ) | ( ~w16652 & w17287 ) ;
  assign w17289 = w5710 | w17288 ;
  assign w17290 = ( w16654 & w17288 ) | ( w16654 & w17289 ) | ( w17288 & w17289 ) ;
  assign w17291 = w17287 | w17290 ;
  assign w17292 = w16652 ^ w16712 ;
  assign w17293 = w16654 ^ w17292 ;
  assign w17294 = w5497 & ~w17293 ;
  assign w17295 = ( w5497 & w17291 ) | ( w5497 & ~w17294 ) | ( w17291 & ~w17294 ) ;
  assign w17296 = \pi17 ^ w17295 ;
  assign w17297 = w17083 ^ w17189 ;
  assign w17298 = w17085 ^ w17297 ;
  assign w17299 = w5494 & ~w16658 ;
  assign w17300 = ( w5948 & w16654 ) | ( w5948 & w17299 ) | ( w16654 & w17299 ) ;
  assign w17301 = w5710 | w17300 ;
  assign w17302 = ( ~w16656 & w17300 ) | ( ~w16656 & w17301 ) | ( w17300 & w17301 ) ;
  assign w17303 = w17299 | w17302 ;
  assign w17304 = ~w5497 & w17266 ;
  assign w17305 = ( w17266 & w17303 ) | ( w17266 & ~w17304 ) | ( w17303 & ~w17304 ) ;
  assign w17306 = \pi17 ^ w17305 ;
  assign w17307 = w5710 | w16658 ;
  assign w17308 = w5494 & w16660 ;
  assign w17309 = ( ~w16658 & w17307 ) | ( ~w16658 & w17308 ) | ( w17307 & w17308 ) ;
  assign w17310 = w5948 | w16656 ;
  assign w17311 = w17057 | w17309 ;
  assign w17312 = ( w5497 & w17309 ) | ( w5497 & w17311 ) | ( w17309 & w17311 ) ;
  assign w17313 = ( ~w16656 & w17310 ) | ( ~w16656 & w17312 ) | ( w17310 & w17312 ) ;
  assign w17314 = \pi17 ^ w17313 ;
  assign w17315 = w17095 ^ w17188 ;
  assign w17316 = w17087 ^ w17315 ;
  assign w17317 = ~w5710 & w16660 ;
  assign w17318 = w5494 & ~w16662 ;
  assign w17319 = ( w16660 & ~w17317 ) | ( w16660 & w17318 ) | ( ~w17317 & w17318 ) ;
  assign w17320 = w5948 | w16658 ;
  assign w17321 = w17065 & ~w17319 ;
  assign w17322 = ( w5497 & w17319 ) | ( w5497 & ~w17321 ) | ( w17319 & ~w17321 ) ;
  assign w17323 = ( ~w16658 & w17320 ) | ( ~w16658 & w17322 ) | ( w17320 & w17322 ) ;
  assign w17324 = \pi17 ^ w17323 ;
  assign w17325 = w17105 ^ w17187 ;
  assign w17326 = w17097 ^ w17325 ;
  assign w17327 = w5710 | w16662 ;
  assign w17328 = w5494 & w16665 ;
  assign w17329 = ( ~w16662 & w17327 ) | ( ~w16662 & w17328 ) | ( w17327 & w17328 ) ;
  assign w17330 = ~w5948 & w16660 ;
  assign w17331 = w17078 & ~w17329 ;
  assign w17332 = ( w5497 & w17329 ) | ( w5497 & ~w17331 ) | ( w17329 & ~w17331 ) ;
  assign w17333 = ( w16660 & ~w17330 ) | ( w16660 & w17332 ) | ( ~w17330 & w17332 ) ;
  assign w17334 = \pi17 ^ w17333 ;
  assign w17335 = w17115 ^ w17186 ;
  assign w17336 = w17107 ^ w17335 ;
  assign w17337 = w17123 ^ w17185 ;
  assign w17338 = w17125 ^ w17337 ;
  assign w17339 = w5494 & w16670 ;
  assign w17340 = ( w5948 & ~w16662 ) | ( w5948 & w17339 ) | ( ~w16662 & w17339 ) ;
  assign w17341 = w5710 | w17340 ;
  assign w17342 = ( w16665 & w17340 ) | ( w16665 & w17341 ) | ( w17340 & w17341 ) ;
  assign w17343 = w17339 | w17342 ;
  assign w17344 = w5497 | w16762 ;
  assign w17345 = ( ~w16762 & w17343 ) | ( ~w16762 & w17344 ) | ( w17343 & w17344 ) ;
  assign w17346 = \pi17 ^ w17345 ;
  assign w17347 = w17135 ^ w17184 ;
  assign w17348 = w17127 ^ w17347 ;
  assign w17349 = w5494 & w16675 ;
  assign w17350 = ( w5948 & w16665 ) | ( w5948 & w17349 ) | ( w16665 & w17349 ) ;
  assign w17351 = w5710 | w17350 ;
  assign w17352 = ( w16670 & w17350 ) | ( w16670 & w17351 ) | ( w17350 & w17351 ) ;
  assign w17353 = w17349 | w17352 ;
  assign w17354 = ~w5497 & w16960 ;
  assign w17355 = ( w16960 & w17353 ) | ( w16960 & ~w17354 ) | ( w17353 & ~w17354 ) ;
  assign w17356 = \pi17 ^ w17355 ;
  assign w17357 = w17143 ^ w17183 ;
  assign w17358 = w17144 ^ w17357 ;
  assign w17359 = w5494 & w16680 ;
  assign w17360 = ( w5948 & w16670 ) | ( w5948 & w17359 ) | ( w16670 & w17359 ) ;
  assign w17361 = w5710 | w17360 ;
  assign w17362 = ( w16675 & w17360 ) | ( w16675 & w17361 ) | ( w17360 & w17361 ) ;
  assign w17363 = w17359 | w17362 ;
  assign w17364 = ~w5497 & w16972 ;
  assign w17365 = ( w16972 & w17363 ) | ( w16972 & ~w17364 ) | ( w17363 & ~w17364 ) ;
  assign w17366 = \pi17 ^ w17365 ;
  assign w17367 = ~w5710 & w16680 ;
  assign w17368 = w5494 & w16685 ;
  assign w17369 = ( w16680 & ~w17367 ) | ( w16680 & w17368 ) | ( ~w17367 & w17368 ) ;
  assign w17370 = ~w5948 & w16675 ;
  assign w17371 = w16946 | w17369 ;
  assign w17372 = ( w5497 & w17369 ) | ( w5497 & w17371 ) | ( w17369 & w17371 ) ;
  assign w17373 = ( w16675 & ~w17370 ) | ( w16675 & w17372 ) | ( ~w17370 & w17372 ) ;
  assign w17374 = \pi17 ^ w17373 ;
  assign w17375 = w17157 ^ w17182 ;
  assign w17376 = w17149 ^ w17375 ;
  assign w17377 = w17172 ^ w17180 ;
  assign w17378 = w17181 ^ w17377 ;
  assign w17379 = w5494 & ~w16690 ;
  assign w17380 = ( w5948 & w16680 ) | ( w5948 & w17379 ) | ( w16680 & w17379 ) ;
  assign w17381 = w5710 | w17380 ;
  assign w17382 = ( w16685 & w17380 ) | ( w16685 & w17381 ) | ( w17380 & w17381 ) ;
  assign w17383 = w17379 | w17382 ;
  assign w17384 = w5497 | w16772 ;
  assign w17385 = ( ~w16772 & w17383 ) | ( ~w16772 & w17384 ) | ( w17383 & w17384 ) ;
  assign w17386 = \pi17 ^ w17385 ;
  assign w17387 = w5710 | w16690 ;
  assign w17388 = w5494 & ~w16692 ;
  assign w17389 = ( ~w16690 & w17387 ) | ( ~w16690 & w17388 ) | ( w17387 & w17388 ) ;
  assign w17390 = ~w5948 & w16685 ;
  assign w17391 = w16818 | w17389 ;
  assign w17392 = ( w5497 & w17389 ) | ( w5497 & w17391 ) | ( w17389 & w17391 ) ;
  assign w17393 = ( w16685 & ~w17390 ) | ( w16685 & w17392 ) | ( ~w17390 & w17392 ) ;
  assign w17394 = \pi17 ^ w17393 ;
  assign w17395 = w17163 ^ w17171 ;
  assign w17396 = ( \pi17 & \pi18 ) | ( \pi17 & ~w16696 ) | ( \pi18 & ~w16696 ) ;
  assign w17397 = ( \pi17 & \pi18 ) | ( \pi17 & ~w16698 ) | ( \pi18 & ~w16698 ) ;
  assign w17398 = \pi19 ^ w16698 ;
  assign w17399 = ( \pi19 & w17397 ) | ( \pi19 & w17398 ) | ( w17397 & w17398 ) ;
  assign w17400 = w17396 ^ w17399 ;
  assign w17401 = w5494 & w16694 ;
  assign w17402 = ( w5948 & ~w16690 ) | ( w5948 & w17401 ) | ( ~w16690 & w17401 ) ;
  assign w17403 = w5710 | w17402 ;
  assign w17404 = ( ~w16692 & w17402 ) | ( ~w16692 & w17403 ) | ( w17402 & w17403 ) ;
  assign w17405 = w17401 | w17404 ;
  assign w17406 = w5497 | w16839 ;
  assign w17407 = ( ~w16839 & w17405 ) | ( ~w16839 & w17406 ) | ( w17405 & w17406 ) ;
  assign w17408 = \pi17 ^ w17407 ;
  assign w17409 = \pi17 & w16698 ;
  assign w17410 = w16696 & w17409 ;
  assign w17411 = ( \pi14 & \pi15 ) | ( \pi14 & ~w17410 ) | ( \pi15 & ~w17410 ) ;
  assign w17412 = ( \pi16 & \pi17 ) | ( \pi16 & ~w17411 ) | ( \pi17 & ~w17411 ) ;
  assign w17413 = ( \pi16 & ~w17409 ) | ( \pi16 & w17411 ) | ( ~w17409 & w17411 ) ;
  assign w17414 = ( w7879 & w17412 ) | ( w7879 & ~w17413 ) | ( w17412 & ~w17413 ) ;
  assign w17415 = w5494 & ~w16698 ;
  assign w17416 = ( w5948 & w16694 ) | ( w5948 & w17415 ) | ( w16694 & w17415 ) ;
  assign w17417 = w5710 | w17416 ;
  assign w17418 = ( ~w16696 & w17416 ) | ( ~w16696 & w17417 ) | ( w17416 & w17417 ) ;
  assign w17419 = w17415 | w17418 ;
  assign w17420 = ~w5497 & w16802 ;
  assign w17421 = ( w16802 & w17419 ) | ( w16802 & ~w17420 ) | ( w17419 & ~w17420 ) ;
  assign w17422 = \pi17 ^ w17421 ;
  assign w17423 = w17414 & w17422 ;
  assign w17424 = ~w5710 & w16694 ;
  assign w17425 = w5494 & ~w16696 ;
  assign w17426 = ( w16694 & ~w17424 ) | ( w16694 & w17425 ) | ( ~w17424 & w17425 ) ;
  assign w17427 = w5948 | w16692 ;
  assign w17428 = w16784 | w17426 ;
  assign w17429 = ( w5497 & w17426 ) | ( w5497 & w17428 ) | ( w17426 & w17428 ) ;
  assign w17430 = ( ~w16692 & w17427 ) | ( ~w16692 & w17429 ) | ( w17427 & w17429 ) ;
  assign w17431 = \pi17 ^ w17430 ;
  assign w17432 = w4907 & ~w16698 ;
  assign w17433 = ( w17423 & w17431 ) | ( w17423 & w17432 ) | ( w17431 & w17432 ) ;
  assign w17434 = ( w17400 & w17408 ) | ( w17400 & w17433 ) | ( w17408 & w17433 ) ;
  assign w17435 = ( w17394 & w17395 ) | ( w17394 & w17434 ) | ( w17395 & w17434 ) ;
  assign w17436 = ( w17378 & w17386 ) | ( w17378 & w17435 ) | ( w17386 & w17435 ) ;
  assign w17437 = ( w17374 & w17376 ) | ( w17374 & w17436 ) | ( w17376 & w17436 ) ;
  assign w17438 = ( w17358 & w17366 ) | ( w17358 & w17437 ) | ( w17366 & w17437 ) ;
  assign w17439 = ( w17348 & w17356 ) | ( w17348 & w17438 ) | ( w17356 & w17438 ) ;
  assign w17440 = ( w17338 & w17346 ) | ( w17338 & w17439 ) | ( w17346 & w17439 ) ;
  assign w17441 = ( w17334 & w17336 ) | ( w17334 & w17440 ) | ( w17336 & w17440 ) ;
  assign w17442 = ( w17324 & w17326 ) | ( w17324 & w17441 ) | ( w17326 & w17441 ) ;
  assign w17443 = ( w17314 & w17316 ) | ( w17314 & w17442 ) | ( w17316 & w17442 ) ;
  assign w17444 = ( w17298 & w17306 ) | ( w17298 & w17443 ) | ( w17306 & w17443 ) ;
  assign w17445 = ( w17286 & w17296 ) | ( w17286 & w17444 ) | ( w17296 & w17444 ) ;
  assign w17446 = ( w17282 & ~w17284 ) | ( w17282 & w17445 ) | ( ~w17284 & w17445 ) ;
  assign w17447 = w16757 ^ w17446 ;
  assign w17448 = w17271 ^ w17447 ;
  assign w17449 = w6048 & ~w16646 ;
  assign w17450 = ( w6637 & w16642 ) | ( w6637 & w17449 ) | ( w16642 & w17449 ) ;
  assign w17451 = w6549 | w17450 ;
  assign w17452 = ( ~w16644 & w17450 ) | ( ~w16644 & w17451 ) | ( w17450 & w17451 ) ;
  assign w17453 = w17449 | w17452 ;
  assign w17454 = w16642 ^ w16717 ;
  assign w17455 = w16644 ^ w17454 ;
  assign w17456 = w6045 & ~w17455 ;
  assign w17457 = ( w6045 & w17453 ) | ( w6045 & ~w17456 ) | ( w17453 & ~w17456 ) ;
  assign w17458 = \pi14 ^ w17457 ;
  assign w17459 = w17282 ^ w17445 ;
  assign w17460 = w17284 ^ w17459 ;
  assign w17461 = w6048 & ~w16648 ;
  assign w17462 = ( w6637 & ~w16644 ) | ( w6637 & w17461 ) | ( ~w16644 & w17461 ) ;
  assign w17463 = w6549 | w17462 ;
  assign w17464 = ( ~w16646 & w17462 ) | ( ~w16646 & w17463 ) | ( w17462 & w17463 ) ;
  assign w17465 = w17461 | w17464 ;
  assign w17466 = ( w16646 & w16648 ) | ( w16646 & w16715 ) | ( w16648 & w16715 ) ;
  assign w17467 = w16646 ^ w17466 ;
  assign w17468 = w16644 ^ w17467 ;
  assign w17469 = w6045 & w17468 ;
  assign w17470 = ( w6045 & w17465 ) | ( w6045 & ~w17469 ) | ( w17465 & ~w17469 ) ;
  assign w17471 = \pi14 ^ w17470 ;
  assign w17472 = w6549 | w16648 ;
  assign w17473 = w6048 & ~w16650 ;
  assign w17474 = ( ~w16648 & w17472 ) | ( ~w16648 & w17473 ) | ( w17472 & w17473 ) ;
  assign w17475 = w16646 ^ w16715 ;
  assign w17476 = w16648 ^ w17475 ;
  assign w17477 = w6637 | w16646 ;
  assign w17478 = ~w17474 & w17476 ;
  assign w17479 = ( w6045 & w17474 ) | ( w6045 & ~w17478 ) | ( w17474 & ~w17478 ) ;
  assign w17480 = ( ~w16646 & w17477 ) | ( ~w16646 & w17479 ) | ( w17477 & w17479 ) ;
  assign w17481 = \pi14 ^ w17480 ;
  assign w17482 = w17296 ^ w17444 ;
  assign w17483 = w17286 ^ w17482 ;
  assign w17484 = w6549 | w16650 ;
  assign w17485 = w6048 & ~w16652 ;
  assign w17486 = ( ~w16650 & w17484 ) | ( ~w16650 & w17485 ) | ( w17484 & w17485 ) ;
  assign w17487 = w6637 | w16648 ;
  assign w17488 = w16752 & ~w17486 ;
  assign w17489 = ( w6045 & w17486 ) | ( w6045 & ~w17488 ) | ( w17486 & ~w17488 ) ;
  assign w17490 = ( ~w16648 & w17487 ) | ( ~w16648 & w17489 ) | ( w17487 & w17489 ) ;
  assign w17491 = \pi14 ^ w17490 ;
  assign w17492 = w17306 ^ w17443 ;
  assign w17493 = w17298 ^ w17492 ;
  assign w17494 = w17314 ^ w17442 ;
  assign w17495 = w17316 ^ w17494 ;
  assign w17496 = w6048 & w16654 ;
  assign w17497 = ( w6637 & ~w16650 ) | ( w6637 & w17496 ) | ( ~w16650 & w17496 ) ;
  assign w17498 = w6549 | w17497 ;
  assign w17499 = ( ~w16652 & w17497 ) | ( ~w16652 & w17498 ) | ( w17497 & w17498 ) ;
  assign w17500 = w17496 | w17499 ;
  assign w17501 = w6045 | w17277 ;
  assign w17502 = ( ~w17277 & w17500 ) | ( ~w17277 & w17501 ) | ( w17500 & w17501 ) ;
  assign w17503 = \pi14 ^ w17502 ;
  assign w17504 = w17324 ^ w17441 ;
  assign w17505 = w17326 ^ w17504 ;
  assign w17506 = w6048 & ~w16656 ;
  assign w17507 = ( w6637 & ~w16652 ) | ( w6637 & w17506 ) | ( ~w16652 & w17506 ) ;
  assign w17508 = w6549 | w17507 ;
  assign w17509 = ( w16654 & w17507 ) | ( w16654 & w17508 ) | ( w17507 & w17508 ) ;
  assign w17510 = w17506 | w17509 ;
  assign w17511 = ~w6045 & w17293 ;
  assign w17512 = ( w17293 & w17510 ) | ( w17293 & ~w17511 ) | ( w17510 & ~w17511 ) ;
  assign w17513 = \pi14 ^ w17512 ;
  assign w17514 = w17334 ^ w17440 ;
  assign w17515 = w17336 ^ w17514 ;
  assign w17516 = w6048 & ~w16658 ;
  assign w17517 = ( w6637 & w16654 ) | ( w6637 & w17516 ) | ( w16654 & w17516 ) ;
  assign w17518 = w6549 | w17517 ;
  assign w17519 = ( ~w16656 & w17517 ) | ( ~w16656 & w17518 ) | ( w17517 & w17518 ) ;
  assign w17520 = w17516 | w17519 ;
  assign w17521 = ~w6045 & w17266 ;
  assign w17522 = ( w17266 & w17520 ) | ( w17266 & ~w17521 ) | ( w17520 & ~w17521 ) ;
  assign w17523 = \pi14 ^ w17522 ;
  assign w17524 = w6549 | w16658 ;
  assign w17525 = w6048 & w16660 ;
  assign w17526 = ( ~w16658 & w17524 ) | ( ~w16658 & w17525 ) | ( w17524 & w17525 ) ;
  assign w17527 = w6637 | w16656 ;
  assign w17528 = w17057 | w17526 ;
  assign w17529 = ( w6045 & w17526 ) | ( w6045 & w17528 ) | ( w17526 & w17528 ) ;
  assign w17530 = ( ~w16656 & w17527 ) | ( ~w16656 & w17529 ) | ( w17527 & w17529 ) ;
  assign w17531 = \pi14 ^ w17530 ;
  assign w17532 = w17346 ^ w17439 ;
  assign w17533 = w17338 ^ w17532 ;
  assign w17534 = ~w6549 & w16660 ;
  assign w17535 = w6048 & ~w16662 ;
  assign w17536 = ( w16660 & ~w17534 ) | ( w16660 & w17535 ) | ( ~w17534 & w17535 ) ;
  assign w17537 = w6637 | w16658 ;
  assign w17538 = w17065 & ~w17536 ;
  assign w17539 = ( w6045 & w17536 ) | ( w6045 & ~w17538 ) | ( w17536 & ~w17538 ) ;
  assign w17540 = ( ~w16658 & w17537 ) | ( ~w16658 & w17539 ) | ( w17537 & w17539 ) ;
  assign w17541 = \pi14 ^ w17540 ;
  assign w17542 = w17356 ^ w17438 ;
  assign w17543 = w17348 ^ w17542 ;
  assign w17544 = w6549 | w16662 ;
  assign w17545 = w6048 & w16665 ;
  assign w17546 = ( ~w16662 & w17544 ) | ( ~w16662 & w17545 ) | ( w17544 & w17545 ) ;
  assign w17547 = ~w6637 & w16660 ;
  assign w17548 = w17078 & ~w17546 ;
  assign w17549 = ( w6045 & w17546 ) | ( w6045 & ~w17548 ) | ( w17546 & ~w17548 ) ;
  assign w17550 = ( w16660 & ~w17547 ) | ( w16660 & w17549 ) | ( ~w17547 & w17549 ) ;
  assign w17551 = \pi14 ^ w17550 ;
  assign w17552 = w17366 ^ w17437 ;
  assign w17553 = w17358 ^ w17552 ;
  assign w17554 = w17374 ^ w17436 ;
  assign w17555 = w17376 ^ w17554 ;
  assign w17556 = w6048 & w16670 ;
  assign w17557 = ( w6637 & ~w16662 ) | ( w6637 & w17556 ) | ( ~w16662 & w17556 ) ;
  assign w17558 = w6549 | w17557 ;
  assign w17559 = ( w16665 & w17557 ) | ( w16665 & w17558 ) | ( w17557 & w17558 ) ;
  assign w17560 = w17556 | w17559 ;
  assign w17561 = w6045 | w16762 ;
  assign w17562 = ( ~w16762 & w17560 ) | ( ~w16762 & w17561 ) | ( w17560 & w17561 ) ;
  assign w17563 = \pi14 ^ w17562 ;
  assign w17564 = w17386 ^ w17435 ;
  assign w17565 = w17378 ^ w17564 ;
  assign w17566 = w6048 & w16675 ;
  assign w17567 = ( w6637 & w16665 ) | ( w6637 & w17566 ) | ( w16665 & w17566 ) ;
  assign w17568 = w6549 | w17567 ;
  assign w17569 = ( w16670 & w17567 ) | ( w16670 & w17568 ) | ( w17567 & w17568 ) ;
  assign w17570 = w17566 | w17569 ;
  assign w17571 = ~w6045 & w16960 ;
  assign w17572 = ( w16960 & w17570 ) | ( w16960 & ~w17571 ) | ( w17570 & ~w17571 ) ;
  assign w17573 = \pi14 ^ w17572 ;
  assign w17574 = w17394 ^ w17434 ;
  assign w17575 = w17395 ^ w17574 ;
  assign w17576 = w6048 & w16680 ;
  assign w17577 = ( w6637 & w16670 ) | ( w6637 & w17576 ) | ( w16670 & w17576 ) ;
  assign w17578 = w6549 | w17577 ;
  assign w17579 = ( w16675 & w17577 ) | ( w16675 & w17578 ) | ( w17577 & w17578 ) ;
  assign w17580 = w17576 | w17579 ;
  assign w17581 = ~w6045 & w16972 ;
  assign w17582 = ( w16972 & w17580 ) | ( w16972 & ~w17581 ) | ( w17580 & ~w17581 ) ;
  assign w17583 = \pi14 ^ w17582 ;
  assign w17584 = ~w6549 & w16680 ;
  assign w17585 = w6048 & w16685 ;
  assign w17586 = ( w16680 & ~w17584 ) | ( w16680 & w17585 ) | ( ~w17584 & w17585 ) ;
  assign w17587 = ~w6637 & w16675 ;
  assign w17588 = w16946 | w17586 ;
  assign w17589 = ( w6045 & w17586 ) | ( w6045 & w17588 ) | ( w17586 & w17588 ) ;
  assign w17590 = ( w16675 & ~w17587 ) | ( w16675 & w17589 ) | ( ~w17587 & w17589 ) ;
  assign w17591 = \pi14 ^ w17590 ;
  assign w17592 = w17408 ^ w17433 ;
  assign w17593 = w17400 ^ w17592 ;
  assign w17594 = w17423 ^ w17431 ;
  assign w17595 = w17432 ^ w17594 ;
  assign w17596 = w6048 & ~w16690 ;
  assign w17597 = ( w6637 & w16680 ) | ( w6637 & w17596 ) | ( w16680 & w17596 ) ;
  assign w17598 = w6549 | w17597 ;
  assign w17599 = ( w16685 & w17597 ) | ( w16685 & w17598 ) | ( w17597 & w17598 ) ;
  assign w17600 = w17596 | w17599 ;
  assign w17601 = w6045 | w16772 ;
  assign w17602 = ( ~w16772 & w17600 ) | ( ~w16772 & w17601 ) | ( w17600 & w17601 ) ;
  assign w17603 = \pi14 ^ w17602 ;
  assign w17604 = w6549 | w16690 ;
  assign w17605 = w6048 & ~w16692 ;
  assign w17606 = ( ~w16690 & w17604 ) | ( ~w16690 & w17605 ) | ( w17604 & w17605 ) ;
  assign w17607 = ~w6637 & w16685 ;
  assign w17608 = w16818 | w17606 ;
  assign w17609 = ( w6045 & w17606 ) | ( w6045 & w17608 ) | ( w17606 & w17608 ) ;
  assign w17610 = ( w16685 & ~w17607 ) | ( w16685 & w17609 ) | ( ~w17607 & w17609 ) ;
  assign w17611 = \pi14 ^ w17610 ;
  assign w17612 = w17414 ^ w17422 ;
  assign w17613 = ( \pi14 & \pi15 ) | ( \pi14 & ~w16696 ) | ( \pi15 & ~w16696 ) ;
  assign w17614 = ( \pi14 & \pi15 ) | ( \pi14 & ~w16698 ) | ( \pi15 & ~w16698 ) ;
  assign w17615 = \pi16 ^ w16698 ;
  assign w17616 = ( \pi16 & w17614 ) | ( \pi16 & w17615 ) | ( w17614 & w17615 ) ;
  assign w17617 = w17613 ^ w17616 ;
  assign w17618 = w6048 & w16694 ;
  assign w17619 = ( w6637 & ~w16690 ) | ( w6637 & w17618 ) | ( ~w16690 & w17618 ) ;
  assign w17620 = w6549 | w17619 ;
  assign w17621 = ( ~w16692 & w17619 ) | ( ~w16692 & w17620 ) | ( w17619 & w17620 ) ;
  assign w17622 = w17618 | w17621 ;
  assign w17623 = w6045 | w16839 ;
  assign w17624 = ( ~w16839 & w17622 ) | ( ~w16839 & w17623 ) | ( w17622 & w17623 ) ;
  assign w17625 = \pi14 ^ w17624 ;
  assign w17626 = \pi14 & w16698 ;
  assign w17627 = w16696 & w17626 ;
  assign w17628 = ( \pi11 & \pi12 ) | ( \pi11 & ~w17627 ) | ( \pi12 & ~w17627 ) ;
  assign w17629 = ( \pi13 & \pi14 ) | ( \pi13 & ~w17628 ) | ( \pi14 & ~w17628 ) ;
  assign w17630 = ( \pi13 & ~w17626 ) | ( \pi13 & w17628 ) | ( ~w17626 & w17628 ) ;
  assign w17631 = ( w8192 & w17629 ) | ( w8192 & ~w17630 ) | ( w17629 & ~w17630 ) ;
  assign w17632 = w6048 & ~w16698 ;
  assign w17633 = ( w6637 & w16694 ) | ( w6637 & w17632 ) | ( w16694 & w17632 ) ;
  assign w17634 = w6549 | w17633 ;
  assign w17635 = ( ~w16696 & w17633 ) | ( ~w16696 & w17634 ) | ( w17633 & w17634 ) ;
  assign w17636 = w17632 | w17635 ;
  assign w17637 = ~w6045 & w16802 ;
  assign w17638 = ( w16802 & w17636 ) | ( w16802 & ~w17637 ) | ( w17636 & ~w17637 ) ;
  assign w17639 = \pi14 ^ w17638 ;
  assign w17640 = w17631 & w17639 ;
  assign w17641 = ~w6549 & w16694 ;
  assign w17642 = w6048 & ~w16696 ;
  assign w17643 = ( w16694 & ~w17641 ) | ( w16694 & w17642 ) | ( ~w17641 & w17642 ) ;
  assign w17644 = w6637 | w16692 ;
  assign w17645 = w16784 | w17643 ;
  assign w17646 = ( w6045 & w17643 ) | ( w6045 & w17645 ) | ( w17643 & w17645 ) ;
  assign w17647 = ( ~w16692 & w17644 ) | ( ~w16692 & w17646 ) | ( w17644 & w17646 ) ;
  assign w17648 = \pi14 ^ w17647 ;
  assign w17649 = w5496 & ~w16698 ;
  assign w17650 = ( w17640 & w17648 ) | ( w17640 & w17649 ) | ( w17648 & w17649 ) ;
  assign w17651 = ( w17617 & w17625 ) | ( w17617 & w17650 ) | ( w17625 & w17650 ) ;
  assign w17652 = ( w17611 & w17612 ) | ( w17611 & w17651 ) | ( w17612 & w17651 ) ;
  assign w17653 = ( w17595 & w17603 ) | ( w17595 & w17652 ) | ( w17603 & w17652 ) ;
  assign w17654 = ( w17591 & w17593 ) | ( w17591 & w17653 ) | ( w17593 & w17653 ) ;
  assign w17655 = ( w17575 & w17583 ) | ( w17575 & w17654 ) | ( w17583 & w17654 ) ;
  assign w17656 = ( w17565 & w17573 ) | ( w17565 & w17655 ) | ( w17573 & w17655 ) ;
  assign w17657 = ( w17555 & w17563 ) | ( w17555 & w17656 ) | ( w17563 & w17656 ) ;
  assign w17658 = ( w17551 & w17553 ) | ( w17551 & w17657 ) | ( w17553 & w17657 ) ;
  assign w17659 = ( w17541 & w17543 ) | ( w17541 & w17658 ) | ( w17543 & w17658 ) ;
  assign w17660 = ( w17531 & w17533 ) | ( w17531 & w17659 ) | ( w17533 & w17659 ) ;
  assign w17661 = ( w17515 & w17523 ) | ( w17515 & w17660 ) | ( w17523 & w17660 ) ;
  assign w17662 = ( w17505 & w17513 ) | ( w17505 & w17661 ) | ( w17513 & w17661 ) ;
  assign w17663 = ( w17495 & w17503 ) | ( w17495 & w17662 ) | ( w17503 & w17662 ) ;
  assign w17664 = ( w17491 & w17493 ) | ( w17491 & w17663 ) | ( w17493 & w17663 ) ;
  assign w17665 = ( w17481 & w17483 ) | ( w17481 & w17664 ) | ( w17483 & w17664 ) ;
  assign w17666 = ( ~w17460 & w17471 ) | ( ~w17460 & w17665 ) | ( w17471 & w17665 ) ;
  assign w17667 = ( ~w17448 & w17458 ) | ( ~w17448 & w17666 ) | ( w17458 & w17666 ) ;
  assign w17668 = w5710 | w16648 ;
  assign w17669 = w5494 & ~w16650 ;
  assign w17670 = ( ~w16648 & w17668 ) | ( ~w16648 & w17669 ) | ( w17668 & w17669 ) ;
  assign w17671 = w5948 | w16646 ;
  assign w17672 = w17476 & ~w17670 ;
  assign w17673 = ( w5497 & w17670 ) | ( w5497 & ~w17672 ) | ( w17670 & ~w17672 ) ;
  assign w17674 = ( ~w16646 & w17671 ) | ( ~w16646 & w17673 ) | ( w17671 & w17673 ) ;
  assign w17675 = \pi17 ^ w17674 ;
  assign w17676 = ( w17192 & ~w17259 ) | ( w17192 & w17269 ) | ( ~w17259 & w17269 ) ;
  assign w17677 = ~w4651 & w16660 ;
  assign w17678 = w4606 & ~w16662 ;
  assign w17679 = ( w16660 & ~w17677 ) | ( w16660 & w17678 ) | ( ~w17677 & w17678 ) ;
  assign w17680 = w4706 | w16658 ;
  assign w17681 = w17065 & ~w17679 ;
  assign w17682 = ( w4609 & w17679 ) | ( w4609 & ~w17681 ) | ( w17679 & ~w17681 ) ;
  assign w17683 = ( ~w16658 & w17680 ) | ( ~w16658 & w17682 ) | ( w17680 & w17682 ) ;
  assign w17684 = \pi23 ^ w17683 ;
  assign w17685 = ( w17201 & ~w17246 ) | ( w17201 & w17254 ) | ( ~w17246 & w17254 ) ;
  assign w17686 = ~w3717 & w16685 ;
  assign w17687 = w3649 & ~w16690 ;
  assign w17688 = ( w16685 & ~w17686 ) | ( w16685 & w17687 ) | ( ~w17686 & w17687 ) ;
  assign w17689 = ~w3549 & w16680 ;
  assign w17690 = w16772 & ~w17688 ;
  assign w17691 = ( w3448 & w17688 ) | ( w3448 & ~w17690 ) | ( w17688 & ~w17690 ) ;
  assign w17692 = ( w16680 & ~w17689 ) | ( w16680 & w17691 ) | ( ~w17689 & w17691 ) ;
  assign w17693 = \pi29 ^ w17692 ;
  assign w17694 = ( w16935 & w17219 ) | ( w16935 & ~w17241 ) | ( w17219 & ~w17241 ) ;
  assign w17695 = ( w384 & w511 ) | ( w384 & ~w513 ) | ( w511 & ~w513 ) ;
  assign w17696 = w82 | w2037 ;
  assign w17697 = ( ~w82 & w513 ) | ( ~w82 & w1086 ) | ( w513 & w1086 ) ;
  assign w17698 = w17696 | w17697 ;
  assign w17699 = w17695 | w17698 ;
  assign w17700 = w424 | w1663 ;
  assign w17701 = ( w386 & ~w1663 ) | ( w386 & w17699 ) | ( ~w1663 & w17699 ) ;
  assign w17702 = w17700 | w17701 ;
  assign w17703 = ( ~w273 & w3379 ) | ( ~w273 & w5266 ) | ( w3379 & w5266 ) ;
  assign w17704 = w933 | w17702 ;
  assign w17705 = ( w273 & ~w933 ) | ( w273 & w2452 ) | ( ~w933 & w2452 ) ;
  assign w17706 = w17704 | w17705 ;
  assign w17707 = w17703 | w17706 ;
  assign w17708 = w84 | w1566 ;
  assign w17709 = w468 | w17708 ;
  assign w17710 = ( ~w468 & w517 ) | ( ~w468 & w17707 ) | ( w517 & w17707 ) ;
  assign w17711 = w17709 | w17710 ;
  assign w17712 = w68 | w802 ;
  assign w17713 = ( ~w68 & w202 ) | ( ~w68 & w17711 ) | ( w202 & w17711 ) ;
  assign w17714 = w17712 | w17713 ;
  assign w17715 = ~w37 & w16784 ;
  assign w17716 = w3098 & ~w16696 ;
  assign w17717 = ( w16784 & ~w17715 ) | ( w16784 & w17716 ) | ( ~w17715 & w17716 ) ;
  assign w17718 = ( \pi29 & \pi30 ) | ( \pi29 & ~w16692 ) | ( \pi30 & ~w16692 ) ;
  assign w17719 = \pi31 | w17718 ;
  assign w17720 = ( \pi29 & ~\pi30 ) | ( \pi29 & w16694 ) | ( ~\pi30 & w16694 ) ;
  assign w17721 = ( \pi29 & \pi31 ) | ( \pi29 & ~w17720 ) | ( \pi31 & ~w17720 ) ;
  assign w17722 = ( w17717 & w17719 ) | ( w17717 & ~w17721 ) | ( w17719 & ~w17721 ) ;
  assign w17723 = w17694 ^ w17722 ;
  assign w17724 = w17714 ^ w17723 ;
  assign w17725 = ( w17209 & ~w17243 ) | ( w17209 & w17244 ) | ( ~w17243 & w17244 ) ;
  assign w17726 = w17693 ^ w17725 ;
  assign w17727 = w17724 ^ w17726 ;
  assign w17728 = w3964 & w16665 ;
  assign w17729 = ( w4143 & w16670 ) | ( w4143 & w17728 ) | ( w16670 & w17728 ) ;
  assign w17730 = w4052 | w17729 ;
  assign w17731 = ( w16675 & w17729 ) | ( w16675 & w17730 ) | ( w17729 & w17730 ) ;
  assign w17732 = w17728 | w17731 ;
  assign w17733 = ~w4147 & w16960 ;
  assign w17734 = ( w16960 & w17732 ) | ( w16960 & ~w17733 ) | ( w17732 & ~w17733 ) ;
  assign w17735 = \pi26 ^ w17734 ;
  assign w17736 = w17685 ^ w17735 ;
  assign w17737 = w17727 ^ w17736 ;
  assign w17738 = ( w17200 & ~w17256 ) | ( w17200 & w17257 ) | ( ~w17256 & w17257 ) ;
  assign w17739 = w17684 ^ w17738 ;
  assign w17740 = w17737 ^ w17739 ;
  assign w17741 = w4905 & ~w16656 ;
  assign w17742 = ( w5395 & ~w16652 ) | ( w5395 & w17741 ) | ( ~w16652 & w17741 ) ;
  assign w17743 = w5343 | w17742 ;
  assign w17744 = ( w16654 & w17742 ) | ( w16654 & w17743 ) | ( w17742 & w17743 ) ;
  assign w17745 = w17741 | w17744 ;
  assign w17746 = ~w4908 & w17293 ;
  assign w17747 = ( w17293 & w17745 ) | ( w17293 & ~w17746 ) | ( w17745 & ~w17746 ) ;
  assign w17748 = \pi20 ^ w17747 ;
  assign w17749 = w17676 ^ w17748 ;
  assign w17750 = w17740 ^ w17749 ;
  assign w17751 = ( w16757 & ~w17271 ) | ( w16757 & w17446 ) | ( ~w17271 & w17446 ) ;
  assign w17752 = w17675 ^ w17751 ;
  assign w17753 = w17750 ^ w17752 ;
  assign w17754 = w6048 & ~w16644 ;
  assign w17755 = ( w6637 & w16640 ) | ( w6637 & w17754 ) | ( w16640 & w17754 ) ;
  assign w17756 = w6549 | w17755 ;
  assign w17757 = ( w16642 & w17755 ) | ( w16642 & w17756 ) | ( w17755 & w17756 ) ;
  assign w17758 = w17754 | w17757 ;
  assign w17759 = w16640 ^ w16718 ;
  assign w17760 = w16642 ^ w17759 ;
  assign w17761 = w6045 & w17760 ;
  assign w17762 = ( w6045 & w17758 ) | ( w6045 & ~w17761 ) | ( w17758 & ~w17761 ) ;
  assign w17763 = \pi14 ^ w17762 ;
  assign w17764 = w17667 ^ w17763 ;
  assign w17765 = w17753 ^ w17764 ;
  assign w17766 = w6949 | w16638 ;
  assign w17767 = w6748 & w16640 ;
  assign w17768 = ( ~w16638 & w17766 ) | ( ~w16638 & w17767 ) | ( w17766 & w17767 ) ;
  assign w17769 = w16636 ^ w16720 ;
  assign w17770 = w16638 ^ w17769 ;
  assign w17771 = ~w7154 & w16636 ;
  assign w17772 = ~w17768 & w17770 ;
  assign w17773 = ( w6751 & w17768 ) | ( w6751 & ~w17772 ) | ( w17768 & ~w17772 ) ;
  assign w17774 = ( w16636 & ~w17771 ) | ( w16636 & w17773 ) | ( ~w17771 & w17773 ) ;
  assign w17775 = \pi11 ^ w17774 ;
  assign w17776 = w17458 ^ w17666 ;
  assign w17777 = w17448 ^ w17776 ;
  assign w17778 = ~w6949 & w16640 ;
  assign w17779 = w6748 & w16642 ;
  assign w17780 = ( w16640 & ~w17778 ) | ( w16640 & w17779 ) | ( ~w17778 & w17779 ) ;
  assign w17781 = ( w16640 & w16642 ) | ( w16640 & ~w16718 ) | ( w16642 & ~w16718 ) ;
  assign w17782 = w16640 ^ w17781 ;
  assign w17783 = w16638 ^ w17782 ;
  assign w17784 = w7154 | w16638 ;
  assign w17785 = ~w17780 & w17783 ;
  assign w17786 = ( w6751 & w17780 ) | ( w6751 & ~w17785 ) | ( w17780 & ~w17785 ) ;
  assign w17787 = ( ~w16638 & w17784 ) | ( ~w16638 & w17786 ) | ( w17784 & w17786 ) ;
  assign w17788 = \pi11 ^ w17787 ;
  assign w17789 = w17471 ^ w17665 ;
  assign w17790 = w17460 ^ w17789 ;
  assign w17791 = w17481 ^ w17664 ;
  assign w17792 = w17483 ^ w17791 ;
  assign w17793 = w6748 & ~w16644 ;
  assign w17794 = ( w7154 & w16640 ) | ( w7154 & w17793 ) | ( w16640 & w17793 ) ;
  assign w17795 = w6949 | w17794 ;
  assign w17796 = ( w16642 & w17794 ) | ( w16642 & w17795 ) | ( w17794 & w17795 ) ;
  assign w17797 = w17793 | w17796 ;
  assign w17798 = w6751 | w17760 ;
  assign w17799 = ( ~w17760 & w17797 ) | ( ~w17760 & w17798 ) | ( w17797 & w17798 ) ;
  assign w17800 = \pi11 ^ w17799 ;
  assign w17801 = w17491 ^ w17663 ;
  assign w17802 = w17493 ^ w17801 ;
  assign w17803 = w6748 & ~w16646 ;
  assign w17804 = ( w7154 & w16642 ) | ( w7154 & w17803 ) | ( w16642 & w17803 ) ;
  assign w17805 = w6949 | w17804 ;
  assign w17806 = ( ~w16644 & w17804 ) | ( ~w16644 & w17805 ) | ( w17804 & w17805 ) ;
  assign w17807 = w17803 | w17806 ;
  assign w17808 = ~w6751 & w17455 ;
  assign w17809 = ( w17455 & w17807 ) | ( w17455 & ~w17808 ) | ( w17807 & ~w17808 ) ;
  assign w17810 = \pi11 ^ w17809 ;
  assign w17811 = w6949 | w16646 ;
  assign w17812 = w6748 & ~w16648 ;
  assign w17813 = ( ~w16646 & w17811 ) | ( ~w16646 & w17812 ) | ( w17811 & w17812 ) ;
  assign w17814 = w7154 | w16644 ;
  assign w17815 = w17468 & ~w17813 ;
  assign w17816 = ( w6751 & w17813 ) | ( w6751 & ~w17815 ) | ( w17813 & ~w17815 ) ;
  assign w17817 = ( ~w16644 & w17814 ) | ( ~w16644 & w17816 ) | ( w17814 & w17816 ) ;
  assign w17818 = \pi11 ^ w17817 ;
  assign w17819 = w17503 ^ w17662 ;
  assign w17820 = w17495 ^ w17819 ;
  assign w17821 = w6949 | w16648 ;
  assign w17822 = w6748 & ~w16650 ;
  assign w17823 = ( ~w16648 & w17821 ) | ( ~w16648 & w17822 ) | ( w17821 & w17822 ) ;
  assign w17824 = w7154 | w16646 ;
  assign w17825 = w17476 & ~w17823 ;
  assign w17826 = ( w6751 & w17823 ) | ( w6751 & ~w17825 ) | ( w17823 & ~w17825 ) ;
  assign w17827 = ( ~w16646 & w17824 ) | ( ~w16646 & w17826 ) | ( w17824 & w17826 ) ;
  assign w17828 = \pi11 ^ w17827 ;
  assign w17829 = w17513 ^ w17661 ;
  assign w17830 = w17505 ^ w17829 ;
  assign w17831 = w6949 | w16650 ;
  assign w17832 = w6748 & ~w16652 ;
  assign w17833 = ( ~w16650 & w17831 ) | ( ~w16650 & w17832 ) | ( w17831 & w17832 ) ;
  assign w17834 = w7154 | w16648 ;
  assign w17835 = w16752 & ~w17833 ;
  assign w17836 = ( w6751 & w17833 ) | ( w6751 & ~w17835 ) | ( w17833 & ~w17835 ) ;
  assign w17837 = ( ~w16648 & w17834 ) | ( ~w16648 & w17836 ) | ( w17834 & w17836 ) ;
  assign w17838 = \pi11 ^ w17837 ;
  assign w17839 = w17523 ^ w17660 ;
  assign w17840 = w17515 ^ w17839 ;
  assign w17841 = w17531 ^ w17659 ;
  assign w17842 = w17533 ^ w17841 ;
  assign w17843 = w6748 & w16654 ;
  assign w17844 = ( w7154 & ~w16650 ) | ( w7154 & w17843 ) | ( ~w16650 & w17843 ) ;
  assign w17845 = w6949 | w17844 ;
  assign w17846 = ( ~w16652 & w17844 ) | ( ~w16652 & w17845 ) | ( w17844 & w17845 ) ;
  assign w17847 = w17843 | w17846 ;
  assign w17848 = w6751 | w17277 ;
  assign w17849 = ( ~w17277 & w17847 ) | ( ~w17277 & w17848 ) | ( w17847 & w17848 ) ;
  assign w17850 = \pi11 ^ w17849 ;
  assign w17851 = w17541 ^ w17658 ;
  assign w17852 = w17543 ^ w17851 ;
  assign w17853 = w6748 & ~w16656 ;
  assign w17854 = ( w7154 & ~w16652 ) | ( w7154 & w17853 ) | ( ~w16652 & w17853 ) ;
  assign w17855 = w6949 | w17854 ;
  assign w17856 = ( w16654 & w17854 ) | ( w16654 & w17855 ) | ( w17854 & w17855 ) ;
  assign w17857 = w17853 | w17856 ;
  assign w17858 = ~w6751 & w17293 ;
  assign w17859 = ( w17293 & w17857 ) | ( w17293 & ~w17858 ) | ( w17857 & ~w17858 ) ;
  assign w17860 = \pi11 ^ w17859 ;
  assign w17861 = w17551 ^ w17657 ;
  assign w17862 = w17553 ^ w17861 ;
  assign w17863 = w6748 & ~w16658 ;
  assign w17864 = ( w7154 & w16654 ) | ( w7154 & w17863 ) | ( w16654 & w17863 ) ;
  assign w17865 = w6949 | w17864 ;
  assign w17866 = ( ~w16656 & w17864 ) | ( ~w16656 & w17865 ) | ( w17864 & w17865 ) ;
  assign w17867 = w17863 | w17866 ;
  assign w17868 = ~w6751 & w17266 ;
  assign w17869 = ( w17266 & w17867 ) | ( w17266 & ~w17868 ) | ( w17867 & ~w17868 ) ;
  assign w17870 = \pi11 ^ w17869 ;
  assign w17871 = w6949 | w16658 ;
  assign w17872 = w6748 & w16660 ;
  assign w17873 = ( ~w16658 & w17871 ) | ( ~w16658 & w17872 ) | ( w17871 & w17872 ) ;
  assign w17874 = w7154 | w16656 ;
  assign w17875 = w17057 | w17873 ;
  assign w17876 = ( w6751 & w17873 ) | ( w6751 & w17875 ) | ( w17873 & w17875 ) ;
  assign w17877 = ( ~w16656 & w17874 ) | ( ~w16656 & w17876 ) | ( w17874 & w17876 ) ;
  assign w17878 = \pi11 ^ w17877 ;
  assign w17879 = w17563 ^ w17656 ;
  assign w17880 = w17555 ^ w17879 ;
  assign w17881 = ~w6949 & w16660 ;
  assign w17882 = w6748 & ~w16662 ;
  assign w17883 = ( w16660 & ~w17881 ) | ( w16660 & w17882 ) | ( ~w17881 & w17882 ) ;
  assign w17884 = w7154 | w16658 ;
  assign w17885 = w17065 & ~w17883 ;
  assign w17886 = ( w6751 & w17883 ) | ( w6751 & ~w17885 ) | ( w17883 & ~w17885 ) ;
  assign w17887 = ( ~w16658 & w17884 ) | ( ~w16658 & w17886 ) | ( w17884 & w17886 ) ;
  assign w17888 = \pi11 ^ w17887 ;
  assign w17889 = w17573 ^ w17655 ;
  assign w17890 = w17565 ^ w17889 ;
  assign w17891 = w6949 | w16662 ;
  assign w17892 = w6748 & w16665 ;
  assign w17893 = ( ~w16662 & w17891 ) | ( ~w16662 & w17892 ) | ( w17891 & w17892 ) ;
  assign w17894 = ~w7154 & w16660 ;
  assign w17895 = w17078 & ~w17893 ;
  assign w17896 = ( w6751 & w17893 ) | ( w6751 & ~w17895 ) | ( w17893 & ~w17895 ) ;
  assign w17897 = ( w16660 & ~w17894 ) | ( w16660 & w17896 ) | ( ~w17894 & w17896 ) ;
  assign w17898 = \pi11 ^ w17897 ;
  assign w17899 = w17583 ^ w17654 ;
  assign w17900 = w17575 ^ w17899 ;
  assign w17901 = w17591 ^ w17653 ;
  assign w17902 = w17593 ^ w17901 ;
  assign w17903 = w6748 & w16670 ;
  assign w17904 = ( w7154 & ~w16662 ) | ( w7154 & w17903 ) | ( ~w16662 & w17903 ) ;
  assign w17905 = w6949 | w17904 ;
  assign w17906 = ( w16665 & w17904 ) | ( w16665 & w17905 ) | ( w17904 & w17905 ) ;
  assign w17907 = w17903 | w17906 ;
  assign w17908 = w6751 | w16762 ;
  assign w17909 = ( ~w16762 & w17907 ) | ( ~w16762 & w17908 ) | ( w17907 & w17908 ) ;
  assign w17910 = \pi11 ^ w17909 ;
  assign w17911 = w17603 ^ w17652 ;
  assign w17912 = w17595 ^ w17911 ;
  assign w17913 = w6748 & w16675 ;
  assign w17914 = ( w7154 & w16665 ) | ( w7154 & w17913 ) | ( w16665 & w17913 ) ;
  assign w17915 = w6949 | w17914 ;
  assign w17916 = ( w16670 & w17914 ) | ( w16670 & w17915 ) | ( w17914 & w17915 ) ;
  assign w17917 = w17913 | w17916 ;
  assign w17918 = ~w6751 & w16960 ;
  assign w17919 = ( w16960 & w17917 ) | ( w16960 & ~w17918 ) | ( w17917 & ~w17918 ) ;
  assign w17920 = \pi11 ^ w17919 ;
  assign w17921 = w17611 ^ w17651 ;
  assign w17922 = w17612 ^ w17921 ;
  assign w17923 = w6748 & w16680 ;
  assign w17924 = ( w7154 & w16670 ) | ( w7154 & w17923 ) | ( w16670 & w17923 ) ;
  assign w17925 = w6949 | w17924 ;
  assign w17926 = ( w16675 & w17924 ) | ( w16675 & w17925 ) | ( w17924 & w17925 ) ;
  assign w17927 = w17923 | w17926 ;
  assign w17928 = ~w6751 & w16972 ;
  assign w17929 = ( w16972 & w17927 ) | ( w16972 & ~w17928 ) | ( w17927 & ~w17928 ) ;
  assign w17930 = \pi11 ^ w17929 ;
  assign w17931 = ~w6949 & w16680 ;
  assign w17932 = w6748 & w16685 ;
  assign w17933 = ( w16680 & ~w17931 ) | ( w16680 & w17932 ) | ( ~w17931 & w17932 ) ;
  assign w17934 = ~w7154 & w16675 ;
  assign w17935 = w16946 | w17933 ;
  assign w17936 = ( w6751 & w17933 ) | ( w6751 & w17935 ) | ( w17933 & w17935 ) ;
  assign w17937 = ( w16675 & ~w17934 ) | ( w16675 & w17936 ) | ( ~w17934 & w17936 ) ;
  assign w17938 = \pi11 ^ w17937 ;
  assign w17939 = w17625 ^ w17650 ;
  assign w17940 = w17617 ^ w17939 ;
  assign w17941 = w17640 ^ w17648 ;
  assign w17942 = w17649 ^ w17941 ;
  assign w17943 = w6748 & ~w16690 ;
  assign w17944 = ( w7154 & w16680 ) | ( w7154 & w17943 ) | ( w16680 & w17943 ) ;
  assign w17945 = w6949 | w17944 ;
  assign w17946 = ( w16685 & w17944 ) | ( w16685 & w17945 ) | ( w17944 & w17945 ) ;
  assign w17947 = w17943 | w17946 ;
  assign w17948 = w6751 | w16772 ;
  assign w17949 = ( ~w16772 & w17947 ) | ( ~w16772 & w17948 ) | ( w17947 & w17948 ) ;
  assign w17950 = \pi11 ^ w17949 ;
  assign w17951 = w6949 | w16690 ;
  assign w17952 = w6748 & ~w16692 ;
  assign w17953 = ( ~w16690 & w17951 ) | ( ~w16690 & w17952 ) | ( w17951 & w17952 ) ;
  assign w17954 = ~w7154 & w16685 ;
  assign w17955 = w16818 | w17953 ;
  assign w17956 = ( w6751 & w17953 ) | ( w6751 & w17955 ) | ( w17953 & w17955 ) ;
  assign w17957 = ( w16685 & ~w17954 ) | ( w16685 & w17956 ) | ( ~w17954 & w17956 ) ;
  assign w17958 = \pi11 ^ w17957 ;
  assign w17959 = w17631 ^ w17639 ;
  assign w17960 = ( \pi11 & \pi12 ) | ( \pi11 & ~w16696 ) | ( \pi12 & ~w16696 ) ;
  assign w17961 = ( \pi11 & \pi12 ) | ( \pi11 & ~w16698 ) | ( \pi12 & ~w16698 ) ;
  assign w17962 = \pi13 ^ w16698 ;
  assign w17963 = ( \pi13 & w17961 ) | ( \pi13 & w17962 ) | ( w17961 & w17962 ) ;
  assign w17964 = w17960 ^ w17963 ;
  assign w17965 = w6748 & w16694 ;
  assign w17966 = ( w7154 & ~w16690 ) | ( w7154 & w17965 ) | ( ~w16690 & w17965 ) ;
  assign w17967 = w6949 | w17966 ;
  assign w17968 = ( ~w16692 & w17966 ) | ( ~w16692 & w17967 ) | ( w17966 & w17967 ) ;
  assign w17969 = w17965 | w17968 ;
  assign w17970 = w6751 | w16839 ;
  assign w17971 = ( ~w16839 & w17969 ) | ( ~w16839 & w17970 ) | ( w17969 & w17970 ) ;
  assign w17972 = \pi11 ^ w17971 ;
  assign w17973 = \pi11 & w16698 ;
  assign w17974 = w16696 & w17973 ;
  assign w17975 = ( \pi08 & \pi09 ) | ( \pi08 & ~w17974 ) | ( \pi09 & ~w17974 ) ;
  assign w17976 = ( \pi10 & \pi11 ) | ( \pi10 & ~w17975 ) | ( \pi11 & ~w17975 ) ;
  assign w17977 = ( \pi10 & ~w17973 ) | ( \pi10 & w17975 ) | ( ~w17973 & w17975 ) ;
  assign w17978 = ( w8530 & w17976 ) | ( w8530 & ~w17977 ) | ( w17976 & ~w17977 ) ;
  assign w17979 = w6748 & ~w16698 ;
  assign w17980 = ( w7154 & w16694 ) | ( w7154 & w17979 ) | ( w16694 & w17979 ) ;
  assign w17981 = w6949 | w17980 ;
  assign w17982 = ( ~w16696 & w17980 ) | ( ~w16696 & w17981 ) | ( w17980 & w17981 ) ;
  assign w17983 = w17979 | w17982 ;
  assign w17984 = ~w6751 & w16802 ;
  assign w17985 = ( w16802 & w17983 ) | ( w16802 & ~w17984 ) | ( w17983 & ~w17984 ) ;
  assign w17986 = \pi11 ^ w17985 ;
  assign w17987 = w17978 & w17986 ;
  assign w17988 = ~w6949 & w16694 ;
  assign w17989 = w6748 & ~w16696 ;
  assign w17990 = ( w16694 & ~w17988 ) | ( w16694 & w17989 ) | ( ~w17988 & w17989 ) ;
  assign w17991 = w7154 | w16692 ;
  assign w17992 = w16784 | w17990 ;
  assign w17993 = ( w6751 & w17990 ) | ( w6751 & w17992 ) | ( w17990 & w17992 ) ;
  assign w17994 = ( ~w16692 & w17991 ) | ( ~w16692 & w17993 ) | ( w17991 & w17993 ) ;
  assign w17995 = \pi11 ^ w17994 ;
  assign w17996 = w6044 & ~w16698 ;
  assign w17997 = ( w17987 & w17995 ) | ( w17987 & w17996 ) | ( w17995 & w17996 ) ;
  assign w17998 = ( w17964 & w17972 ) | ( w17964 & w17997 ) | ( w17972 & w17997 ) ;
  assign w17999 = ( w17958 & w17959 ) | ( w17958 & w17998 ) | ( w17959 & w17998 ) ;
  assign w18000 = ( w17942 & w17950 ) | ( w17942 & w17999 ) | ( w17950 & w17999 ) ;
  assign w18001 = ( w17938 & w17940 ) | ( w17938 & w18000 ) | ( w17940 & w18000 ) ;
  assign w18002 = ( w17922 & w17930 ) | ( w17922 & w18001 ) | ( w17930 & w18001 ) ;
  assign w18003 = ( w17912 & w17920 ) | ( w17912 & w18002 ) | ( w17920 & w18002 ) ;
  assign w18004 = ( w17902 & w17910 ) | ( w17902 & w18003 ) | ( w17910 & w18003 ) ;
  assign w18005 = ( w17898 & w17900 ) | ( w17898 & w18004 ) | ( w17900 & w18004 ) ;
  assign w18006 = ( w17888 & w17890 ) | ( w17888 & w18005 ) | ( w17890 & w18005 ) ;
  assign w18007 = ( w17878 & w17880 ) | ( w17878 & w18006 ) | ( w17880 & w18006 ) ;
  assign w18008 = ( w17862 & w17870 ) | ( w17862 & w18007 ) | ( w17870 & w18007 ) ;
  assign w18009 = ( w17852 & w17860 ) | ( w17852 & w18008 ) | ( w17860 & w18008 ) ;
  assign w18010 = ( w17842 & w17850 ) | ( w17842 & w18009 ) | ( w17850 & w18009 ) ;
  assign w18011 = ( w17838 & w17840 ) | ( w17838 & w18010 ) | ( w17840 & w18010 ) ;
  assign w18012 = ( w17828 & w17830 ) | ( w17828 & w18011 ) | ( w17830 & w18011 ) ;
  assign w18013 = ( w17818 & w17820 ) | ( w17818 & w18012 ) | ( w17820 & w18012 ) ;
  assign w18014 = ( w17802 & w17810 ) | ( w17802 & w18013 ) | ( w17810 & w18013 ) ;
  assign w18015 = ( w17792 & w17800 ) | ( w17792 & w18014 ) | ( w17800 & w18014 ) ;
  assign w18016 = ( w17788 & ~w17790 ) | ( w17788 & w18015 ) | ( ~w17790 & w18015 ) ;
  assign w18017 = ( w17775 & ~w17777 ) | ( w17775 & w18016 ) | ( ~w17777 & w18016 ) ;
  assign w18018 = w16747 ^ w18017 ;
  assign w18019 = w17765 ^ w18018 ;
  assign w18020 = w7411 & w16632 ;
  assign w18021 = ( w7944 & ~w16628 ) | ( w7944 & w18020 ) | ( ~w16628 & w18020 ) ;
  assign w18022 = w7673 | w18021 ;
  assign w18023 = ( ~w16630 & w18021 ) | ( ~w16630 & w18022 ) | ( w18021 & w18022 ) ;
  assign w18024 = w18020 | w18023 ;
  assign w18025 = w16628 ^ w16724 ;
  assign w18026 = w16630 ^ w18025 ;
  assign w18027 = w7414 & ~w18026 ;
  assign w18028 = ( w7414 & w18024 ) | ( w7414 & ~w18027 ) | ( w18024 & ~w18027 ) ;
  assign w18029 = \pi08 ^ w18028 ;
  assign w18030 = w17775 ^ w18016 ;
  assign w18031 = w17777 ^ w18030 ;
  assign w18032 = w7411 & ~w16634 ;
  assign w18033 = ( w7944 & ~w16630 ) | ( w7944 & w18032 ) | ( ~w16630 & w18032 ) ;
  assign w18034 = w7673 | w18033 ;
  assign w18035 = ( w16632 & w18033 ) | ( w16632 & w18034 ) | ( w18033 & w18034 ) ;
  assign w18036 = w18032 | w18035 ;
  assign w18037 = w16630 ^ w16723 ;
  assign w18038 = w16632 ^ w18037 ;
  assign w18039 = w7414 & w18038 ;
  assign w18040 = ( w7414 & w18036 ) | ( w7414 & ~w18039 ) | ( w18036 & ~w18039 ) ;
  assign w18041 = \pi08 ^ w18040 ;
  assign w18042 = w17788 ^ w18015 ;
  assign w18043 = w17790 ^ w18042 ;
  assign w18044 = w7411 & w16636 ;
  assign w18045 = ( w7944 & w16632 ) | ( w7944 & w18044 ) | ( w16632 & w18044 ) ;
  assign w18046 = w7673 | w18045 ;
  assign w18047 = ( ~w16634 & w18045 ) | ( ~w16634 & w18046 ) | ( w18045 & w18046 ) ;
  assign w18048 = w18044 | w18047 ;
  assign w18049 = ( ~w16634 & w16636 ) | ( ~w16634 & w16721 ) | ( w16636 & w16721 ) ;
  assign w18050 = w16634 ^ w18049 ;
  assign w18051 = w16632 ^ w18050 ;
  assign w18052 = w7414 & w18051 ;
  assign w18053 = ( w7414 & w18048 ) | ( w7414 & ~w18052 ) | ( w18048 & ~w18052 ) ;
  assign w18054 = \pi08 ^ w18053 ;
  assign w18055 = ~w7673 & w16636 ;
  assign w18056 = w7411 & ~w16638 ;
  assign w18057 = ( w16636 & ~w18055 ) | ( w16636 & w18056 ) | ( ~w18055 & w18056 ) ;
  assign w18058 = w7944 | w16634 ;
  assign w18059 = w16742 & ~w18057 ;
  assign w18060 = ( w7414 & w18057 ) | ( w7414 & ~w18059 ) | ( w18057 & ~w18059 ) ;
  assign w18061 = ( ~w16634 & w18058 ) | ( ~w16634 & w18060 ) | ( w18058 & w18060 ) ;
  assign w18062 = \pi08 ^ w18061 ;
  assign w18063 = w17800 ^ w18014 ;
  assign w18064 = w17792 ^ w18063 ;
  assign w18065 = w7673 | w16638 ;
  assign w18066 = w7411 & w16640 ;
  assign w18067 = ( ~w16638 & w18065 ) | ( ~w16638 & w18066 ) | ( w18065 & w18066 ) ;
  assign w18068 = ~w7944 & w16636 ;
  assign w18069 = w17770 & ~w18067 ;
  assign w18070 = ( w7414 & w18067 ) | ( w7414 & ~w18069 ) | ( w18067 & ~w18069 ) ;
  assign w18071 = ( w16636 & ~w18068 ) | ( w16636 & w18070 ) | ( ~w18068 & w18070 ) ;
  assign w18072 = \pi08 ^ w18071 ;
  assign w18073 = w17810 ^ w18013 ;
  assign w18074 = w17802 ^ w18073 ;
  assign w18075 = w17818 ^ w18012 ;
  assign w18076 = w17820 ^ w18075 ;
  assign w18077 = w7411 & w16642 ;
  assign w18078 = ( w7944 & ~w16638 ) | ( w7944 & w18077 ) | ( ~w16638 & w18077 ) ;
  assign w18079 = w7673 | w18078 ;
  assign w18080 = ( w16640 & w18078 ) | ( w16640 & w18079 ) | ( w18078 & w18079 ) ;
  assign w18081 = w18077 | w18080 ;
  assign w18082 = w7414 | w17783 ;
  assign w18083 = ( ~w17783 & w18081 ) | ( ~w17783 & w18082 ) | ( w18081 & w18082 ) ;
  assign w18084 = \pi08 ^ w18083 ;
  assign w18085 = w17828 ^ w18011 ;
  assign w18086 = w17830 ^ w18085 ;
  assign w18087 = w7411 & ~w16644 ;
  assign w18088 = ( w7944 & w16640 ) | ( w7944 & w18087 ) | ( w16640 & w18087 ) ;
  assign w18089 = w7673 | w18088 ;
  assign w18090 = ( w16642 & w18088 ) | ( w16642 & w18089 ) | ( w18088 & w18089 ) ;
  assign w18091 = w18087 | w18090 ;
  assign w18092 = w7414 | w17760 ;
  assign w18093 = ( ~w17760 & w18091 ) | ( ~w17760 & w18092 ) | ( w18091 & w18092 ) ;
  assign w18094 = \pi08 ^ w18093 ;
  assign w18095 = w17838 ^ w18010 ;
  assign w18096 = w17840 ^ w18095 ;
  assign w18097 = w7411 & ~w16646 ;
  assign w18098 = ( w7944 & w16642 ) | ( w7944 & w18097 ) | ( w16642 & w18097 ) ;
  assign w18099 = w7673 | w18098 ;
  assign w18100 = ( ~w16644 & w18098 ) | ( ~w16644 & w18099 ) | ( w18098 & w18099 ) ;
  assign w18101 = w18097 | w18100 ;
  assign w18102 = ~w7414 & w17455 ;
  assign w18103 = ( w17455 & w18101 ) | ( w17455 & ~w18102 ) | ( w18101 & ~w18102 ) ;
  assign w18104 = \pi08 ^ w18103 ;
  assign w18105 = w7673 | w16646 ;
  assign w18106 = w7411 & ~w16648 ;
  assign w18107 = ( ~w16646 & w18105 ) | ( ~w16646 & w18106 ) | ( w18105 & w18106 ) ;
  assign w18108 = w7944 | w16644 ;
  assign w18109 = w17468 & ~w18107 ;
  assign w18110 = ( w7414 & w18107 ) | ( w7414 & ~w18109 ) | ( w18107 & ~w18109 ) ;
  assign w18111 = ( ~w16644 & w18108 ) | ( ~w16644 & w18110 ) | ( w18108 & w18110 ) ;
  assign w18112 = \pi08 ^ w18111 ;
  assign w18113 = w17850 ^ w18009 ;
  assign w18114 = w17842 ^ w18113 ;
  assign w18115 = w7673 | w16648 ;
  assign w18116 = w7411 & ~w16650 ;
  assign w18117 = ( ~w16648 & w18115 ) | ( ~w16648 & w18116 ) | ( w18115 & w18116 ) ;
  assign w18118 = w7944 | w16646 ;
  assign w18119 = w17476 & ~w18117 ;
  assign w18120 = ( w7414 & w18117 ) | ( w7414 & ~w18119 ) | ( w18117 & ~w18119 ) ;
  assign w18121 = ( ~w16646 & w18118 ) | ( ~w16646 & w18120 ) | ( w18118 & w18120 ) ;
  assign w18122 = \pi08 ^ w18121 ;
  assign w18123 = w17860 ^ w18008 ;
  assign w18124 = w17852 ^ w18123 ;
  assign w18125 = w7673 | w16650 ;
  assign w18126 = w7411 & ~w16652 ;
  assign w18127 = ( ~w16650 & w18125 ) | ( ~w16650 & w18126 ) | ( w18125 & w18126 ) ;
  assign w18128 = w7944 | w16648 ;
  assign w18129 = w16752 & ~w18127 ;
  assign w18130 = ( w7414 & w18127 ) | ( w7414 & ~w18129 ) | ( w18127 & ~w18129 ) ;
  assign w18131 = ( ~w16648 & w18128 ) | ( ~w16648 & w18130 ) | ( w18128 & w18130 ) ;
  assign w18132 = \pi08 ^ w18131 ;
  assign w18133 = w17870 ^ w18007 ;
  assign w18134 = w17862 ^ w18133 ;
  assign w18135 = w17878 ^ w18006 ;
  assign w18136 = w17880 ^ w18135 ;
  assign w18137 = w7411 & w16654 ;
  assign w18138 = ( w7944 & ~w16650 ) | ( w7944 & w18137 ) | ( ~w16650 & w18137 ) ;
  assign w18139 = w7673 | w18138 ;
  assign w18140 = ( ~w16652 & w18138 ) | ( ~w16652 & w18139 ) | ( w18138 & w18139 ) ;
  assign w18141 = w18137 | w18140 ;
  assign w18142 = w7414 | w17277 ;
  assign w18143 = ( ~w17277 & w18141 ) | ( ~w17277 & w18142 ) | ( w18141 & w18142 ) ;
  assign w18144 = \pi08 ^ w18143 ;
  assign w18145 = w17888 ^ w18005 ;
  assign w18146 = w17890 ^ w18145 ;
  assign w18147 = w7411 & ~w16656 ;
  assign w18148 = ( w7944 & ~w16652 ) | ( w7944 & w18147 ) | ( ~w16652 & w18147 ) ;
  assign w18149 = w7673 | w18148 ;
  assign w18150 = ( w16654 & w18148 ) | ( w16654 & w18149 ) | ( w18148 & w18149 ) ;
  assign w18151 = w18147 | w18150 ;
  assign w18152 = ~w7414 & w17293 ;
  assign w18153 = ( w17293 & w18151 ) | ( w17293 & ~w18152 ) | ( w18151 & ~w18152 ) ;
  assign w18154 = \pi08 ^ w18153 ;
  assign w18155 = w17898 ^ w18004 ;
  assign w18156 = w17900 ^ w18155 ;
  assign w18157 = w7411 & ~w16658 ;
  assign w18158 = ( w7944 & w16654 ) | ( w7944 & w18157 ) | ( w16654 & w18157 ) ;
  assign w18159 = w7673 | w18158 ;
  assign w18160 = ( ~w16656 & w18158 ) | ( ~w16656 & w18159 ) | ( w18158 & w18159 ) ;
  assign w18161 = w18157 | w18160 ;
  assign w18162 = ~w7414 & w17266 ;
  assign w18163 = ( w17266 & w18161 ) | ( w17266 & ~w18162 ) | ( w18161 & ~w18162 ) ;
  assign w18164 = \pi08 ^ w18163 ;
  assign w18165 = w7673 | w16658 ;
  assign w18166 = w7411 & w16660 ;
  assign w18167 = ( ~w16658 & w18165 ) | ( ~w16658 & w18166 ) | ( w18165 & w18166 ) ;
  assign w18168 = w7944 | w16656 ;
  assign w18169 = w17057 | w18167 ;
  assign w18170 = ( w7414 & w18167 ) | ( w7414 & w18169 ) | ( w18167 & w18169 ) ;
  assign w18171 = ( ~w16656 & w18168 ) | ( ~w16656 & w18170 ) | ( w18168 & w18170 ) ;
  assign w18172 = \pi08 ^ w18171 ;
  assign w18173 = w17910 ^ w18003 ;
  assign w18174 = w17902 ^ w18173 ;
  assign w18175 = ~w7673 & w16660 ;
  assign w18176 = w7411 & ~w16662 ;
  assign w18177 = ( w16660 & ~w18175 ) | ( w16660 & w18176 ) | ( ~w18175 & w18176 ) ;
  assign w18178 = w7944 | w16658 ;
  assign w18179 = w17065 & ~w18177 ;
  assign w18180 = ( w7414 & w18177 ) | ( w7414 & ~w18179 ) | ( w18177 & ~w18179 ) ;
  assign w18181 = ( ~w16658 & w18178 ) | ( ~w16658 & w18180 ) | ( w18178 & w18180 ) ;
  assign w18182 = \pi08 ^ w18181 ;
  assign w18183 = w17920 ^ w18002 ;
  assign w18184 = w17912 ^ w18183 ;
  assign w18185 = w7673 | w16662 ;
  assign w18186 = w7411 & w16665 ;
  assign w18187 = ( ~w16662 & w18185 ) | ( ~w16662 & w18186 ) | ( w18185 & w18186 ) ;
  assign w18188 = ~w7944 & w16660 ;
  assign w18189 = w17078 & ~w18187 ;
  assign w18190 = ( w7414 & w18187 ) | ( w7414 & ~w18189 ) | ( w18187 & ~w18189 ) ;
  assign w18191 = ( w16660 & ~w18188 ) | ( w16660 & w18190 ) | ( ~w18188 & w18190 ) ;
  assign w18192 = \pi08 ^ w18191 ;
  assign w18193 = w17930 ^ w18001 ;
  assign w18194 = w17922 ^ w18193 ;
  assign w18195 = w17938 ^ w18000 ;
  assign w18196 = w17940 ^ w18195 ;
  assign w18197 = w7411 & w16670 ;
  assign w18198 = ( w7944 & ~w16662 ) | ( w7944 & w18197 ) | ( ~w16662 & w18197 ) ;
  assign w18199 = w7673 | w18198 ;
  assign w18200 = ( w16665 & w18198 ) | ( w16665 & w18199 ) | ( w18198 & w18199 ) ;
  assign w18201 = w18197 | w18200 ;
  assign w18202 = w7414 | w16762 ;
  assign w18203 = ( ~w16762 & w18201 ) | ( ~w16762 & w18202 ) | ( w18201 & w18202 ) ;
  assign w18204 = \pi08 ^ w18203 ;
  assign w18205 = w17950 ^ w17999 ;
  assign w18206 = w17942 ^ w18205 ;
  assign w18207 = w7411 & w16675 ;
  assign w18208 = ( w7944 & w16665 ) | ( w7944 & w18207 ) | ( w16665 & w18207 ) ;
  assign w18209 = w7673 | w18208 ;
  assign w18210 = ( w16670 & w18208 ) | ( w16670 & w18209 ) | ( w18208 & w18209 ) ;
  assign w18211 = w18207 | w18210 ;
  assign w18212 = ~w7414 & w16960 ;
  assign w18213 = ( w16960 & w18211 ) | ( w16960 & ~w18212 ) | ( w18211 & ~w18212 ) ;
  assign w18214 = \pi08 ^ w18213 ;
  assign w18215 = w17958 ^ w17998 ;
  assign w18216 = w17959 ^ w18215 ;
  assign w18217 = w7411 & w16680 ;
  assign w18218 = ( w7944 & w16670 ) | ( w7944 & w18217 ) | ( w16670 & w18217 ) ;
  assign w18219 = w7673 | w18218 ;
  assign w18220 = ( w16675 & w18218 ) | ( w16675 & w18219 ) | ( w18218 & w18219 ) ;
  assign w18221 = w18217 | w18220 ;
  assign w18222 = ~w7414 & w16972 ;
  assign w18223 = ( w16972 & w18221 ) | ( w16972 & ~w18222 ) | ( w18221 & ~w18222 ) ;
  assign w18224 = \pi08 ^ w18223 ;
  assign w18225 = ~w7673 & w16680 ;
  assign w18226 = w7411 & w16685 ;
  assign w18227 = ( w16680 & ~w18225 ) | ( w16680 & w18226 ) | ( ~w18225 & w18226 ) ;
  assign w18228 = ~w7944 & w16675 ;
  assign w18229 = w16946 | w18227 ;
  assign w18230 = ( w7414 & w18227 ) | ( w7414 & w18229 ) | ( w18227 & w18229 ) ;
  assign w18231 = ( w16675 & ~w18228 ) | ( w16675 & w18230 ) | ( ~w18228 & w18230 ) ;
  assign w18232 = \pi08 ^ w18231 ;
  assign w18233 = w17972 ^ w17997 ;
  assign w18234 = w17964 ^ w18233 ;
  assign w18235 = w17987 ^ w17995 ;
  assign w18236 = w17996 ^ w18235 ;
  assign w18237 = w7411 & ~w16690 ;
  assign w18238 = ( w7944 & w16680 ) | ( w7944 & w18237 ) | ( w16680 & w18237 ) ;
  assign w18239 = w7673 | w18238 ;
  assign w18240 = ( w16685 & w18238 ) | ( w16685 & w18239 ) | ( w18238 & w18239 ) ;
  assign w18241 = w18237 | w18240 ;
  assign w18242 = w7414 | w16772 ;
  assign w18243 = ( ~w16772 & w18241 ) | ( ~w16772 & w18242 ) | ( w18241 & w18242 ) ;
  assign w18244 = \pi08 ^ w18243 ;
  assign w18245 = w7673 | w16690 ;
  assign w18246 = w7411 & ~w16692 ;
  assign w18247 = ( ~w16690 & w18245 ) | ( ~w16690 & w18246 ) | ( w18245 & w18246 ) ;
  assign w18248 = ~w7944 & w16685 ;
  assign w18249 = w16818 | w18247 ;
  assign w18250 = ( w7414 & w18247 ) | ( w7414 & w18249 ) | ( w18247 & w18249 ) ;
  assign w18251 = ( w16685 & ~w18248 ) | ( w16685 & w18250 ) | ( ~w18248 & w18250 ) ;
  assign w18252 = \pi08 ^ w18251 ;
  assign w18253 = w17978 ^ w17986 ;
  assign w18254 = ( \pi08 & \pi09 ) | ( \pi08 & ~w16696 ) | ( \pi09 & ~w16696 ) ;
  assign w18255 = ( \pi08 & \pi09 ) | ( \pi08 & ~w16698 ) | ( \pi09 & ~w16698 ) ;
  assign w18256 = \pi10 ^ w16698 ;
  assign w18257 = ( \pi10 & w18255 ) | ( \pi10 & w18256 ) | ( w18255 & w18256 ) ;
  assign w18258 = w18254 ^ w18257 ;
  assign w18259 = w7411 & w16694 ;
  assign w18260 = ( w7944 & ~w16690 ) | ( w7944 & w18259 ) | ( ~w16690 & w18259 ) ;
  assign w18261 = w7673 | w18260 ;
  assign w18262 = ( ~w16692 & w18260 ) | ( ~w16692 & w18261 ) | ( w18260 & w18261 ) ;
  assign w18263 = w18259 | w18262 ;
  assign w18264 = w7414 | w16839 ;
  assign w18265 = ( ~w16839 & w18263 ) | ( ~w16839 & w18264 ) | ( w18263 & w18264 ) ;
  assign w18266 = \pi08 ^ w18265 ;
  assign w18267 = \pi08 & w16698 ;
  assign w18268 = w16696 & w18267 ;
  assign w18269 = ( \pi05 & \pi06 ) | ( \pi05 & ~w18268 ) | ( \pi06 & ~w18268 ) ;
  assign w18270 = ( \pi07 & \pi08 ) | ( \pi07 & ~w18269 ) | ( \pi08 & ~w18269 ) ;
  assign w18271 = ( \pi07 & ~w18267 ) | ( \pi07 & w18269 ) | ( ~w18267 & w18269 ) ;
  assign w18272 = ( w8885 & w18270 ) | ( w8885 & ~w18271 ) | ( w18270 & ~w18271 ) ;
  assign w18273 = w7411 & ~w16698 ;
  assign w18274 = ( w7944 & w16694 ) | ( w7944 & w18273 ) | ( w16694 & w18273 ) ;
  assign w18275 = w7673 | w18274 ;
  assign w18276 = ( ~w16696 & w18274 ) | ( ~w16696 & w18275 ) | ( w18274 & w18275 ) ;
  assign w18277 = w18273 | w18276 ;
  assign w18278 = ~w7414 & w16802 ;
  assign w18279 = ( w16802 & w18277 ) | ( w16802 & ~w18278 ) | ( w18277 & ~w18278 ) ;
  assign w18280 = \pi08 ^ w18279 ;
  assign w18281 = w18272 & w18280 ;
  assign w18282 = ~w7673 & w16694 ;
  assign w18283 = w7411 & ~w16696 ;
  assign w18284 = ( w16694 & ~w18282 ) | ( w16694 & w18283 ) | ( ~w18282 & w18283 ) ;
  assign w18285 = w7944 | w16692 ;
  assign w18286 = w16784 | w18284 ;
  assign w18287 = ( w7414 & w18284 ) | ( w7414 & w18286 ) | ( w18284 & w18286 ) ;
  assign w18288 = ( ~w16692 & w18285 ) | ( ~w16692 & w18287 ) | ( w18285 & w18287 ) ;
  assign w18289 = \pi08 ^ w18288 ;
  assign w18290 = w6750 & ~w16698 ;
  assign w18291 = ( w18281 & w18289 ) | ( w18281 & w18290 ) | ( w18289 & w18290 ) ;
  assign w18292 = ( w18258 & w18266 ) | ( w18258 & w18291 ) | ( w18266 & w18291 ) ;
  assign w18293 = ( w18252 & w18253 ) | ( w18252 & w18292 ) | ( w18253 & w18292 ) ;
  assign w18294 = ( w18236 & w18244 ) | ( w18236 & w18293 ) | ( w18244 & w18293 ) ;
  assign w18295 = ( w18232 & w18234 ) | ( w18232 & w18294 ) | ( w18234 & w18294 ) ;
  assign w18296 = ( w18216 & w18224 ) | ( w18216 & w18295 ) | ( w18224 & w18295 ) ;
  assign w18297 = ( w18206 & w18214 ) | ( w18206 & w18296 ) | ( w18214 & w18296 ) ;
  assign w18298 = ( w18196 & w18204 ) | ( w18196 & w18297 ) | ( w18204 & w18297 ) ;
  assign w18299 = ( w18192 & w18194 ) | ( w18192 & w18298 ) | ( w18194 & w18298 ) ;
  assign w18300 = ( w18182 & w18184 ) | ( w18182 & w18299 ) | ( w18184 & w18299 ) ;
  assign w18301 = ( w18172 & w18174 ) | ( w18172 & w18300 ) | ( w18174 & w18300 ) ;
  assign w18302 = ( w18156 & w18164 ) | ( w18156 & w18301 ) | ( w18164 & w18301 ) ;
  assign w18303 = ( w18146 & w18154 ) | ( w18146 & w18302 ) | ( w18154 & w18302 ) ;
  assign w18304 = ( w18136 & w18144 ) | ( w18136 & w18303 ) | ( w18144 & w18303 ) ;
  assign w18305 = ( w18132 & w18134 ) | ( w18132 & w18304 ) | ( w18134 & w18304 ) ;
  assign w18306 = ( w18122 & w18124 ) | ( w18122 & w18305 ) | ( w18124 & w18305 ) ;
  assign w18307 = ( w18112 & w18114 ) | ( w18112 & w18306 ) | ( w18114 & w18306 ) ;
  assign w18308 = ( w18096 & w18104 ) | ( w18096 & w18307 ) | ( w18104 & w18307 ) ;
  assign w18309 = ( w18086 & w18094 ) | ( w18086 & w18308 ) | ( w18094 & w18308 ) ;
  assign w18310 = ( w18076 & w18084 ) | ( w18076 & w18309 ) | ( w18084 & w18309 ) ;
  assign w18311 = ( w18072 & w18074 ) | ( w18072 & w18310 ) | ( w18074 & w18310 ) ;
  assign w18312 = ( w18062 & w18064 ) | ( w18062 & w18311 ) | ( w18064 & w18311 ) ;
  assign w18313 = ( ~w18043 & w18054 ) | ( ~w18043 & w18312 ) | ( w18054 & w18312 ) ;
  assign w18314 = ( ~w18031 & w18041 ) | ( ~w18031 & w18313 ) | ( w18041 & w18313 ) ;
  assign w18315 = ( w18019 & w18029 ) | ( w18019 & w18314 ) | ( w18029 & w18314 ) ;
  assign w18316 = w6949 | w16634 ;
  assign w18317 = w6748 & w16636 ;
  assign w18318 = ( ~w16634 & w18316 ) | ( ~w16634 & w18317 ) | ( w18316 & w18317 ) ;
  assign w18319 = ~w7154 & w16632 ;
  assign w18320 = w18051 & ~w18318 ;
  assign w18321 = ( w6751 & w18318 ) | ( w6751 & ~w18320 ) | ( w18318 & ~w18320 ) ;
  assign w18322 = ( w16632 & ~w18319 ) | ( w16632 & w18321 ) | ( ~w18319 & w18321 ) ;
  assign w18323 = \pi11 ^ w18322 ;
  assign w18324 = ( w17667 & w17753 ) | ( w17667 & w17763 ) | ( w17753 & w17763 ) ;
  assign w18325 = w5710 | w16646 ;
  assign w18326 = w5494 & ~w16648 ;
  assign w18327 = ( ~w16646 & w18325 ) | ( ~w16646 & w18326 ) | ( w18325 & w18326 ) ;
  assign w18328 = w5948 | w16644 ;
  assign w18329 = w17468 & ~w18327 ;
  assign w18330 = ( w5497 & w18327 ) | ( w5497 & ~w18329 ) | ( w18327 & ~w18329 ) ;
  assign w18331 = ( ~w16644 & w18328 ) | ( ~w16644 & w18330 ) | ( w18328 & w18330 ) ;
  assign w18332 = \pi17 ^ w18331 ;
  assign w18333 = ( w17676 & w17740 ) | ( w17676 & w17748 ) | ( w17740 & w17748 ) ;
  assign w18334 = w4651 | w16658 ;
  assign w18335 = w4606 & w16660 ;
  assign w18336 = ( ~w16658 & w18334 ) | ( ~w16658 & w18335 ) | ( w18334 & w18335 ) ;
  assign w18337 = w4706 | w16656 ;
  assign w18338 = w17057 | w18336 ;
  assign w18339 = ( w4609 & w18336 ) | ( w4609 & w18338 ) | ( w18336 & w18338 ) ;
  assign w18340 = ( ~w16656 & w18337 ) | ( ~w16656 & w18339 ) | ( w18337 & w18339 ) ;
  assign w18341 = \pi23 ^ w18340 ;
  assign w18342 = ( w17685 & w17727 ) | ( w17685 & w17735 ) | ( w17727 & w17735 ) ;
  assign w18343 = ~w3717 & w16680 ;
  assign w18344 = w3649 & w16685 ;
  assign w18345 = ( w16680 & ~w18343 ) | ( w16680 & w18344 ) | ( ~w18343 & w18344 ) ;
  assign w18346 = ~w3549 & w16675 ;
  assign w18347 = w16946 | w18345 ;
  assign w18348 = ( w3448 & w18345 ) | ( w3448 & w18347 ) | ( w18345 & w18347 ) ;
  assign w18349 = ( w16675 & ~w18346 ) | ( w16675 & w18348 ) | ( ~w18346 & w18348 ) ;
  assign w18350 = \pi29 ^ w18349 ;
  assign w18351 = ( w17694 & w17714 ) | ( w17694 & w17722 ) | ( w17714 & w17722 ) ;
  assign w18352 = ( w271 & w351 ) | ( w271 & ~w491 ) | ( w351 & ~w491 ) ;
  assign w18353 = w269 | w4352 ;
  assign w18354 = ( ~w269 & w491 ) | ( ~w269 & w1030 ) | ( w491 & w1030 ) ;
  assign w18355 = w18353 | w18354 ;
  assign w18356 = w18352 | w18355 ;
  assign w18357 = w178 | w698 ;
  assign w18358 = w18356 | w18357 ;
  assign w18359 = ( w177 & w10835 ) | ( w177 & ~w18356 ) | ( w10835 & ~w18356 ) ;
  assign w18360 = w18358 | w18359 ;
  assign w18361 = ( ~w514 & w10230 ) | ( ~w514 & w10257 ) | ( w10230 & w10257 ) ;
  assign w18362 = w12670 & ~w18360 ;
  assign w18363 = ( w260 & w514 ) | ( w260 & ~w18360 ) | ( w514 & ~w18360 ) ;
  assign w18364 = w18362 & ~w18363 ;
  assign w18365 = ~w18361 & w18364 ;
  assign w18366 = w315 | w570 ;
  assign w18367 = w103 | w18366 ;
  assign w18368 = ( w103 & ~w202 ) | ( w103 & w18365 ) | ( ~w202 & w18365 ) ;
  assign w18369 = ~w18367 & w18368 ;
  assign w18370 = w37 | w16839 ;
  assign w18371 = w3098 & w16694 ;
  assign w18372 = ( ~w16839 & w18370 ) | ( ~w16839 & w18371 ) | ( w18370 & w18371 ) ;
  assign w18373 = ( \pi29 & \pi30 ) | ( \pi29 & ~w16690 ) | ( \pi30 & ~w16690 ) ;
  assign w18374 = \pi31 | w18373 ;
  assign w18375 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w16692 ) | ( \pi30 & w16692 ) ;
  assign w18376 = ( \pi29 & \pi31 ) | ( \pi29 & w18375 ) | ( \pi31 & w18375 ) ;
  assign w18377 = ( w18372 & w18374 ) | ( w18372 & ~w18376 ) | ( w18374 & ~w18376 ) ;
  assign w18378 = w18351 ^ w18377 ;
  assign w18379 = w18369 ^ w18378 ;
  assign w18380 = ( w17693 & w17724 ) | ( w17693 & w17725 ) | ( w17724 & w17725 ) ;
  assign w18381 = w18350 ^ w18380 ;
  assign w18382 = w18379 ^ w18381 ;
  assign w18383 = w3964 & ~w16662 ;
  assign w18384 = ( w4143 & w16665 ) | ( w4143 & w18383 ) | ( w16665 & w18383 ) ;
  assign w18385 = w4052 | w18384 ;
  assign w18386 = ( w16670 & w18384 ) | ( w16670 & w18385 ) | ( w18384 & w18385 ) ;
  assign w18387 = w18383 | w18386 ;
  assign w18388 = w4147 | w16762 ;
  assign w18389 = ( ~w16762 & w18387 ) | ( ~w16762 & w18388 ) | ( w18387 & w18388 ) ;
  assign w18390 = \pi26 ^ w18389 ;
  assign w18391 = w18342 ^ w18390 ;
  assign w18392 = w18382 ^ w18391 ;
  assign w18393 = ( w17684 & w17737 ) | ( w17684 & w17738 ) | ( w17737 & w17738 ) ;
  assign w18394 = w18341 ^ w18393 ;
  assign w18395 = w18392 ^ w18394 ;
  assign w18396 = w4905 & w16654 ;
  assign w18397 = ( w5395 & ~w16650 ) | ( w5395 & w18396 ) | ( ~w16650 & w18396 ) ;
  assign w18398 = w5343 | w18397 ;
  assign w18399 = ( ~w16652 & w18397 ) | ( ~w16652 & w18398 ) | ( w18397 & w18398 ) ;
  assign w18400 = w18396 | w18399 ;
  assign w18401 = w4908 | w17277 ;
  assign w18402 = ( ~w17277 & w18400 ) | ( ~w17277 & w18401 ) | ( w18400 & w18401 ) ;
  assign w18403 = \pi20 ^ w18402 ;
  assign w18404 = w18333 ^ w18403 ;
  assign w18405 = w18395 ^ w18404 ;
  assign w18406 = ( w17675 & w17750 ) | ( w17675 & w17751 ) | ( w17750 & w17751 ) ;
  assign w18407 = w18332 ^ w18406 ;
  assign w18408 = w18405 ^ w18407 ;
  assign w18409 = w6048 & w16642 ;
  assign w18410 = ( w6637 & ~w16638 ) | ( w6637 & w18409 ) | ( ~w16638 & w18409 ) ;
  assign w18411 = w6549 | w18410 ;
  assign w18412 = ( w16640 & w18410 ) | ( w16640 & w18411 ) | ( w18410 & w18411 ) ;
  assign w18413 = w18409 | w18412 ;
  assign w18414 = w6045 | w17783 ;
  assign w18415 = ( ~w17783 & w18413 ) | ( ~w17783 & w18414 ) | ( w18413 & w18414 ) ;
  assign w18416 = \pi14 ^ w18415 ;
  assign w18417 = w18324 ^ w18416 ;
  assign w18418 = w18408 ^ w18417 ;
  assign w18419 = ( w16747 & w17765 ) | ( w16747 & w18017 ) | ( w17765 & w18017 ) ;
  assign w18420 = w18323 ^ w18419 ;
  assign w18421 = w18418 ^ w18420 ;
  assign w18422 = w7411 & ~w16630 ;
  assign w18423 = ( w7944 & ~w16626 ) | ( w7944 & w18422 ) | ( ~w16626 & w18422 ) ;
  assign w18424 = w7673 | w18423 ;
  assign w18425 = ( ~w16628 & w18423 ) | ( ~w16628 & w18424 ) | ( w18423 & w18424 ) ;
  assign w18426 = w18422 | w18425 ;
  assign w18427 = ( w16628 & w16630 ) | ( w16628 & ~w16724 ) | ( w16630 & ~w16724 ) ;
  assign w18428 = w16628 ^ w18427 ;
  assign w18429 = w16626 ^ w18428 ;
  assign w18430 = w7414 & w18429 ;
  assign w18431 = ( w7414 & w18426 ) | ( w7414 & ~w18430 ) | ( w18426 & ~w18430 ) ;
  assign w18432 = \pi08 ^ w18431 ;
  assign w18433 = w18315 ^ w18432 ;
  assign w18434 = w18421 ^ w18433 ;
  assign w18435 = ~w8593 & w16619 ;
  assign w18436 = w8262 & ~w16626 ;
  assign w18437 = ( w16619 & ~w18435 ) | ( w16619 & w18436 ) | ( ~w18435 & w18436 ) ;
  assign w18438 = w16621 ^ w16727 ;
  assign w18439 = w16619 ^ w18438 ;
  assign w18440 = w8263 | w18439 ;
  assign w18441 = w16621 | w18437 ;
  assign w18442 = ( w35 & w18437 ) | ( w35 & w18441 ) | ( w18437 & w18441 ) ;
  assign w18443 = ( ~w18439 & w18440 ) | ( ~w18439 & w18442 ) | ( w18440 & w18442 ) ;
  assign w18444 = \pi05 ^ w18443 ;
  assign w18445 = w18029 ^ w18314 ;
  assign w18446 = w18019 ^ w18445 ;
  assign w18447 = w8593 | w16626 ;
  assign w18448 = w8262 & ~w16628 ;
  assign w18449 = ( ~w16626 & w18447 ) | ( ~w16626 & w18448 ) | ( w18447 & w18448 ) ;
  assign w18450 = w16619 ^ w16726 ;
  assign w18451 = w16626 ^ w18450 ;
  assign w18452 = ~w8263 & w18451 ;
  assign w18453 = w16619 | w18449 ;
  assign w18454 = ( w35 & w18449 ) | ( w35 & w18453 ) | ( w18449 & w18453 ) ;
  assign w18455 = ( w18451 & ~w18452 ) | ( w18451 & w18454 ) | ( ~w18452 & w18454 ) ;
  assign w18456 = \pi05 ^ w18455 ;
  assign w18457 = w18041 ^ w18313 ;
  assign w18458 = w18031 ^ w18457 ;
  assign w18459 = w8593 | w16628 ;
  assign w18460 = w8262 & ~w16630 ;
  assign w18461 = ( ~w16628 & w18459 ) | ( ~w16628 & w18460 ) | ( w18459 & w18460 ) ;
  assign w18462 = w8263 | w18429 ;
  assign w18463 = w16626 & ~w18461 ;
  assign w18464 = ( w35 & w18461 ) | ( w35 & ~w18463 ) | ( w18461 & ~w18463 ) ;
  assign w18465 = ( ~w18429 & w18462 ) | ( ~w18429 & w18464 ) | ( w18462 & w18464 ) ;
  assign w18466 = \pi05 ^ w18465 ;
  assign w18467 = w18054 ^ w18312 ;
  assign w18468 = w18043 ^ w18467 ;
  assign w18469 = w18062 ^ w18311 ;
  assign w18470 = w18064 ^ w18469 ;
  assign w18471 = w35 & ~w16628 ;
  assign w18472 = ( w8593 & ~w16630 ) | ( w8593 & w18471 ) | ( ~w16630 & w18471 ) ;
  assign w18473 = w8262 | w18472 ;
  assign w18474 = ( w16632 & w18472 ) | ( w16632 & w18473 ) | ( w18472 & w18473 ) ;
  assign w18475 = w18471 | w18474 ;
  assign w18476 = ~w8263 & w18026 ;
  assign w18477 = ( w18026 & w18475 ) | ( w18026 & ~w18476 ) | ( w18475 & ~w18476 ) ;
  assign w18478 = \pi05 ^ w18477 ;
  assign w18479 = w18072 ^ w18310 ;
  assign w18480 = w18074 ^ w18479 ;
  assign w18481 = w35 & ~w16630 ;
  assign w18482 = ( w8593 & w16632 ) | ( w8593 & w18481 ) | ( w16632 & w18481 ) ;
  assign w18483 = w8262 | w18482 ;
  assign w18484 = ( ~w16634 & w18482 ) | ( ~w16634 & w18483 ) | ( w18482 & w18483 ) ;
  assign w18485 = w18481 | w18484 ;
  assign w18486 = w8263 | w18038 ;
  assign w18487 = ( ~w18038 & w18485 ) | ( ~w18038 & w18486 ) | ( w18485 & w18486 ) ;
  assign w18488 = \pi05 ^ w18487 ;
  assign w18489 = w8593 | w16634 ;
  assign w18490 = w8262 & w16636 ;
  assign w18491 = ( ~w16634 & w18489 ) | ( ~w16634 & w18490 ) | ( w18489 & w18490 ) ;
  assign w18492 = w8263 | w18051 ;
  assign w18493 = w16632 | w18491 ;
  assign w18494 = ( w35 & w18491 ) | ( w35 & w18493 ) | ( w18491 & w18493 ) ;
  assign w18495 = ( ~w18051 & w18492 ) | ( ~w18051 & w18494 ) | ( w18492 & w18494 ) ;
  assign w18496 = \pi05 ^ w18495 ;
  assign w18497 = w18084 ^ w18309 ;
  assign w18498 = w18076 ^ w18497 ;
  assign w18499 = ~w8593 & w16636 ;
  assign w18500 = w8262 & ~w16638 ;
  assign w18501 = ( w16636 & ~w18499 ) | ( w16636 & w18500 ) | ( ~w18499 & w18500 ) ;
  assign w18502 = w8263 | w16742 ;
  assign w18503 = w16634 & ~w18501 ;
  assign w18504 = ( w35 & w18501 ) | ( w35 & ~w18503 ) | ( w18501 & ~w18503 ) ;
  assign w18505 = ( ~w16742 & w18502 ) | ( ~w16742 & w18504 ) | ( w18502 & w18504 ) ;
  assign w18506 = \pi05 ^ w18505 ;
  assign w18507 = w18094 ^ w18308 ;
  assign w18508 = w18086 ^ w18507 ;
  assign w18509 = w8593 | w16638 ;
  assign w18510 = w8262 & w16640 ;
  assign w18511 = ( ~w16638 & w18509 ) | ( ~w16638 & w18510 ) | ( w18509 & w18510 ) ;
  assign w18512 = w8263 | w17770 ;
  assign w18513 = w16636 | w18511 ;
  assign w18514 = ( w35 & w18511 ) | ( w35 & w18513 ) | ( w18511 & w18513 ) ;
  assign w18515 = ( ~w17770 & w18512 ) | ( ~w17770 & w18514 ) | ( w18512 & w18514 ) ;
  assign w18516 = \pi05 ^ w18515 ;
  assign w18517 = w18104 ^ w18307 ;
  assign w18518 = w18096 ^ w18517 ;
  assign w18519 = w18112 ^ w18306 ;
  assign w18520 = w18114 ^ w18519 ;
  assign w18521 = w35 & ~w16638 ;
  assign w18522 = ( w8593 & w16640 ) | ( w8593 & w18521 ) | ( w16640 & w18521 ) ;
  assign w18523 = w8262 | w18522 ;
  assign w18524 = ( w16642 & w18522 ) | ( w16642 & w18523 ) | ( w18522 & w18523 ) ;
  assign w18525 = w18521 | w18524 ;
  assign w18526 = w8263 | w17783 ;
  assign w18527 = ( ~w17783 & w18525 ) | ( ~w17783 & w18526 ) | ( w18525 & w18526 ) ;
  assign w18528 = \pi05 ^ w18527 ;
  assign w18529 = w18122 ^ w18305 ;
  assign w18530 = w18124 ^ w18529 ;
  assign w18531 = w35 & w16640 ;
  assign w18532 = ( w8593 & w16642 ) | ( w8593 & w18531 ) | ( w16642 & w18531 ) ;
  assign w18533 = w8262 | w18532 ;
  assign w18534 = ( ~w16644 & w18532 ) | ( ~w16644 & w18533 ) | ( w18532 & w18533 ) ;
  assign w18535 = w18531 | w18534 ;
  assign w18536 = w8263 | w17760 ;
  assign w18537 = ( ~w17760 & w18535 ) | ( ~w17760 & w18536 ) | ( w18535 & w18536 ) ;
  assign w18538 = \pi05 ^ w18537 ;
  assign w18539 = w18132 ^ w18304 ;
  assign w18540 = w18134 ^ w18539 ;
  assign w18541 = w35 & w16642 ;
  assign w18542 = ( w8593 & ~w16644 ) | ( w8593 & w18541 ) | ( ~w16644 & w18541 ) ;
  assign w18543 = w8262 | w18542 ;
  assign w18544 = ( ~w16646 & w18542 ) | ( ~w16646 & w18543 ) | ( w18542 & w18543 ) ;
  assign w18545 = w18541 | w18544 ;
  assign w18546 = ~w8263 & w17455 ;
  assign w18547 = ( w17455 & w18545 ) | ( w17455 & ~w18546 ) | ( w18545 & ~w18546 ) ;
  assign w18548 = \pi05 ^ w18547 ;
  assign w18549 = w8593 | w16646 ;
  assign w18550 = w8262 & ~w16648 ;
  assign w18551 = ( ~w16646 & w18549 ) | ( ~w16646 & w18550 ) | ( w18549 & w18550 ) ;
  assign w18552 = w8263 | w17468 ;
  assign w18553 = w16644 & ~w18551 ;
  assign w18554 = ( w35 & w18551 ) | ( w35 & ~w18553 ) | ( w18551 & ~w18553 ) ;
  assign w18555 = ( ~w17468 & w18552 ) | ( ~w17468 & w18554 ) | ( w18552 & w18554 ) ;
  assign w18556 = \pi05 ^ w18555 ;
  assign w18557 = w18144 ^ w18303 ;
  assign w18558 = w18136 ^ w18557 ;
  assign w18559 = w8593 | w16648 ;
  assign w18560 = w8262 & ~w16650 ;
  assign w18561 = ( ~w16648 & w18559 ) | ( ~w16648 & w18560 ) | ( w18559 & w18560 ) ;
  assign w18562 = w8263 | w17476 ;
  assign w18563 = w16646 & ~w18561 ;
  assign w18564 = ( w35 & w18561 ) | ( w35 & ~w18563 ) | ( w18561 & ~w18563 ) ;
  assign w18565 = ( ~w17476 & w18562 ) | ( ~w17476 & w18564 ) | ( w18562 & w18564 ) ;
  assign w18566 = \pi05 ^ w18565 ;
  assign w18567 = w18154 ^ w18302 ;
  assign w18568 = w18146 ^ w18567 ;
  assign w18569 = w8593 | w16650 ;
  assign w18570 = w8262 & ~w16652 ;
  assign w18571 = ( ~w16650 & w18569 ) | ( ~w16650 & w18570 ) | ( w18569 & w18570 ) ;
  assign w18572 = w8263 | w16752 ;
  assign w18573 = w16648 & ~w18571 ;
  assign w18574 = ( w35 & w18571 ) | ( w35 & ~w18573 ) | ( w18571 & ~w18573 ) ;
  assign w18575 = ( ~w16752 & w18572 ) | ( ~w16752 & w18574 ) | ( w18572 & w18574 ) ;
  assign w18576 = \pi05 ^ w18575 ;
  assign w18577 = w18164 ^ w18301 ;
  assign w18578 = w18156 ^ w18577 ;
  assign w18579 = w18172 ^ w18300 ;
  assign w18580 = w18174 ^ w18579 ;
  assign w18581 = w35 & ~w16650 ;
  assign w18582 = ( w8593 & ~w16652 ) | ( w8593 & w18581 ) | ( ~w16652 & w18581 ) ;
  assign w18583 = w8262 | w18582 ;
  assign w18584 = ( w16654 & w18582 ) | ( w16654 & w18583 ) | ( w18582 & w18583 ) ;
  assign w18585 = w18581 | w18584 ;
  assign w18586 = w8263 | w17277 ;
  assign w18587 = ( ~w17277 & w18585 ) | ( ~w17277 & w18586 ) | ( w18585 & w18586 ) ;
  assign w18588 = \pi05 ^ w18587 ;
  assign w18589 = w18182 ^ w18299 ;
  assign w18590 = w18184 ^ w18589 ;
  assign w18591 = w35 & ~w16652 ;
  assign w18592 = ( w8593 & w16654 ) | ( w8593 & w18591 ) | ( w16654 & w18591 ) ;
  assign w18593 = w8262 | w18592 ;
  assign w18594 = ( ~w16656 & w18592 ) | ( ~w16656 & w18593 ) | ( w18592 & w18593 ) ;
  assign w18595 = w18591 | w18594 ;
  assign w18596 = ~w8263 & w17293 ;
  assign w18597 = ( w17293 & w18595 ) | ( w17293 & ~w18596 ) | ( w18595 & ~w18596 ) ;
  assign w18598 = \pi05 ^ w18597 ;
  assign w18599 = w18192 ^ w18298 ;
  assign w18600 = w18194 ^ w18599 ;
  assign w18601 = w35 & w16654 ;
  assign w18602 = ( w8593 & ~w16656 ) | ( w8593 & w18601 ) | ( ~w16656 & w18601 ) ;
  assign w18603 = w8262 | w18602 ;
  assign w18604 = ( ~w16658 & w18602 ) | ( ~w16658 & w18603 ) | ( w18602 & w18603 ) ;
  assign w18605 = w18601 | w18604 ;
  assign w18606 = ~w8263 & w17266 ;
  assign w18607 = ( w17266 & w18605 ) | ( w17266 & ~w18606 ) | ( w18605 & ~w18606 ) ;
  assign w18608 = \pi05 ^ w18607 ;
  assign w18609 = w8593 | w16658 ;
  assign w18610 = w8262 & w16660 ;
  assign w18611 = ( ~w16658 & w18609 ) | ( ~w16658 & w18610 ) | ( w18609 & w18610 ) ;
  assign w18612 = ~w8263 & w17057 ;
  assign w18613 = w16656 & ~w18611 ;
  assign w18614 = ( w35 & w18611 ) | ( w35 & ~w18613 ) | ( w18611 & ~w18613 ) ;
  assign w18615 = ( w17057 & ~w18612 ) | ( w17057 & w18614 ) | ( ~w18612 & w18614 ) ;
  assign w18616 = \pi05 ^ w18615 ;
  assign w18617 = w18204 ^ w18297 ;
  assign w18618 = w18196 ^ w18617 ;
  assign w18619 = ~w8593 & w16660 ;
  assign w18620 = w8262 & ~w16662 ;
  assign w18621 = ( w16660 & ~w18619 ) | ( w16660 & w18620 ) | ( ~w18619 & w18620 ) ;
  assign w18622 = w8263 | w17065 ;
  assign w18623 = w16658 & ~w18621 ;
  assign w18624 = ( w35 & w18621 ) | ( w35 & ~w18623 ) | ( w18621 & ~w18623 ) ;
  assign w18625 = ( ~w17065 & w18622 ) | ( ~w17065 & w18624 ) | ( w18622 & w18624 ) ;
  assign w18626 = \pi05 ^ w18625 ;
  assign w18627 = w18214 ^ w18296 ;
  assign w18628 = w18206 ^ w18627 ;
  assign w18629 = w8593 | w16662 ;
  assign w18630 = w8262 & w16665 ;
  assign w18631 = ( ~w16662 & w18629 ) | ( ~w16662 & w18630 ) | ( w18629 & w18630 ) ;
  assign w18632 = w8263 | w17078 ;
  assign w18633 = w16660 | w18631 ;
  assign w18634 = ( w35 & w18631 ) | ( w35 & w18633 ) | ( w18631 & w18633 ) ;
  assign w18635 = ( ~w17078 & w18632 ) | ( ~w17078 & w18634 ) | ( w18632 & w18634 ) ;
  assign w18636 = \pi05 ^ w18635 ;
  assign w18637 = w18224 ^ w18295 ;
  assign w18638 = w18216 ^ w18637 ;
  assign w18639 = w18232 ^ w18294 ;
  assign w18640 = w18234 ^ w18639 ;
  assign w18641 = w35 & ~w16662 ;
  assign w18642 = ( w8593 & w16665 ) | ( w8593 & w18641 ) | ( w16665 & w18641 ) ;
  assign w18643 = w8262 | w18642 ;
  assign w18644 = ( w16670 & w18642 ) | ( w16670 & w18643 ) | ( w18642 & w18643 ) ;
  assign w18645 = w18641 | w18644 ;
  assign w18646 = w8263 | w16762 ;
  assign w18647 = ( ~w16762 & w18645 ) | ( ~w16762 & w18646 ) | ( w18645 & w18646 ) ;
  assign w18648 = \pi05 ^ w18647 ;
  assign w18649 = w18244 ^ w18293 ;
  assign w18650 = w18236 ^ w18649 ;
  assign w18651 = w35 & w16665 ;
  assign w18652 = ( w8593 & w16670 ) | ( w8593 & w18651 ) | ( w16670 & w18651 ) ;
  assign w18653 = w8262 | w18652 ;
  assign w18654 = ( w16675 & w18652 ) | ( w16675 & w18653 ) | ( w18652 & w18653 ) ;
  assign w18655 = w18651 | w18654 ;
  assign w18656 = ~w8263 & w16960 ;
  assign w18657 = ( w16960 & w18655 ) | ( w16960 & ~w18656 ) | ( w18655 & ~w18656 ) ;
  assign w18658 = \pi05 ^ w18657 ;
  assign w18659 = w18252 ^ w18292 ;
  assign w18660 = w18253 ^ w18659 ;
  assign w18661 = w35 & w16670 ;
  assign w18662 = ( w8593 & w16675 ) | ( w8593 & w18661 ) | ( w16675 & w18661 ) ;
  assign w18663 = w8262 | w18662 ;
  assign w18664 = ( w16680 & w18662 ) | ( w16680 & w18663 ) | ( w18662 & w18663 ) ;
  assign w18665 = w18661 | w18664 ;
  assign w18666 = ~w8263 & w16972 ;
  assign w18667 = ( w16972 & w18665 ) | ( w16972 & ~w18666 ) | ( w18665 & ~w18666 ) ;
  assign w18668 = \pi05 ^ w18667 ;
  assign w18669 = ~w8593 & w16680 ;
  assign w18670 = w8262 & w16685 ;
  assign w18671 = ( w16680 & ~w18669 ) | ( w16680 & w18670 ) | ( ~w18669 & w18670 ) ;
  assign w18672 = ~w8263 & w16946 ;
  assign w18673 = w16675 | w18671 ;
  assign w18674 = ( w35 & w18671 ) | ( w35 & w18673 ) | ( w18671 & w18673 ) ;
  assign w18675 = ( w16946 & ~w18672 ) | ( w16946 & w18674 ) | ( ~w18672 & w18674 ) ;
  assign w18676 = \pi05 ^ w18675 ;
  assign w18677 = w18266 ^ w18291 ;
  assign w18678 = w18258 ^ w18677 ;
  assign w18679 = w18281 ^ w18289 ;
  assign w18680 = w18290 ^ w18679 ;
  assign w18681 = w35 & w16680 ;
  assign w18682 = ( w8593 & w16685 ) | ( w8593 & w18681 ) | ( w16685 & w18681 ) ;
  assign w18683 = w8262 | w18682 ;
  assign w18684 = ( ~w16690 & w18682 ) | ( ~w16690 & w18683 ) | ( w18682 & w18683 ) ;
  assign w18685 = w18681 | w18684 ;
  assign w18686 = w8263 | w16772 ;
  assign w18687 = ( ~w16772 & w18685 ) | ( ~w16772 & w18686 ) | ( w18685 & w18686 ) ;
  assign w18688 = \pi05 ^ w18687 ;
  assign w18689 = w8593 | w16690 ;
  assign w18690 = w8262 & ~w16692 ;
  assign w18691 = ( ~w16690 & w18689 ) | ( ~w16690 & w18690 ) | ( w18689 & w18690 ) ;
  assign w18692 = ~w8263 & w16818 ;
  assign w18693 = w16685 | w18691 ;
  assign w18694 = ( w35 & w18691 ) | ( w35 & w18693 ) | ( w18691 & w18693 ) ;
  assign w18695 = ( w16818 & ~w18692 ) | ( w16818 & w18694 ) | ( ~w18692 & w18694 ) ;
  assign w18696 = \pi05 ^ w18695 ;
  assign w18697 = w18272 ^ w18280 ;
  assign w18698 = ( \pi05 & \pi06 ) | ( \pi05 & ~w16696 ) | ( \pi06 & ~w16696 ) ;
  assign w18699 = ( \pi05 & \pi06 ) | ( \pi05 & ~w16698 ) | ( \pi06 & ~w16698 ) ;
  assign w18700 = \pi07 ^ w16698 ;
  assign w18701 = ( \pi07 & w18699 ) | ( \pi07 & w18700 ) | ( w18699 & w18700 ) ;
  assign w18702 = w18698 ^ w18701 ;
  assign w18703 = w35 & ~w16690 ;
  assign w18704 = ( w8593 & ~w16692 ) | ( w8593 & w18703 ) | ( ~w16692 & w18703 ) ;
  assign w18705 = w8262 | w18704 ;
  assign w18706 = ( w16694 & w18704 ) | ( w16694 & w18705 ) | ( w18704 & w18705 ) ;
  assign w18707 = w18703 | w18706 ;
  assign w18708 = w8263 | w16839 ;
  assign w18709 = ( ~w16839 & w18707 ) | ( ~w16839 & w18708 ) | ( w18707 & w18708 ) ;
  assign w18710 = \pi05 ^ w18709 ;
  assign w18711 = w16696 ^ w16698 ;
  assign w18712 = ( w8593 & ~w16696 ) | ( w8593 & w18711 ) | ( ~w16696 & w18711 ) ;
  assign w18713 = ( ~w8263 & w16696 ) | ( ~w8263 & w16698 ) | ( w16696 & w16698 ) ;
  assign w18714 = w35 | w16696 ;
  assign w18715 = ( w18712 & ~w18713 ) | ( w18712 & w18714 ) | ( ~w18713 & w18714 ) ;
  assign w18716 = w34 & ~w16698 ;
  assign w18717 = ( \pi05 & ~w18715 ) | ( \pi05 & w18716 ) | ( ~w18715 & w18716 ) ;
  assign w18718 = ~w18716 & w18717 ;
  assign w18719 = w35 & w16694 ;
  assign w18720 = ( w8593 & ~w16696 ) | ( w8593 & w18719 ) | ( ~w16696 & w18719 ) ;
  assign w18721 = w8262 | w18720 ;
  assign w18722 = ( ~w16698 & w18720 ) | ( ~w16698 & w18721 ) | ( w18720 & w18721 ) ;
  assign w18723 = w18719 | w18722 ;
  assign w18724 = ~w8263 & w16802 ;
  assign w18725 = ( w16802 & w18723 ) | ( w16802 & ~w18724 ) | ( w18723 & ~w18724 ) ;
  assign w18726 = \pi05 ^ w18725 ;
  assign w18727 = w18718 & w18726 ;
  assign w18728 = ~w8593 & w16694 ;
  assign w18729 = w8262 & ~w16696 ;
  assign w18730 = ( w16694 & ~w18728 ) | ( w16694 & w18729 ) | ( ~w18728 & w18729 ) ;
  assign w18731 = ~w8263 & w16784 ;
  assign w18732 = w16692 & ~w18730 ;
  assign w18733 = ( w35 & w18730 ) | ( w35 & ~w18732 ) | ( w18730 & ~w18732 ) ;
  assign w18734 = ( w16784 & ~w18731 ) | ( w16784 & w18733 ) | ( ~w18731 & w18733 ) ;
  assign w18735 = \pi05 ^ w18734 ;
  assign w18736 = w7413 & ~w16698 ;
  assign w18737 = ( w18727 & w18735 ) | ( w18727 & w18736 ) | ( w18735 & w18736 ) ;
  assign w18738 = ( w18702 & w18710 ) | ( w18702 & w18737 ) | ( w18710 & w18737 ) ;
  assign w18739 = ( w18696 & w18697 ) | ( w18696 & w18738 ) | ( w18697 & w18738 ) ;
  assign w18740 = ( w18680 & w18688 ) | ( w18680 & w18739 ) | ( w18688 & w18739 ) ;
  assign w18741 = ( w18676 & w18678 ) | ( w18676 & w18740 ) | ( w18678 & w18740 ) ;
  assign w18742 = ( w18660 & w18668 ) | ( w18660 & w18741 ) | ( w18668 & w18741 ) ;
  assign w18743 = ( w18650 & w18658 ) | ( w18650 & w18742 ) | ( w18658 & w18742 ) ;
  assign w18744 = ( w18640 & w18648 ) | ( w18640 & w18743 ) | ( w18648 & w18743 ) ;
  assign w18745 = ( w18636 & w18638 ) | ( w18636 & w18744 ) | ( w18638 & w18744 ) ;
  assign w18746 = ( w18626 & w18628 ) | ( w18626 & w18745 ) | ( w18628 & w18745 ) ;
  assign w18747 = ( w18616 & w18618 ) | ( w18616 & w18746 ) | ( w18618 & w18746 ) ;
  assign w18748 = ( w18600 & w18608 ) | ( w18600 & w18747 ) | ( w18608 & w18747 ) ;
  assign w18749 = ( w18590 & w18598 ) | ( w18590 & w18748 ) | ( w18598 & w18748 ) ;
  assign w18750 = ( w18580 & w18588 ) | ( w18580 & w18749 ) | ( w18588 & w18749 ) ;
  assign w18751 = ( w18576 & w18578 ) | ( w18576 & w18750 ) | ( w18578 & w18750 ) ;
  assign w18752 = ( w18566 & w18568 ) | ( w18566 & w18751 ) | ( w18568 & w18751 ) ;
  assign w18753 = ( w18556 & w18558 ) | ( w18556 & w18752 ) | ( w18558 & w18752 ) ;
  assign w18754 = ( w18540 & w18548 ) | ( w18540 & w18753 ) | ( w18548 & w18753 ) ;
  assign w18755 = ( w18530 & w18538 ) | ( w18530 & w18754 ) | ( w18538 & w18754 ) ;
  assign w18756 = ( w18520 & w18528 ) | ( w18520 & w18755 ) | ( w18528 & w18755 ) ;
  assign w18757 = ( w18516 & w18518 ) | ( w18516 & w18756 ) | ( w18518 & w18756 ) ;
  assign w18758 = ( w18506 & w18508 ) | ( w18506 & w18757 ) | ( w18508 & w18757 ) ;
  assign w18759 = ( w18496 & w18498 ) | ( w18496 & w18758 ) | ( w18498 & w18758 ) ;
  assign w18760 = ( w18480 & w18488 ) | ( w18480 & w18759 ) | ( w18488 & w18759 ) ;
  assign w18761 = ( w18470 & w18478 ) | ( w18470 & w18760 ) | ( w18478 & w18760 ) ;
  assign w18762 = ( w18466 & ~w18468 ) | ( w18466 & w18761 ) | ( ~w18468 & w18761 ) ;
  assign w18763 = ( w18456 & ~w18458 ) | ( w18456 & w18762 ) | ( ~w18458 & w18762 ) ;
  assign w18764 = ( w18444 & w18446 ) | ( w18444 & w18763 ) | ( w18446 & w18763 ) ;
  assign w18765 = w16737 ^ w18764 ;
  assign w18766 = w18434 ^ w18765 ;
  assign w18767 = ( w16602 & w16603 ) | ( w16602 & w16611 ) | ( w16603 & w16611 ) ;
  assign w18768 = ( w10851 & ~w16574 ) | ( w10851 & w16600 ) | ( ~w16574 & w16600 ) ;
  assign w18769 = ( w10850 & ~w16578 ) | ( w10850 & w16598 ) | ( ~w16578 & w16598 ) ;
  assign w18770 = ( w785 & ~w1881 ) | ( w785 & w6365 ) | ( ~w1881 & w6365 ) ;
  assign w18771 = w1881 | w18770 ;
  assign w18772 = ( w215 & w447 ) | ( w215 & ~w625 ) | ( w447 & ~w625 ) ;
  assign w18773 = w3965 | w18771 ;
  assign w18774 = ( w625 & w1229 ) | ( w625 & ~w3965 ) | ( w1229 & ~w3965 ) ;
  assign w18775 = w18773 | w18774 ;
  assign w18776 = w18772 | w18775 ;
  assign w18777 = ( ~w139 & w3861 ) | ( ~w139 & w10407 ) | ( w3861 & w10407 ) ;
  assign w18778 = w3490 & ~w3522 ;
  assign w18779 = ( w139 & w802 ) | ( w139 & w3490 ) | ( w802 & w3490 ) ;
  assign w18780 = w18778 & ~w18779 ;
  assign w18781 = ~w18777 & w18780 ;
  assign w18782 = w149 | w214 ;
  assign w18783 = w18776 | w18782 ;
  assign w18784 = ( ~w2374 & w18776 ) | ( ~w2374 & w18781 ) | ( w18776 & w18781 ) ;
  assign w18785 = ~w18783 & w18784 ;
  assign w18786 = w351 | w495 ;
  assign w18787 = w1401 | w18786 ;
  assign w18788 = ( ~w278 & w1401 ) | ( ~w278 & w18785 ) | ( w1401 & w18785 ) ;
  assign w18789 = ~w18787 & w18788 ;
  assign w18790 = ~w37 & w10814 ;
  assign w18791 = w3098 & ~w10805 ;
  assign w18792 = ( w10814 & ~w18790 ) | ( w10814 & w18791 ) | ( ~w18790 & w18791 ) ;
  assign w18793 = ( \pi29 & \pi30 ) | ( \pi29 & w10801 ) | ( \pi30 & w10801 ) ;
  assign w18794 = \pi31 | w18793 ;
  assign w18795 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w10807 ) | ( \pi30 & w10807 ) ;
  assign w18796 = ( \pi29 & \pi31 ) | ( \pi29 & w18795 ) | ( \pi31 & w18795 ) ;
  assign w18797 = ( w18792 & w18794 ) | ( w18792 & ~w18796 ) | ( w18794 & ~w18796 ) ;
  assign w18798 = w18769 ^ w18797 ;
  assign w18799 = w18789 ^ w18798 ;
  assign w18800 = w3717 | w10885 ;
  assign w18801 = w3649 & ~w10866 ;
  assign w18802 = ( ~w10885 & w18800 ) | ( ~w10885 & w18801 ) | ( w18800 & w18801 ) ;
  assign w18803 = w3549 | w10887 ;
  assign w18804 = w11131 & ~w18802 ;
  assign w18805 = ( w3448 & w18802 ) | ( w3448 & ~w18804 ) | ( w18802 & ~w18804 ) ;
  assign w18806 = ( ~w10887 & w18803 ) | ( ~w10887 & w18805 ) | ( w18803 & w18805 ) ;
  assign w18807 = \pi29 ^ w18806 ;
  assign w18808 = w18768 ^ w18799 ;
  assign w18809 = w18807 ^ w18808 ;
  assign w18810 = w4143 | w11139 ;
  assign w18811 = w4052 & w10883 ;
  assign w18812 = ( ~w11139 & w18810 ) | ( ~w11139 & w18811 ) | ( w18810 & w18811 ) ;
  assign w18813 = w4147 | w11145 ;
  assign w18814 = w10738 & ~w18812 ;
  assign w18815 = ( w3964 & w18812 ) | ( w3964 & ~w18814 ) | ( w18812 & ~w18814 ) ;
  assign w18816 = ( ~w11145 & w18813 ) | ( ~w11145 & w18815 ) | ( w18813 & w18815 ) ;
  assign w18817 = \pi26 ^ w18816 ;
  assign w18818 = ( w18767 & ~w18809 ) | ( w18767 & w18817 ) | ( ~w18809 & w18817 ) ;
  assign w18819 = ( \pi29 & \pi31 ) | ( \pi29 & w10801 ) | ( \pi31 & w10801 ) ;
  assign w18820 = ( \pi29 & ~\pi30 ) | ( \pi29 & w18819 ) | ( ~\pi30 & w18819 ) ;
  assign w18821 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w18819 ) | ( \pi30 & w18819 ) ;
  assign w18822 = ( \pi29 & w10807 ) | ( \pi29 & ~w18821 ) | ( w10807 & ~w18821 ) ;
  assign w18823 = ( ~w10866 & w18821 ) | ( ~w10866 & w18822 ) | ( w18821 & w18822 ) ;
  assign w18824 = ~\pi31 & w18823 ;
  assign w18825 = ( w18820 & ~w18822 ) | ( w18820 & w18824 ) | ( ~w18822 & w18824 ) ;
  assign w18826 = ( w37 & w10874 ) | ( w37 & w18825 ) | ( w10874 & w18825 ) ;
  assign w18827 = w18825 | w18826 ;
  assign w18828 = ( w133 & ~w465 ) | ( w133 & w1069 ) | ( ~w465 & w1069 ) ;
  assign w18829 = w468 | w4066 ;
  assign w18830 = ( w465 & w466 ) | ( w465 & ~w468 ) | ( w466 & ~w468 ) ;
  assign w18831 = w18829 | w18830 ;
  assign w18832 = w18828 | w18831 ;
  assign w18833 = w1783 | w2253 ;
  assign w18834 = w18832 | w18833 ;
  assign w18835 = ( w3881 & w10407 ) | ( w3881 & ~w18832 ) | ( w10407 & ~w18832 ) ;
  assign w18836 = w18834 | w18835 ;
  assign w18837 = ( w144 & w278 ) | ( w144 & ~w605 ) | ( w278 & ~w605 ) ;
  assign w18838 = w3853 | w18836 ;
  assign w18839 = ( w605 & w758 ) | ( w605 & ~w18836 ) | ( w758 & ~w18836 ) ;
  assign w18840 = w18838 | w18839 ;
  assign w18841 = w18837 | w18840 ;
  assign w18842 = ( ~w111 & w223 ) | ( ~w111 & w18841 ) | ( w223 & w18841 ) ;
  assign w18843 = w111 | w18842 ;
  assign w18844 = ( w18789 & w18827 ) | ( w18789 & w18843 ) | ( w18827 & w18843 ) ;
  assign w18845 = w18789 ^ w18827 ;
  assign w18846 = w18843 ^ w18845 ;
  assign w18847 = ( w18769 & w18789 ) | ( w18769 & w18797 ) | ( w18789 & w18797 ) ;
  assign w18848 = ( ~w18768 & w18799 ) | ( ~w18768 & w18807 ) | ( w18799 & w18807 ) ;
  assign w18849 = w18847 ^ w18848 ;
  assign w18850 = w18846 ^ w18849 ;
  assign w18851 = w3964 | w4143 ;
  assign w18852 = w4147 & ~w11138 ;
  assign w18853 = ( w4147 & w11144 ) | ( w4147 & w18852 ) | ( w11144 & w18852 ) ;
  assign w18854 = ( w4052 & ~w11138 ) | ( w4052 & w18852 ) | ( ~w11138 & w18852 ) ;
  assign w18855 = w18851 & ~w18854 ;
  assign w18856 = ( ~w10738 & w18854 ) | ( ~w10738 & w18855 ) | ( w18854 & w18855 ) ;
  assign w18857 = ( w4147 & ~w18853 ) | ( w4147 & w18856 ) | ( ~w18853 & w18856 ) ;
  assign w18858 = w3717 | w10887 ;
  assign w18859 = w3649 & ~w10885 ;
  assign w18860 = ( ~w10887 & w18858 ) | ( ~w10887 & w18859 ) | ( w18858 & w18859 ) ;
  assign w18861 = ~w3549 & w10883 ;
  assign w18862 = w10895 | w18860 ;
  assign w18863 = ( w3448 & w18860 ) | ( w3448 & w18862 ) | ( w18860 & w18862 ) ;
  assign w18864 = ( w10883 & ~w18861 ) | ( w10883 & w18863 ) | ( ~w18861 & w18863 ) ;
  assign w18865 = \pi29 ^ w18864 ;
  assign w18866 = \pi26 ^ w18865 ;
  assign w18867 = w18850 ^ w18866 ;
  assign w18868 = w18857 ^ w18867 ;
  assign w18869 = w18767 ^ w18809 ;
  assign w18870 = w18817 ^ w18869 ;
  assign w18871 = ( w16557 & w16565 ) | ( w16557 & w16613 ) | ( w16565 & w16613 ) ;
  assign w18872 = ( w16552 & w16556 ) | ( w16552 & w16615 ) | ( w16556 & w16615 ) ;
  assign w18873 = ( ~w18870 & w18871 ) | ( ~w18870 & w18872 ) | ( w18871 & w18872 ) ;
  assign w18874 = ( w18818 & w18868 ) | ( w18818 & w18873 ) | ( w18868 & w18873 ) ;
  assign w18875 = ( \pi29 & \pi31 ) | ( \pi29 & ~w10866 ) | ( \pi31 & ~w10866 ) ;
  assign w18876 = ( \pi29 & ~\pi30 ) | ( \pi29 & w18875 ) | ( ~\pi30 & w18875 ) ;
  assign w18877 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w18875 ) | ( \pi30 & w18875 ) ;
  assign w18878 = ( ~\pi29 & w10801 ) | ( ~\pi29 & w18877 ) | ( w10801 & w18877 ) ;
  assign w18879 = ( w10885 & ~w18877 ) | ( w10885 & w18878 ) | ( ~w18877 & w18878 ) ;
  assign w18880 = \pi31 | w18879 ;
  assign w18881 = ( w18876 & w18878 ) | ( w18876 & ~w18880 ) | ( w18878 & ~w18880 ) ;
  assign w18882 = ( w37 & ~w11160 ) | ( w37 & w18881 ) | ( ~w11160 & w18881 ) ;
  assign w18883 = w18881 | w18882 ;
  assign w18884 = ( \pi25 & ~\pi26 ) | ( \pi25 & w99 ) | ( ~\pi26 & w99 ) ;
  assign w18885 = w10738 ^ w18884 ;
  assign w18886 = ( \pi26 & w18884 ) | ( \pi26 & w18885 ) | ( w18884 & w18885 ) ;
  assign w18887 = ( w278 & ~w3958 ) | ( w278 & w4057 ) | ( ~w3958 & w4057 ) ;
  assign w18888 = w3958 | w18887 ;
  assign w18889 = ( ~w312 & w2873 ) | ( ~w312 & w18888 ) | ( w2873 & w18888 ) ;
  assign w18890 = w4110 & ~w4137 ;
  assign w18891 = ( w312 & w605 ) | ( w312 & ~w4137 ) | ( w605 & ~w4137 ) ;
  assign w18892 = w18890 & ~w18891 ;
  assign w18893 = ~w18889 & w18892 ;
  assign w18894 = w18789 ^ w18886 ;
  assign w18895 = w18893 ^ w18894 ;
  assign w18896 = w18844 ^ w18895 ;
  assign w18897 = w18883 ^ w18896 ;
  assign w18898 = ~w3717 & w10883 ;
  assign w18899 = w3649 & ~w10887 ;
  assign w18900 = ( w10883 & ~w18898 ) | ( w10883 & w18899 ) | ( ~w18898 & w18899 ) ;
  assign w18901 = w3549 | w11139 ;
  assign w18902 = w11256 | w18900 ;
  assign w18903 = ( w3448 & w18900 ) | ( w3448 & w18902 ) | ( w18900 & w18902 ) ;
  assign w18904 = ( ~w11139 & w18901 ) | ( ~w11139 & w18903 ) | ( w18901 & w18903 ) ;
  assign w18905 = \pi29 ^ w18904 ;
  assign w18906 = ( w18846 & w18847 ) | ( w18846 & w18848 ) | ( w18847 & w18848 ) ;
  assign w18907 = w18897 ^ w18906 ;
  assign w18908 = w18905 ^ w18907 ;
  assign w18909 = \pi26 ^ w18857 ;
  assign w18910 = ( w18850 & w18865 ) | ( w18850 & w18909 ) | ( w18865 & w18909 ) ;
  assign w18911 = w18874 ^ w18908 ;
  assign w18912 = w18910 ^ w18911 ;
  assign w18913 = w18870 ^ w18872 ;
  assign w18914 = w18871 ^ w18913 ;
  assign w18915 = w18868 ^ w18873 ;
  assign w18916 = w18818 ^ w18915 ;
  assign w18917 = ( \pi02 & w18912 ) | ( \pi02 & ~w18916 ) | ( w18912 & ~w18916 ) ;
  assign w18918 = \pi00 ^ w18917 ;
  assign w18919 = ( \pi02 & ~w18912 ) | ( \pi02 & w18918 ) | ( ~w18912 & w18918 ) ;
  assign w18920 = ( \pi02 & w18916 ) | ( \pi02 & ~w18918 ) | ( w18916 & ~w18918 ) ;
  assign w18921 = \pi01 & w18920 ;
  assign w18922 = ( \pi00 & w18914 ) | ( \pi00 & ~w18921 ) | ( w18914 & ~w18921 ) ;
  assign w18923 = ( \pi01 & \pi02 ) | ( \pi01 & w18922 ) | ( \pi02 & w18922 ) ;
  assign w18924 = ( w18919 & w18921 ) | ( w18919 & ~w18923 ) | ( w18921 & ~w18923 ) ;
  assign w18925 = ( w16617 & w16729 ) | ( w16617 & ~w18914 ) | ( w16729 & ~w18914 ) ;
  assign w18926 = ( ~w18914 & w18916 ) | ( ~w18914 & w18925 ) | ( w18916 & w18925 ) ;
  assign w18927 = ( ~w18912 & w18916 ) | ( ~w18912 & w18926 ) | ( w18916 & w18926 ) ;
  assign w18928 = w18912 ^ w18926 ;
  assign w18929 = w18916 ^ w18928 ;
  assign w18930 = w8954 & w18929 ;
  assign w18931 = ( w8954 & w18924 ) | ( w8954 & ~w18930 ) | ( w18924 & ~w18930 ) ;
  assign w18932 = \pi02 ^ w18931 ;
  assign w18933 = \pi00 ^ w16694 ;
  assign w18934 = ( \pi01 & w16694 ) | ( \pi01 & ~w18933 ) | ( w16694 & ~w18933 ) ;
  assign w18935 = ( \pi00 & ~w16696 ) | ( \pi00 & w18934 ) | ( ~w16696 & w18934 ) ;
  assign w18936 = ( \pi02 & ~w16698 ) | ( \pi02 & w18935 ) | ( ~w16698 & w18935 ) ;
  assign w18937 = \pi02 & ~w18936 ;
  assign w18938 = ( \pi02 & w16692 ) | ( \pi02 & ~w16694 ) | ( w16692 & ~w16694 ) ;
  assign w18939 = \pi00 ^ w18938 ;
  assign w18940 = ( \pi02 & ~w16692 ) | ( \pi02 & w18939 ) | ( ~w16692 & w18939 ) ;
  assign w18941 = ( \pi02 & w16694 ) | ( \pi02 & ~w18939 ) | ( w16694 & ~w18939 ) ;
  assign w18942 = \pi01 & w18941 ;
  assign w18943 = ( \pi00 & w16696 ) | ( \pi00 & ~w18942 ) | ( w16696 & ~w18942 ) ;
  assign w18944 = ( \pi01 & \pi02 ) | ( \pi01 & w18943 ) | ( \pi02 & w18943 ) ;
  assign w18945 = ( w18940 & w18942 ) | ( w18940 & ~w18944 ) | ( w18942 & ~w18944 ) ;
  assign w18946 = w16784 | w18945 ;
  assign w18947 = ( w8954 & w18945 ) | ( w8954 & w18946 ) | ( w18945 & w18946 ) ;
  assign w18948 = \pi02 ^ w18947 ;
  assign w18949 = ( w18716 & w18937 ) | ( w18716 & w18948 ) | ( w18937 & w18948 ) ;
  assign w18950 = ( \pi02 & w16690 ) | ( \pi02 & w16692 ) | ( w16690 & w16692 ) ;
  assign w18951 = \pi00 ^ w18950 ;
  assign w18952 = ( \pi02 & ~w16690 ) | ( \pi02 & w18951 ) | ( ~w16690 & w18951 ) ;
  assign w18953 = ( ~\pi02 & w16692 ) | ( ~\pi02 & w18951 ) | ( w16692 & w18951 ) ;
  assign w18954 = \pi01 & ~w18953 ;
  assign w18955 = ( ~\pi00 & w16694 ) | ( ~\pi00 & w18954 ) | ( w16694 & w18954 ) ;
  assign w18956 = ( \pi01 & \pi02 ) | ( \pi01 & ~w18955 ) | ( \pi02 & ~w18955 ) ;
  assign w18957 = ( w18952 & w18954 ) | ( w18952 & ~w18956 ) | ( w18954 & ~w18956 ) ;
  assign w18958 = w8954 | w16839 ;
  assign w18959 = ( ~w16839 & w18957 ) | ( ~w16839 & w18958 ) | ( w18957 & w18958 ) ;
  assign w18960 = \pi02 ^ w18959 ;
  assign w18961 = \pi05 & w18716 ;
  assign w18962 = w18715 ^ w18961 ;
  assign w18963 = ( w18949 & w18960 ) | ( w18949 & w18962 ) | ( w18960 & w18962 ) ;
  assign w18964 = ( \pi02 & ~w16685 ) | ( \pi02 & w16690 ) | ( ~w16685 & w16690 ) ;
  assign w18965 = \pi00 ^ w18964 ;
  assign w18966 = ( \pi02 & w16685 ) | ( \pi02 & w18965 ) | ( w16685 & w18965 ) ;
  assign w18967 = ( ~\pi02 & w16690 ) | ( ~\pi02 & w18965 ) | ( w16690 & w18965 ) ;
  assign w18968 = \pi01 & ~w18967 ;
  assign w18969 = ( \pi00 & w16692 ) | ( \pi00 & ~w18968 ) | ( w16692 & ~w18968 ) ;
  assign w18970 = ( \pi01 & \pi02 ) | ( \pi01 & w18969 ) | ( \pi02 & w18969 ) ;
  assign w18971 = ( w18966 & w18968 ) | ( w18966 & ~w18970 ) | ( w18968 & ~w18970 ) ;
  assign w18972 = ~w8954 & w16818 ;
  assign w18973 = ( w16818 & w18971 ) | ( w16818 & ~w18972 ) | ( w18971 & ~w18972 ) ;
  assign w18974 = \pi02 ^ w18973 ;
  assign w18975 = w18718 ^ w18726 ;
  assign w18976 = ( w18963 & w18974 ) | ( w18963 & w18975 ) | ( w18974 & w18975 ) ;
  assign w18977 = ( ~\pi02 & w16680 ) | ( ~\pi02 & w16685 ) | ( w16680 & w16685 ) ;
  assign w18978 = \pi00 ^ w18977 ;
  assign w18979 = ( \pi02 & w16680 ) | ( \pi02 & ~w18978 ) | ( w16680 & ~w18978 ) ;
  assign w18980 = ( \pi02 & w16685 ) | ( \pi02 & w18978 ) | ( w16685 & w18978 ) ;
  assign w18981 = \pi01 & w18980 ;
  assign w18982 = ( \pi00 & w16690 ) | ( \pi00 & ~w18981 ) | ( w16690 & ~w18981 ) ;
  assign w18983 = ( \pi01 & \pi02 ) | ( \pi01 & w18982 ) | ( \pi02 & w18982 ) ;
  assign w18984 = ( w18979 & w18981 ) | ( w18979 & ~w18983 ) | ( w18981 & ~w18983 ) ;
  assign w18985 = w18727 ^ w18735 ;
  assign w18986 = w18736 ^ w18985 ;
  assign w18987 = w16772 & ~w18984 ;
  assign w18988 = ( w8954 & w18984 ) | ( w8954 & ~w18987 ) | ( w18984 & ~w18987 ) ;
  assign w18989 = \pi02 ^ w18988 ;
  assign w18990 = ( w18976 & w18986 ) | ( w18976 & w18989 ) | ( w18986 & w18989 ) ;
  assign w18991 = ( ~\pi02 & w16675 ) | ( ~\pi02 & w16680 ) | ( w16675 & w16680 ) ;
  assign w18992 = \pi00 ^ w18991 ;
  assign w18993 = ( \pi02 & w16675 ) | ( \pi02 & ~w18992 ) | ( w16675 & ~w18992 ) ;
  assign w18994 = ( \pi02 & w16680 ) | ( \pi02 & w18992 ) | ( w16680 & w18992 ) ;
  assign w18995 = \pi01 & w18994 ;
  assign w18996 = ( ~\pi00 & w16685 ) | ( ~\pi00 & w18995 ) | ( w16685 & w18995 ) ;
  assign w18997 = ( \pi01 & \pi02 ) | ( \pi01 & ~w18996 ) | ( \pi02 & ~w18996 ) ;
  assign w18998 = ( w18993 & w18995 ) | ( w18993 & ~w18997 ) | ( w18995 & ~w18997 ) ;
  assign w18999 = ~w8954 & w16946 ;
  assign w19000 = ( w16946 & w18998 ) | ( w16946 & ~w18999 ) | ( w18998 & ~w18999 ) ;
  assign w19001 = \pi02 ^ w19000 ;
  assign w19002 = w18710 ^ w18737 ;
  assign w19003 = w18702 ^ w19002 ;
  assign w19004 = ( w18990 & w19001 ) | ( w18990 & w19003 ) | ( w19001 & w19003 ) ;
  assign w19005 = ( ~\pi02 & w16670 ) | ( ~\pi02 & w16675 ) | ( w16670 & w16675 ) ;
  assign w19006 = \pi00 ^ w19005 ;
  assign w19007 = ( \pi02 & w16670 ) | ( \pi02 & ~w19006 ) | ( w16670 & ~w19006 ) ;
  assign w19008 = ( \pi02 & w16675 ) | ( \pi02 & w19006 ) | ( w16675 & w19006 ) ;
  assign w19009 = \pi01 & w19008 ;
  assign w19010 = ( ~\pi00 & w16680 ) | ( ~\pi00 & w19009 ) | ( w16680 & w19009 ) ;
  assign w19011 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19010 ) | ( \pi02 & ~w19010 ) ;
  assign w19012 = ( w19007 & w19009 ) | ( w19007 & ~w19011 ) | ( w19009 & ~w19011 ) ;
  assign w19013 = ~w8954 & w16972 ;
  assign w19014 = ( w16972 & w19012 ) | ( w16972 & ~w19013 ) | ( w19012 & ~w19013 ) ;
  assign w19015 = \pi02 ^ w19014 ;
  assign w19016 = w18696 ^ w18738 ;
  assign w19017 = w18697 ^ w19016 ;
  assign w19018 = ( w19004 & w19015 ) | ( w19004 & w19017 ) | ( w19015 & w19017 ) ;
  assign w19019 = ( ~\pi02 & w16665 ) | ( ~\pi02 & w16670 ) | ( w16665 & w16670 ) ;
  assign w19020 = \pi00 ^ w19019 ;
  assign w19021 = ( \pi02 & w16665 ) | ( \pi02 & ~w19020 ) | ( w16665 & ~w19020 ) ;
  assign w19022 = ( \pi02 & w16670 ) | ( \pi02 & w19020 ) | ( w16670 & w19020 ) ;
  assign w19023 = \pi01 & w19022 ;
  assign w19024 = ( ~\pi00 & w16675 ) | ( ~\pi00 & w19023 ) | ( w16675 & w19023 ) ;
  assign w19025 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19024 ) | ( \pi02 & ~w19024 ) ;
  assign w19026 = ( w19021 & w19023 ) | ( w19021 & ~w19025 ) | ( w19023 & ~w19025 ) ;
  assign w19027 = ~w8954 & w16960 ;
  assign w19028 = ( w16960 & w19026 ) | ( w16960 & ~w19027 ) | ( w19026 & ~w19027 ) ;
  assign w19029 = \pi02 ^ w19028 ;
  assign w19030 = w18688 ^ w18739 ;
  assign w19031 = w18680 ^ w19030 ;
  assign w19032 = ( w19018 & w19029 ) | ( w19018 & w19031 ) | ( w19029 & w19031 ) ;
  assign w19033 = ( \pi02 & w16662 ) | ( \pi02 & ~w16665 ) | ( w16662 & ~w16665 ) ;
  assign w19034 = \pi00 ^ w19033 ;
  assign w19035 = ( \pi02 & ~w16662 ) | ( \pi02 & w19034 ) | ( ~w16662 & w19034 ) ;
  assign w19036 = ( \pi02 & w16665 ) | ( \pi02 & ~w19034 ) | ( w16665 & ~w19034 ) ;
  assign w19037 = \pi01 & w19036 ;
  assign w19038 = ( ~\pi00 & w16670 ) | ( ~\pi00 & w19037 ) | ( w16670 & w19037 ) ;
  assign w19039 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19038 ) | ( \pi02 & ~w19038 ) ;
  assign w19040 = ( w19035 & w19037 ) | ( w19035 & ~w19039 ) | ( w19037 & ~w19039 ) ;
  assign w19041 = w8954 | w16762 ;
  assign w19042 = ( ~w16762 & w19040 ) | ( ~w16762 & w19041 ) | ( w19040 & w19041 ) ;
  assign w19043 = \pi02 ^ w19042 ;
  assign w19044 = w18676 ^ w18740 ;
  assign w19045 = w18678 ^ w19044 ;
  assign w19046 = ( w19032 & w19043 ) | ( w19032 & w19045 ) | ( w19043 & w19045 ) ;
  assign w19047 = ( \pi02 & ~w16660 ) | ( \pi02 & w16662 ) | ( ~w16660 & w16662 ) ;
  assign w19048 = \pi00 ^ w19047 ;
  assign w19049 = ( \pi02 & w16660 ) | ( \pi02 & w19048 ) | ( w16660 & w19048 ) ;
  assign w19050 = ( ~\pi02 & w16662 ) | ( ~\pi02 & w19048 ) | ( w16662 & w19048 ) ;
  assign w19051 = \pi01 & ~w19050 ;
  assign w19052 = ( ~\pi00 & w16665 ) | ( ~\pi00 & w19051 ) | ( w16665 & w19051 ) ;
  assign w19053 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19052 ) | ( \pi02 & ~w19052 ) ;
  assign w19054 = ( w19049 & w19051 ) | ( w19049 & ~w19053 ) | ( w19051 & ~w19053 ) ;
  assign w19055 = w8954 | w17078 ;
  assign w19056 = ( ~w17078 & w19054 ) | ( ~w17078 & w19055 ) | ( w19054 & w19055 ) ;
  assign w19057 = \pi02 ^ w19056 ;
  assign w19058 = w18668 ^ w18741 ;
  assign w19059 = w18660 ^ w19058 ;
  assign w19060 = ( w19046 & w19057 ) | ( w19046 & w19059 ) | ( w19057 & w19059 ) ;
  assign w19061 = ( \pi02 & w16658 ) | ( \pi02 & ~w16660 ) | ( w16658 & ~w16660 ) ;
  assign w19062 = \pi00 ^ w19061 ;
  assign w19063 = ( \pi02 & ~w16658 ) | ( \pi02 & w19062 ) | ( ~w16658 & w19062 ) ;
  assign w19064 = ( \pi02 & w16660 ) | ( \pi02 & ~w19062 ) | ( w16660 & ~w19062 ) ;
  assign w19065 = \pi01 & w19064 ;
  assign w19066 = ( \pi00 & w16662 ) | ( \pi00 & ~w19065 ) | ( w16662 & ~w19065 ) ;
  assign w19067 = ( \pi01 & \pi02 ) | ( \pi01 & w19066 ) | ( \pi02 & w19066 ) ;
  assign w19068 = ( w19063 & w19065 ) | ( w19063 & ~w19067 ) | ( w19065 & ~w19067 ) ;
  assign w19069 = w8954 | w17065 ;
  assign w19070 = ( ~w17065 & w19068 ) | ( ~w17065 & w19069 ) | ( w19068 & w19069 ) ;
  assign w19071 = \pi02 ^ w19070 ;
  assign w19072 = w18658 ^ w18742 ;
  assign w19073 = w18650 ^ w19072 ;
  assign w19074 = ( w19060 & w19071 ) | ( w19060 & w19073 ) | ( w19071 & w19073 ) ;
  assign w19075 = ( \pi02 & w16656 ) | ( \pi02 & w16658 ) | ( w16656 & w16658 ) ;
  assign w19076 = \pi00 ^ w19075 ;
  assign w19077 = ( \pi02 & ~w16656 ) | ( \pi02 & w19076 ) | ( ~w16656 & w19076 ) ;
  assign w19078 = ( ~\pi02 & w16658 ) | ( ~\pi02 & w19076 ) | ( w16658 & w19076 ) ;
  assign w19079 = \pi01 & ~w19078 ;
  assign w19080 = ( ~\pi00 & w16660 ) | ( ~\pi00 & w19079 ) | ( w16660 & w19079 ) ;
  assign w19081 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19080 ) | ( \pi02 & ~w19080 ) ;
  assign w19082 = ( w19077 & w19079 ) | ( w19077 & ~w19081 ) | ( w19079 & ~w19081 ) ;
  assign w19083 = ~w8954 & w17057 ;
  assign w19084 = ( w17057 & w19082 ) | ( w17057 & ~w19083 ) | ( w19082 & ~w19083 ) ;
  assign w19085 = \pi02 ^ w19084 ;
  assign w19086 = w18648 ^ w18743 ;
  assign w19087 = w18640 ^ w19086 ;
  assign w19088 = ( w19074 & w19085 ) | ( w19074 & w19087 ) | ( w19085 & w19087 ) ;
  assign w19089 = ( \pi02 & ~w16654 ) | ( \pi02 & w16656 ) | ( ~w16654 & w16656 ) ;
  assign w19090 = \pi00 ^ w19089 ;
  assign w19091 = ( \pi02 & w16654 ) | ( \pi02 & w19090 ) | ( w16654 & w19090 ) ;
  assign w19092 = ( ~\pi02 & w16656 ) | ( ~\pi02 & w19090 ) | ( w16656 & w19090 ) ;
  assign w19093 = \pi01 & ~w19092 ;
  assign w19094 = ( \pi00 & w16658 ) | ( \pi00 & ~w19093 ) | ( w16658 & ~w19093 ) ;
  assign w19095 = ( \pi01 & \pi02 ) | ( \pi01 & w19094 ) | ( \pi02 & w19094 ) ;
  assign w19096 = ( w19091 & w19093 ) | ( w19091 & ~w19095 ) | ( w19093 & ~w19095 ) ;
  assign w19097 = ~w8954 & w17266 ;
  assign w19098 = ( w17266 & w19096 ) | ( w17266 & ~w19097 ) | ( w19096 & ~w19097 ) ;
  assign w19099 = \pi02 ^ w19098 ;
  assign w19100 = w18636 ^ w18744 ;
  assign w19101 = w18638 ^ w19100 ;
  assign w19102 = ( w19088 & w19099 ) | ( w19088 & w19101 ) | ( w19099 & w19101 ) ;
  assign w19103 = ( \pi02 & w16652 ) | ( \pi02 & ~w16654 ) | ( w16652 & ~w16654 ) ;
  assign w19104 = \pi00 ^ w19103 ;
  assign w19105 = ( \pi02 & ~w16652 ) | ( \pi02 & w19104 ) | ( ~w16652 & w19104 ) ;
  assign w19106 = ( \pi02 & w16654 ) | ( \pi02 & ~w19104 ) | ( w16654 & ~w19104 ) ;
  assign w19107 = \pi01 & w19106 ;
  assign w19108 = ( \pi00 & w16656 ) | ( \pi00 & ~w19107 ) | ( w16656 & ~w19107 ) ;
  assign w19109 = ( \pi01 & \pi02 ) | ( \pi01 & w19108 ) | ( \pi02 & w19108 ) ;
  assign w19110 = ( w19105 & w19107 ) | ( w19105 & ~w19109 ) | ( w19107 & ~w19109 ) ;
  assign w19111 = ~w8954 & w17293 ;
  assign w19112 = ( w17293 & w19110 ) | ( w17293 & ~w19111 ) | ( w19110 & ~w19111 ) ;
  assign w19113 = \pi02 ^ w19112 ;
  assign w19114 = w18626 ^ w18745 ;
  assign w19115 = w18628 ^ w19114 ;
  assign w19116 = ( w19102 & w19113 ) | ( w19102 & w19115 ) | ( w19113 & w19115 ) ;
  assign w19117 = ( \pi02 & w16650 ) | ( \pi02 & w16652 ) | ( w16650 & w16652 ) ;
  assign w19118 = \pi00 ^ w19117 ;
  assign w19119 = ( \pi02 & ~w16650 ) | ( \pi02 & w19118 ) | ( ~w16650 & w19118 ) ;
  assign w19120 = ( ~\pi02 & w16652 ) | ( ~\pi02 & w19118 ) | ( w16652 & w19118 ) ;
  assign w19121 = \pi01 & ~w19120 ;
  assign w19122 = ( ~\pi00 & w16654 ) | ( ~\pi00 & w19121 ) | ( w16654 & w19121 ) ;
  assign w19123 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19122 ) | ( \pi02 & ~w19122 ) ;
  assign w19124 = ( w19119 & w19121 ) | ( w19119 & ~w19123 ) | ( w19121 & ~w19123 ) ;
  assign w19125 = w8954 | w17277 ;
  assign w19126 = ( ~w17277 & w19124 ) | ( ~w17277 & w19125 ) | ( w19124 & w19125 ) ;
  assign w19127 = \pi02 ^ w19126 ;
  assign w19128 = w18616 ^ w18746 ;
  assign w19129 = w18618 ^ w19128 ;
  assign w19130 = ( w19116 & w19127 ) | ( w19116 & w19129 ) | ( w19127 & w19129 ) ;
  assign w19131 = ( \pi02 & w16648 ) | ( \pi02 & w16650 ) | ( w16648 & w16650 ) ;
  assign w19132 = \pi00 ^ w19131 ;
  assign w19133 = ( \pi02 & ~w16648 ) | ( \pi02 & w19132 ) | ( ~w16648 & w19132 ) ;
  assign w19134 = ( ~\pi02 & w16650 ) | ( ~\pi02 & w19132 ) | ( w16650 & w19132 ) ;
  assign w19135 = \pi01 & ~w19134 ;
  assign w19136 = ( \pi00 & w16652 ) | ( \pi00 & ~w19135 ) | ( w16652 & ~w19135 ) ;
  assign w19137 = ( \pi01 & \pi02 ) | ( \pi01 & w19136 ) | ( \pi02 & w19136 ) ;
  assign w19138 = ( w19133 & w19135 ) | ( w19133 & ~w19137 ) | ( w19135 & ~w19137 ) ;
  assign w19139 = w8954 | w16752 ;
  assign w19140 = ( ~w16752 & w19138 ) | ( ~w16752 & w19139 ) | ( w19138 & w19139 ) ;
  assign w19141 = \pi02 ^ w19140 ;
  assign w19142 = w18608 ^ w18747 ;
  assign w19143 = w18600 ^ w19142 ;
  assign w19144 = ( w19130 & w19141 ) | ( w19130 & w19143 ) | ( w19141 & w19143 ) ;
  assign w19145 = ( \pi02 & w16646 ) | ( \pi02 & w16648 ) | ( w16646 & w16648 ) ;
  assign w19146 = \pi00 ^ w19145 ;
  assign w19147 = ( \pi02 & ~w16646 ) | ( \pi02 & w19146 ) | ( ~w16646 & w19146 ) ;
  assign w19148 = ( ~\pi02 & w16648 ) | ( ~\pi02 & w19146 ) | ( w16648 & w19146 ) ;
  assign w19149 = \pi01 & ~w19148 ;
  assign w19150 = ( \pi00 & w16650 ) | ( \pi00 & ~w19149 ) | ( w16650 & ~w19149 ) ;
  assign w19151 = ( \pi01 & \pi02 ) | ( \pi01 & w19150 ) | ( \pi02 & w19150 ) ;
  assign w19152 = ( w19147 & w19149 ) | ( w19147 & ~w19151 ) | ( w19149 & ~w19151 ) ;
  assign w19153 = w8954 | w17476 ;
  assign w19154 = ( ~w17476 & w19152 ) | ( ~w17476 & w19153 ) | ( w19152 & w19153 ) ;
  assign w19155 = \pi02 ^ w19154 ;
  assign w19156 = w18598 ^ w18748 ;
  assign w19157 = w18590 ^ w19156 ;
  assign w19158 = ( w19144 & w19155 ) | ( w19144 & w19157 ) | ( w19155 & w19157 ) ;
  assign w19159 = ( \pi02 & w16644 ) | ( \pi02 & w16646 ) | ( w16644 & w16646 ) ;
  assign w19160 = \pi00 ^ w19159 ;
  assign w19161 = ( \pi02 & ~w16644 ) | ( \pi02 & w19160 ) | ( ~w16644 & w19160 ) ;
  assign w19162 = ( ~\pi02 & w16646 ) | ( ~\pi02 & w19160 ) | ( w16646 & w19160 ) ;
  assign w19163 = \pi01 & ~w19162 ;
  assign w19164 = ( \pi00 & w16648 ) | ( \pi00 & ~w19163 ) | ( w16648 & ~w19163 ) ;
  assign w19165 = ( \pi01 & \pi02 ) | ( \pi01 & w19164 ) | ( \pi02 & w19164 ) ;
  assign w19166 = ( w19161 & w19163 ) | ( w19161 & ~w19165 ) | ( w19163 & ~w19165 ) ;
  assign w19167 = w8954 | w17468 ;
  assign w19168 = ( ~w17468 & w19166 ) | ( ~w17468 & w19167 ) | ( w19166 & w19167 ) ;
  assign w19169 = \pi02 ^ w19168 ;
  assign w19170 = w18588 ^ w18749 ;
  assign w19171 = w18580 ^ w19170 ;
  assign w19172 = ( w19158 & w19169 ) | ( w19158 & w19171 ) | ( w19169 & w19171 ) ;
  assign w19173 = ( \pi02 & ~w16642 ) | ( \pi02 & w16644 ) | ( ~w16642 & w16644 ) ;
  assign w19174 = \pi00 ^ w19173 ;
  assign w19175 = ( \pi02 & w16642 ) | ( \pi02 & w19174 ) | ( w16642 & w19174 ) ;
  assign w19176 = ( ~\pi02 & w16644 ) | ( ~\pi02 & w19174 ) | ( w16644 & w19174 ) ;
  assign w19177 = \pi01 & ~w19176 ;
  assign w19178 = ( \pi00 & w16646 ) | ( \pi00 & ~w19177 ) | ( w16646 & ~w19177 ) ;
  assign w19179 = ( \pi01 & \pi02 ) | ( \pi01 & w19178 ) | ( \pi02 & w19178 ) ;
  assign w19180 = ( w19175 & w19177 ) | ( w19175 & ~w19179 ) | ( w19177 & ~w19179 ) ;
  assign w19181 = ~w8954 & w17455 ;
  assign w19182 = ( w17455 & w19180 ) | ( w17455 & ~w19181 ) | ( w19180 & ~w19181 ) ;
  assign w19183 = \pi02 ^ w19182 ;
  assign w19184 = w18576 ^ w18750 ;
  assign w19185 = w18578 ^ w19184 ;
  assign w19186 = ( w19172 & w19183 ) | ( w19172 & w19185 ) | ( w19183 & w19185 ) ;
  assign w19187 = ( ~\pi02 & w16640 ) | ( ~\pi02 & w16642 ) | ( w16640 & w16642 ) ;
  assign w19188 = \pi00 ^ w19187 ;
  assign w19189 = ( \pi02 & w16640 ) | ( \pi02 & ~w19188 ) | ( w16640 & ~w19188 ) ;
  assign w19190 = ( \pi02 & w16642 ) | ( \pi02 & w19188 ) | ( w16642 & w19188 ) ;
  assign w19191 = \pi01 & w19190 ;
  assign w19192 = ( \pi00 & w16644 ) | ( \pi00 & ~w19191 ) | ( w16644 & ~w19191 ) ;
  assign w19193 = ( \pi01 & \pi02 ) | ( \pi01 & w19192 ) | ( \pi02 & w19192 ) ;
  assign w19194 = ( w19189 & w19191 ) | ( w19189 & ~w19193 ) | ( w19191 & ~w19193 ) ;
  assign w19195 = w8954 | w17760 ;
  assign w19196 = ( ~w17760 & w19194 ) | ( ~w17760 & w19195 ) | ( w19194 & w19195 ) ;
  assign w19197 = \pi02 ^ w19196 ;
  assign w19198 = w18566 ^ w18751 ;
  assign w19199 = w18568 ^ w19198 ;
  assign w19200 = ( w19186 & w19197 ) | ( w19186 & w19199 ) | ( w19197 & w19199 ) ;
  assign w19201 = ( \pi02 & w16638 ) | ( \pi02 & ~w16640 ) | ( w16638 & ~w16640 ) ;
  assign w19202 = \pi00 ^ w19201 ;
  assign w19203 = ( \pi02 & ~w16638 ) | ( \pi02 & w19202 ) | ( ~w16638 & w19202 ) ;
  assign w19204 = ( \pi02 & w16640 ) | ( \pi02 & ~w19202 ) | ( w16640 & ~w19202 ) ;
  assign w19205 = \pi01 & w19204 ;
  assign w19206 = ( ~\pi00 & w16642 ) | ( ~\pi00 & w19205 ) | ( w16642 & w19205 ) ;
  assign w19207 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19206 ) | ( \pi02 & ~w19206 ) ;
  assign w19208 = ( w19203 & w19205 ) | ( w19203 & ~w19207 ) | ( w19205 & ~w19207 ) ;
  assign w19209 = w8954 | w17783 ;
  assign w19210 = ( ~w17783 & w19208 ) | ( ~w17783 & w19209 ) | ( w19208 & w19209 ) ;
  assign w19211 = \pi02 ^ w19210 ;
  assign w19212 = w18556 ^ w18752 ;
  assign w19213 = w18558 ^ w19212 ;
  assign w19214 = ( w19200 & w19211 ) | ( w19200 & w19213 ) | ( w19211 & w19213 ) ;
  assign w19215 = ( \pi02 & ~w16636 ) | ( \pi02 & w16638 ) | ( ~w16636 & w16638 ) ;
  assign w19216 = \pi00 ^ w19215 ;
  assign w19217 = ( \pi02 & w16636 ) | ( \pi02 & w19216 ) | ( w16636 & w19216 ) ;
  assign w19218 = ( ~\pi02 & w16638 ) | ( ~\pi02 & w19216 ) | ( w16638 & w19216 ) ;
  assign w19219 = \pi01 & ~w19218 ;
  assign w19220 = ( ~\pi00 & w16640 ) | ( ~\pi00 & w19219 ) | ( w16640 & w19219 ) ;
  assign w19221 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19220 ) | ( \pi02 & ~w19220 ) ;
  assign w19222 = ( w19217 & w19219 ) | ( w19217 & ~w19221 ) | ( w19219 & ~w19221 ) ;
  assign w19223 = w8954 | w17770 ;
  assign w19224 = ( ~w17770 & w19222 ) | ( ~w17770 & w19223 ) | ( w19222 & w19223 ) ;
  assign w19225 = \pi02 ^ w19224 ;
  assign w19226 = w18548 ^ w18753 ;
  assign w19227 = w18540 ^ w19226 ;
  assign w19228 = ( w19214 & w19225 ) | ( w19214 & w19227 ) | ( w19225 & w19227 ) ;
  assign w19229 = ( \pi02 & w16634 ) | ( \pi02 & ~w16636 ) | ( w16634 & ~w16636 ) ;
  assign w19230 = \pi00 ^ w19229 ;
  assign w19231 = ( \pi02 & ~w16634 ) | ( \pi02 & w19230 ) | ( ~w16634 & w19230 ) ;
  assign w19232 = ( \pi02 & w16636 ) | ( \pi02 & ~w19230 ) | ( w16636 & ~w19230 ) ;
  assign w19233 = \pi01 & w19232 ;
  assign w19234 = ( \pi00 & w16638 ) | ( \pi00 & ~w19233 ) | ( w16638 & ~w19233 ) ;
  assign w19235 = ( \pi01 & \pi02 ) | ( \pi01 & w19234 ) | ( \pi02 & w19234 ) ;
  assign w19236 = ( w19231 & w19233 ) | ( w19231 & ~w19235 ) | ( w19233 & ~w19235 ) ;
  assign w19237 = w8954 | w16742 ;
  assign w19238 = ( ~w16742 & w19236 ) | ( ~w16742 & w19237 ) | ( w19236 & w19237 ) ;
  assign w19239 = \pi02 ^ w19238 ;
  assign w19240 = w18538 ^ w18754 ;
  assign w19241 = w18530 ^ w19240 ;
  assign w19242 = ( w19228 & w19239 ) | ( w19228 & w19241 ) | ( w19239 & w19241 ) ;
  assign w19243 = ( \pi02 & ~w16632 ) | ( \pi02 & w16634 ) | ( ~w16632 & w16634 ) ;
  assign w19244 = \pi00 ^ w19243 ;
  assign w19245 = ( \pi02 & w16632 ) | ( \pi02 & w19244 ) | ( w16632 & w19244 ) ;
  assign w19246 = ( ~\pi02 & w16634 ) | ( ~\pi02 & w19244 ) | ( w16634 & w19244 ) ;
  assign w19247 = \pi01 & ~w19246 ;
  assign w19248 = ( ~\pi00 & w16636 ) | ( ~\pi00 & w19247 ) | ( w16636 & w19247 ) ;
  assign w19249 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19248 ) | ( \pi02 & ~w19248 ) ;
  assign w19250 = ( w19245 & w19247 ) | ( w19245 & ~w19249 ) | ( w19247 & ~w19249 ) ;
  assign w19251 = w8954 | w18051 ;
  assign w19252 = ( ~w18051 & w19250 ) | ( ~w18051 & w19251 ) | ( w19250 & w19251 ) ;
  assign w19253 = \pi02 ^ w19252 ;
  assign w19254 = w18528 ^ w18755 ;
  assign w19255 = w18520 ^ w19254 ;
  assign w19256 = ( w19242 & w19253 ) | ( w19242 & w19255 ) | ( w19253 & w19255 ) ;
  assign w19257 = ( \pi02 & w16630 ) | ( \pi02 & ~w16632 ) | ( w16630 & ~w16632 ) ;
  assign w19258 = \pi00 ^ w19257 ;
  assign w19259 = ( \pi02 & ~w16630 ) | ( \pi02 & w19258 ) | ( ~w16630 & w19258 ) ;
  assign w19260 = ( \pi02 & w16632 ) | ( \pi02 & ~w19258 ) | ( w16632 & ~w19258 ) ;
  assign w19261 = \pi01 & w19260 ;
  assign w19262 = ( \pi00 & w16634 ) | ( \pi00 & ~w19261 ) | ( w16634 & ~w19261 ) ;
  assign w19263 = ( \pi01 & \pi02 ) | ( \pi01 & w19262 ) | ( \pi02 & w19262 ) ;
  assign w19264 = ( w19259 & w19261 ) | ( w19259 & ~w19263 ) | ( w19261 & ~w19263 ) ;
  assign w19265 = w8954 | w18038 ;
  assign w19266 = ( ~w18038 & w19264 ) | ( ~w18038 & w19265 ) | ( w19264 & w19265 ) ;
  assign w19267 = \pi02 ^ w19266 ;
  assign w19268 = w18516 ^ w18756 ;
  assign w19269 = w18518 ^ w19268 ;
  assign w19270 = ( w19256 & w19267 ) | ( w19256 & w19269 ) | ( w19267 & w19269 ) ;
  assign w19271 = ( \pi02 & w16628 ) | ( \pi02 & w16630 ) | ( w16628 & w16630 ) ;
  assign w19272 = \pi00 ^ w19271 ;
  assign w19273 = ( \pi02 & ~w16628 ) | ( \pi02 & w19272 ) | ( ~w16628 & w19272 ) ;
  assign w19274 = ( ~\pi02 & w16630 ) | ( ~\pi02 & w19272 ) | ( w16630 & w19272 ) ;
  assign w19275 = \pi01 & ~w19274 ;
  assign w19276 = ( ~\pi00 & w16632 ) | ( ~\pi00 & w19275 ) | ( w16632 & w19275 ) ;
  assign w19277 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19276 ) | ( \pi02 & ~w19276 ) ;
  assign w19278 = ( w19273 & w19275 ) | ( w19273 & ~w19277 ) | ( w19275 & ~w19277 ) ;
  assign w19279 = ~w8954 & w18026 ;
  assign w19280 = ( w18026 & w19278 ) | ( w18026 & ~w19279 ) | ( w19278 & ~w19279 ) ;
  assign w19281 = \pi02 ^ w19280 ;
  assign w19282 = w18506 ^ w18757 ;
  assign w19283 = w18508 ^ w19282 ;
  assign w19284 = ( w19270 & w19281 ) | ( w19270 & w19283 ) | ( w19281 & w19283 ) ;
  assign w19285 = ( \pi02 & w16626 ) | ( \pi02 & w16628 ) | ( w16626 & w16628 ) ;
  assign w19286 = \pi00 ^ w19285 ;
  assign w19287 = ( \pi02 & ~w16626 ) | ( \pi02 & w19286 ) | ( ~w16626 & w19286 ) ;
  assign w19288 = ( ~\pi02 & w16628 ) | ( ~\pi02 & w19286 ) | ( w16628 & w19286 ) ;
  assign w19289 = \pi01 & ~w19288 ;
  assign w19290 = ( \pi00 & w16630 ) | ( \pi00 & ~w19289 ) | ( w16630 & ~w19289 ) ;
  assign w19291 = ( \pi01 & \pi02 ) | ( \pi01 & w19290 ) | ( \pi02 & w19290 ) ;
  assign w19292 = ( w19287 & w19289 ) | ( w19287 & ~w19291 ) | ( w19289 & ~w19291 ) ;
  assign w19293 = w8954 | w18429 ;
  assign w19294 = ( ~w18429 & w19292 ) | ( ~w18429 & w19293 ) | ( w19292 & w19293 ) ;
  assign w19295 = \pi02 ^ w19294 ;
  assign w19296 = w18496 ^ w18758 ;
  assign w19297 = w18498 ^ w19296 ;
  assign w19298 = ( w19284 & w19295 ) | ( w19284 & w19297 ) | ( w19295 & w19297 ) ;
  assign w19299 = ( \pi02 & ~w16619 ) | ( \pi02 & w16626 ) | ( ~w16619 & w16626 ) ;
  assign w19300 = \pi00 ^ w19299 ;
  assign w19301 = ( \pi02 & w16619 ) | ( \pi02 & w19300 ) | ( w16619 & w19300 ) ;
  assign w19302 = ( ~\pi02 & w16626 ) | ( ~\pi02 & w19300 ) | ( w16626 & w19300 ) ;
  assign w19303 = \pi01 & ~w19302 ;
  assign w19304 = ( \pi00 & w16628 ) | ( \pi00 & ~w19303 ) | ( w16628 & ~w19303 ) ;
  assign w19305 = ( \pi01 & \pi02 ) | ( \pi01 & w19304 ) | ( \pi02 & w19304 ) ;
  assign w19306 = ( w19301 & w19303 ) | ( w19301 & ~w19305 ) | ( w19303 & ~w19305 ) ;
  assign w19307 = ~w8954 & w18451 ;
  assign w19308 = ( w18451 & w19306 ) | ( w18451 & ~w19307 ) | ( w19306 & ~w19307 ) ;
  assign w19309 = \pi02 ^ w19308 ;
  assign w19310 = w18488 ^ w18759 ;
  assign w19311 = w18480 ^ w19310 ;
  assign w19312 = ( w19298 & w19309 ) | ( w19298 & w19311 ) | ( w19309 & w19311 ) ;
  assign w19313 = ( ~\pi02 & w16619 ) | ( ~\pi02 & w16621 ) | ( w16619 & w16621 ) ;
  assign w19314 = \pi00 ^ w19313 ;
  assign w19315 = ( \pi02 & w16621 ) | ( \pi02 & ~w19314 ) | ( w16621 & ~w19314 ) ;
  assign w19316 = ( \pi02 & w16619 ) | ( \pi02 & w19314 ) | ( w16619 & w19314 ) ;
  assign w19317 = \pi01 & w19316 ;
  assign w19318 = ( \pi00 & w16626 ) | ( \pi00 & ~w19317 ) | ( w16626 & ~w19317 ) ;
  assign w19319 = ( \pi01 & \pi02 ) | ( \pi01 & w19318 ) | ( \pi02 & w19318 ) ;
  assign w19320 = ( w19315 & w19317 ) | ( w19315 & ~w19319 ) | ( w19317 & ~w19319 ) ;
  assign w19321 = w8954 | w18439 ;
  assign w19322 = ( ~w18439 & w19320 ) | ( ~w18439 & w19321 ) | ( w19320 & w19321 ) ;
  assign w19323 = \pi02 ^ w19322 ;
  assign w19324 = w18478 ^ w18760 ;
  assign w19325 = w18470 ^ w19324 ;
  assign w19326 = ( w19312 & w19323 ) | ( w19312 & w19325 ) | ( w19323 & w19325 ) ;
  assign w19327 = ( ~\pi02 & w16617 ) | ( ~\pi02 & w16621 ) | ( w16617 & w16621 ) ;
  assign w19328 = \pi00 ^ w19327 ;
  assign w19329 = ( \pi02 & w16617 ) | ( \pi02 & ~w19328 ) | ( w16617 & ~w19328 ) ;
  assign w19330 = ( \pi02 & w16621 ) | ( \pi02 & w19328 ) | ( w16621 & w19328 ) ;
  assign w19331 = \pi01 & w19330 ;
  assign w19332 = ( ~\pi00 & w16619 ) | ( ~\pi00 & w19331 ) | ( w16619 & w19331 ) ;
  assign w19333 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19332 ) | ( \pi02 & ~w19332 ) ;
  assign w19334 = ( w19329 & w19331 ) | ( w19329 & ~w19333 ) | ( w19331 & ~w19333 ) ;
  assign w19335 = ~w8954 & w16732 ;
  assign w19336 = ( w16732 & w19334 ) | ( w16732 & ~w19335 ) | ( w19334 & ~w19335 ) ;
  assign w19337 = \pi02 ^ w19336 ;
  assign w19338 = w18466 ^ w18761 ;
  assign w19339 = w18468 ^ w19338 ;
  assign w19340 = ( w19326 & w19337 ) | ( w19326 & ~w19339 ) | ( w19337 & ~w19339 ) ;
  assign w19341 = ( \pi02 & ~w16617 ) | ( \pi02 & w18914 ) | ( ~w16617 & w18914 ) ;
  assign w19342 = \pi00 ^ w19341 ;
  assign w19343 = ( \pi02 & ~w18914 ) | ( \pi02 & w19342 ) | ( ~w18914 & w19342 ) ;
  assign w19344 = ( \pi02 & w16617 ) | ( \pi02 & ~w19342 ) | ( w16617 & ~w19342 ) ;
  assign w19345 = \pi01 & w19344 ;
  assign w19346 = ( ~\pi00 & w16621 ) | ( ~\pi00 & w19345 ) | ( w16621 & w19345 ) ;
  assign w19347 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19346 ) | ( \pi02 & ~w19346 ) ;
  assign w19348 = ( w19343 & w19345 ) | ( w19343 & ~w19347 ) | ( w19345 & ~w19347 ) ;
  assign w19349 = w16729 ^ w18914 ;
  assign w19350 = w16617 ^ w19349 ;
  assign w19351 = w8954 & w19350 ;
  assign w19352 = ( w8954 & w19348 ) | ( w8954 & ~w19351 ) | ( w19348 & ~w19351 ) ;
  assign w19353 = \pi02 ^ w19352 ;
  assign w19354 = w18456 ^ w18762 ;
  assign w19355 = w18458 ^ w19354 ;
  assign w19356 = ( w19340 & w19353 ) | ( w19340 & ~w19355 ) | ( w19353 & ~w19355 ) ;
  assign w19357 = ( \pi02 & w18914 ) | ( \pi02 & ~w18916 ) | ( w18914 & ~w18916 ) ;
  assign w19358 = \pi00 ^ w19357 ;
  assign w19359 = ( \pi02 & w18916 ) | ( \pi02 & w19358 ) | ( w18916 & w19358 ) ;
  assign w19360 = ( ~\pi02 & w18914 ) | ( ~\pi02 & w19358 ) | ( w18914 & w19358 ) ;
  assign w19361 = \pi01 & ~w19360 ;
  assign w19362 = ( ~\pi00 & w16617 ) | ( ~\pi00 & w19361 ) | ( w16617 & w19361 ) ;
  assign w19363 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19362 ) | ( \pi02 & ~w19362 ) ;
  assign w19364 = ( w19359 & w19361 ) | ( w19359 & ~w19363 ) | ( w19361 & ~w19363 ) ;
  assign w19365 = w18916 ^ w18925 ;
  assign w19366 = w18914 ^ w19365 ;
  assign w19367 = w8954 & w19366 ;
  assign w19368 = ( w8954 & w19364 ) | ( w8954 & ~w19367 ) | ( w19364 & ~w19367 ) ;
  assign w19369 = \pi02 ^ w19368 ;
  assign w19370 = w18444 ^ w18763 ;
  assign w19371 = w18446 ^ w19370 ;
  assign w19372 = ( w19356 & w19369 ) | ( w19356 & w19371 ) | ( w19369 & w19371 ) ;
  assign w19373 = ( ~w18766 & w18932 ) | ( ~w18766 & w19372 ) | ( w18932 & w19372 ) ;
  assign w19374 = ~w8593 & w16617 ;
  assign w19375 = w8262 & w16621 ;
  assign w19376 = ( w16617 & ~w19374 ) | ( w16617 & w19375 ) | ( ~w19374 & w19375 ) ;
  assign w19377 = w8263 | w19350 ;
  assign w19378 = w18914 & ~w19376 ;
  assign w19379 = ( w35 & w19376 ) | ( w35 & ~w19378 ) | ( w19376 & ~w19378 ) ;
  assign w19380 = ( ~w19350 & w19377 ) | ( ~w19350 & w19379 ) | ( w19377 & w19379 ) ;
  assign w19381 = \pi05 ^ w19380 ;
  assign w19382 = ( w18315 & ~w18421 ) | ( w18315 & w18432 ) | ( ~w18421 & w18432 ) ;
  assign w19383 = ~w6949 & w16632 ;
  assign w19384 = w6748 & ~w16634 ;
  assign w19385 = ( w16632 & ~w19383 ) | ( w16632 & w19384 ) | ( ~w19383 & w19384 ) ;
  assign w19386 = w7154 | w16630 ;
  assign w19387 = w18038 & ~w19385 ;
  assign w19388 = ( w6751 & w19385 ) | ( w6751 & ~w19387 ) | ( w19385 & ~w19387 ) ;
  assign w19389 = ( ~w16630 & w19386 ) | ( ~w16630 & w19388 ) | ( w19386 & w19388 ) ;
  assign w19390 = \pi11 ^ w19389 ;
  assign w19391 = ( w18324 & ~w18408 ) | ( w18324 & w18416 ) | ( ~w18408 & w18416 ) ;
  assign w19392 = w5710 | w16644 ;
  assign w19393 = w5494 & ~w16646 ;
  assign w19394 = ( ~w16644 & w19392 ) | ( ~w16644 & w19393 ) | ( w19392 & w19393 ) ;
  assign w19395 = ~w5948 & w16642 ;
  assign w19396 = w17455 | w19394 ;
  assign w19397 = ( w5497 & w19394 ) | ( w5497 & w19396 ) | ( w19394 & w19396 ) ;
  assign w19398 = ( w16642 & ~w19395 ) | ( w16642 & w19397 ) | ( ~w19395 & w19397 ) ;
  assign w19399 = \pi17 ^ w19398 ;
  assign w19400 = ( w18333 & ~w18395 ) | ( w18333 & w18403 ) | ( ~w18395 & w18403 ) ;
  assign w19401 = w4651 | w16656 ;
  assign w19402 = w4606 & ~w16658 ;
  assign w19403 = ( ~w16656 & w19401 ) | ( ~w16656 & w19402 ) | ( w19401 & w19402 ) ;
  assign w19404 = ~w4706 & w16654 ;
  assign w19405 = w17266 | w19403 ;
  assign w19406 = ( w4609 & w19403 ) | ( w4609 & w19405 ) | ( w19403 & w19405 ) ;
  assign w19407 = ( w16654 & ~w19404 ) | ( w16654 & w19406 ) | ( ~w19404 & w19406 ) ;
  assign w19408 = \pi23 ^ w19407 ;
  assign w19409 = ( w18342 & ~w18382 ) | ( w18342 & w18390 ) | ( ~w18382 & w18390 ) ;
  assign w19410 = ~w3717 & w16675 ;
  assign w19411 = w3649 & w16680 ;
  assign w19412 = ( w16675 & ~w19410 ) | ( w16675 & w19411 ) | ( ~w19410 & w19411 ) ;
  assign w19413 = ~w3549 & w16670 ;
  assign w19414 = w16972 | w19412 ;
  assign w19415 = ( w3448 & w19412 ) | ( w3448 & w19414 ) | ( w19412 & w19414 ) ;
  assign w19416 = ( w16670 & ~w19413 ) | ( w16670 & w19415 ) | ( ~w19413 & w19415 ) ;
  assign w19417 = \pi29 ^ w19416 ;
  assign w19418 = ( w18351 & ~w18369 ) | ( w18351 & w18377 ) | ( ~w18369 & w18377 ) ;
  assign w19419 = ( ~w390 & w800 ) | ( ~w390 & w1948 ) | ( w800 & w1948 ) ;
  assign w19420 = w4764 | w11021 ;
  assign w19421 = ( w390 & w1229 ) | ( w390 & ~w4764 ) | ( w1229 & ~w4764 ) ;
  assign w19422 = w19420 | w19421 ;
  assign w19423 = w19419 | w19422 ;
  assign w19424 = ~w222 & w10912 ;
  assign w19425 = ~w4400 & w19424 ;
  assign w19426 = ( w3244 & ~w4400 ) | ( w3244 & w19423 ) | ( ~w4400 & w19423 ) ;
  assign w19427 = w19425 & ~w19426 ;
  assign w19428 = w1126 | w1265 ;
  assign w19429 = w82 | w19428 ;
  assign w19430 = ( w82 & ~w952 ) | ( w82 & w19427 ) | ( ~w952 & w19427 ) ;
  assign w19431 = ~w19429 & w19430 ;
  assign w19432 = w415 | w492 ;
  assign w19433 = ( w415 & ~w422 ) | ( w415 & w19431 ) | ( ~w422 & w19431 ) ;
  assign w19434 = ~w19432 & w19433 ;
  assign w19435 = ~w37 & w16818 ;
  assign w19436 = w3098 & ~w16692 ;
  assign w19437 = ( w16818 & ~w19435 ) | ( w16818 & w19436 ) | ( ~w19435 & w19436 ) ;
  assign w19438 = ( \pi29 & \pi30 ) | ( \pi29 & w16685 ) | ( \pi30 & w16685 ) ;
  assign w19439 = \pi31 | w19438 ;
  assign w19440 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w16690 ) | ( \pi30 & w16690 ) ;
  assign w19441 = ( \pi29 & \pi31 ) | ( \pi29 & w19440 ) | ( \pi31 & w19440 ) ;
  assign w19442 = ( w19437 & w19439 ) | ( w19437 & ~w19441 ) | ( w19439 & ~w19441 ) ;
  assign w19443 = w19418 ^ w19442 ;
  assign w19444 = w19434 ^ w19443 ;
  assign w19445 = ( w18350 & ~w18379 ) | ( w18350 & w18380 ) | ( ~w18379 & w18380 ) ;
  assign w19446 = w19417 ^ w19445 ;
  assign w19447 = w19444 ^ w19446 ;
  assign w19448 = w3964 & w16660 ;
  assign w19449 = ( w4143 & ~w16662 ) | ( w4143 & w19448 ) | ( ~w16662 & w19448 ) ;
  assign w19450 = w4052 | w19449 ;
  assign w19451 = ( w16665 & w19449 ) | ( w16665 & w19450 ) | ( w19449 & w19450 ) ;
  assign w19452 = w19448 | w19451 ;
  assign w19453 = w4147 | w17078 ;
  assign w19454 = ( ~w17078 & w19452 ) | ( ~w17078 & w19453 ) | ( w19452 & w19453 ) ;
  assign w19455 = \pi26 ^ w19454 ;
  assign w19456 = w19409 ^ w19455 ;
  assign w19457 = w19447 ^ w19456 ;
  assign w19458 = ( w18341 & ~w18392 ) | ( w18341 & w18393 ) | ( ~w18392 & w18393 ) ;
  assign w19459 = w19408 ^ w19458 ;
  assign w19460 = w19457 ^ w19459 ;
  assign w19461 = w4905 & ~w16652 ;
  assign w19462 = ( w5395 & ~w16648 ) | ( w5395 & w19461 ) | ( ~w16648 & w19461 ) ;
  assign w19463 = w5343 | w19462 ;
  assign w19464 = ( ~w16650 & w19462 ) | ( ~w16650 & w19463 ) | ( w19462 & w19463 ) ;
  assign w19465 = w19461 | w19464 ;
  assign w19466 = w4908 | w16752 ;
  assign w19467 = ( ~w16752 & w19465 ) | ( ~w16752 & w19466 ) | ( w19465 & w19466 ) ;
  assign w19468 = \pi20 ^ w19467 ;
  assign w19469 = w19400 ^ w19468 ;
  assign w19470 = w19460 ^ w19469 ;
  assign w19471 = ( w18332 & ~w18405 ) | ( w18332 & w18406 ) | ( ~w18405 & w18406 ) ;
  assign w19472 = w19399 ^ w19471 ;
  assign w19473 = w19470 ^ w19472 ;
  assign w19474 = w6048 & w16640 ;
  assign w19475 = ( w6637 & w16636 ) | ( w6637 & w19474 ) | ( w16636 & w19474 ) ;
  assign w19476 = w6549 | w19475 ;
  assign w19477 = ( ~w16638 & w19475 ) | ( ~w16638 & w19476 ) | ( w19475 & w19476 ) ;
  assign w19478 = w19474 | w19477 ;
  assign w19479 = w6045 | w17770 ;
  assign w19480 = ( ~w17770 & w19478 ) | ( ~w17770 & w19479 ) | ( w19478 & w19479 ) ;
  assign w19481 = \pi14 ^ w19480 ;
  assign w19482 = w19391 ^ w19481 ;
  assign w19483 = w19473 ^ w19482 ;
  assign w19484 = ( w18323 & ~w18418 ) | ( w18323 & w18419 ) | ( ~w18418 & w18419 ) ;
  assign w19485 = w19390 ^ w19484 ;
  assign w19486 = w19483 ^ w19485 ;
  assign w19487 = w7411 & ~w16628 ;
  assign w19488 = ( w7944 & w16619 ) | ( w7944 & w19487 ) | ( w16619 & w19487 ) ;
  assign w19489 = w7673 | w19488 ;
  assign w19490 = ( ~w16626 & w19488 ) | ( ~w16626 & w19489 ) | ( w19488 & w19489 ) ;
  assign w19491 = w19487 | w19490 ;
  assign w19492 = ~w7414 & w18451 ;
  assign w19493 = ( w18451 & w19491 ) | ( w18451 & ~w19492 ) | ( w19491 & ~w19492 ) ;
  assign w19494 = \pi08 ^ w19493 ;
  assign w19495 = w19382 ^ w19494 ;
  assign w19496 = w19486 ^ w19495 ;
  assign w19497 = ( w16737 & ~w18434 ) | ( w16737 & w18764 ) | ( ~w18434 & w18764 ) ;
  assign w19498 = w19381 ^ w19497 ;
  assign w19499 = w19496 ^ w19498 ;
  assign w19500 = ( w18874 & ~w18908 ) | ( w18874 & w18910 ) | ( ~w18908 & w18910 ) ;
  assign w19501 = ( ~w18897 & w18905 ) | ( ~w18897 & w18906 ) | ( w18905 & w18906 ) ;
  assign w19502 = ( \pi29 & \pi31 ) | ( \pi29 & ~w10885 ) | ( \pi31 & ~w10885 ) ;
  assign w19503 = ( \pi29 & ~\pi30 ) | ( \pi29 & w19502 ) | ( ~\pi30 & w19502 ) ;
  assign w19504 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w19502 ) | ( \pi30 & w19502 ) ;
  assign w19505 = ( \pi29 & w10866 ) | ( \pi29 & ~w19504 ) | ( w10866 & ~w19504 ) ;
  assign w19506 = ( ~w10887 & w19504 ) | ( ~w10887 & w19505 ) | ( w19504 & w19505 ) ;
  assign w19507 = ~\pi31 & w19506 ;
  assign w19508 = ( w19503 & ~w19505 ) | ( w19503 & w19507 ) | ( ~w19505 & w19507 ) ;
  assign w19509 = ( w37 & ~w11131 ) | ( w37 & w19508 ) | ( ~w11131 & w19508 ) ;
  assign w19510 = w19508 | w19509 ;
  assign w19511 = ( w18789 & w18886 ) | ( w18789 & w18893 ) | ( w18886 & w18893 ) ;
  assign w19512 = w312 | w4596 ;
  assign w19513 = ( w4126 & ~w4596 ) | ( w4126 & w18888 ) | ( ~w4596 & w18888 ) ;
  assign w19514 = w19512 | w19513 ;
  assign w19515 = w19510 ^ w19511 ;
  assign w19516 = w19514 ^ w19515 ;
  assign w19517 = ( w18844 & w18883 ) | ( w18844 & ~w18895 ) | ( w18883 & ~w18895 ) ;
  assign w19518 = w3717 | w11139 ;
  assign w19519 = w3649 & w10883 ;
  assign w19520 = ( ~w11139 & w19518 ) | ( ~w11139 & w19519 ) | ( w19518 & w19519 ) ;
  assign w19521 = w3549 | w10738 ;
  assign w19522 = w11145 & ~w19520 ;
  assign w19523 = ( w3448 & w19520 ) | ( w3448 & ~w19522 ) | ( w19520 & ~w19522 ) ;
  assign w19524 = ( ~w10738 & w19521 ) | ( ~w10738 & w19523 ) | ( w19521 & w19523 ) ;
  assign w19525 = \pi29 ^ w19524 ;
  assign w19526 = w19516 ^ w19525 ;
  assign w19527 = w19517 ^ w19526 ;
  assign w19528 = w19500 ^ w19501 ;
  assign w19529 = w19527 ^ w19528 ;
  assign w19530 = ( \pi02 & w18912 ) | ( \pi02 & ~w19529 ) | ( w18912 & ~w19529 ) ;
  assign w19531 = \pi00 ^ w19530 ;
  assign w19532 = ( \pi02 & w19529 ) | ( \pi02 & w19531 ) | ( w19529 & w19531 ) ;
  assign w19533 = ( ~\pi02 & w18912 ) | ( ~\pi02 & w19531 ) | ( w18912 & w19531 ) ;
  assign w19534 = \pi01 & ~w19533 ;
  assign w19535 = ( ~\pi00 & w18916 ) | ( ~\pi00 & w19534 ) | ( w18916 & w19534 ) ;
  assign w19536 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19535 ) | ( \pi02 & ~w19535 ) ;
  assign w19537 = ( w19532 & w19534 ) | ( w19532 & ~w19536 ) | ( w19534 & ~w19536 ) ;
  assign w19538 = ( ~w18912 & w18927 ) | ( ~w18912 & w19529 ) | ( w18927 & w19529 ) ;
  assign w19539 = w18927 ^ w19529 ;
  assign w19540 = w18912 ^ w19539 ;
  assign w19541 = w8954 & w19540 ;
  assign w19542 = ( w8954 & w19537 ) | ( w8954 & ~w19541 ) | ( w19537 & ~w19541 ) ;
  assign w19543 = w19373 ^ w19542 ;
  assign w19544 = \pi02 ^ w19499 ;
  assign w19545 = w19543 ^ w19544 ;
  assign w19546 = w18932 ^ w19372 ;
  assign w19547 = w18766 ^ w19546 ;
  assign w19548 = w19545 ^ w19547 ;
  assign w19549 = w19545 | w19547 ;
  assign w19550 = ~w19537 & w19540 ;
  assign w19551 = ( w8954 & w19537 ) | ( w8954 & ~w19550 ) | ( w19537 & ~w19550 ) ;
  assign w19552 = \pi02 ^ w19551 ;
  assign w19553 = ( w19373 & ~w19499 ) | ( w19373 & w19552 ) | ( ~w19499 & w19552 ) ;
  assign w19554 = w8593 | w18914 ;
  assign w19555 = w8262 & w16617 ;
  assign w19556 = ( ~w18914 & w19554 ) | ( ~w18914 & w19555 ) | ( w19554 & w19555 ) ;
  assign w19557 = w8263 | w19366 ;
  assign w19558 = w18916 | w19556 ;
  assign w19559 = ( w35 & w19556 ) | ( w35 & w19558 ) | ( w19556 & w19558 ) ;
  assign w19560 = ( ~w19366 & w19557 ) | ( ~w19366 & w19559 ) | ( w19557 & w19559 ) ;
  assign w19561 = \pi05 ^ w19560 ;
  assign w19562 = ( w19382 & ~w19486 ) | ( w19382 & w19494 ) | ( ~w19486 & w19494 ) ;
  assign w19563 = w6949 | w16630 ;
  assign w19564 = w6748 & w16632 ;
  assign w19565 = ( ~w16630 & w19563 ) | ( ~w16630 & w19564 ) | ( w19563 & w19564 ) ;
  assign w19566 = w7154 | w16628 ;
  assign w19567 = w18026 | w19565 ;
  assign w19568 = ( w6751 & w19565 ) | ( w6751 & w19567 ) | ( w19565 & w19567 ) ;
  assign w19569 = ( ~w16628 & w19566 ) | ( ~w16628 & w19568 ) | ( w19566 & w19568 ) ;
  assign w19570 = \pi11 ^ w19569 ;
  assign w19571 = ( w19391 & ~w19473 ) | ( w19391 & w19481 ) | ( ~w19473 & w19481 ) ;
  assign w19572 = ~w5710 & w16642 ;
  assign w19573 = w5494 & ~w16644 ;
  assign w19574 = ( w16642 & ~w19572 ) | ( w16642 & w19573 ) | ( ~w19572 & w19573 ) ;
  assign w19575 = ~w5948 & w16640 ;
  assign w19576 = w17760 & ~w19574 ;
  assign w19577 = ( w5497 & w19574 ) | ( w5497 & ~w19576 ) | ( w19574 & ~w19576 ) ;
  assign w19578 = ( w16640 & ~w19575 ) | ( w16640 & w19577 ) | ( ~w19575 & w19577 ) ;
  assign w19579 = \pi17 ^ w19578 ;
  assign w19580 = ( w19400 & ~w19460 ) | ( w19400 & w19468 ) | ( ~w19460 & w19468 ) ;
  assign w19581 = ~w4651 & w16654 ;
  assign w19582 = w4606 & ~w16656 ;
  assign w19583 = ( w16654 & ~w19581 ) | ( w16654 & w19582 ) | ( ~w19581 & w19582 ) ;
  assign w19584 = w4706 | w16652 ;
  assign w19585 = w17293 | w19583 ;
  assign w19586 = ( w4609 & w19583 ) | ( w4609 & w19585 ) | ( w19583 & w19585 ) ;
  assign w19587 = ( ~w16652 & w19584 ) | ( ~w16652 & w19586 ) | ( w19584 & w19586 ) ;
  assign w19588 = \pi23 ^ w19587 ;
  assign w19589 = ( w19409 & ~w19447 ) | ( w19409 & w19455 ) | ( ~w19447 & w19455 ) ;
  assign w19590 = ( w19417 & ~w19444 ) | ( w19417 & w19445 ) | ( ~w19444 & w19445 ) ;
  assign w19591 = ( w19418 & ~w19434 ) | ( w19418 & w19442 ) | ( ~w19434 & w19442 ) ;
  assign w19592 = ( w164 & w262 ) | ( w164 & ~w419 ) | ( w262 & ~w419 ) ;
  assign w19593 = w988 | w2095 ;
  assign w19594 = ( w419 & w1086 ) | ( w419 & ~w2095 ) | ( w1086 & ~w2095 ) ;
  assign w19595 = w19593 | w19594 ;
  assign w19596 = w19592 | w19595 ;
  assign w19597 = w6265 | w19596 ;
  assign w19598 = w11614 | w19597 ;
  assign w19599 = ( w3059 & w6409 ) | ( w3059 & ~w11614 ) | ( w6409 & ~w11614 ) ;
  assign w19600 = w19598 | w19599 ;
  assign w19601 = ( ~w210 & w1616 ) | ( ~w210 & w2705 ) | ( w1616 & w2705 ) ;
  assign w19602 = w1265 | w19600 ;
  assign w19603 = ( w210 & w899 ) | ( w210 & ~w1265 ) | ( w899 & ~w1265 ) ;
  assign w19604 = w19602 | w19603 ;
  assign w19605 = w19601 | w19604 ;
  assign w19606 = w565 | w1274 ;
  assign w19607 = w2517 | w19606 ;
  assign w19608 = ( w199 & ~w2517 ) | ( w199 & w19605 ) | ( ~w2517 & w19605 ) ;
  assign w19609 = w19607 | w19608 ;
  assign w19610 = ( ~w314 & w359 ) | ( ~w314 & w783 ) | ( w359 & w783 ) ;
  assign w19611 = w278 | w19609 ;
  assign w19612 = ( ~w278 & w783 ) | ( ~w278 & w951 ) | ( w783 & w951 ) ;
  assign w19613 = w19611 | w19612 ;
  assign w19614 = w19610 & ~w19613 ;
  assign w19615 = w37 | w16772 ;
  assign w19616 = w3098 & ~w16690 ;
  assign w19617 = ( ~w16772 & w19615 ) | ( ~w16772 & w19616 ) | ( w19615 & w19616 ) ;
  assign w19618 = ( \pi29 & \pi30 ) | ( \pi29 & w16680 ) | ( \pi30 & w16680 ) ;
  assign w19619 = \pi31 | w19618 ;
  assign w19620 = ( \pi29 & ~\pi30 ) | ( \pi29 & w16685 ) | ( ~\pi30 & w16685 ) ;
  assign w19621 = ( \pi29 & \pi31 ) | ( \pi29 & ~w19620 ) | ( \pi31 & ~w19620 ) ;
  assign w19622 = ( w19617 & w19619 ) | ( w19617 & ~w19621 ) | ( w19619 & ~w19621 ) ;
  assign w19623 = w19591 ^ w19622 ;
  assign w19624 = w19614 ^ w19623 ;
  assign w19625 = w3549 & w16665 ;
  assign w19626 = ( w3717 & w16670 ) | ( w3717 & w19625 ) | ( w16670 & w19625 ) ;
  assign w19627 = w3649 | w19626 ;
  assign w19628 = ( w16675 & w19626 ) | ( w16675 & w19627 ) | ( w19626 & w19627 ) ;
  assign w19629 = w19625 | w19628 ;
  assign w19630 = ~w3448 & w16960 ;
  assign w19631 = ( w16960 & w19629 ) | ( w16960 & ~w19630 ) | ( w19629 & ~w19630 ) ;
  assign w19632 = \pi29 ^ w19631 ;
  assign w19633 = w19590 ^ w19632 ;
  assign w19634 = w19624 ^ w19633 ;
  assign w19635 = w3964 & ~w16658 ;
  assign w19636 = ( w4143 & w16660 ) | ( w4143 & w19635 ) | ( w16660 & w19635 ) ;
  assign w19637 = w4052 | w19636 ;
  assign w19638 = ( ~w16662 & w19636 ) | ( ~w16662 & w19637 ) | ( w19636 & w19637 ) ;
  assign w19639 = w19635 | w19638 ;
  assign w19640 = w4147 | w17065 ;
  assign w19641 = ( ~w17065 & w19639 ) | ( ~w17065 & w19640 ) | ( w19639 & w19640 ) ;
  assign w19642 = \pi26 ^ w19641 ;
  assign w19643 = w19589 ^ w19642 ;
  assign w19644 = w19634 ^ w19643 ;
  assign w19645 = ( w19408 & ~w19457 ) | ( w19408 & w19458 ) | ( ~w19457 & w19458 ) ;
  assign w19646 = w19588 ^ w19645 ;
  assign w19647 = w19644 ^ w19646 ;
  assign w19648 = w4905 & ~w16650 ;
  assign w19649 = ( w5395 & ~w16646 ) | ( w5395 & w19648 ) | ( ~w16646 & w19648 ) ;
  assign w19650 = w5343 | w19649 ;
  assign w19651 = ( ~w16648 & w19649 ) | ( ~w16648 & w19650 ) | ( w19649 & w19650 ) ;
  assign w19652 = w19648 | w19651 ;
  assign w19653 = w4908 | w17476 ;
  assign w19654 = ( ~w17476 & w19652 ) | ( ~w17476 & w19653 ) | ( w19652 & w19653 ) ;
  assign w19655 = \pi20 ^ w19654 ;
  assign w19656 = w19580 ^ w19655 ;
  assign w19657 = w19647 ^ w19656 ;
  assign w19658 = ( w19399 & ~w19470 ) | ( w19399 & w19471 ) | ( ~w19470 & w19471 ) ;
  assign w19659 = w19579 ^ w19658 ;
  assign w19660 = w19657 ^ w19659 ;
  assign w19661 = w6048 & ~w16638 ;
  assign w19662 = ( w6637 & ~w16634 ) | ( w6637 & w19661 ) | ( ~w16634 & w19661 ) ;
  assign w19663 = w6549 | w19662 ;
  assign w19664 = ( w16636 & w19662 ) | ( w16636 & w19663 ) | ( w19662 & w19663 ) ;
  assign w19665 = w19661 | w19664 ;
  assign w19666 = w6045 | w16742 ;
  assign w19667 = ( ~w16742 & w19665 ) | ( ~w16742 & w19666 ) | ( w19665 & w19666 ) ;
  assign w19668 = \pi14 ^ w19667 ;
  assign w19669 = w19571 ^ w19668 ;
  assign w19670 = w19660 ^ w19669 ;
  assign w19671 = ( w19390 & ~w19483 ) | ( w19390 & w19484 ) | ( ~w19483 & w19484 ) ;
  assign w19672 = w19570 ^ w19671 ;
  assign w19673 = w19670 ^ w19672 ;
  assign w19674 = w7411 & ~w16626 ;
  assign w19675 = ( w7944 & w16621 ) | ( w7944 & w19674 ) | ( w16621 & w19674 ) ;
  assign w19676 = w7673 | w19675 ;
  assign w19677 = ( w16619 & w19675 ) | ( w16619 & w19676 ) | ( w19675 & w19676 ) ;
  assign w19678 = w19674 | w19677 ;
  assign w19679 = w7414 | w18439 ;
  assign w19680 = ( ~w18439 & w19678 ) | ( ~w18439 & w19679 ) | ( w19678 & w19679 ) ;
  assign w19681 = \pi08 ^ w19680 ;
  assign w19682 = w19562 ^ w19681 ;
  assign w19683 = w19673 ^ w19682 ;
  assign w19684 = ( w19381 & ~w19496 ) | ( w19381 & w19497 ) | ( ~w19496 & w19497 ) ;
  assign w19685 = w19561 ^ w19684 ;
  assign w19686 = w19683 ^ w19685 ;
  assign w19687 = ( w19500 & w19501 ) | ( w19500 & w19527 ) | ( w19501 & w19527 ) ;
  assign w19688 = ( w19516 & w19517 ) | ( w19516 & w19525 ) | ( w19517 & w19525 ) ;
  assign w19689 = ( ~w19510 & w19511 ) | ( ~w19510 & w19514 ) | ( w19511 & w19514 ) ;
  assign w19690 = w3945 | w4599 ;
  assign w19691 = ( ~w19514 & w19689 ) | ( ~w19514 & w19690 ) | ( w19689 & w19690 ) ;
  assign w19692 = w19514 ^ w19689 ;
  assign w19693 = w19690 ^ w19692 ;
  assign w19694 = ( w3549 & w3649 ) | ( w3549 & ~w11138 ) | ( w3649 & ~w11138 ) ;
  assign w19695 = w3549 & ~w19694 ;
  assign w19696 = ( w3717 & ~w19694 ) | ( w3717 & w19695 ) | ( ~w19694 & w19695 ) ;
  assign w19697 = ( ~w10738 & w19694 ) | ( ~w10738 & w19696 ) | ( w19694 & w19696 ) ;
  assign w19698 = w3448 | w11146 ;
  assign w19699 = ( ~w11146 & w19697 ) | ( ~w11146 & w19698 ) | ( w19697 & w19698 ) ;
  assign w19700 = \pi29 ^ w19699 ;
  assign w19701 = ( \pi29 & \pi31 ) | ( \pi29 & ~w10887 ) | ( \pi31 & ~w10887 ) ;
  assign w19702 = ( \pi29 & ~\pi30 ) | ( \pi29 & w19701 ) | ( ~\pi30 & w19701 ) ;
  assign w19703 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w19701 ) | ( \pi30 & w19701 ) ;
  assign w19704 = ( \pi29 & w10885 ) | ( \pi29 & ~w19703 ) | ( w10885 & ~w19703 ) ;
  assign w19705 = ( w10883 & w19703 ) | ( w10883 & w19704 ) | ( w19703 & w19704 ) ;
  assign w19706 = ~\pi31 & w19705 ;
  assign w19707 = ( w19702 & ~w19704 ) | ( w19702 & w19706 ) | ( ~w19704 & w19706 ) ;
  assign w19708 = ( w37 & w10895 ) | ( w37 & w19707 ) | ( w10895 & w19707 ) ;
  assign w19709 = w19707 | w19708 ;
  assign w19710 = w19693 ^ w19700 ;
  assign w19711 = w19709 ^ w19710 ;
  assign w19712 = w19687 ^ w19688 ;
  assign w19713 = w19711 ^ w19712 ;
  assign w19714 = ( ~\pi02 & w19529 ) | ( ~\pi02 & w19713 ) | ( w19529 & w19713 ) ;
  assign w19715 = \pi00 ^ w19714 ;
  assign w19716 = ( \pi02 & w19713 ) | ( \pi02 & ~w19715 ) | ( w19713 & ~w19715 ) ;
  assign w19717 = ( \pi02 & w19529 ) | ( \pi02 & w19715 ) | ( w19529 & w19715 ) ;
  assign w19718 = \pi01 & w19717 ;
  assign w19719 = ( \pi00 & w18912 ) | ( \pi00 & ~w19718 ) | ( w18912 & ~w19718 ) ;
  assign w19720 = ( \pi01 & \pi02 ) | ( \pi01 & w19719 ) | ( \pi02 & w19719 ) ;
  assign w19721 = ( w19716 & w19718 ) | ( w19716 & ~w19720 ) | ( w19718 & ~w19720 ) ;
  assign w19722 = w19538 ^ w19713 ;
  assign w19723 = w19529 ^ w19722 ;
  assign w19724 = w8954 & ~w19723 ;
  assign w19725 = ( w8954 & w19721 ) | ( w8954 & ~w19724 ) | ( w19721 & ~w19724 ) ;
  assign w19726 = w19553 ^ w19725 ;
  assign w19727 = \pi02 ^ w19686 ;
  assign w19728 = w19726 ^ w19727 ;
  assign w19729 = w19549 | w19728 ;
  assign w19730 = w19549 ^ w19728 ;
  assign w19731 = w19721 | w19723 ;
  assign w19732 = ( w8954 & w19721 ) | ( w8954 & w19731 ) | ( w19721 & w19731 ) ;
  assign w19733 = \pi02 ^ w19732 ;
  assign w19734 = ( w19553 & ~w19686 ) | ( w19553 & w19733 ) | ( ~w19686 & w19733 ) ;
  assign w19735 = ~w8593 & w18916 ;
  assign w19736 = w8262 & ~w18914 ;
  assign w19737 = ( w18916 & ~w19735 ) | ( w18916 & w19736 ) | ( ~w19735 & w19736 ) ;
  assign w19738 = w8263 | w18929 ;
  assign w19739 = w18912 & ~w19737 ;
  assign w19740 = ( w35 & w19737 ) | ( w35 & ~w19739 ) | ( w19737 & ~w19739 ) ;
  assign w19741 = ( ~w18929 & w19738 ) | ( ~w18929 & w19740 ) | ( w19738 & w19740 ) ;
  assign w19742 = \pi05 ^ w19741 ;
  assign w19743 = ( w19562 & ~w19673 ) | ( w19562 & w19681 ) | ( ~w19673 & w19681 ) ;
  assign w19744 = w6949 | w16628 ;
  assign w19745 = w6748 & ~w16630 ;
  assign w19746 = ( ~w16628 & w19744 ) | ( ~w16628 & w19745 ) | ( w19744 & w19745 ) ;
  assign w19747 = w7154 | w16626 ;
  assign w19748 = w18429 & ~w19746 ;
  assign w19749 = ( w6751 & w19746 ) | ( w6751 & ~w19748 ) | ( w19746 & ~w19748 ) ;
  assign w19750 = ( ~w16626 & w19747 ) | ( ~w16626 & w19749 ) | ( w19747 & w19749 ) ;
  assign w19751 = \pi11 ^ w19750 ;
  assign w19752 = ( w19571 & ~w19660 ) | ( w19571 & w19668 ) | ( ~w19660 & w19668 ) ;
  assign w19753 = ~w5710 & w16640 ;
  assign w19754 = w5494 & w16642 ;
  assign w19755 = ( w16640 & ~w19753 ) | ( w16640 & w19754 ) | ( ~w19753 & w19754 ) ;
  assign w19756 = w5948 | w16638 ;
  assign w19757 = w17783 & ~w19755 ;
  assign w19758 = ( w5497 & w19755 ) | ( w5497 & ~w19757 ) | ( w19755 & ~w19757 ) ;
  assign w19759 = ( ~w16638 & w19756 ) | ( ~w16638 & w19758 ) | ( w19756 & w19758 ) ;
  assign w19760 = \pi17 ^ w19759 ;
  assign w19761 = ( w19580 & ~w19647 ) | ( w19580 & w19655 ) | ( ~w19647 & w19655 ) ;
  assign w19762 = w4651 | w16652 ;
  assign w19763 = w4606 & w16654 ;
  assign w19764 = ( ~w16652 & w19762 ) | ( ~w16652 & w19763 ) | ( w19762 & w19763 ) ;
  assign w19765 = w4706 | w16650 ;
  assign w19766 = w17277 & ~w19764 ;
  assign w19767 = ( w4609 & w19764 ) | ( w4609 & ~w19766 ) | ( w19764 & ~w19766 ) ;
  assign w19768 = ( ~w16650 & w19765 ) | ( ~w16650 & w19767 ) | ( w19765 & w19767 ) ;
  assign w19769 = \pi23 ^ w19768 ;
  assign w19770 = ( w19589 & ~w19634 ) | ( w19589 & w19642 ) | ( ~w19634 & w19642 ) ;
  assign w19771 = ( w19590 & ~w19624 ) | ( w19590 & w19632 ) | ( ~w19624 & w19632 ) ;
  assign w19772 = ( w19591 & ~w19614 ) | ( w19591 & w19622 ) | ( ~w19614 & w19622 ) ;
  assign w19773 = w596 | w726 ;
  assign w19774 = w1565 | w19773 ;
  assign w19775 = ( w315 & w784 ) | ( w315 & ~w1565 ) | ( w784 & ~w1565 ) ;
  assign w19776 = w19774 | w19775 ;
  assign w19777 = w1155 | w6366 ;
  assign w19778 = ( ~w1155 & w2522 ) | ( ~w1155 & w19776 ) | ( w2522 & w19776 ) ;
  assign w19779 = w19777 | w19778 ;
  assign w19780 = ( ~w622 & w3285 ) | ( ~w622 & w19779 ) | ( w3285 & w19779 ) ;
  assign w19781 = w1645 | w3273 ;
  assign w19782 = ( w622 & w1513 ) | ( w622 & ~w3273 ) | ( w1513 & ~w3273 ) ;
  assign w19783 = w19781 | w19782 ;
  assign w19784 = w19780 | w19783 ;
  assign w19785 = ( ~w147 & w514 ) | ( ~w147 & w1302 ) | ( w514 & w1302 ) ;
  assign w19786 = w1903 | w19784 ;
  assign w19787 = ( w147 & w205 ) | ( w147 & ~w1903 ) | ( w205 & ~w1903 ) ;
  assign w19788 = w19786 | w19787 ;
  assign w19789 = w19785 | w19788 ;
  assign w19790 = ( w223 & w268 ) | ( w223 & ~w467 ) | ( w268 & ~w467 ) ;
  assign w19791 = w74 | w19789 ;
  assign w19792 = ( ~w74 & w467 ) | ( ~w74 & w490 ) | ( w467 & w490 ) ;
  assign w19793 = w19791 | w19792 ;
  assign w19794 = w19790 | w19793 ;
  assign w19795 = ~w37 & w16946 ;
  assign w19796 = w3098 & w16685 ;
  assign w19797 = ( w16946 & ~w19795 ) | ( w16946 & w19796 ) | ( ~w19795 & w19796 ) ;
  assign w19798 = ( \pi29 & \pi30 ) | ( \pi29 & w16675 ) | ( \pi30 & w16675 ) ;
  assign w19799 = \pi31 | w19798 ;
  assign w19800 = ( \pi29 & ~\pi30 ) | ( \pi29 & w16680 ) | ( ~\pi30 & w16680 ) ;
  assign w19801 = ( \pi29 & \pi31 ) | ( \pi29 & ~w19800 ) | ( \pi31 & ~w19800 ) ;
  assign w19802 = ( w19797 & w19799 ) | ( w19797 & ~w19801 ) | ( w19799 & ~w19801 ) ;
  assign w19803 = w19772 ^ w19802 ;
  assign w19804 = w19794 ^ w19803 ;
  assign w19805 = w3549 & ~w16662 ;
  assign w19806 = ( w3717 & w16665 ) | ( w3717 & w19805 ) | ( w16665 & w19805 ) ;
  assign w19807 = w3649 | w19806 ;
  assign w19808 = ( w16670 & w19806 ) | ( w16670 & w19807 ) | ( w19806 & w19807 ) ;
  assign w19809 = w19805 | w19808 ;
  assign w19810 = w3448 | w16762 ;
  assign w19811 = ( ~w16762 & w19809 ) | ( ~w16762 & w19810 ) | ( w19809 & w19810 ) ;
  assign w19812 = \pi29 ^ w19811 ;
  assign w19813 = w19771 ^ w19812 ;
  assign w19814 = w19804 ^ w19813 ;
  assign w19815 = w3964 & ~w16656 ;
  assign w19816 = ( w4143 & ~w16658 ) | ( w4143 & w19815 ) | ( ~w16658 & w19815 ) ;
  assign w19817 = w4052 | w19816 ;
  assign w19818 = ( w16660 & w19816 ) | ( w16660 & w19817 ) | ( w19816 & w19817 ) ;
  assign w19819 = w19815 | w19818 ;
  assign w19820 = ~w4147 & w17057 ;
  assign w19821 = ( w17057 & w19819 ) | ( w17057 & ~w19820 ) | ( w19819 & ~w19820 ) ;
  assign w19822 = \pi26 ^ w19821 ;
  assign w19823 = w19770 ^ w19822 ;
  assign w19824 = w19814 ^ w19823 ;
  assign w19825 = ( w19588 & ~w19644 ) | ( w19588 & w19645 ) | ( ~w19644 & w19645 ) ;
  assign w19826 = w19769 ^ w19825 ;
  assign w19827 = w19824 ^ w19826 ;
  assign w19828 = w4905 & ~w16648 ;
  assign w19829 = ( w5395 & ~w16644 ) | ( w5395 & w19828 ) | ( ~w16644 & w19828 ) ;
  assign w19830 = w5343 | w19829 ;
  assign w19831 = ( ~w16646 & w19829 ) | ( ~w16646 & w19830 ) | ( w19829 & w19830 ) ;
  assign w19832 = w19828 | w19831 ;
  assign w19833 = w4908 | w17468 ;
  assign w19834 = ( ~w17468 & w19832 ) | ( ~w17468 & w19833 ) | ( w19832 & w19833 ) ;
  assign w19835 = \pi20 ^ w19834 ;
  assign w19836 = w19761 ^ w19835 ;
  assign w19837 = w19827 ^ w19836 ;
  assign w19838 = ( w19579 & ~w19657 ) | ( w19579 & w19658 ) | ( ~w19657 & w19658 ) ;
  assign w19839 = w19760 ^ w19838 ;
  assign w19840 = w19837 ^ w19839 ;
  assign w19841 = w6048 & w16636 ;
  assign w19842 = ( w6637 & w16632 ) | ( w6637 & w19841 ) | ( w16632 & w19841 ) ;
  assign w19843 = w6549 | w19842 ;
  assign w19844 = ( ~w16634 & w19842 ) | ( ~w16634 & w19843 ) | ( w19842 & w19843 ) ;
  assign w19845 = w19841 | w19844 ;
  assign w19846 = w6045 | w18051 ;
  assign w19847 = ( ~w18051 & w19845 ) | ( ~w18051 & w19846 ) | ( w19845 & w19846 ) ;
  assign w19848 = \pi14 ^ w19847 ;
  assign w19849 = w19752 ^ w19848 ;
  assign w19850 = w19840 ^ w19849 ;
  assign w19851 = ( w19570 & ~w19670 ) | ( w19570 & w19671 ) | ( ~w19670 & w19671 ) ;
  assign w19852 = w19751 ^ w19851 ;
  assign w19853 = w19850 ^ w19852 ;
  assign w19854 = ~w7673 & w16621 ;
  assign w19855 = w7411 & w16619 ;
  assign w19856 = ( w16621 & ~w19854 ) | ( w16621 & w19855 ) | ( ~w19854 & w19855 ) ;
  assign w19857 = ~w7944 & w16617 ;
  assign w19858 = w16732 | w19856 ;
  assign w19859 = ( w7414 & w19856 ) | ( w7414 & w19858 ) | ( w19856 & w19858 ) ;
  assign w19860 = ( w16617 & ~w19857 ) | ( w16617 & w19859 ) | ( ~w19857 & w19859 ) ;
  assign w19861 = \pi08 ^ w19860 ;
  assign w19862 = w19743 ^ w19861 ;
  assign w19863 = w19853 ^ w19862 ;
  assign w19864 = ( w19561 & ~w19683 ) | ( w19561 & w19684 ) | ( ~w19683 & w19684 ) ;
  assign w19865 = w19742 ^ w19864 ;
  assign w19866 = w19863 ^ w19865 ;
  assign w19867 = ( w19687 & w19688 ) | ( w19687 & w19711 ) | ( w19688 & w19711 ) ;
  assign w19868 = ( w19693 & w19700 ) | ( w19693 & w19709 ) | ( w19700 & w19709 ) ;
  assign w19869 = ( \pi29 & \pi31 ) | ( \pi29 & w10883 ) | ( \pi31 & w10883 ) ;
  assign w19870 = ( \pi29 & ~\pi30 ) | ( \pi29 & w19869 ) | ( ~\pi30 & w19869 ) ;
  assign w19871 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w19869 ) | ( \pi30 & w19869 ) ;
  assign w19872 = ( \pi29 & w10887 ) | ( \pi29 & ~w19871 ) | ( w10887 & ~w19871 ) ;
  assign w19873 = ( ~w11139 & w19871 ) | ( ~w11139 & w19872 ) | ( w19871 & w19872 ) ;
  assign w19874 = ~\pi31 & w19873 ;
  assign w19875 = ( w19870 & ~w19872 ) | ( w19870 & w19874 ) | ( ~w19872 & w19874 ) ;
  assign w19876 = ( w37 & w11256 ) | ( w37 & w19875 ) | ( w11256 & w19875 ) ;
  assign w19877 = w19875 | w19876 ;
  assign w19878 = ( \pi26 & \pi27 ) | ( \pi26 & ~\pi28 ) | ( \pi27 & ~\pi28 ) ;
  assign w19879 = ( \pi28 & ~\pi29 ) | ( \pi28 & w19878 ) | ( ~\pi29 & w19878 ) ;
  assign w19880 = w10738 ^ w19879 ;
  assign w19881 = ( \pi29 & w19879 ) | ( \pi29 & w19880 ) | ( w19879 & w19880 ) ;
  assign w19882 = w10399 ^ w19881 ;
  assign w19883 = w19690 ^ w19882 ;
  assign w19884 = w19691 ^ w19877 ;
  assign w19885 = w19883 ^ w19884 ;
  assign w19886 = w19867 ^ w19868 ;
  assign w19887 = w19885 ^ w19886 ;
  assign w19888 = ( ~\pi02 & w19713 ) | ( ~\pi02 & w19887 ) | ( w19713 & w19887 ) ;
  assign w19889 = \pi00 ^ w19888 ;
  assign w19890 = ( \pi02 & w19887 ) | ( \pi02 & ~w19889 ) | ( w19887 & ~w19889 ) ;
  assign w19891 = ( \pi02 & w19713 ) | ( \pi02 & w19889 ) | ( w19713 & w19889 ) ;
  assign w19892 = \pi01 & w19891 ;
  assign w19893 = ( ~\pi00 & w19529 ) | ( ~\pi00 & w19892 ) | ( w19529 & w19892 ) ;
  assign w19894 = ( \pi01 & \pi02 ) | ( \pi01 & ~w19893 ) | ( \pi02 & ~w19893 ) ;
  assign w19895 = ( w19890 & w19892 ) | ( w19890 & ~w19894 ) | ( w19892 & ~w19894 ) ;
  assign w19896 = ( ~w19529 & w19538 ) | ( ~w19529 & w19713 ) | ( w19538 & w19713 ) ;
  assign w19897 = w19538 ^ w19896 ;
  assign w19898 = w19887 ^ w19897 ;
  assign w19899 = w8954 & ~w19898 ;
  assign w19900 = ( w8954 & w19895 ) | ( w8954 & ~w19899 ) | ( w19895 & ~w19899 ) ;
  assign w19901 = w19734 ^ w19900 ;
  assign w19902 = \pi02 ^ w19866 ;
  assign w19903 = w19901 ^ w19902 ;
  assign w19904 = ~w19729 & w19903 ;
  assign w19905 = w19729 ^ w19903 ;
  assign w19906 = w19895 | w19898 ;
  assign w19907 = ( w8954 & w19895 ) | ( w8954 & w19906 ) | ( w19895 & w19906 ) ;
  assign w19908 = \pi02 ^ w19907 ;
  assign w19909 = ( w19734 & w19866 ) | ( w19734 & w19908 ) | ( w19866 & w19908 ) ;
  assign w19910 = w8593 | w18912 ;
  assign w19911 = w8262 & w18916 ;
  assign w19912 = ( ~w18912 & w19910 ) | ( ~w18912 & w19911 ) | ( w19910 & w19911 ) ;
  assign w19913 = w8263 | w19540 ;
  assign w19914 = w19529 | w19912 ;
  assign w19915 = ( w35 & w19912 ) | ( w35 & w19914 ) | ( w19912 & w19914 ) ;
  assign w19916 = ( ~w19540 & w19913 ) | ( ~w19540 & w19915 ) | ( w19913 & w19915 ) ;
  assign w19917 = \pi05 ^ w19916 ;
  assign w19918 = ( w19743 & w19853 ) | ( w19743 & w19861 ) | ( w19853 & w19861 ) ;
  assign w19919 = w6949 | w16626 ;
  assign w19920 = w6748 & ~w16628 ;
  assign w19921 = ( ~w16626 & w19919 ) | ( ~w16626 & w19920 ) | ( w19919 & w19920 ) ;
  assign w19922 = ~w7154 & w16619 ;
  assign w19923 = w18451 | w19921 ;
  assign w19924 = ( w6751 & w19921 ) | ( w6751 & w19923 ) | ( w19921 & w19923 ) ;
  assign w19925 = ( w16619 & ~w19922 ) | ( w16619 & w19924 ) | ( ~w19922 & w19924 ) ;
  assign w19926 = \pi11 ^ w19925 ;
  assign w19927 = ( w19752 & w19840 ) | ( w19752 & w19848 ) | ( w19840 & w19848 ) ;
  assign w19928 = w5710 | w16638 ;
  assign w19929 = w5494 & w16640 ;
  assign w19930 = ( ~w16638 & w19928 ) | ( ~w16638 & w19929 ) | ( w19928 & w19929 ) ;
  assign w19931 = ~w5948 & w16636 ;
  assign w19932 = w17770 & ~w19930 ;
  assign w19933 = ( w5497 & w19930 ) | ( w5497 & ~w19932 ) | ( w19930 & ~w19932 ) ;
  assign w19934 = ( w16636 & ~w19931 ) | ( w16636 & w19933 ) | ( ~w19931 & w19933 ) ;
  assign w19935 = \pi17 ^ w19934 ;
  assign w19936 = ( w19761 & w19827 ) | ( w19761 & w19835 ) | ( w19827 & w19835 ) ;
  assign w19937 = w4651 | w16650 ;
  assign w19938 = w4606 & ~w16652 ;
  assign w19939 = ( ~w16650 & w19937 ) | ( ~w16650 & w19938 ) | ( w19937 & w19938 ) ;
  assign w19940 = w4706 | w16648 ;
  assign w19941 = w16752 & ~w19939 ;
  assign w19942 = ( w4609 & w19939 ) | ( w4609 & ~w19941 ) | ( w19939 & ~w19941 ) ;
  assign w19943 = ( ~w16648 & w19940 ) | ( ~w16648 & w19942 ) | ( w19940 & w19942 ) ;
  assign w19944 = \pi23 ^ w19943 ;
  assign w19945 = ( w19770 & w19814 ) | ( w19770 & w19822 ) | ( w19814 & w19822 ) ;
  assign w19946 = ( w19771 & w19804 ) | ( w19771 & w19812 ) | ( w19804 & w19812 ) ;
  assign w19947 = ( w19772 & w19794 ) | ( w19772 & w19802 ) | ( w19794 & w19802 ) ;
  assign w19948 = w88 | w10501 ;
  assign w19949 = ( ~w88 & w126 ) | ( ~w88 & w149 ) | ( w126 & w149 ) ;
  assign w19950 = w19948 | w19949 ;
  assign w19951 = w447 | w516 ;
  assign w19952 = w1790 | w19951 ;
  assign w19953 = ( w175 & ~w1790 ) | ( w175 & w19950 ) | ( ~w1790 & w19950 ) ;
  assign w19954 = w19952 | w19953 ;
  assign w19955 = w2522 | w19954 ;
  assign w19956 = ( w573 & w901 ) | ( w573 & ~w2522 ) | ( w901 & ~w2522 ) ;
  assign w19957 = w19955 | w19956 ;
  assign w19958 = w4765 | w19957 ;
  assign w19959 = ( w6429 & ~w12462 ) | ( w6429 & w19958 ) | ( ~w12462 & w19958 ) ;
  assign w19960 = ~w2318 & w6385 ;
  assign w19961 = ( w510 & ~w2318 ) | ( w510 & w12462 ) | ( ~w2318 & w12462 ) ;
  assign w19962 = w19960 & ~w19961 ;
  assign w19963 = ~w19959 & w19962 ;
  assign w19964 = w165 | w325 ;
  assign w19965 = w1207 | w19964 ;
  assign w19966 = ( w1207 & ~w1883 ) | ( w1207 & w19963 ) | ( ~w1883 & w19963 ) ;
  assign w19967 = ~w19965 & w19966 ;
  assign w19968 = ~w37 & w16972 ;
  assign w19969 = w3098 & w16680 ;
  assign w19970 = ( w16972 & ~w19968 ) | ( w16972 & w19969 ) | ( ~w19968 & w19969 ) ;
  assign w19971 = ( \pi29 & \pi30 ) | ( \pi29 & w16670 ) | ( \pi30 & w16670 ) ;
  assign w19972 = \pi31 | w19971 ;
  assign w19973 = ( \pi29 & ~\pi30 ) | ( \pi29 & w16675 ) | ( ~\pi30 & w16675 ) ;
  assign w19974 = ( \pi29 & \pi31 ) | ( \pi29 & ~w19973 ) | ( \pi31 & ~w19973 ) ;
  assign w19975 = ( w19970 & w19972 ) | ( w19970 & ~w19974 ) | ( w19972 & ~w19974 ) ;
  assign w19976 = w19947 ^ w19975 ;
  assign w19977 = w19967 ^ w19976 ;
  assign w19978 = w3549 & w16660 ;
  assign w19979 = ( w3717 & ~w16662 ) | ( w3717 & w19978 ) | ( ~w16662 & w19978 ) ;
  assign w19980 = w3649 | w19979 ;
  assign w19981 = ( w16665 & w19979 ) | ( w16665 & w19980 ) | ( w19979 & w19980 ) ;
  assign w19982 = w19978 | w19981 ;
  assign w19983 = w3448 | w17078 ;
  assign w19984 = ( ~w17078 & w19982 ) | ( ~w17078 & w19983 ) | ( w19982 & w19983 ) ;
  assign w19985 = \pi29 ^ w19984 ;
  assign w19986 = w19946 ^ w19985 ;
  assign w19987 = w19977 ^ w19986 ;
  assign w19988 = w3964 & w16654 ;
  assign w19989 = ( w4143 & ~w16656 ) | ( w4143 & w19988 ) | ( ~w16656 & w19988 ) ;
  assign w19990 = w4052 | w19989 ;
  assign w19991 = ( ~w16658 & w19989 ) | ( ~w16658 & w19990 ) | ( w19989 & w19990 ) ;
  assign w19992 = w19988 | w19991 ;
  assign w19993 = ~w4147 & w17266 ;
  assign w19994 = ( w17266 & w19992 ) | ( w17266 & ~w19993 ) | ( w19992 & ~w19993 ) ;
  assign w19995 = \pi26 ^ w19994 ;
  assign w19996 = w19945 ^ w19995 ;
  assign w19997 = w19987 ^ w19996 ;
  assign w19998 = ( w19769 & w19824 ) | ( w19769 & w19825 ) | ( w19824 & w19825 ) ;
  assign w19999 = w19944 ^ w19998 ;
  assign w20000 = w19997 ^ w19999 ;
  assign w20001 = w4905 & ~w16646 ;
  assign w20002 = ( w5395 & w16642 ) | ( w5395 & w20001 ) | ( w16642 & w20001 ) ;
  assign w20003 = w5343 | w20002 ;
  assign w20004 = ( ~w16644 & w20002 ) | ( ~w16644 & w20003 ) | ( w20002 & w20003 ) ;
  assign w20005 = w20001 | w20004 ;
  assign w20006 = ~w4908 & w17455 ;
  assign w20007 = ( w17455 & w20005 ) | ( w17455 & ~w20006 ) | ( w20005 & ~w20006 ) ;
  assign w20008 = \pi20 ^ w20007 ;
  assign w20009 = w19936 ^ w20008 ;
  assign w20010 = w20000 ^ w20009 ;
  assign w20011 = ( w19760 & w19837 ) | ( w19760 & w19838 ) | ( w19837 & w19838 ) ;
  assign w20012 = w19935 ^ w20011 ;
  assign w20013 = w20010 ^ w20012 ;
  assign w20014 = w6048 & ~w16634 ;
  assign w20015 = ( w6637 & ~w16630 ) | ( w6637 & w20014 ) | ( ~w16630 & w20014 ) ;
  assign w20016 = w6549 | w20015 ;
  assign w20017 = ( w16632 & w20015 ) | ( w16632 & w20016 ) | ( w20015 & w20016 ) ;
  assign w20018 = w20014 | w20017 ;
  assign w20019 = w6045 | w18038 ;
  assign w20020 = ( ~w18038 & w20018 ) | ( ~w18038 & w20019 ) | ( w20018 & w20019 ) ;
  assign w20021 = \pi14 ^ w20020 ;
  assign w20022 = w19927 ^ w20021 ;
  assign w20023 = w20013 ^ w20022 ;
  assign w20024 = ( w19751 & w19850 ) | ( w19751 & w19851 ) | ( w19850 & w19851 ) ;
  assign w20025 = w19926 ^ w20024 ;
  assign w20026 = w20023 ^ w20025 ;
  assign w20027 = ~w7673 & w16617 ;
  assign w20028 = w7411 & w16621 ;
  assign w20029 = ( w16617 & ~w20027 ) | ( w16617 & w20028 ) | ( ~w20027 & w20028 ) ;
  assign w20030 = w7944 | w18914 ;
  assign w20031 = w19350 & ~w20029 ;
  assign w20032 = ( w7414 & w20029 ) | ( w7414 & ~w20031 ) | ( w20029 & ~w20031 ) ;
  assign w20033 = ( ~w18914 & w20030 ) | ( ~w18914 & w20032 ) | ( w20030 & w20032 ) ;
  assign w20034 = \pi08 ^ w20033 ;
  assign w20035 = w19918 ^ w20034 ;
  assign w20036 = w20026 ^ w20035 ;
  assign w20037 = ( w19742 & w19863 ) | ( w19742 & w19864 ) | ( w19863 & w19864 ) ;
  assign w20038 = w19917 ^ w20037 ;
  assign w20039 = w20036 ^ w20038 ;
  assign w20040 = w6462 & w10431 ;
  assign w20041 = w10736 ^ w20040 ;
  assign w20042 = ~w16009 & w20041 ;
  assign w20043 = w10431 & ~w10736 ;
  assign w20044 = ~w10402 & w20043 ;
  assign w20045 = ~\pi31 & w20044 ;
  assign w20046 = \pi30 ^ w20045 ;
  assign w20047 = ( \pi29 & \pi30 ) | ( \pi29 & \pi31 ) | ( \pi30 & \pi31 ) ;
  assign w20048 = ~w20046 & w20047 ;
  assign w20049 = w20042 | w20048 ;
  assign w20050 = ( w10402 & ~w10431 ) | ( w10402 & w10736 ) | ( ~w10431 & w10736 ) ;
  assign w20051 = ( w6462 & ~w10431 ) | ( w6462 & w10736 ) | ( ~w10431 & w10736 ) ;
  assign w20052 = ~w20050 & w20051 ;
  assign w20053 = \pi30 ^ \pi31 ;
  assign w20054 = \pi31 & w20043 ;
  assign w20055 = ( w10402 & w20053 ) | ( w10402 & ~w20054 ) | ( w20053 & ~w20054 ) ;
  assign w20056 = w20053 & w20055 ;
  assign w20057 = ( \pi29 & ~w20049 ) | ( \pi29 & w20056 ) | ( ~w20049 & w20056 ) ;
  assign w20058 = ( w20049 & ~w20052 ) | ( w20049 & w20057 ) | ( ~w20052 & w20057 ) ;
  assign w20059 = ~w20049 & w20058 ;
  assign w20060 = ( w37 & ~w11145 ) | ( w37 & w20059 ) | ( ~w11145 & w20059 ) ;
  assign w20061 = w20059 | w20060 ;
  assign w20062 = ( w10399 & w19690 ) | ( w10399 & ~w19881 ) | ( w19690 & ~w19881 ) ;
  assign w20063 = w20061 ^ w20062 ;
  assign w20064 = w3927 ^ w20063 ;
  assign w20065 = ( w19691 & ~w19877 ) | ( w19691 & w19883 ) | ( ~w19877 & w19883 ) ;
  assign w20066 = ( w19867 & w19868 ) | ( w19867 & w19885 ) | ( w19868 & w19885 ) ;
  assign w20067 = w20064 ^ w20066 ;
  assign w20068 = w20065 ^ w20067 ;
  assign w20069 = ( \pi02 & ~w19887 ) | ( \pi02 & w20068 ) | ( ~w19887 & w20068 ) ;
  assign w20070 = \pi00 ^ w20069 ;
  assign w20071 = ( \pi02 & ~w20068 ) | ( \pi02 & w20070 ) | ( ~w20068 & w20070 ) ;
  assign w20072 = ( \pi02 & w19887 ) | ( \pi02 & ~w20070 ) | ( w19887 & ~w20070 ) ;
  assign w20073 = \pi01 & w20072 ;
  assign w20074 = ( ~\pi00 & w19713 ) | ( ~\pi00 & w20073 ) | ( w19713 & w20073 ) ;
  assign w20075 = ( \pi01 & \pi02 ) | ( \pi01 & ~w20074 ) | ( \pi02 & ~w20074 ) ;
  assign w20076 = ( w20071 & w20073 ) | ( w20071 & ~w20075 ) | ( w20073 & ~w20075 ) ;
  assign w20077 = ( w19529 & w19538 ) | ( w19529 & w19713 ) | ( w19538 & w19713 ) ;
  assign w20078 = ( w19713 & w19887 ) | ( w19713 & w20077 ) | ( w19887 & w20077 ) ;
  assign w20079 = ( w19887 & ~w20068 ) | ( w19887 & w20078 ) | ( ~w20068 & w20078 ) ;
  assign w20080 = w20068 ^ w20078 ;
  assign w20081 = w19887 ^ w20080 ;
  assign w20082 = w8954 & w20081 ;
  assign w20083 = ( w8954 & w20076 ) | ( w8954 & ~w20082 ) | ( w20076 & ~w20082 ) ;
  assign w20084 = w19909 ^ w20083 ;
  assign w20085 = \pi02 ^ w20039 ;
  assign w20086 = w20084 ^ w20085 ;
  assign w20087 = w19904 & ~w20086 ;
  assign w20088 = w19904 ^ w20086 ;
  assign w20089 = ~w20076 & w20081 ;
  assign w20090 = ( w8954 & w20076 ) | ( w8954 & ~w20089 ) | ( w20076 & ~w20089 ) ;
  assign w20091 = \pi02 ^ w20090 ;
  assign w20092 = ( w19909 & ~w20039 ) | ( w19909 & w20091 ) | ( ~w20039 & w20091 ) ;
  assign w20093 = ~w8593 & w19529 ;
  assign w20094 = w8262 & ~w18912 ;
  assign w20095 = ( w19529 & ~w20093 ) | ( w19529 & w20094 ) | ( ~w20093 & w20094 ) ;
  assign w20096 = ~w8263 & w19723 ;
  assign w20097 = w19713 | w20095 ;
  assign w20098 = ( w35 & w20095 ) | ( w35 & w20097 ) | ( w20095 & w20097 ) ;
  assign w20099 = ( w19723 & ~w20096 ) | ( w19723 & w20098 ) | ( ~w20096 & w20098 ) ;
  assign w20100 = \pi05 ^ w20099 ;
  assign w20101 = ( w19918 & ~w20026 ) | ( w19918 & w20034 ) | ( ~w20026 & w20034 ) ;
  assign w20102 = ~w6949 & w16619 ;
  assign w20103 = w6748 & ~w16626 ;
  assign w20104 = ( w16619 & ~w20102 ) | ( w16619 & w20103 ) | ( ~w20102 & w20103 ) ;
  assign w20105 = ~w7154 & w16621 ;
  assign w20106 = w18439 & ~w20104 ;
  assign w20107 = ( w6751 & w20104 ) | ( w6751 & ~w20106 ) | ( w20104 & ~w20106 ) ;
  assign w20108 = ( w16621 & ~w20105 ) | ( w16621 & w20107 ) | ( ~w20105 & w20107 ) ;
  assign w20109 = \pi11 ^ w20108 ;
  assign w20110 = ( w19927 & ~w20013 ) | ( w19927 & w20021 ) | ( ~w20013 & w20021 ) ;
  assign w20111 = ~w5710 & w16636 ;
  assign w20112 = w5494 & ~w16638 ;
  assign w20113 = ( w16636 & ~w20111 ) | ( w16636 & w20112 ) | ( ~w20111 & w20112 ) ;
  assign w20114 = w5948 | w16634 ;
  assign w20115 = w16742 & ~w20113 ;
  assign w20116 = ( w5497 & w20113 ) | ( w5497 & ~w20115 ) | ( w20113 & ~w20115 ) ;
  assign w20117 = ( ~w16634 & w20114 ) | ( ~w16634 & w20116 ) | ( w20114 & w20116 ) ;
  assign w20118 = \pi17 ^ w20117 ;
  assign w20119 = ( w19936 & ~w20000 ) | ( w19936 & w20008 ) | ( ~w20000 & w20008 ) ;
  assign w20120 = w4651 | w16648 ;
  assign w20121 = w4606 & ~w16650 ;
  assign w20122 = ( ~w16648 & w20120 ) | ( ~w16648 & w20121 ) | ( w20120 & w20121 ) ;
  assign w20123 = w4706 | w16646 ;
  assign w20124 = w17476 & ~w20122 ;
  assign w20125 = ( w4609 & w20122 ) | ( w4609 & ~w20124 ) | ( w20122 & ~w20124 ) ;
  assign w20126 = ( ~w16646 & w20123 ) | ( ~w16646 & w20125 ) | ( w20123 & w20125 ) ;
  assign w20127 = \pi23 ^ w20126 ;
  assign w20128 = ( w19945 & ~w19987 ) | ( w19945 & w19995 ) | ( ~w19987 & w19995 ) ;
  assign w20129 = ( w19946 & ~w19977 ) | ( w19946 & w19985 ) | ( ~w19977 & w19985 ) ;
  assign w20130 = ( w19947 & ~w19967 ) | ( w19947 & w19975 ) | ( ~w19967 & w19975 ) ;
  assign w20131 = w63 | w3659 ;
  assign w20132 = ( ~w63 & w199 ) | ( ~w63 & w1460 ) | ( w199 & w1460 ) ;
  assign w20133 = w20131 | w20132 ;
  assign w20134 = w203 | w390 ;
  assign w20135 = w1616 | w20134 ;
  assign w20136 = ( w76 & ~w1616 ) | ( w76 & w20133 ) | ( ~w1616 & w20133 ) ;
  assign w20137 = w20135 | w20136 ;
  assign w20138 = ( w180 & w490 ) | ( w180 & ~w802 ) | ( w490 & ~w802 ) ;
  assign w20139 = w136 | w20137 ;
  assign w20140 = ( ~w136 & w802 ) | ( ~w136 & w901 ) | ( w802 & w901 ) ;
  assign w20141 = w20139 | w20140 ;
  assign w20142 = w20138 | w20141 ;
  assign w20143 = w568 | w2170 ;
  assign w20144 = w1268 | w20143 ;
  assign w20145 = ( w1165 & ~w1268 ) | ( w1165 & w1729 ) | ( ~w1268 & w1729 ) ;
  assign w20146 = w20144 | w20145 ;
  assign w20147 = w449 | w524 ;
  assign w20148 = w254 | w20147 ;
  assign w20149 = ( ~w254 & w268 ) | ( ~w254 & w20146 ) | ( w268 & w20146 ) ;
  assign w20150 = w20148 | w20149 ;
  assign w20151 = ~w1759 & w2082 ;
  assign w20152 = ~w4489 & w20151 ;
  assign w20153 = ( w3212 & ~w4489 ) | ( w3212 & w20150 ) | ( ~w4489 & w20150 ) ;
  assign w20154 = w20152 & ~w20153 ;
  assign w20155 = w572 | w998 ;
  assign w20156 = w20142 | w20155 ;
  assign w20157 = ( ~w87 & w20142 ) | ( ~w87 & w20154 ) | ( w20142 & w20154 ) ;
  assign w20158 = ~w20156 & w20157 ;
  assign w20159 = ( w223 & w314 ) | ( w223 & ~w423 ) | ( w314 & ~w423 ) ;
  assign w20160 = ~w74 & w20158 ;
  assign w20161 = ( ~w74 & w423 ) | ( ~w74 & w606 ) | ( w423 & w606 ) ;
  assign w20162 = w20160 & ~w20161 ;
  assign w20163 = ~w20159 & w20162 ;
  assign w20164 = ~w37 & w16960 ;
  assign w20165 = w3098 & w16675 ;
  assign w20166 = ( w16960 & ~w20164 ) | ( w16960 & w20165 ) | ( ~w20164 & w20165 ) ;
  assign w20167 = ( \pi29 & \pi30 ) | ( \pi29 & w16665 ) | ( \pi30 & w16665 ) ;
  assign w20168 = \pi31 | w20167 ;
  assign w20169 = ( \pi29 & ~\pi30 ) | ( \pi29 & w16670 ) | ( ~\pi30 & w16670 ) ;
  assign w20170 = ( \pi29 & \pi31 ) | ( \pi29 & ~w20169 ) | ( \pi31 & ~w20169 ) ;
  assign w20171 = ( w20166 & w20168 ) | ( w20166 & ~w20170 ) | ( w20168 & ~w20170 ) ;
  assign w20172 = w20130 ^ w20171 ;
  assign w20173 = w20163 ^ w20172 ;
  assign w20174 = w3549 & ~w16658 ;
  assign w20175 = ( w3717 & w16660 ) | ( w3717 & w20174 ) | ( w16660 & w20174 ) ;
  assign w20176 = w3649 | w20175 ;
  assign w20177 = ( ~w16662 & w20175 ) | ( ~w16662 & w20176 ) | ( w20175 & w20176 ) ;
  assign w20178 = w20174 | w20177 ;
  assign w20179 = w3448 | w17065 ;
  assign w20180 = ( ~w17065 & w20178 ) | ( ~w17065 & w20179 ) | ( w20178 & w20179 ) ;
  assign w20181 = \pi29 ^ w20180 ;
  assign w20182 = w20129 ^ w20181 ;
  assign w20183 = w20173 ^ w20182 ;
  assign w20184 = w3964 & ~w16652 ;
  assign w20185 = ( w4143 & w16654 ) | ( w4143 & w20184 ) | ( w16654 & w20184 ) ;
  assign w20186 = w4052 | w20185 ;
  assign w20187 = ( ~w16656 & w20185 ) | ( ~w16656 & w20186 ) | ( w20185 & w20186 ) ;
  assign w20188 = w20184 | w20187 ;
  assign w20189 = ~w4147 & w17293 ;
  assign w20190 = ( w17293 & w20188 ) | ( w17293 & ~w20189 ) | ( w20188 & ~w20189 ) ;
  assign w20191 = \pi26 ^ w20190 ;
  assign w20192 = w20128 ^ w20191 ;
  assign w20193 = w20183 ^ w20192 ;
  assign w20194 = ( w19944 & ~w19997 ) | ( w19944 & w19998 ) | ( ~w19997 & w19998 ) ;
  assign w20195 = w20127 ^ w20194 ;
  assign w20196 = w20193 ^ w20195 ;
  assign w20197 = w4905 & ~w16644 ;
  assign w20198 = ( w5395 & w16640 ) | ( w5395 & w20197 ) | ( w16640 & w20197 ) ;
  assign w20199 = w5343 | w20198 ;
  assign w20200 = ( w16642 & w20198 ) | ( w16642 & w20199 ) | ( w20198 & w20199 ) ;
  assign w20201 = w20197 | w20200 ;
  assign w20202 = w4908 | w17760 ;
  assign w20203 = ( ~w17760 & w20201 ) | ( ~w17760 & w20202 ) | ( w20201 & w20202 ) ;
  assign w20204 = \pi20 ^ w20203 ;
  assign w20205 = w20119 ^ w20204 ;
  assign w20206 = w20196 ^ w20205 ;
  assign w20207 = ( w19935 & ~w20010 ) | ( w19935 & w20011 ) | ( ~w20010 & w20011 ) ;
  assign w20208 = w20118 ^ w20207 ;
  assign w20209 = w20206 ^ w20208 ;
  assign w20210 = w6048 & w16632 ;
  assign w20211 = ( w6637 & ~w16628 ) | ( w6637 & w20210 ) | ( ~w16628 & w20210 ) ;
  assign w20212 = w6549 | w20211 ;
  assign w20213 = ( ~w16630 & w20211 ) | ( ~w16630 & w20212 ) | ( w20211 & w20212 ) ;
  assign w20214 = w20210 | w20213 ;
  assign w20215 = ~w6045 & w18026 ;
  assign w20216 = ( w18026 & w20214 ) | ( w18026 & ~w20215 ) | ( w20214 & ~w20215 ) ;
  assign w20217 = \pi14 ^ w20216 ;
  assign w20218 = w20110 ^ w20217 ;
  assign w20219 = w20209 ^ w20218 ;
  assign w20220 = ( w19926 & ~w20023 ) | ( w19926 & w20024 ) | ( ~w20023 & w20024 ) ;
  assign w20221 = w20109 ^ w20220 ;
  assign w20222 = w20219 ^ w20221 ;
  assign w20223 = w7673 | w18914 ;
  assign w20224 = w7411 & w16617 ;
  assign w20225 = ( ~w18914 & w20223 ) | ( ~w18914 & w20224 ) | ( w20223 & w20224 ) ;
  assign w20226 = ~w7944 & w18916 ;
  assign w20227 = w19366 & ~w20225 ;
  assign w20228 = ( w7414 & w20225 ) | ( w7414 & ~w20227 ) | ( w20225 & ~w20227 ) ;
  assign w20229 = ( w18916 & ~w20226 ) | ( w18916 & w20228 ) | ( ~w20226 & w20228 ) ;
  assign w20230 = \pi08 ^ w20229 ;
  assign w20231 = w20101 ^ w20230 ;
  assign w20232 = w20222 ^ w20231 ;
  assign w20233 = ( w19917 & ~w20036 ) | ( w19917 & w20037 ) | ( ~w20036 & w20037 ) ;
  assign w20234 = w20100 ^ w20233 ;
  assign w20235 = w20232 ^ w20234 ;
  assign w20236 = \pi31 ^ w10738 ;
  assign w20237 = ( \pi29 & \pi30 ) | ( \pi29 & w11146 ) | ( \pi30 & w11146 ) ;
  assign w20238 = ( w10738 & w20236 ) | ( w10738 & w20237 ) | ( w20236 & w20237 ) ;
  assign w20239 = ( \pi29 & w10738 ) | ( \pi29 & w11138 ) | ( w10738 & w11138 ) ;
  assign w20240 = w20236 & ~w20239 ;
  assign w20241 = ( \pi29 & ~\pi30 ) | ( \pi29 & w20240 ) | ( ~\pi30 & w20240 ) ;
  assign w20242 = ( \pi30 & ~w20238 ) | ( \pi30 & w20241 ) | ( ~w20238 & w20241 ) ;
  assign w20243 = ( w3927 & w20061 ) | ( w3927 & w20062 ) | ( w20061 & w20062 ) ;
  assign w20244 = ( w20064 & ~w20065 ) | ( w20064 & w20066 ) | ( ~w20065 & w20066 ) ;
  assign w20245 = w3927 ^ w20242 ;
  assign w20246 = w20244 ^ w20245 ;
  assign w20247 = w20243 ^ w20246 ;
  assign w20248 = ( \pi02 & w20068 ) | ( \pi02 & ~w20247 ) | ( w20068 & ~w20247 ) ;
  assign w20249 = \pi00 ^ w20248 ;
  assign w20250 = ( \pi02 & w20247 ) | ( \pi02 & w20249 ) | ( w20247 & w20249 ) ;
  assign w20251 = ( ~\pi02 & w20068 ) | ( ~\pi02 & w20249 ) | ( w20068 & w20249 ) ;
  assign w20252 = \pi01 & ~w20251 ;
  assign w20253 = ( ~\pi00 & w19887 ) | ( ~\pi00 & w20252 ) | ( w19887 & w20252 ) ;
  assign w20254 = ( \pi01 & \pi02 ) | ( \pi01 & ~w20253 ) | ( \pi02 & ~w20253 ) ;
  assign w20255 = ( w20250 & w20252 ) | ( w20250 & ~w20254 ) | ( w20252 & ~w20254 ) ;
  assign w20256 = w20079 ^ w20247 ;
  assign w20257 = w20068 ^ w20256 ;
  assign w20258 = w8954 & w20257 ;
  assign w20259 = ( w8954 & w20255 ) | ( w8954 & ~w20258 ) | ( w20255 & ~w20258 ) ;
  assign w20260 = w20092 ^ w20259 ;
  assign w20261 = \pi02 ^ w20235 ;
  assign w20262 = w20260 ^ w20261 ;
  assign w20263 = w20087 & ~w20262 ;
  assign w20264 = w20087 ^ w20262 ;
  assign w20265 = ~w20255 & w20257 ;
  assign w20266 = ( w8954 & w20255 ) | ( w8954 & ~w20265 ) | ( w20255 & ~w20265 ) ;
  assign w20267 = \pi02 ^ w20266 ;
  assign w20268 = ( w20092 & ~w20235 ) | ( w20092 & w20267 ) | ( ~w20235 & w20267 ) ;
  assign w20269 = ~w8593 & w19713 ;
  assign w20270 = w8262 & w19529 ;
  assign w20271 = ( w19713 & ~w20269 ) | ( w19713 & w20270 ) | ( ~w20269 & w20270 ) ;
  assign w20272 = ~w8263 & w19898 ;
  assign w20273 = w19887 | w20271 ;
  assign w20274 = ( w35 & w20271 ) | ( w35 & w20273 ) | ( w20271 & w20273 ) ;
  assign w20275 = ( w19898 & ~w20272 ) | ( w19898 & w20274 ) | ( ~w20272 & w20274 ) ;
  assign w20276 = \pi05 ^ w20275 ;
  assign w20277 = ( w20101 & ~w20222 ) | ( w20101 & w20230 ) | ( ~w20222 & w20230 ) ;
  assign w20278 = ~w6949 & w16621 ;
  assign w20279 = w6748 & w16619 ;
  assign w20280 = ( w16621 & ~w20278 ) | ( w16621 & w20279 ) | ( ~w20278 & w20279 ) ;
  assign w20281 = ~w7154 & w16617 ;
  assign w20282 = w16732 | w20280 ;
  assign w20283 = ( w6751 & w20280 ) | ( w6751 & w20282 ) | ( w20280 & w20282 ) ;
  assign w20284 = ( w16617 & ~w20281 ) | ( w16617 & w20283 ) | ( ~w20281 & w20283 ) ;
  assign w20285 = \pi11 ^ w20284 ;
  assign w20286 = ( w20110 & ~w20209 ) | ( w20110 & w20217 ) | ( ~w20209 & w20217 ) ;
  assign w20287 = w5710 | w16634 ;
  assign w20288 = w5494 & w16636 ;
  assign w20289 = ( ~w16634 & w20287 ) | ( ~w16634 & w20288 ) | ( w20287 & w20288 ) ;
  assign w20290 = ~w5948 & w16632 ;
  assign w20291 = w18051 & ~w20289 ;
  assign w20292 = ( w5497 & w20289 ) | ( w5497 & ~w20291 ) | ( w20289 & ~w20291 ) ;
  assign w20293 = ( w16632 & ~w20290 ) | ( w16632 & w20292 ) | ( ~w20290 & w20292 ) ;
  assign w20294 = \pi17 ^ w20293 ;
  assign w20295 = ( w20119 & ~w20196 ) | ( w20119 & w20204 ) | ( ~w20196 & w20204 ) ;
  assign w20296 = w4651 | w16646 ;
  assign w20297 = w4606 & ~w16648 ;
  assign w20298 = ( ~w16646 & w20296 ) | ( ~w16646 & w20297 ) | ( w20296 & w20297 ) ;
  assign w20299 = w4706 | w16644 ;
  assign w20300 = w17468 & ~w20298 ;
  assign w20301 = ( w4609 & w20298 ) | ( w4609 & ~w20300 ) | ( w20298 & ~w20300 ) ;
  assign w20302 = ( ~w16644 & w20299 ) | ( ~w16644 & w20301 ) | ( w20299 & w20301 ) ;
  assign w20303 = \pi23 ^ w20302 ;
  assign w20304 = ( w20128 & ~w20183 ) | ( w20128 & w20191 ) | ( ~w20183 & w20191 ) ;
  assign w20305 = ( w20129 & ~w20173 ) | ( w20129 & w20181 ) | ( ~w20173 & w20181 ) ;
  assign w20306 = ( w20130 & ~w20163 ) | ( w20130 & w20171 ) | ( ~w20163 & w20171 ) ;
  assign w20307 = w3697 | w12586 ;
  assign w20308 = ( w181 & ~w3697 ) | ( w181 & w9881 ) | ( ~w3697 & w9881 ) ;
  assign w20309 = w20307 | w20308 ;
  assign w20310 = ( ~w1069 & w3741 ) | ( ~w1069 & w20309 ) | ( w3741 & w20309 ) ;
  assign w20311 = ~w5255 & w12725 ;
  assign w20312 = ( w466 & w1069 ) | ( w466 & w12725 ) | ( w1069 & w12725 ) ;
  assign w20313 = w20311 & ~w20312 ;
  assign w20314 = ~w20310 & w20313 ;
  assign w20315 = ( w143 & w220 ) | ( w143 & ~w362 ) | ( w220 & ~w362 ) ;
  assign w20316 = ~w76 & w20314 ;
  assign w20317 = ( ~w76 & w362 ) | ( ~w76 & w605 ) | ( w362 & w605 ) ;
  assign w20318 = w20316 & ~w20317 ;
  assign w20319 = ~w20315 & w20318 ;
  assign w20320 = ( w131 & w198 ) | ( w131 & ~w227 ) | ( w198 & ~w227 ) ;
  assign w20321 = ~w128 & w20319 ;
  assign w20322 = ( ~w128 & w227 ) | ( ~w128 & w492 ) | ( w227 & w492 ) ;
  assign w20323 = w20321 & ~w20322 ;
  assign w20324 = ~w20320 & w20323 ;
  assign w20325 = w37 | w16762 ;
  assign w20326 = w3098 & w16670 ;
  assign w20327 = ( ~w16762 & w20325 ) | ( ~w16762 & w20326 ) | ( w20325 & w20326 ) ;
  assign w20328 = ( \pi29 & \pi30 ) | ( \pi29 & ~w16662 ) | ( \pi30 & ~w16662 ) ;
  assign w20329 = \pi31 | w20328 ;
  assign w20330 = ( \pi29 & ~\pi30 ) | ( \pi29 & w16665 ) | ( ~\pi30 & w16665 ) ;
  assign w20331 = ( \pi29 & \pi31 ) | ( \pi29 & ~w20330 ) | ( \pi31 & ~w20330 ) ;
  assign w20332 = ( w20327 & w20329 ) | ( w20327 & ~w20331 ) | ( w20329 & ~w20331 ) ;
  assign w20333 = w20306 ^ w20332 ;
  assign w20334 = w20324 ^ w20333 ;
  assign w20335 = w3549 & ~w16656 ;
  assign w20336 = ( w3717 & ~w16658 ) | ( w3717 & w20335 ) | ( ~w16658 & w20335 ) ;
  assign w20337 = w3649 | w20336 ;
  assign w20338 = ( w16660 & w20336 ) | ( w16660 & w20337 ) | ( w20336 & w20337 ) ;
  assign w20339 = w20335 | w20338 ;
  assign w20340 = ~w3448 & w17057 ;
  assign w20341 = ( w17057 & w20339 ) | ( w17057 & ~w20340 ) | ( w20339 & ~w20340 ) ;
  assign w20342 = \pi29 ^ w20341 ;
  assign w20343 = w20305 ^ w20342 ;
  assign w20344 = w20334 ^ w20343 ;
  assign w20345 = w3964 & ~w16650 ;
  assign w20346 = ( w4143 & ~w16652 ) | ( w4143 & w20345 ) | ( ~w16652 & w20345 ) ;
  assign w20347 = w4052 | w20346 ;
  assign w20348 = ( w16654 & w20346 ) | ( w16654 & w20347 ) | ( w20346 & w20347 ) ;
  assign w20349 = w20345 | w20348 ;
  assign w20350 = w4147 | w17277 ;
  assign w20351 = ( ~w17277 & w20349 ) | ( ~w17277 & w20350 ) | ( w20349 & w20350 ) ;
  assign w20352 = \pi26 ^ w20351 ;
  assign w20353 = w20304 ^ w20352 ;
  assign w20354 = w20344 ^ w20353 ;
  assign w20355 = ( w20127 & ~w20193 ) | ( w20127 & w20194 ) | ( ~w20193 & w20194 ) ;
  assign w20356 = w20303 ^ w20355 ;
  assign w20357 = w20354 ^ w20356 ;
  assign w20358 = w4905 & w16642 ;
  assign w20359 = ( w5395 & ~w16638 ) | ( w5395 & w20358 ) | ( ~w16638 & w20358 ) ;
  assign w20360 = w5343 | w20359 ;
  assign w20361 = ( w16640 & w20359 ) | ( w16640 & w20360 ) | ( w20359 & w20360 ) ;
  assign w20362 = w20358 | w20361 ;
  assign w20363 = w4908 | w17783 ;
  assign w20364 = ( ~w17783 & w20362 ) | ( ~w17783 & w20363 ) | ( w20362 & w20363 ) ;
  assign w20365 = \pi20 ^ w20364 ;
  assign w20366 = w20295 ^ w20365 ;
  assign w20367 = w20357 ^ w20366 ;
  assign w20368 = ( w20118 & ~w20206 ) | ( w20118 & w20207 ) | ( ~w20206 & w20207 ) ;
  assign w20369 = w20294 ^ w20368 ;
  assign w20370 = w20367 ^ w20369 ;
  assign w20371 = w6048 & ~w16630 ;
  assign w20372 = ( w6637 & ~w16626 ) | ( w6637 & w20371 ) | ( ~w16626 & w20371 ) ;
  assign w20373 = w6549 | w20372 ;
  assign w20374 = ( ~w16628 & w20372 ) | ( ~w16628 & w20373 ) | ( w20372 & w20373 ) ;
  assign w20375 = w20371 | w20374 ;
  assign w20376 = w6045 | w18429 ;
  assign w20377 = ( ~w18429 & w20375 ) | ( ~w18429 & w20376 ) | ( w20375 & w20376 ) ;
  assign w20378 = \pi14 ^ w20377 ;
  assign w20379 = w20286 ^ w20378 ;
  assign w20380 = w20370 ^ w20379 ;
  assign w20381 = ( w20109 & ~w20219 ) | ( w20109 & w20220 ) | ( ~w20219 & w20220 ) ;
  assign w20382 = w20285 ^ w20381 ;
  assign w20383 = w20380 ^ w20382 ;
  assign w20384 = ~w7673 & w18916 ;
  assign w20385 = w7411 & ~w18914 ;
  assign w20386 = ( w18916 & ~w20384 ) | ( w18916 & w20385 ) | ( ~w20384 & w20385 ) ;
  assign w20387 = w7944 | w18912 ;
  assign w20388 = w18929 & ~w20386 ;
  assign w20389 = ( w7414 & w20386 ) | ( w7414 & ~w20388 ) | ( w20386 & ~w20388 ) ;
  assign w20390 = ( ~w18912 & w20387 ) | ( ~w18912 & w20389 ) | ( w20387 & w20389 ) ;
  assign w20391 = \pi08 ^ w20390 ;
  assign w20392 = w20277 ^ w20391 ;
  assign w20393 = w20383 ^ w20392 ;
  assign w20394 = ( w20100 & ~w20232 ) | ( w20100 & w20233 ) | ( ~w20232 & w20233 ) ;
  assign w20395 = w20276 ^ w20394 ;
  assign w20396 = w20393 ^ w20395 ;
  assign w20397 = ~\pi30 & \pi31 ;
  assign w20398 = ( \pi29 & \pi30 ) | ( \pi29 & ~w20397 ) | ( \pi30 & ~w20397 ) ;
  assign w20399 = ( ~w10738 & w20397 ) | ( ~w10738 & w20398 ) | ( w20397 & w20398 ) ;
  assign w20400 = w20243 ^ w20244 ;
  assign w20401 = ( w20243 & w20244 ) | ( w20243 & w20400 ) | ( w20244 & w20400 ) ;
  assign w20402 = w20399 ^ w20401 ;
  assign w20403 = ( w3927 & ~w20242 ) | ( w3927 & w20400 ) | ( ~w20242 & w20400 ) ;
  assign w20404 = w20402 ^ w20403 ;
  assign w20405 = ( ~\pi02 & w20247 ) | ( ~\pi02 & w20404 ) | ( w20247 & w20404 ) ;
  assign w20406 = \pi00 ^ w20405 ;
  assign w20407 = ( \pi02 & w20404 ) | ( \pi02 & ~w20406 ) | ( w20404 & ~w20406 ) ;
  assign w20408 = ( \pi02 & w20247 ) | ( \pi02 & w20406 ) | ( w20247 & w20406 ) ;
  assign w20409 = \pi01 & w20408 ;
  assign w20410 = ( \pi00 & w20068 ) | ( \pi00 & ~w20409 ) | ( w20068 & ~w20409 ) ;
  assign w20411 = ( \pi01 & \pi02 ) | ( \pi01 & w20410 ) | ( \pi02 & w20410 ) ;
  assign w20412 = ( w20407 & w20409 ) | ( w20407 & ~w20411 ) | ( w20409 & ~w20411 ) ;
  assign w20413 = ( w20079 & w20247 ) | ( w20079 & w20404 ) | ( w20247 & w20404 ) ;
  assign w20414 = ( ~w20068 & w20247 ) | ( ~w20068 & w20413 ) | ( w20247 & w20413 ) ;
  assign w20415 = ( ~w20068 & w20079 ) | ( ~w20068 & w20247 ) | ( w20079 & w20247 ) ;
  assign w20416 = w20247 ^ w20415 ;
  assign w20417 = w20404 ^ w20416 ;
  assign w20418 = w8954 & ~w20417 ;
  assign w20419 = ( w8954 & w20412 ) | ( w8954 & ~w20418 ) | ( w20412 & ~w20418 ) ;
  assign w20420 = w20268 ^ w20419 ;
  assign w20421 = \pi02 ^ w20396 ;
  assign w20422 = w20420 ^ w20421 ;
  assign w20423 = w20263 & ~w20422 ;
  assign w20424 = w20263 ^ w20422 ;
  assign w20425 = ~w8593 & w19887 ;
  assign w20426 = w8262 & w19713 ;
  assign w20427 = ( w19887 & ~w20425 ) | ( w19887 & w20426 ) | ( ~w20425 & w20426 ) ;
  assign w20428 = w8263 | w20081 ;
  assign w20429 = w20068 & ~w20427 ;
  assign w20430 = ( w35 & w20427 ) | ( w35 & ~w20429 ) | ( w20427 & ~w20429 ) ;
  assign w20431 = ( ~w20081 & w20428 ) | ( ~w20081 & w20430 ) | ( w20428 & w20430 ) ;
  assign w20432 = \pi05 ^ w20431 ;
  assign w20433 = ( w20277 & ~w20383 ) | ( w20277 & w20391 ) | ( ~w20383 & w20391 ) ;
  assign w20434 = ~w6949 & w16617 ;
  assign w20435 = w6748 & w16621 ;
  assign w20436 = ( w16617 & ~w20434 ) | ( w16617 & w20435 ) | ( ~w20434 & w20435 ) ;
  assign w20437 = w7154 | w18914 ;
  assign w20438 = w19350 & ~w20436 ;
  assign w20439 = ( w6751 & w20436 ) | ( w6751 & ~w20438 ) | ( w20436 & ~w20438 ) ;
  assign w20440 = ( ~w18914 & w20437 ) | ( ~w18914 & w20439 ) | ( w20437 & w20439 ) ;
  assign w20441 = \pi11 ^ w20440 ;
  assign w20442 = ( w20286 & ~w20370 ) | ( w20286 & w20378 ) | ( ~w20370 & w20378 ) ;
  assign w20443 = ~w5710 & w16632 ;
  assign w20444 = w5494 & ~w16634 ;
  assign w20445 = ( w16632 & ~w20443 ) | ( w16632 & w20444 ) | ( ~w20443 & w20444 ) ;
  assign w20446 = w5948 | w16630 ;
  assign w20447 = w18038 & ~w20445 ;
  assign w20448 = ( w5497 & w20445 ) | ( w5497 & ~w20447 ) | ( w20445 & ~w20447 ) ;
  assign w20449 = ( ~w16630 & w20446 ) | ( ~w16630 & w20448 ) | ( w20446 & w20448 ) ;
  assign w20450 = \pi17 ^ w20449 ;
  assign w20451 = ( w20295 & ~w20357 ) | ( w20295 & w20365 ) | ( ~w20357 & w20365 ) ;
  assign w20452 = w4651 | w16644 ;
  assign w20453 = w4606 & ~w16646 ;
  assign w20454 = ( ~w16644 & w20452 ) | ( ~w16644 & w20453 ) | ( w20452 & w20453 ) ;
  assign w20455 = ~w4706 & w16642 ;
  assign w20456 = w17455 | w20454 ;
  assign w20457 = ( w4609 & w20454 ) | ( w4609 & w20456 ) | ( w20454 & w20456 ) ;
  assign w20458 = ( w16642 & ~w20455 ) | ( w16642 & w20457 ) | ( ~w20455 & w20457 ) ;
  assign w20459 = \pi23 ^ w20458 ;
  assign w20460 = ( w20304 & ~w20344 ) | ( w20304 & w20352 ) | ( ~w20344 & w20352 ) ;
  assign w20461 = ( w20305 & ~w20334 ) | ( w20305 & w20342 ) | ( ~w20334 & w20342 ) ;
  assign w20462 = ( w20306 & ~w20324 ) | ( w20306 & w20332 ) | ( ~w20324 & w20332 ) ;
  assign w20463 = w205 | w281 ;
  assign w20464 = w104 | w20463 ;
  assign w20465 = ( ~w104 & w141 ) | ( ~w104 & w1590 ) | ( w141 & w1590 ) ;
  assign w20466 = w20464 | w20465 ;
  assign w20467 = w309 | w569 ;
  assign w20468 = w128 | w20467 ;
  assign w20469 = ( ~w128 & w165 ) | ( ~w128 & w20466 ) | ( w165 & w20466 ) ;
  assign w20470 = w20468 | w20469 ;
  assign w20471 = w279 | w430 ;
  assign w20472 = ( ~w279 & w429 ) | ( ~w279 & w19950 ) | ( w429 & w19950 ) ;
  assign w20473 = w20471 | w20472 ;
  assign w20474 = ( ~w268 & w11635 ) | ( ~w268 & w20473 ) | ( w11635 & w20473 ) ;
  assign w20475 = w4959 | w20470 ;
  assign w20476 = ( w268 & w449 ) | ( w268 & ~w20470 ) | ( w449 & ~w20470 ) ;
  assign w20477 = w20475 | w20476 ;
  assign w20478 = w20474 | w20477 ;
  assign w20479 = w507 | w998 ;
  assign w20480 = w11965 | w20479 ;
  assign w20481 = ( w204 & ~w11965 ) | ( w204 & w20478 ) | ( ~w11965 & w20478 ) ;
  assign w20482 = w20480 | w20481 ;
  assign w20483 = ( w82 & w224 ) | ( w82 & w359 ) | ( w224 & w359 ) ;
  assign w20484 = w2517 | w20482 ;
  assign w20485 = ( w359 & ~w663 ) | ( w359 & w20482 ) | ( ~w663 & w20482 ) ;
  assign w20486 = ~w20484 & w20485 ;
  assign w20487 = ~w20483 & w20486 ;
  assign w20488 = ( w422 & w664 ) | ( w422 & ~w722 ) | ( w664 & ~w722 ) ;
  assign w20489 = ~w59 & w20487 ;
  assign w20490 = ( ~w59 & w722 ) | ( ~w59 & w901 ) | ( w722 & w901 ) ;
  assign w20491 = w20489 & ~w20490 ;
  assign w20492 = ~w20488 & w20491 ;
  assign w20493 = w37 | w17078 ;
  assign w20494 = w3098 & w16665 ;
  assign w20495 = ( ~w17078 & w20493 ) | ( ~w17078 & w20494 ) | ( w20493 & w20494 ) ;
  assign w20496 = ( \pi29 & \pi30 ) | ( \pi29 & w16660 ) | ( \pi30 & w16660 ) ;
  assign w20497 = \pi31 | w20496 ;
  assign w20498 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w16662 ) | ( \pi30 & w16662 ) ;
  assign w20499 = ( \pi29 & \pi31 ) | ( \pi29 & w20498 ) | ( \pi31 & w20498 ) ;
  assign w20500 = ( w20495 & w20497 ) | ( w20495 & ~w20499 ) | ( w20497 & ~w20499 ) ;
  assign w20501 = w20462 ^ w20500 ;
  assign w20502 = w20492 ^ w20501 ;
  assign w20503 = w3549 & w16654 ;
  assign w20504 = ( w3717 & ~w16656 ) | ( w3717 & w20503 ) | ( ~w16656 & w20503 ) ;
  assign w20505 = w3649 | w20504 ;
  assign w20506 = ( ~w16658 & w20504 ) | ( ~w16658 & w20505 ) | ( w20504 & w20505 ) ;
  assign w20507 = w20503 | w20506 ;
  assign w20508 = ~w3448 & w17266 ;
  assign w20509 = ( w17266 & w20507 ) | ( w17266 & ~w20508 ) | ( w20507 & ~w20508 ) ;
  assign w20510 = \pi29 ^ w20509 ;
  assign w20511 = w20461 ^ w20510 ;
  assign w20512 = w20502 ^ w20511 ;
  assign w20513 = w3964 & ~w16648 ;
  assign w20514 = ( w4143 & ~w16650 ) | ( w4143 & w20513 ) | ( ~w16650 & w20513 ) ;
  assign w20515 = w4052 | w20514 ;
  assign w20516 = ( ~w16652 & w20514 ) | ( ~w16652 & w20515 ) | ( w20514 & w20515 ) ;
  assign w20517 = w20513 | w20516 ;
  assign w20518 = w4147 | w16752 ;
  assign w20519 = ( ~w16752 & w20517 ) | ( ~w16752 & w20518 ) | ( w20517 & w20518 ) ;
  assign w20520 = \pi26 ^ w20519 ;
  assign w20521 = w20460 ^ w20520 ;
  assign w20522 = w20512 ^ w20521 ;
  assign w20523 = ( w20303 & ~w20354 ) | ( w20303 & w20355 ) | ( ~w20354 & w20355 ) ;
  assign w20524 = w20459 ^ w20523 ;
  assign w20525 = w20522 ^ w20524 ;
  assign w20526 = w4905 & w16640 ;
  assign w20527 = ( w5395 & w16636 ) | ( w5395 & w20526 ) | ( w16636 & w20526 ) ;
  assign w20528 = w5343 | w20527 ;
  assign w20529 = ( ~w16638 & w20527 ) | ( ~w16638 & w20528 ) | ( w20527 & w20528 ) ;
  assign w20530 = w20526 | w20529 ;
  assign w20531 = w4908 | w17770 ;
  assign w20532 = ( ~w17770 & w20530 ) | ( ~w17770 & w20531 ) | ( w20530 & w20531 ) ;
  assign w20533 = \pi20 ^ w20532 ;
  assign w20534 = w20451 ^ w20533 ;
  assign w20535 = w20525 ^ w20534 ;
  assign w20536 = ( w20294 & ~w20367 ) | ( w20294 & w20368 ) | ( ~w20367 & w20368 ) ;
  assign w20537 = w20450 ^ w20536 ;
  assign w20538 = w20535 ^ w20537 ;
  assign w20539 = w6048 & ~w16628 ;
  assign w20540 = ( w6637 & w16619 ) | ( w6637 & w20539 ) | ( w16619 & w20539 ) ;
  assign w20541 = w6549 | w20540 ;
  assign w20542 = ( ~w16626 & w20540 ) | ( ~w16626 & w20541 ) | ( w20540 & w20541 ) ;
  assign w20543 = w20539 | w20542 ;
  assign w20544 = ~w6045 & w18451 ;
  assign w20545 = ( w18451 & w20543 ) | ( w18451 & ~w20544 ) | ( w20543 & ~w20544 ) ;
  assign w20546 = \pi14 ^ w20545 ;
  assign w20547 = w20442 ^ w20546 ;
  assign w20548 = w20538 ^ w20547 ;
  assign w20549 = ( w20285 & ~w20380 ) | ( w20285 & w20381 ) | ( ~w20380 & w20381 ) ;
  assign w20550 = w20441 ^ w20549 ;
  assign w20551 = w20548 ^ w20550 ;
  assign w20552 = w7673 | w18912 ;
  assign w20553 = w7411 & w18916 ;
  assign w20554 = ( ~w18912 & w20552 ) | ( ~w18912 & w20553 ) | ( w20552 & w20553 ) ;
  assign w20555 = ~w7944 & w19529 ;
  assign w20556 = w19540 & ~w20554 ;
  assign w20557 = ( w7414 & w20554 ) | ( w7414 & ~w20556 ) | ( w20554 & ~w20556 ) ;
  assign w20558 = ( w19529 & ~w20555 ) | ( w19529 & w20557 ) | ( ~w20555 & w20557 ) ;
  assign w20559 = \pi08 ^ w20558 ;
  assign w20560 = w20433 ^ w20559 ;
  assign w20561 = w20551 ^ w20560 ;
  assign w20562 = \pi00 & ~\pi02 ;
  assign w20563 = ( \pi01 & w20404 ) | ( \pi01 & w20562 ) | ( w20404 & w20562 ) ;
  assign w20564 = ( \pi01 & \pi02 ) | ( \pi01 & w20562 ) | ( \pi02 & w20562 ) ;
  assign w20565 = \pi00 ^ w20414 ;
  assign w20566 = ( w20247 & w20414 ) | ( w20247 & ~w20565 ) | ( w20414 & ~w20565 ) ;
  assign w20567 = ( \pi02 & w20564 ) | ( \pi02 & ~w20566 ) | ( w20564 & ~w20566 ) ;
  assign w20568 = w20563 ^ w20567 ;
  assign w20569 = w20432 ^ w20568 ;
  assign w20570 = w20561 ^ w20569 ;
  assign w20571 = ( w20276 & ~w20393 ) | ( w20276 & w20394 ) | ( ~w20393 & w20394 ) ;
  assign w20572 = w20412 | w20417 ;
  assign w20573 = ( w8954 & w20412 ) | ( w8954 & w20572 ) | ( w20412 & w20572 ) ;
  assign w20574 = \pi02 ^ w20573 ;
  assign w20575 = ( w20268 & ~w20396 ) | ( w20268 & w20574 ) | ( ~w20396 & w20574 ) ;
  assign w20576 = w20570 ^ w20575 ;
  assign w20577 = w20571 ^ w20576 ;
  assign w20578 = w20423 & ~w20577 ;
  assign w20579 = w20423 ^ w20577 ;
  assign w20580 = ( w20461 & ~w20502 ) | ( w20461 & w20510 ) | ( ~w20502 & w20510 ) ;
  assign w20581 = ( \pi29 & \pi31 ) | ( \pi29 & w16660 ) | ( \pi31 & w16660 ) ;
  assign w20582 = ( \pi29 & ~\pi30 ) | ( \pi29 & w20581 ) | ( ~\pi30 & w20581 ) ;
  assign w20583 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w20581 ) | ( \pi30 & w20581 ) ;
  assign w20584 = ( \pi29 & w16662 ) | ( \pi29 & ~w20583 ) | ( w16662 & ~w20583 ) ;
  assign w20585 = ( ~w16658 & w20583 ) | ( ~w16658 & w20584 ) | ( w20583 & w20584 ) ;
  assign w20586 = ~\pi31 & w20585 ;
  assign w20587 = ( w20582 & ~w20584 ) | ( w20582 & w20586 ) | ( ~w20584 & w20586 ) ;
  assign w20588 = ( w37 & ~w17065 ) | ( w37 & w20587 ) | ( ~w17065 & w20587 ) ;
  assign w20589 = w20587 | w20588 ;
  assign w20590 = w115 | w1094 ;
  assign w20591 = w1154 | w20590 ;
  assign w20592 = ( ~w1154 & w2536 ) | ( ~w1154 & w6387 ) | ( w2536 & w6387 ) ;
  assign w20593 = w20591 | w20592 ;
  assign w20594 = w2092 | w20593 ;
  assign w20595 = ( w663 & w821 ) | ( w663 & ~w2092 ) | ( w821 & ~w2092 ) ;
  assign w20596 = w20594 | w20595 ;
  assign w20597 = w10944 | w20596 ;
  assign w20598 = ( w1615 & ~w1945 ) | ( w1615 & w10272 ) | ( ~w1945 & w10272 ) ;
  assign w20599 = w3853 | w20597 ;
  assign w20600 = ( w1615 & w1618 ) | ( w1615 & ~w20597 ) | ( w1618 & ~w20597 ) ;
  assign w20601 = w20599 | w20600 ;
  assign w20602 = w20598 & ~w20601 ;
  assign w20603 = ( w625 & ~w860 ) | ( w625 & w1421 ) | ( ~w860 & w1421 ) ;
  assign w20604 = ~w2600 & w20602 ;
  assign w20605 = ( w860 & ~w2600 ) | ( w860 & w4073 ) | ( ~w2600 & w4073 ) ;
  assign w20606 = w20604 & ~w20605 ;
  assign w20607 = ~w20603 & w20606 ;
  assign w20608 = w534 | w605 ;
  assign w20609 = w127 | w20608 ;
  assign w20610 = ( w127 & ~w530 ) | ( w127 & w20607 ) | ( ~w530 & w20607 ) ;
  assign w20611 = ~w20609 & w20610 ;
  assign w20612 = \pi02 ^ w20404 ;
  assign w20613 = ~\pi01 & w20404 ;
  assign w20614 = ( \pi00 & w20612 ) | ( \pi00 & ~w20613 ) | ( w20612 & ~w20613 ) ;
  assign w20615 = w20612 & w20614 ;
  assign w20616 = ( w20589 & ~w20611 ) | ( w20589 & w20615 ) | ( ~w20611 & w20615 ) ;
  assign w20617 = w20589 ^ w20615 ;
  assign w20618 = w20611 ^ w20617 ;
  assign w20619 = ( w20462 & ~w20492 ) | ( w20462 & w20500 ) | ( ~w20492 & w20500 ) ;
  assign w20620 = w3549 & ~w16652 ;
  assign w20621 = ( w3717 & w16654 ) | ( w3717 & w20620 ) | ( w16654 & w20620 ) ;
  assign w20622 = w3649 | w20621 ;
  assign w20623 = ( ~w16656 & w20621 ) | ( ~w16656 & w20622 ) | ( w20621 & w20622 ) ;
  assign w20624 = w20620 | w20623 ;
  assign w20625 = ~w3448 & w17293 ;
  assign w20626 = ( w17293 & w20624 ) | ( w17293 & ~w20625 ) | ( w20624 & ~w20625 ) ;
  assign w20627 = \pi29 ^ w20626 ;
  assign w20628 = w20618 ^ w20627 ;
  assign w20629 = w20619 ^ w20628 ;
  assign w20630 = w4143 | w16648 ;
  assign w20631 = w4052 & ~w16650 ;
  assign w20632 = ( ~w16648 & w20630 ) | ( ~w16648 & w20631 ) | ( w20630 & w20631 ) ;
  assign w20633 = w4147 | w17476 ;
  assign w20634 = w16646 & ~w20632 ;
  assign w20635 = ( w3964 & w20632 ) | ( w3964 & ~w20634 ) | ( w20632 & ~w20634 ) ;
  assign w20636 = ( ~w17476 & w20633 ) | ( ~w17476 & w20635 ) | ( w20633 & w20635 ) ;
  assign w20637 = \pi26 ^ w20636 ;
  assign w20638 = w20629 ^ w20637 ;
  assign w20639 = w20580 ^ w20638 ;
  assign w20640 = ( w20460 & ~w20512 ) | ( w20460 & w20520 ) | ( ~w20512 & w20520 ) ;
  assign w20641 = ~w4651 & w16642 ;
  assign w20642 = w4606 & ~w16644 ;
  assign w20643 = ( w16642 & ~w20641 ) | ( w16642 & w20642 ) | ( ~w20641 & w20642 ) ;
  assign w20644 = ~w4706 & w16640 ;
  assign w20645 = w17760 & ~w20643 ;
  assign w20646 = ( w4609 & w20643 ) | ( w4609 & ~w20645 ) | ( w20643 & ~w20645 ) ;
  assign w20647 = ( w16640 & ~w20644 ) | ( w16640 & w20646 ) | ( ~w20644 & w20646 ) ;
  assign w20648 = \pi23 ^ w20647 ;
  assign w20649 = w20639 ^ w20648 ;
  assign w20650 = w20640 ^ w20649 ;
  assign w20651 = ( w20459 & ~w20522 ) | ( w20459 & w20523 ) | ( ~w20522 & w20523 ) ;
  assign w20652 = ~w5343 & w16636 ;
  assign w20653 = w4905 & ~w16638 ;
  assign w20654 = ( w16636 & ~w20652 ) | ( w16636 & w20653 ) | ( ~w20652 & w20653 ) ;
  assign w20655 = w5395 | w16634 ;
  assign w20656 = w16742 & ~w20654 ;
  assign w20657 = ( w4908 & w20654 ) | ( w4908 & ~w20656 ) | ( w20654 & ~w20656 ) ;
  assign w20658 = ( ~w16634 & w20655 ) | ( ~w16634 & w20657 ) | ( w20655 & w20657 ) ;
  assign w20659 = \pi20 ^ w20658 ;
  assign w20660 = w20650 ^ w20659 ;
  assign w20661 = w20651 ^ w20660 ;
  assign w20662 = ( w20451 & ~w20525 ) | ( w20451 & w20533 ) | ( ~w20525 & w20533 ) ;
  assign w20663 = w5710 | w16630 ;
  assign w20664 = w5494 & w16632 ;
  assign w20665 = ( ~w16630 & w20663 ) | ( ~w16630 & w20664 ) | ( w20663 & w20664 ) ;
  assign w20666 = w5948 | w16628 ;
  assign w20667 = w18026 | w20665 ;
  assign w20668 = ( w5497 & w20665 ) | ( w5497 & w20667 ) | ( w20665 & w20667 ) ;
  assign w20669 = ( ~w16628 & w20666 ) | ( ~w16628 & w20668 ) | ( w20666 & w20668 ) ;
  assign w20670 = \pi17 ^ w20669 ;
  assign w20671 = w20661 ^ w20670 ;
  assign w20672 = w20662 ^ w20671 ;
  assign w20673 = ( w20450 & ~w20535 ) | ( w20450 & w20536 ) | ( ~w20535 & w20536 ) ;
  assign w20674 = ~w6549 & w16619 ;
  assign w20675 = w6048 & ~w16626 ;
  assign w20676 = ( w16619 & ~w20674 ) | ( w16619 & w20675 ) | ( ~w20674 & w20675 ) ;
  assign w20677 = ~w6637 & w16621 ;
  assign w20678 = w18439 & ~w20676 ;
  assign w20679 = ( w6045 & w20676 ) | ( w6045 & ~w20678 ) | ( w20676 & ~w20678 ) ;
  assign w20680 = ( w16621 & ~w20677 ) | ( w16621 & w20679 ) | ( ~w20677 & w20679 ) ;
  assign w20681 = \pi14 ^ w20680 ;
  assign w20682 = w20672 ^ w20681 ;
  assign w20683 = w20673 ^ w20682 ;
  assign w20684 = ( w20442 & ~w20538 ) | ( w20442 & w20546 ) | ( ~w20538 & w20546 ) ;
  assign w20685 = w6949 | w18914 ;
  assign w20686 = w6748 & w16617 ;
  assign w20687 = ( ~w18914 & w20685 ) | ( ~w18914 & w20686 ) | ( w20685 & w20686 ) ;
  assign w20688 = ~w7154 & w18916 ;
  assign w20689 = w19366 & ~w20687 ;
  assign w20690 = ( w6751 & w20687 ) | ( w6751 & ~w20689 ) | ( w20687 & ~w20689 ) ;
  assign w20691 = ( w18916 & ~w20688 ) | ( w18916 & w20690 ) | ( ~w20688 & w20690 ) ;
  assign w20692 = \pi11 ^ w20691 ;
  assign w20693 = w20683 ^ w20692 ;
  assign w20694 = w20684 ^ w20693 ;
  assign w20695 = ( w20441 & ~w20548 ) | ( w20441 & w20549 ) | ( ~w20548 & w20549 ) ;
  assign w20696 = ~w7673 & w19529 ;
  assign w20697 = w7411 & ~w18912 ;
  assign w20698 = ( w19529 & ~w20696 ) | ( w19529 & w20697 ) | ( ~w20696 & w20697 ) ;
  assign w20699 = ~w7944 & w19713 ;
  assign w20700 = w19723 | w20698 ;
  assign w20701 = ( w7414 & w20698 ) | ( w7414 & w20700 ) | ( w20698 & w20700 ) ;
  assign w20702 = ( w19713 & ~w20699 ) | ( w19713 & w20701 ) | ( ~w20699 & w20701 ) ;
  assign w20703 = \pi08 ^ w20702 ;
  assign w20704 = w20694 ^ w20703 ;
  assign w20705 = w20695 ^ w20704 ;
  assign w20706 = ( w20433 & ~w20551 ) | ( w20433 & w20559 ) | ( ~w20551 & w20559 ) ;
  assign w20707 = w8593 | w20068 ;
  assign w20708 = w8262 & w19887 ;
  assign w20709 = ( ~w20068 & w20707 ) | ( ~w20068 & w20708 ) | ( w20707 & w20708 ) ;
  assign w20710 = w8263 | w20257 ;
  assign w20711 = w20247 | w20709 ;
  assign w20712 = ( w35 & w20709 ) | ( w35 & w20711 ) | ( w20709 & w20711 ) ;
  assign w20713 = ( ~w20257 & w20710 ) | ( ~w20257 & w20712 ) | ( w20710 & w20712 ) ;
  assign w20714 = \pi05 ^ w20713 ;
  assign w20715 = w20705 ^ w20714 ;
  assign w20716 = w20706 ^ w20715 ;
  assign w20717 = ( w20432 & ~w20561 ) | ( w20432 & w20568 ) | ( ~w20561 & w20568 ) ;
  assign w20718 = ( ~w20570 & w20571 ) | ( ~w20570 & w20575 ) | ( w20571 & w20575 ) ;
  assign w20719 = w20716 ^ w20718 ;
  assign w20720 = w20717 ^ w20719 ;
  assign w20721 = w20578 & ~w20720 ;
  assign w20722 = w20578 ^ w20720 ;
  assign w20723 = ( w283 & w573 ) | ( w283 & ~w593 ) | ( w573 & ~w593 ) ;
  assign w20724 = w119 | w731 ;
  assign w20725 = ( ~w119 & w593 ) | ( ~w119 & w723 ) | ( w593 & w723 ) ;
  assign w20726 = w20724 | w20725 ;
  assign w20727 = w20723 | w20726 ;
  assign w20728 = w901 | w20727 ;
  assign w20729 = w353 | w390 ;
  assign w20730 = w210 | w20729 ;
  assign w20731 = ( w51 & ~w210 ) | ( w51 & w316 ) | ( ~w210 & w316 ) ;
  assign w20732 = w20730 | w20731 ;
  assign w20733 = w136 | w495 ;
  assign w20734 = w2522 | w20733 ;
  assign w20735 = ( ~w2522 & w20728 ) | ( ~w2522 & w20732 ) | ( w20728 & w20732 ) ;
  assign w20736 = w20734 | w20735 ;
  assign w20737 = ( ~w201 & w1347 ) | ( ~w201 & w1836 ) | ( w1347 & w1836 ) ;
  assign w20738 = w12844 | w20736 ;
  assign w20739 = ( w201 & w221 ) | ( w201 & ~w20736 ) | ( w221 & ~w20736 ) ;
  assign w20740 = w20738 | w20739 ;
  assign w20741 = w20737 | w20740 ;
  assign w20742 = ( ~w311 & w999 ) | ( ~w311 & w2705 ) | ( w999 & w2705 ) ;
  assign w20743 = w2167 | w20741 ;
  assign w20744 = ( w311 & w389 ) | ( w311 & ~w20741 ) | ( w389 & ~w20741 ) ;
  assign w20745 = w20743 | w20744 ;
  assign w20746 = w20742 | w20745 ;
  assign w20747 = w3251 | w10639 ;
  assign w20748 = ( w88 & ~w3251 ) | ( w88 & w20746 ) | ( ~w3251 & w20746 ) ;
  assign w20749 = w20747 | w20748 ;
  assign w20750 = w265 | w673 ;
  assign w20751 = ( ~w265 & w350 ) | ( ~w265 & w20749 ) | ( w350 & w20749 ) ;
  assign w20752 = w20750 | w20751 ;
  assign w20753 = ( w20615 & w20616 ) | ( w20615 & w20752 ) | ( w20616 & w20752 ) ;
  assign w20754 = w20615 ^ w20616 ;
  assign w20755 = w20752 ^ w20754 ;
  assign w20756 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16658 ) | ( \pi31 & ~w16658 ) ;
  assign w20757 = ( \pi29 & ~\pi30 ) | ( \pi29 & w20756 ) | ( ~\pi30 & w20756 ) ;
  assign w20758 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w20756 ) | ( \pi30 & w20756 ) ;
  assign w20759 = ( ~\pi29 & w16660 ) | ( ~\pi29 & w20758 ) | ( w16660 & w20758 ) ;
  assign w20760 = ( w16656 & ~w20758 ) | ( w16656 & w20759 ) | ( ~w20758 & w20759 ) ;
  assign w20761 = \pi31 | w20760 ;
  assign w20762 = ( w20757 & w20759 ) | ( w20757 & ~w20761 ) | ( w20759 & ~w20761 ) ;
  assign w20763 = ( w37 & w17057 ) | ( w37 & w20762 ) | ( w17057 & w20762 ) ;
  assign w20764 = w20762 | w20763 ;
  assign w20765 = ( ~w20618 & w20619 ) | ( ~w20618 & w20627 ) | ( w20619 & w20627 ) ;
  assign w20766 = w20755 ^ w20765 ;
  assign w20767 = w20764 ^ w20766 ;
  assign w20768 = w3717 | w16652 ;
  assign w20769 = w3649 & w16654 ;
  assign w20770 = ( ~w16652 & w20768 ) | ( ~w16652 & w20769 ) | ( w20768 & w20769 ) ;
  assign w20771 = w3549 | w16650 ;
  assign w20772 = w17277 & ~w20770 ;
  assign w20773 = ( w3448 & w20770 ) | ( w3448 & ~w20772 ) | ( w20770 & ~w20772 ) ;
  assign w20774 = ( ~w16650 & w20771 ) | ( ~w16650 & w20773 ) | ( w20771 & w20773 ) ;
  assign w20775 = \pi29 ^ w20774 ;
  assign w20776 = w4143 | w16646 ;
  assign w20777 = w4052 & ~w16648 ;
  assign w20778 = ( ~w16646 & w20776 ) | ( ~w16646 & w20777 ) | ( w20776 & w20777 ) ;
  assign w20779 = w4147 | w17468 ;
  assign w20780 = w16644 & ~w20778 ;
  assign w20781 = ( w3964 & w20778 ) | ( w3964 & ~w20780 ) | ( w20778 & ~w20780 ) ;
  assign w20782 = ( ~w17468 & w20779 ) | ( ~w17468 & w20781 ) | ( w20779 & w20781 ) ;
  assign w20783 = \pi26 ^ w20782 ;
  assign w20784 = w20767 ^ w20783 ;
  assign w20785 = w20775 ^ w20784 ;
  assign w20786 = ( w20580 & ~w20629 ) | ( w20580 & w20637 ) | ( ~w20629 & w20637 ) ;
  assign w20787 = ~w4651 & w16640 ;
  assign w20788 = w4606 & w16642 ;
  assign w20789 = ( w16640 & ~w20787 ) | ( w16640 & w20788 ) | ( ~w20787 & w20788 ) ;
  assign w20790 = w4706 | w16638 ;
  assign w20791 = w17783 & ~w20789 ;
  assign w20792 = ( w4609 & w20789 ) | ( w4609 & ~w20791 ) | ( w20789 & ~w20791 ) ;
  assign w20793 = ( ~w16638 & w20790 ) | ( ~w16638 & w20792 ) | ( w20790 & w20792 ) ;
  assign w20794 = \pi23 ^ w20793 ;
  assign w20795 = w20785 ^ w20786 ;
  assign w20796 = w20794 ^ w20795 ;
  assign w20797 = ( ~w20639 & w20640 ) | ( ~w20639 & w20648 ) | ( w20640 & w20648 ) ;
  assign w20798 = w5343 | w16634 ;
  assign w20799 = w4905 & w16636 ;
  assign w20800 = ( ~w16634 & w20798 ) | ( ~w16634 & w20799 ) | ( w20798 & w20799 ) ;
  assign w20801 = ~w5395 & w16632 ;
  assign w20802 = w18051 & ~w20800 ;
  assign w20803 = ( w4908 & w20800 ) | ( w4908 & ~w20802 ) | ( w20800 & ~w20802 ) ;
  assign w20804 = ( w16632 & ~w20801 ) | ( w16632 & w20803 ) | ( ~w20801 & w20803 ) ;
  assign w20805 = \pi20 ^ w20804 ;
  assign w20806 = w20796 ^ w20797 ;
  assign w20807 = w20805 ^ w20806 ;
  assign w20808 = ( ~w20650 & w20651 ) | ( ~w20650 & w20659 ) | ( w20651 & w20659 ) ;
  assign w20809 = w5710 | w16628 ;
  assign w20810 = w5494 & ~w16630 ;
  assign w20811 = ( ~w16628 & w20809 ) | ( ~w16628 & w20810 ) | ( w20809 & w20810 ) ;
  assign w20812 = w5948 | w16626 ;
  assign w20813 = w18429 & ~w20811 ;
  assign w20814 = ( w5497 & w20811 ) | ( w5497 & ~w20813 ) | ( w20811 & ~w20813 ) ;
  assign w20815 = ( ~w16626 & w20812 ) | ( ~w16626 & w20814 ) | ( w20812 & w20814 ) ;
  assign w20816 = \pi17 ^ w20815 ;
  assign w20817 = w20807 ^ w20808 ;
  assign w20818 = w20816 ^ w20817 ;
  assign w20819 = ( ~w20661 & w20662 ) | ( ~w20661 & w20670 ) | ( w20662 & w20670 ) ;
  assign w20820 = ~w6549 & w16621 ;
  assign w20821 = w6048 & w16619 ;
  assign w20822 = ( w16621 & ~w20820 ) | ( w16621 & w20821 ) | ( ~w20820 & w20821 ) ;
  assign w20823 = ~w6637 & w16617 ;
  assign w20824 = w16732 | w20822 ;
  assign w20825 = ( w6045 & w20822 ) | ( w6045 & w20824 ) | ( w20822 & w20824 ) ;
  assign w20826 = ( w16617 & ~w20823 ) | ( w16617 & w20825 ) | ( ~w20823 & w20825 ) ;
  assign w20827 = \pi14 ^ w20826 ;
  assign w20828 = w20818 ^ w20819 ;
  assign w20829 = w20827 ^ w20828 ;
  assign w20830 = ( ~w20672 & w20673 ) | ( ~w20672 & w20681 ) | ( w20673 & w20681 ) ;
  assign w20831 = ~w6949 & w18916 ;
  assign w20832 = w6748 & ~w18914 ;
  assign w20833 = ( w18916 & ~w20831 ) | ( w18916 & w20832 ) | ( ~w20831 & w20832 ) ;
  assign w20834 = w7154 | w18912 ;
  assign w20835 = w18929 & ~w20833 ;
  assign w20836 = ( w6751 & w20833 ) | ( w6751 & ~w20835 ) | ( w20833 & ~w20835 ) ;
  assign w20837 = ( ~w18912 & w20834 ) | ( ~w18912 & w20836 ) | ( w20834 & w20836 ) ;
  assign w20838 = \pi11 ^ w20837 ;
  assign w20839 = w20829 ^ w20830 ;
  assign w20840 = w20838 ^ w20839 ;
  assign w20841 = ( ~w20683 & w20684 ) | ( ~w20683 & w20692 ) | ( w20684 & w20692 ) ;
  assign w20842 = ~w7673 & w19713 ;
  assign w20843 = w7411 & w19529 ;
  assign w20844 = ( w19713 & ~w20842 ) | ( w19713 & w20843 ) | ( ~w20842 & w20843 ) ;
  assign w20845 = ~w7944 & w19887 ;
  assign w20846 = w19898 | w20844 ;
  assign w20847 = ( w7414 & w20844 ) | ( w7414 & w20846 ) | ( w20844 & w20846 ) ;
  assign w20848 = ( w19887 & ~w20845 ) | ( w19887 & w20847 ) | ( ~w20845 & w20847 ) ;
  assign w20849 = \pi08 ^ w20848 ;
  assign w20850 = w20840 ^ w20841 ;
  assign w20851 = w20849 ^ w20850 ;
  assign w20852 = ( ~w20694 & w20695 ) | ( ~w20694 & w20703 ) | ( w20695 & w20703 ) ;
  assign w20853 = ~w8593 & w20247 ;
  assign w20854 = w8262 & ~w20068 ;
  assign w20855 = ( w20247 & ~w20853 ) | ( w20247 & w20854 ) | ( ~w20853 & w20854 ) ;
  assign w20856 = ~w8263 & w20417 ;
  assign w20857 = w20404 | w20855 ;
  assign w20858 = ( w35 & w20855 ) | ( w35 & w20857 ) | ( w20855 & w20857 ) ;
  assign w20859 = ( w20417 & ~w20856 ) | ( w20417 & w20858 ) | ( ~w20856 & w20858 ) ;
  assign w20860 = \pi05 ^ w20859 ;
  assign w20861 = w20851 ^ w20852 ;
  assign w20862 = w20860 ^ w20861 ;
  assign w20863 = ( ~w20705 & w20706 ) | ( ~w20705 & w20714 ) | ( w20706 & w20714 ) ;
  assign w20864 = ( ~w20716 & w20717 ) | ( ~w20716 & w20718 ) | ( w20717 & w20718 ) ;
  assign w20865 = w20862 ^ w20864 ;
  assign w20866 = w20863 ^ w20865 ;
  assign w20867 = w20721 & w20866 ;
  assign w20868 = w20721 ^ w20866 ;
  assign w20869 = w605 | w889 ;
  assign w20870 = w199 | w20869 ;
  assign w20871 = ( ~w199 & w411 ) | ( ~w199 & w12138 ) | ( w411 & w12138 ) ;
  assign w20872 = w20870 | w20871 ;
  assign w20873 = w1129 | w3786 ;
  assign w20874 = w20872 | w20873 ;
  assign w20875 = ( w782 & w5151 ) | ( w782 & ~w20872 ) | ( w5151 & ~w20872 ) ;
  assign w20876 = w20874 | w20875 ;
  assign w20877 = ( w407 & w956 ) | ( w407 & ~w1207 ) | ( w956 & ~w1207 ) ;
  assign w20878 = w2250 | w20876 ;
  assign w20879 = ( w1207 & ~w2250 ) | ( w1207 & w2556 ) | ( ~w2250 & w2556 ) ;
  assign w20880 = w20878 | w20879 ;
  assign w20881 = w20877 | w20880 ;
  assign w20882 = ( w232 & w258 ) | ( w232 & ~w277 ) | ( w258 & ~w277 ) ;
  assign w20883 = w119 | w20881 ;
  assign w20884 = ( ~w119 & w277 ) | ( ~w119 & w1031 ) | ( w277 & w1031 ) ;
  assign w20885 = w20883 | w20884 ;
  assign w20886 = w20882 | w20885 ;
  assign w20887 = ( w20615 & w20753 ) | ( w20615 & w20886 ) | ( w20753 & w20886 ) ;
  assign w20888 = w20615 ^ w20753 ;
  assign w20889 = w20886 ^ w20888 ;
  assign w20890 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16656 ) | ( \pi31 & ~w16656 ) ;
  assign w20891 = ( \pi29 & ~\pi30 ) | ( \pi29 & w20890 ) | ( ~\pi30 & w20890 ) ;
  assign w20892 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w20890 ) | ( \pi30 & w20890 ) ;
  assign w20893 = ( \pi29 & w16658 ) | ( \pi29 & ~w20892 ) | ( w16658 & ~w20892 ) ;
  assign w20894 = ( w16654 & w20892 ) | ( w16654 & w20893 ) | ( w20892 & w20893 ) ;
  assign w20895 = ~\pi31 & w20894 ;
  assign w20896 = ( w20891 & ~w20893 ) | ( w20891 & w20895 ) | ( ~w20893 & w20895 ) ;
  assign w20897 = ( w37 & w17266 ) | ( w37 & w20896 ) | ( w17266 & w20896 ) ;
  assign w20898 = w20896 | w20897 ;
  assign w20899 = ( w20755 & w20764 ) | ( w20755 & w20765 ) | ( w20764 & w20765 ) ;
  assign w20900 = w20889 ^ w20899 ;
  assign w20901 = w20898 ^ w20900 ;
  assign w20902 = w3717 | w16650 ;
  assign w20903 = w3649 & ~w16652 ;
  assign w20904 = ( ~w16650 & w20902 ) | ( ~w16650 & w20903 ) | ( w20902 & w20903 ) ;
  assign w20905 = w3549 | w16648 ;
  assign w20906 = w16752 & ~w20904 ;
  assign w20907 = ( w3448 & w20904 ) | ( w3448 & ~w20906 ) | ( w20904 & ~w20906 ) ;
  assign w20908 = ( ~w16648 & w20905 ) | ( ~w16648 & w20907 ) | ( w20905 & w20907 ) ;
  assign w20909 = \pi29 ^ w20908 ;
  assign w20910 = w4143 | w16644 ;
  assign w20911 = w4052 & ~w16646 ;
  assign w20912 = ( ~w16644 & w20910 ) | ( ~w16644 & w20911 ) | ( w20910 & w20911 ) ;
  assign w20913 = ~w4147 & w17455 ;
  assign w20914 = w16642 | w20912 ;
  assign w20915 = ( w3964 & w20912 ) | ( w3964 & w20914 ) | ( w20912 & w20914 ) ;
  assign w20916 = ( w17455 & ~w20913 ) | ( w17455 & w20915 ) | ( ~w20913 & w20915 ) ;
  assign w20917 = \pi26 ^ w20916 ;
  assign w20918 = w20901 ^ w20917 ;
  assign w20919 = w20909 ^ w20918 ;
  assign w20920 = ( w20767 & w20775 ) | ( w20767 & w20783 ) | ( w20775 & w20783 ) ;
  assign w20921 = w4651 | w16638 ;
  assign w20922 = w4606 & w16640 ;
  assign w20923 = ( ~w16638 & w20921 ) | ( ~w16638 & w20922 ) | ( w20921 & w20922 ) ;
  assign w20924 = ~w4706 & w16636 ;
  assign w20925 = w17770 & ~w20923 ;
  assign w20926 = ( w4609 & w20923 ) | ( w4609 & ~w20925 ) | ( w20923 & ~w20925 ) ;
  assign w20927 = ( w16636 & ~w20924 ) | ( w16636 & w20926 ) | ( ~w20924 & w20926 ) ;
  assign w20928 = \pi23 ^ w20927 ;
  assign w20929 = w20919 ^ w20920 ;
  assign w20930 = w20928 ^ w20929 ;
  assign w20931 = ( w20785 & w20786 ) | ( w20785 & w20794 ) | ( w20786 & w20794 ) ;
  assign w20932 = ~w5343 & w16632 ;
  assign w20933 = w4905 & ~w16634 ;
  assign w20934 = ( w16632 & ~w20932 ) | ( w16632 & w20933 ) | ( ~w20932 & w20933 ) ;
  assign w20935 = w5395 | w16630 ;
  assign w20936 = w18038 & ~w20934 ;
  assign w20937 = ( w4908 & w20934 ) | ( w4908 & ~w20936 ) | ( w20934 & ~w20936 ) ;
  assign w20938 = ( ~w16630 & w20935 ) | ( ~w16630 & w20937 ) | ( w20935 & w20937 ) ;
  assign w20939 = \pi20 ^ w20938 ;
  assign w20940 = w20930 ^ w20931 ;
  assign w20941 = w20939 ^ w20940 ;
  assign w20942 = ( w20796 & w20797 ) | ( w20796 & w20805 ) | ( w20797 & w20805 ) ;
  assign w20943 = w5710 | w16626 ;
  assign w20944 = w5494 & ~w16628 ;
  assign w20945 = ( ~w16626 & w20943 ) | ( ~w16626 & w20944 ) | ( w20943 & w20944 ) ;
  assign w20946 = ~w5948 & w16619 ;
  assign w20947 = w18451 | w20945 ;
  assign w20948 = ( w5497 & w20945 ) | ( w5497 & w20947 ) | ( w20945 & w20947 ) ;
  assign w20949 = ( w16619 & ~w20946 ) | ( w16619 & w20948 ) | ( ~w20946 & w20948 ) ;
  assign w20950 = \pi17 ^ w20949 ;
  assign w20951 = w20941 ^ w20942 ;
  assign w20952 = w20950 ^ w20951 ;
  assign w20953 = ( w20807 & w20808 ) | ( w20807 & w20816 ) | ( w20808 & w20816 ) ;
  assign w20954 = ~w6549 & w16617 ;
  assign w20955 = w6048 & w16621 ;
  assign w20956 = ( w16617 & ~w20954 ) | ( w16617 & w20955 ) | ( ~w20954 & w20955 ) ;
  assign w20957 = w6637 | w18914 ;
  assign w20958 = w19350 & ~w20956 ;
  assign w20959 = ( w6045 & w20956 ) | ( w6045 & ~w20958 ) | ( w20956 & ~w20958 ) ;
  assign w20960 = ( ~w18914 & w20957 ) | ( ~w18914 & w20959 ) | ( w20957 & w20959 ) ;
  assign w20961 = \pi14 ^ w20960 ;
  assign w20962 = w20952 ^ w20953 ;
  assign w20963 = w20961 ^ w20962 ;
  assign w20964 = ( w20818 & w20819 ) | ( w20818 & w20827 ) | ( w20819 & w20827 ) ;
  assign w20965 = w6949 | w18912 ;
  assign w20966 = w6748 & w18916 ;
  assign w20967 = ( ~w18912 & w20965 ) | ( ~w18912 & w20966 ) | ( w20965 & w20966 ) ;
  assign w20968 = ~w7154 & w19529 ;
  assign w20969 = w19540 & ~w20967 ;
  assign w20970 = ( w6751 & w20967 ) | ( w6751 & ~w20969 ) | ( w20967 & ~w20969 ) ;
  assign w20971 = ( w19529 & ~w20968 ) | ( w19529 & w20970 ) | ( ~w20968 & w20970 ) ;
  assign w20972 = \pi11 ^ w20971 ;
  assign w20973 = w20963 ^ w20964 ;
  assign w20974 = w20972 ^ w20973 ;
  assign w20975 = ( w20829 & w20830 ) | ( w20829 & w20838 ) | ( w20830 & w20838 ) ;
  assign w20976 = ~w7673 & w19887 ;
  assign w20977 = w7411 & w19713 ;
  assign w20978 = ( w19887 & ~w20976 ) | ( w19887 & w20977 ) | ( ~w20976 & w20977 ) ;
  assign w20979 = w7944 | w20068 ;
  assign w20980 = w20081 & ~w20978 ;
  assign w20981 = ( w7414 & w20978 ) | ( w7414 & ~w20980 ) | ( w20978 & ~w20980 ) ;
  assign w20982 = ( ~w20068 & w20979 ) | ( ~w20068 & w20981 ) | ( w20979 & w20981 ) ;
  assign w20983 = \pi08 ^ w20982 ;
  assign w20984 = w20974 ^ w20975 ;
  assign w20985 = w20983 ^ w20984 ;
  assign w20986 = ( w20840 & w20841 ) | ( w20840 & w20849 ) | ( w20841 & w20849 ) ;
  assign w20987 = w8593 & w20404 ;
  assign w20988 = ( w35 & w20404 ) | ( w35 & w20987 ) | ( w20404 & w20987 ) ;
  assign w20989 = w8262 & w20247 ;
  assign w20990 = w20988 | w20989 ;
  assign w20991 = w8263 & ~w20414 ;
  assign w20992 = ( w8263 & w20990 ) | ( w8263 & ~w20991 ) | ( w20990 & ~w20991 ) ;
  assign w20993 = w20985 ^ w20992 ;
  assign w20994 = \pi05 ^ w20986 ;
  assign w20995 = w20993 ^ w20994 ;
  assign w20996 = ( w20851 & w20852 ) | ( w20851 & w20860 ) | ( w20852 & w20860 ) ;
  assign w20997 = ( w20862 & w20863 ) | ( w20862 & w20864 ) | ( w20863 & w20864 ) ;
  assign w20998 = w20995 ^ w20997 ;
  assign w20999 = w20996 ^ w20998 ;
  assign w21000 = w20867 & w20999 ;
  assign w21001 = w20867 ^ w20999 ;
  assign w21002 = ( w20995 & w20996 ) | ( w20995 & w20997 ) | ( w20996 & w20997 ) ;
  assign w21003 = w20414 | w20990 ;
  assign w21004 = ( w8263 & w20990 ) | ( w8263 & w21003 ) | ( w20990 & w21003 ) ;
  assign w21005 = \pi05 ^ w21004 ;
  assign w21006 = ( w20985 & w20986 ) | ( w20985 & w21005 ) | ( w20986 & w21005 ) ;
  assign w21007 = ( w20889 & w20898 ) | ( w20889 & w20899 ) | ( w20898 & w20899 ) ;
  assign w21008 = ( w210 & w681 ) | ( w210 & ~w725 ) | ( w681 & ~w725 ) ;
  assign w21009 = w1095 | w1919 ;
  assign w21010 = ( w725 & ~w1095 ) | ( w725 & w1340 ) | ( ~w1095 & w1340 ) ;
  assign w21011 = w21009 | w21010 ;
  assign w21012 = w21008 | w21011 ;
  assign w21013 = ( w76 & w230 ) | ( w76 & ~w254 ) | ( w230 & ~w254 ) ;
  assign w21014 = w11063 | w21012 ;
  assign w21015 = ( w254 & w524 ) | ( w254 & ~w11063 ) | ( w524 & ~w11063 ) ;
  assign w21016 = w21014 | w21015 ;
  assign w21017 = w21013 | w21016 ;
  assign w21018 = ( ~w286 & w1814 ) | ( ~w286 & w3965 ) | ( w1814 & w3965 ) ;
  assign w21019 = w3132 | w21017 ;
  assign w21020 = ( w286 & w445 ) | ( w286 & ~w3132 ) | ( w445 & ~w3132 ) ;
  assign w21021 = w21019 | w21020 ;
  assign w21022 = w21018 | w21021 ;
  assign w21023 = ( w86 & w262 ) | ( w86 & ~w345 ) | ( w262 & ~w345 ) ;
  assign w21024 = w16891 | w21022 ;
  assign w21025 = ( w345 & w758 ) | ( w345 & ~w16891 ) | ( w758 & ~w16891 ) ;
  assign w21026 = w21024 | w21025 ;
  assign w21027 = w21023 | w21026 ;
  assign w21028 = w20615 ^ w21027 ;
  assign w21029 = w12003 ^ w20404 ;
  assign w21030 = ( \pi05 & w12003 ) | ( \pi05 & ~w21029 ) | ( w12003 & ~w21029 ) ;
  assign w21031 = w21028 | w21030 ;
  assign w21032 = \pi05 ^ w20404 ;
  assign w21033 = ( \pi04 & w12231 ) | ( \pi04 & w21032 ) | ( w12231 & w21032 ) ;
  assign w21034 = w21028 ^ w21033 ;
  assign w21035 = ( \pi29 & \pi31 ) | ( \pi29 & w16654 ) | ( \pi31 & w16654 ) ;
  assign w21036 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21035 ) | ( ~\pi30 & w21035 ) ;
  assign w21037 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21035 ) | ( \pi30 & w21035 ) ;
  assign w21038 = ( \pi29 & w16656 ) | ( \pi29 & ~w21037 ) | ( w16656 & ~w21037 ) ;
  assign w21039 = ( ~w16652 & w21037 ) | ( ~w16652 & w21038 ) | ( w21037 & w21038 ) ;
  assign w21040 = ~\pi31 & w21039 ;
  assign w21041 = ( w21036 & ~w21038 ) | ( w21036 & w21040 ) | ( ~w21038 & w21040 ) ;
  assign w21042 = ( w37 & w17293 ) | ( w37 & w21041 ) | ( w17293 & w21041 ) ;
  assign w21043 = w21041 | w21042 ;
  assign w21044 = w20887 ^ w21034 ;
  assign w21045 = w21043 ^ w21044 ;
  assign w21046 = w3717 | w16648 ;
  assign w21047 = w3649 & ~w16650 ;
  assign w21048 = ( ~w16648 & w21046 ) | ( ~w16648 & w21047 ) | ( w21046 & w21047 ) ;
  assign w21049 = w3549 | w16646 ;
  assign w21050 = w17476 & ~w21048 ;
  assign w21051 = ( w3448 & w21048 ) | ( w3448 & ~w21050 ) | ( w21048 & ~w21050 ) ;
  assign w21052 = ( ~w16646 & w21049 ) | ( ~w16646 & w21051 ) | ( w21049 & w21051 ) ;
  assign w21053 = \pi29 ^ w21052 ;
  assign w21054 = w21007 ^ w21045 ;
  assign w21055 = w21053 ^ w21054 ;
  assign w21056 = ~w4143 & w16642 ;
  assign w21057 = w4052 & ~w16644 ;
  assign w21058 = ( w16642 & ~w21056 ) | ( w16642 & w21057 ) | ( ~w21056 & w21057 ) ;
  assign w21059 = w4147 | w17760 ;
  assign w21060 = w16640 | w21058 ;
  assign w21061 = ( w3964 & w21058 ) | ( w3964 & w21060 ) | ( w21058 & w21060 ) ;
  assign w21062 = ( ~w17760 & w21059 ) | ( ~w17760 & w21061 ) | ( w21059 & w21061 ) ;
  assign w21063 = \pi26 ^ w21062 ;
  assign w21064 = ( w20901 & w20909 ) | ( w20901 & w20917 ) | ( w20909 & w20917 ) ;
  assign w21065 = w21055 ^ w21064 ;
  assign w21066 = w21063 ^ w21065 ;
  assign w21067 = ~w4651 & w16636 ;
  assign w21068 = w4606 & ~w16638 ;
  assign w21069 = ( w16636 & ~w21067 ) | ( w16636 & w21068 ) | ( ~w21067 & w21068 ) ;
  assign w21070 = w4706 | w16634 ;
  assign w21071 = w16742 & ~w21069 ;
  assign w21072 = ( w4609 & w21069 ) | ( w4609 & ~w21071 ) | ( w21069 & ~w21071 ) ;
  assign w21073 = ( ~w16634 & w21070 ) | ( ~w16634 & w21072 ) | ( w21070 & w21072 ) ;
  assign w21074 = \pi23 ^ w21073 ;
  assign w21075 = ( w20919 & w20920 ) | ( w20919 & w20928 ) | ( w20920 & w20928 ) ;
  assign w21076 = w21066 ^ w21075 ;
  assign w21077 = w21074 ^ w21076 ;
  assign w21078 = w5343 | w16630 ;
  assign w21079 = w4905 & w16632 ;
  assign w21080 = ( ~w16630 & w21078 ) | ( ~w16630 & w21079 ) | ( w21078 & w21079 ) ;
  assign w21081 = w5395 | w16628 ;
  assign w21082 = w18026 | w21080 ;
  assign w21083 = ( w4908 & w21080 ) | ( w4908 & w21082 ) | ( w21080 & w21082 ) ;
  assign w21084 = ( ~w16628 & w21081 ) | ( ~w16628 & w21083 ) | ( w21081 & w21083 ) ;
  assign w21085 = \pi20 ^ w21084 ;
  assign w21086 = ( w20930 & w20931 ) | ( w20930 & w20939 ) | ( w20931 & w20939 ) ;
  assign w21087 = w21077 ^ w21086 ;
  assign w21088 = w21085 ^ w21087 ;
  assign w21089 = ~w5710 & w16619 ;
  assign w21090 = w5494 & ~w16626 ;
  assign w21091 = ( w16619 & ~w21089 ) | ( w16619 & w21090 ) | ( ~w21089 & w21090 ) ;
  assign w21092 = ~w5948 & w16621 ;
  assign w21093 = w18439 & ~w21091 ;
  assign w21094 = ( w5497 & w21091 ) | ( w5497 & ~w21093 ) | ( w21091 & ~w21093 ) ;
  assign w21095 = ( w16621 & ~w21092 ) | ( w16621 & w21094 ) | ( ~w21092 & w21094 ) ;
  assign w21096 = \pi17 ^ w21095 ;
  assign w21097 = ( w20941 & w20942 ) | ( w20941 & w20950 ) | ( w20942 & w20950 ) ;
  assign w21098 = w21088 ^ w21097 ;
  assign w21099 = w21096 ^ w21098 ;
  assign w21100 = ( w20952 & w20953 ) | ( w20952 & w20961 ) | ( w20953 & w20961 ) ;
  assign w21101 = w6549 | w18914 ;
  assign w21102 = w6048 & w16617 ;
  assign w21103 = ( ~w18914 & w21101 ) | ( ~w18914 & w21102 ) | ( w21101 & w21102 ) ;
  assign w21104 = ~w6637 & w18916 ;
  assign w21105 = w19366 & ~w21103 ;
  assign w21106 = ( w6045 & w21103 ) | ( w6045 & ~w21105 ) | ( w21103 & ~w21105 ) ;
  assign w21107 = ( w18916 & ~w21104 ) | ( w18916 & w21106 ) | ( ~w21104 & w21106 ) ;
  assign w21108 = \pi14 ^ w21107 ;
  assign w21109 = w21099 ^ w21100 ;
  assign w21110 = w21108 ^ w21109 ;
  assign w21111 = ~w6949 & w19529 ;
  assign w21112 = w6748 & ~w18912 ;
  assign w21113 = ( w19529 & ~w21111 ) | ( w19529 & w21112 ) | ( ~w21111 & w21112 ) ;
  assign w21114 = ~w7154 & w19713 ;
  assign w21115 = w19723 | w21113 ;
  assign w21116 = ( w6751 & w21113 ) | ( w6751 & w21115 ) | ( w21113 & w21115 ) ;
  assign w21117 = ( w19713 & ~w21114 ) | ( w19713 & w21116 ) | ( ~w21114 & w21116 ) ;
  assign w21118 = \pi11 ^ w21117 ;
  assign w21119 = ( w20963 & w20964 ) | ( w20963 & w20972 ) | ( w20964 & w20972 ) ;
  assign w21120 = w21110 ^ w21119 ;
  assign w21121 = w21118 ^ w21120 ;
  assign w21122 = ( w20974 & w20975 ) | ( w20974 & w20983 ) | ( w20975 & w20983 ) ;
  assign w21123 = w7673 | w20068 ;
  assign w21124 = w7411 & w19887 ;
  assign w21125 = ( ~w20068 & w21123 ) | ( ~w20068 & w21124 ) | ( w21123 & w21124 ) ;
  assign w21126 = ~w7944 & w20247 ;
  assign w21127 = w20257 & ~w21125 ;
  assign w21128 = ( w7414 & w21125 ) | ( w7414 & ~w21127 ) | ( w21125 & ~w21127 ) ;
  assign w21129 = ( w20247 & ~w21126 ) | ( w20247 & w21128 ) | ( ~w21126 & w21128 ) ;
  assign w21130 = \pi08 ^ w21129 ;
  assign w21131 = w21121 ^ w21122 ;
  assign w21132 = w21130 ^ w21131 ;
  assign w21133 = w21002 ^ w21006 ;
  assign w21134 = w21132 ^ w21133 ;
  assign w21135 = w21000 & w21134 ;
  assign w21136 = w21000 ^ w21134 ;
  assign w21137 = ( w21007 & w21045 ) | ( w21007 & w21053 ) | ( w21045 & w21053 ) ;
  assign w21138 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16652 ) | ( \pi31 & ~w16652 ) ;
  assign w21139 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21138 ) | ( ~\pi30 & w21138 ) ;
  assign w21140 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21138 ) | ( \pi30 & w21138 ) ;
  assign w21141 = ( ~\pi29 & w16654 ) | ( ~\pi29 & w21140 ) | ( w16654 & w21140 ) ;
  assign w21142 = ( w16650 & ~w21140 ) | ( w16650 & w21141 ) | ( ~w21140 & w21141 ) ;
  assign w21143 = \pi31 | w21142 ;
  assign w21144 = ( w21139 & w21141 ) | ( w21139 & ~w21143 ) | ( w21141 & ~w21143 ) ;
  assign w21145 = ( w37 & ~w17277 ) | ( w37 & w21144 ) | ( ~w17277 & w21144 ) ;
  assign w21146 = w21144 | w21145 ;
  assign w21147 = ( w515 & w525 ) | ( w515 & ~w570 ) | ( w525 & ~w570 ) ;
  assign w21148 = w325 | w5808 ;
  assign w21149 = ( ~w325 & w570 ) | ( ~w325 & w889 ) | ( w570 & w889 ) ;
  assign w21150 = w21148 | w21149 ;
  assign w21151 = w21147 | w21150 ;
  assign w21152 = ( ~w84 & w341 ) | ( ~w84 & w21151 ) | ( w341 & w21151 ) ;
  assign w21153 = w84 | w21152 ;
  assign w21154 = ( ~w201 & w661 ) | ( ~w201 & w6351 ) | ( w661 & w6351 ) ;
  assign w21155 = w3562 | w21153 ;
  assign w21156 = ( w201 & w221 ) | ( w201 & ~w3562 ) | ( w221 & ~w3562 ) ;
  assign w21157 = w21155 | w21156 ;
  assign w21158 = w21154 | w21157 ;
  assign w21159 = ( w88 & w180 ) | ( w88 & ~w206 ) | ( w180 & ~w206 ) ;
  assign w21160 = w1166 | w21158 ;
  assign w21161 = ( w206 & w225 ) | ( w206 & ~w1166 ) | ( w225 & ~w1166 ) ;
  assign w21162 = w21160 | w21161 ;
  assign w21163 = w21159 | w21162 ;
  assign w21164 = ( w758 & w817 ) | ( w758 & ~w821 ) | ( w817 & ~w821 ) ;
  assign w21165 = w309 | w340 ;
  assign w21166 = ( ~w340 & w821 ) | ( ~w340 & w1094 ) | ( w821 & w1094 ) ;
  assign w21167 = w21165 | w21166 ;
  assign w21168 = w21164 | w21167 ;
  assign w21169 = w6432 | w21168 ;
  assign w21170 = ( ~w603 & w1412 ) | ( ~w603 & w21169 ) | ( w1412 & w21169 ) ;
  assign w21171 = w487 | w21163 ;
  assign w21172 = ( ~w487 & w603 ) | ( ~w487 & w2808 ) | ( w603 & w2808 ) ;
  assign w21173 = w21171 | w21172 ;
  assign w21174 = w21170 | w21173 ;
  assign w21175 = ( w119 & w199 ) | ( w119 & ~w229 ) | ( w199 & ~w229 ) ;
  assign w21176 = w1882 | w21174 ;
  assign w21177 = ( w229 & w565 ) | ( w229 & ~w1882 ) | ( w565 & ~w1882 ) ;
  assign w21178 = w21176 | w21177 ;
  assign w21179 = w21175 | w21178 ;
  assign w21180 = ( ~w1031 & w1274 ) | ( ~w1031 & w21179 ) | ( w1274 & w21179 ) ;
  assign w21181 = w1031 | w21180 ;
  assign w21182 = ( w257 & w344 ) | ( w257 & ~w492 ) | ( w344 & ~w492 ) ;
  assign w21183 = w136 | w21181 ;
  assign w21184 = ( ~w136 & w492 ) | ( ~w136 & w662 ) | ( w492 & w662 ) ;
  assign w21185 = w21183 | w21184 ;
  assign w21186 = w21182 | w21185 ;
  assign w21187 = ( w20615 & ~w21027 ) | ( w20615 & w21031 ) | ( ~w21027 & w21031 ) ;
  assign w21188 = w21031 & w21187 ;
  assign w21189 = w21146 ^ w21188 ;
  assign w21190 = w21186 ^ w21189 ;
  assign w21191 = ( w20887 & w21034 ) | ( w20887 & w21043 ) | ( w21034 & w21043 ) ;
  assign w21192 = w3549 & ~w16644 ;
  assign w21193 = ( w3717 & ~w16646 ) | ( w3717 & w21192 ) | ( ~w16646 & w21192 ) ;
  assign w21194 = w3649 | w21193 ;
  assign w21195 = ( ~w16648 & w21193 ) | ( ~w16648 & w21194 ) | ( w21193 & w21194 ) ;
  assign w21196 = w21192 | w21195 ;
  assign w21197 = w3448 | w17468 ;
  assign w21198 = ( ~w17468 & w21196 ) | ( ~w17468 & w21197 ) | ( w21196 & w21197 ) ;
  assign w21199 = \pi29 ^ w21198 ;
  assign w21200 = w21190 ^ w21191 ;
  assign w21201 = w21199 ^ w21200 ;
  assign w21202 = ~w4143 & w16640 ;
  assign w21203 = w4052 & w16642 ;
  assign w21204 = ( w16640 & ~w21202 ) | ( w16640 & w21203 ) | ( ~w21202 & w21203 ) ;
  assign w21205 = w4147 | w17783 ;
  assign w21206 = w16638 & ~w21204 ;
  assign w21207 = ( w3964 & w21204 ) | ( w3964 & ~w21206 ) | ( w21204 & ~w21206 ) ;
  assign w21208 = ( ~w17783 & w21205 ) | ( ~w17783 & w21207 ) | ( w21205 & w21207 ) ;
  assign w21209 = \pi26 ^ w21208 ;
  assign w21210 = w21137 ^ w21201 ;
  assign w21211 = w21209 ^ w21210 ;
  assign w21212 = ( w21055 & w21063 ) | ( w21055 & w21064 ) | ( w21063 & w21064 ) ;
  assign w21213 = w4651 | w16634 ;
  assign w21214 = w4606 & w16636 ;
  assign w21215 = ( ~w16634 & w21213 ) | ( ~w16634 & w21214 ) | ( w21213 & w21214 ) ;
  assign w21216 = ~w4706 & w16632 ;
  assign w21217 = w18051 & ~w21215 ;
  assign w21218 = ( w4609 & w21215 ) | ( w4609 & ~w21217 ) | ( w21215 & ~w21217 ) ;
  assign w21219 = ( w16632 & ~w21216 ) | ( w16632 & w21218 ) | ( ~w21216 & w21218 ) ;
  assign w21220 = \pi23 ^ w21219 ;
  assign w21221 = w21211 ^ w21212 ;
  assign w21222 = w21220 ^ w21221 ;
  assign w21223 = ( w21066 & w21074 ) | ( w21066 & w21075 ) | ( w21074 & w21075 ) ;
  assign w21224 = w5343 | w16628 ;
  assign w21225 = w4905 & ~w16630 ;
  assign w21226 = ( ~w16628 & w21224 ) | ( ~w16628 & w21225 ) | ( w21224 & w21225 ) ;
  assign w21227 = w5395 | w16626 ;
  assign w21228 = w18429 & ~w21226 ;
  assign w21229 = ( w4908 & w21226 ) | ( w4908 & ~w21228 ) | ( w21226 & ~w21228 ) ;
  assign w21230 = ( ~w16626 & w21227 ) | ( ~w16626 & w21229 ) | ( w21227 & w21229 ) ;
  assign w21231 = \pi20 ^ w21230 ;
  assign w21232 = w21222 ^ w21223 ;
  assign w21233 = w21231 ^ w21232 ;
  assign w21234 = ( w21077 & w21085 ) | ( w21077 & w21086 ) | ( w21085 & w21086 ) ;
  assign w21235 = ~w5710 & w16621 ;
  assign w21236 = w5494 & w16619 ;
  assign w21237 = ( w16621 & ~w21235 ) | ( w16621 & w21236 ) | ( ~w21235 & w21236 ) ;
  assign w21238 = ~w5948 & w16617 ;
  assign w21239 = w16732 | w21237 ;
  assign w21240 = ( w5497 & w21237 ) | ( w5497 & w21239 ) | ( w21237 & w21239 ) ;
  assign w21241 = ( w16617 & ~w21238 ) | ( w16617 & w21240 ) | ( ~w21238 & w21240 ) ;
  assign w21242 = \pi17 ^ w21241 ;
  assign w21243 = w21233 ^ w21234 ;
  assign w21244 = w21242 ^ w21243 ;
  assign w21245 = ( w21088 & w21096 ) | ( w21088 & w21097 ) | ( w21096 & w21097 ) ;
  assign w21246 = ~w6549 & w18916 ;
  assign w21247 = w6048 & ~w18914 ;
  assign w21248 = ( w18916 & ~w21246 ) | ( w18916 & w21247 ) | ( ~w21246 & w21247 ) ;
  assign w21249 = w6637 | w18912 ;
  assign w21250 = w18929 & ~w21248 ;
  assign w21251 = ( w6045 & w21248 ) | ( w6045 & ~w21250 ) | ( w21248 & ~w21250 ) ;
  assign w21252 = ( ~w18912 & w21249 ) | ( ~w18912 & w21251 ) | ( w21249 & w21251 ) ;
  assign w21253 = \pi14 ^ w21252 ;
  assign w21254 = w21244 ^ w21245 ;
  assign w21255 = w21253 ^ w21254 ;
  assign w21256 = ( w21099 & w21100 ) | ( w21099 & w21108 ) | ( w21100 & w21108 ) ;
  assign w21257 = ~w6949 & w19713 ;
  assign w21258 = w6748 & w19529 ;
  assign w21259 = ( w19713 & ~w21257 ) | ( w19713 & w21258 ) | ( ~w21257 & w21258 ) ;
  assign w21260 = ~w7154 & w19887 ;
  assign w21261 = w19898 | w21259 ;
  assign w21262 = ( w6751 & w21259 ) | ( w6751 & w21261 ) | ( w21259 & w21261 ) ;
  assign w21263 = ( w19887 & ~w21260 ) | ( w19887 & w21262 ) | ( ~w21260 & w21262 ) ;
  assign w21264 = \pi11 ^ w21263 ;
  assign w21265 = w21255 ^ w21256 ;
  assign w21266 = w21264 ^ w21265 ;
  assign w21267 = ( w21110 & w21118 ) | ( w21110 & w21119 ) | ( w21118 & w21119 ) ;
  assign w21268 = ~w7673 & w20247 ;
  assign w21269 = w7411 & ~w20068 ;
  assign w21270 = ( w20247 & ~w21268 ) | ( w20247 & w21269 ) | ( ~w21268 & w21269 ) ;
  assign w21271 = ~w7944 & w20404 ;
  assign w21272 = w20417 | w21270 ;
  assign w21273 = ( w7414 & w21270 ) | ( w7414 & w21272 ) | ( w21270 & w21272 ) ;
  assign w21274 = ( w20404 & ~w21271 ) | ( w20404 & w21273 ) | ( ~w21271 & w21273 ) ;
  assign w21275 = \pi08 ^ w21274 ;
  assign w21276 = w21266 ^ w21267 ;
  assign w21277 = w21275 ^ w21276 ;
  assign w21278 = ( w21121 & w21122 ) | ( w21121 & w21130 ) | ( w21122 & w21130 ) ;
  assign w21279 = ( w21002 & w21006 ) | ( w21002 & w21132 ) | ( w21006 & w21132 ) ;
  assign w21280 = w21277 ^ w21279 ;
  assign w21281 = w21278 ^ w21280 ;
  assign w21282 = w21135 ^ w21281 ;
  assign w21283 = w21135 & w21281 ;
  assign w21284 = ( ~w21146 & w21186 ) | ( ~w21146 & w21188 ) | ( w21186 & w21188 ) ;
  assign w21285 = ( w232 & w281 ) | ( w232 & ~w286 ) | ( w281 & ~w286 ) ;
  assign w21286 = w136 | w147 ;
  assign w21287 = ( ~w147 & w286 ) | ( ~w147 & w491 ) | ( w286 & w491 ) ;
  assign w21288 = w21286 | w21287 ;
  assign w21289 = w21285 | w21288 ;
  assign w21290 = w252 | w680 ;
  assign w21291 = ( ~w252 & w595 ) | ( ~w252 & w21289 ) | ( w595 & w21289 ) ;
  assign w21292 = w21290 | w21291 ;
  assign w21293 = ( w209 & w283 ) | ( w209 & ~w383 ) | ( w283 & ~w383 ) ;
  assign w21294 = w176 | w959 ;
  assign w21295 = ( ~w176 & w383 ) | ( ~w176 & w722 ) | ( w383 & w722 ) ;
  assign w21296 = w21294 | w21295 ;
  assign w21297 = w21293 | w21296 ;
  assign w21298 = w2518 | w4381 ;
  assign w21299 = w21297 | w21298 ;
  assign w21300 = ( ~w1069 & w2530 ) | ( ~w1069 & w21297 ) | ( w2530 & w21297 ) ;
  assign w21301 = ~w21299 & w21300 ;
  assign w21302 = w135 | w271 ;
  assign w21303 = w900 | w21302 ;
  assign w21304 = ( ~w125 & w900 ) | ( ~w125 & w21301 ) | ( w900 & w21301 ) ;
  assign w21305 = ~w21303 & w21304 ;
  assign w21306 = ( w165 & ~w223 ) | ( w165 & w21305 ) | ( ~w223 & w21305 ) ;
  assign w21307 = ~w165 & w21306 ;
  assign w21308 = ( ~w6174 & w10233 ) | ( ~w6174 & w11042 ) | ( w10233 & w11042 ) ;
  assign w21309 = w6174 | w21308 ;
  assign w21310 = w3140 | w21292 ;
  assign w21311 = w21307 & ~w21310 ;
  assign w21312 = ( w9867 & w21307 ) | ( w9867 & w21309 ) | ( w21307 & w21309 ) ;
  assign w21313 = w21311 & ~w21312 ;
  assign w21314 = ( w221 & w230 ) | ( w221 & ~w429 ) | ( w230 & ~w429 ) ;
  assign w21315 = ~w169 & w21313 ;
  assign w21316 = ( ~w169 & w429 ) | ( ~w169 & w463 ) | ( w429 & w463 ) ;
  assign w21317 = w21315 & ~w21316 ;
  assign w21318 = ~w21314 & w21317 ;
  assign w21319 = w309 | w534 ;
  assign w21320 = ( w309 & ~w316 ) | ( w309 & w21318 ) | ( ~w316 & w21318 ) ;
  assign w21321 = ~w21319 & w21320 ;
  assign w21322 = ( w21186 & w21284 ) | ( w21186 & w21321 ) | ( w21284 & w21321 ) ;
  assign w21323 = w21284 ^ w21321 ;
  assign w21324 = w21186 ^ w21323 ;
  assign w21325 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16650 ) | ( \pi31 & ~w16650 ) ;
  assign w21326 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21325 ) | ( ~\pi30 & w21325 ) ;
  assign w21327 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21325 ) | ( \pi30 & w21325 ) ;
  assign w21328 = ( \pi29 & w16652 ) | ( \pi29 & ~w21327 ) | ( w16652 & ~w21327 ) ;
  assign w21329 = ( ~w16648 & w21327 ) | ( ~w16648 & w21328 ) | ( w21327 & w21328 ) ;
  assign w21330 = ~\pi31 & w21329 ;
  assign w21331 = ( w21326 & ~w21328 ) | ( w21326 & w21330 ) | ( ~w21328 & w21330 ) ;
  assign w21332 = ( w37 & ~w16752 ) | ( w37 & w21331 ) | ( ~w16752 & w21331 ) ;
  assign w21333 = w21331 | w21332 ;
  assign w21334 = ( w21190 & w21191 ) | ( w21190 & w21199 ) | ( w21191 & w21199 ) ;
  assign w21335 = w21324 ^ w21334 ;
  assign w21336 = w21333 ^ w21335 ;
  assign w21337 = w3717 | w16644 ;
  assign w21338 = w3649 & ~w16646 ;
  assign w21339 = ( ~w16644 & w21337 ) | ( ~w16644 & w21338 ) | ( w21337 & w21338 ) ;
  assign w21340 = ~w3549 & w16642 ;
  assign w21341 = w17455 | w21339 ;
  assign w21342 = ( w3448 & w21339 ) | ( w3448 & w21341 ) | ( w21339 & w21341 ) ;
  assign w21343 = ( w16642 & ~w21340 ) | ( w16642 & w21342 ) | ( ~w21340 & w21342 ) ;
  assign w21344 = \pi29 ^ w21343 ;
  assign w21345 = w4143 | w16638 ;
  assign w21346 = w4052 & w16640 ;
  assign w21347 = ( ~w16638 & w21345 ) | ( ~w16638 & w21346 ) | ( w21345 & w21346 ) ;
  assign w21348 = w4147 | w17770 ;
  assign w21349 = w16636 | w21347 ;
  assign w21350 = ( w3964 & w21347 ) | ( w3964 & w21349 ) | ( w21347 & w21349 ) ;
  assign w21351 = ( ~w17770 & w21348 ) | ( ~w17770 & w21350 ) | ( w21348 & w21350 ) ;
  assign w21352 = \pi26 ^ w21351 ;
  assign w21353 = w21336 ^ w21352 ;
  assign w21354 = w21344 ^ w21353 ;
  assign w21355 = ( w21137 & w21201 ) | ( w21137 & w21209 ) | ( w21201 & w21209 ) ;
  assign w21356 = ~w4651 & w16632 ;
  assign w21357 = w4606 & ~w16634 ;
  assign w21358 = ( w16632 & ~w21356 ) | ( w16632 & w21357 ) | ( ~w21356 & w21357 ) ;
  assign w21359 = w4706 | w16630 ;
  assign w21360 = w18038 & ~w21358 ;
  assign w21361 = ( w4609 & w21358 ) | ( w4609 & ~w21360 ) | ( w21358 & ~w21360 ) ;
  assign w21362 = ( ~w16630 & w21359 ) | ( ~w16630 & w21361 ) | ( w21359 & w21361 ) ;
  assign w21363 = \pi23 ^ w21362 ;
  assign w21364 = w21354 ^ w21355 ;
  assign w21365 = w21363 ^ w21364 ;
  assign w21366 = ( w21211 & w21212 ) | ( w21211 & w21220 ) | ( w21212 & w21220 ) ;
  assign w21367 = w5343 | w16626 ;
  assign w21368 = w4905 & ~w16628 ;
  assign w21369 = ( ~w16626 & w21367 ) | ( ~w16626 & w21368 ) | ( w21367 & w21368 ) ;
  assign w21370 = ~w5395 & w16619 ;
  assign w21371 = w18451 | w21369 ;
  assign w21372 = ( w4908 & w21369 ) | ( w4908 & w21371 ) | ( w21369 & w21371 ) ;
  assign w21373 = ( w16619 & ~w21370 ) | ( w16619 & w21372 ) | ( ~w21370 & w21372 ) ;
  assign w21374 = \pi20 ^ w21373 ;
  assign w21375 = w21365 ^ w21366 ;
  assign w21376 = w21374 ^ w21375 ;
  assign w21377 = ( w21222 & w21223 ) | ( w21222 & w21231 ) | ( w21223 & w21231 ) ;
  assign w21378 = ~w5710 & w16617 ;
  assign w21379 = w5494 & w16621 ;
  assign w21380 = ( w16617 & ~w21378 ) | ( w16617 & w21379 ) | ( ~w21378 & w21379 ) ;
  assign w21381 = w5948 | w18914 ;
  assign w21382 = w19350 & ~w21380 ;
  assign w21383 = ( w5497 & w21380 ) | ( w5497 & ~w21382 ) | ( w21380 & ~w21382 ) ;
  assign w21384 = ( ~w18914 & w21381 ) | ( ~w18914 & w21383 ) | ( w21381 & w21383 ) ;
  assign w21385 = \pi17 ^ w21384 ;
  assign w21386 = w21376 ^ w21377 ;
  assign w21387 = w21385 ^ w21386 ;
  assign w21388 = ( w21233 & w21234 ) | ( w21233 & w21242 ) | ( w21234 & w21242 ) ;
  assign w21389 = w6549 | w18912 ;
  assign w21390 = w6048 & w18916 ;
  assign w21391 = ( ~w18912 & w21389 ) | ( ~w18912 & w21390 ) | ( w21389 & w21390 ) ;
  assign w21392 = ~w6637 & w19529 ;
  assign w21393 = w19540 & ~w21391 ;
  assign w21394 = ( w6045 & w21391 ) | ( w6045 & ~w21393 ) | ( w21391 & ~w21393 ) ;
  assign w21395 = ( w19529 & ~w21392 ) | ( w19529 & w21394 ) | ( ~w21392 & w21394 ) ;
  assign w21396 = \pi14 ^ w21395 ;
  assign w21397 = w21387 ^ w21388 ;
  assign w21398 = w21396 ^ w21397 ;
  assign w21399 = ( w21244 & w21245 ) | ( w21244 & w21253 ) | ( w21245 & w21253 ) ;
  assign w21400 = ~w6949 & w19887 ;
  assign w21401 = w6748 & w19713 ;
  assign w21402 = ( w19887 & ~w21400 ) | ( w19887 & w21401 ) | ( ~w21400 & w21401 ) ;
  assign w21403 = w7154 | w20068 ;
  assign w21404 = w20081 & ~w21402 ;
  assign w21405 = ( w6751 & w21402 ) | ( w6751 & ~w21404 ) | ( w21402 & ~w21404 ) ;
  assign w21406 = ( ~w20068 & w21403 ) | ( ~w20068 & w21405 ) | ( w21403 & w21405 ) ;
  assign w21407 = \pi11 ^ w21406 ;
  assign w21408 = w21398 ^ w21399 ;
  assign w21409 = w21407 ^ w21408 ;
  assign w21410 = ( w21255 & w21256 ) | ( w21255 & w21264 ) | ( w21256 & w21264 ) ;
  assign w21411 = w7944 & w20404 ;
  assign w21412 = ( w7673 & w20404 ) | ( w7673 & w21411 ) | ( w20404 & w21411 ) ;
  assign w21413 = w7411 & w20247 ;
  assign w21414 = w21412 | w21413 ;
  assign w21415 = w7414 & ~w20414 ;
  assign w21416 = ( w7414 & w21414 ) | ( w7414 & ~w21415 ) | ( w21414 & ~w21415 ) ;
  assign w21417 = w21409 ^ w21416 ;
  assign w21418 = \pi08 ^ w21410 ;
  assign w21419 = w21417 ^ w21418 ;
  assign w21420 = ( w21266 & w21267 ) | ( w21266 & w21275 ) | ( w21267 & w21275 ) ;
  assign w21421 = ( w21277 & w21278 ) | ( w21277 & w21279 ) | ( w21278 & w21279 ) ;
  assign w21422 = w21419 ^ w21421 ;
  assign w21423 = w21420 ^ w21422 ;
  assign w21424 = w21283 & ~w21423 ;
  assign w21425 = w21283 ^ w21423 ;
  assign w21426 = ( ~w21419 & w21420 ) | ( ~w21419 & w21421 ) | ( w21420 & w21421 ) ;
  assign w21427 = w20414 | w21414 ;
  assign w21428 = ( w7414 & w21414 ) | ( w7414 & w21427 ) | ( w21414 & w21427 ) ;
  assign w21429 = \pi08 ^ w21428 ;
  assign w21430 = ( ~w21409 & w21410 ) | ( ~w21409 & w21429 ) | ( w21410 & w21429 ) ;
  assign w21431 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16648 ) | ( \pi31 & ~w16648 ) ;
  assign w21432 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21431 ) | ( ~\pi30 & w21431 ) ;
  assign w21433 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21431 ) | ( \pi30 & w21431 ) ;
  assign w21434 = ( \pi29 & w16650 ) | ( \pi29 & ~w21433 ) | ( w16650 & ~w21433 ) ;
  assign w21435 = ( ~w16646 & w21433 ) | ( ~w16646 & w21434 ) | ( w21433 & w21434 ) ;
  assign w21436 = ~\pi31 & w21435 ;
  assign w21437 = ( w21432 & ~w21434 ) | ( w21432 & w21436 ) | ( ~w21434 & w21436 ) ;
  assign w21438 = ( w37 & ~w17476 ) | ( w37 & w21437 ) | ( ~w17476 & w21437 ) ;
  assign w21439 = w21437 | w21438 ;
  assign w21440 = w11666 ^ w20404 ;
  assign w21441 = ( \pi08 & w11666 ) | ( \pi08 & ~w21440 ) | ( w11666 & ~w21440 ) ;
  assign w21442 = ( w76 & w230 ) | ( w76 & ~w466 ) | ( w230 & ~w466 ) ;
  assign w21443 = w410 | w1459 ;
  assign w21444 = ( w466 & w470 ) | ( w466 & ~w1459 ) | ( w470 & ~w1459 ) ;
  assign w21445 = w21443 | w21444 ;
  assign w21446 = w21442 | w21445 ;
  assign w21447 = w1616 | w11003 ;
  assign w21448 = w21446 | w21447 ;
  assign w21449 = ( w282 & w2075 ) | ( w282 & ~w21446 ) | ( w2075 & ~w21446 ) ;
  assign w21450 = w21448 | w21449 ;
  assign w21451 = ( ~w138 & w212 ) | ( ~w138 & w21450 ) | ( w212 & w21450 ) ;
  assign w21452 = w2829 & ~w3032 ;
  assign w21453 = ( w138 & w424 ) | ( w138 & w2829 ) | ( w424 & w2829 ) ;
  assign w21454 = w21452 & ~w21453 ;
  assign w21455 = ~w21451 & w21454 ;
  assign w21456 = w354 | w723 ;
  assign w21457 = w126 | w21456 ;
  assign w21458 = ( w126 & ~w2253 ) | ( w126 & w21455 ) | ( ~w2253 & w21455 ) ;
  assign w21459 = ~w21457 & w21458 ;
  assign w21460 = w21186 ^ w21441 ;
  assign w21461 = w21459 ^ w21460 ;
  assign w21462 = w21322 ^ w21461 ;
  assign w21463 = w21439 ^ w21462 ;
  assign w21464 = ~w3717 & w16642 ;
  assign w21465 = w3649 & ~w16644 ;
  assign w21466 = ( w16642 & ~w21464 ) | ( w16642 & w21465 ) | ( ~w21464 & w21465 ) ;
  assign w21467 = ~w3549 & w16640 ;
  assign w21468 = w17760 & ~w21466 ;
  assign w21469 = ( w3448 & w21466 ) | ( w3448 & ~w21468 ) | ( w21466 & ~w21468 ) ;
  assign w21470 = ( w16640 & ~w21467 ) | ( w16640 & w21469 ) | ( ~w21467 & w21469 ) ;
  assign w21471 = \pi29 ^ w21470 ;
  assign w21472 = ( ~w21324 & w21333 ) | ( ~w21324 & w21334 ) | ( w21333 & w21334 ) ;
  assign w21473 = w21463 ^ w21472 ;
  assign w21474 = w21471 ^ w21473 ;
  assign w21475 = ~w4143 & w16636 ;
  assign w21476 = w4052 & ~w16638 ;
  assign w21477 = ( w16636 & ~w21475 ) | ( w16636 & w21476 ) | ( ~w21475 & w21476 ) ;
  assign w21478 = w4147 | w16742 ;
  assign w21479 = w16634 & ~w21477 ;
  assign w21480 = ( w3964 & w21477 ) | ( w3964 & ~w21479 ) | ( w21477 & ~w21479 ) ;
  assign w21481 = ( ~w16742 & w21478 ) | ( ~w16742 & w21480 ) | ( w21478 & w21480 ) ;
  assign w21482 = \pi26 ^ w21481 ;
  assign w21483 = ( ~w21336 & w21344 ) | ( ~w21336 & w21352 ) | ( w21344 & w21352 ) ;
  assign w21484 = w21474 ^ w21483 ;
  assign w21485 = w21482 ^ w21484 ;
  assign w21486 = w4651 | w16630 ;
  assign w21487 = w4606 & w16632 ;
  assign w21488 = ( ~w16630 & w21486 ) | ( ~w16630 & w21487 ) | ( w21486 & w21487 ) ;
  assign w21489 = w4706 | w16628 ;
  assign w21490 = w18026 | w21488 ;
  assign w21491 = ( w4609 & w21488 ) | ( w4609 & w21490 ) | ( w21488 & w21490 ) ;
  assign w21492 = ( ~w16628 & w21489 ) | ( ~w16628 & w21491 ) | ( w21489 & w21491 ) ;
  assign w21493 = \pi23 ^ w21492 ;
  assign w21494 = ( ~w21354 & w21355 ) | ( ~w21354 & w21363 ) | ( w21355 & w21363 ) ;
  assign w21495 = w21485 ^ w21494 ;
  assign w21496 = w21493 ^ w21495 ;
  assign w21497 = ~w5343 & w16619 ;
  assign w21498 = w4905 & ~w16626 ;
  assign w21499 = ( w16619 & ~w21497 ) | ( w16619 & w21498 ) | ( ~w21497 & w21498 ) ;
  assign w21500 = ~w5395 & w16621 ;
  assign w21501 = w18439 & ~w21499 ;
  assign w21502 = ( w4908 & w21499 ) | ( w4908 & ~w21501 ) | ( w21499 & ~w21501 ) ;
  assign w21503 = ( w16621 & ~w21500 ) | ( w16621 & w21502 ) | ( ~w21500 & w21502 ) ;
  assign w21504 = \pi20 ^ w21503 ;
  assign w21505 = ( ~w21365 & w21366 ) | ( ~w21365 & w21374 ) | ( w21366 & w21374 ) ;
  assign w21506 = w21496 ^ w21505 ;
  assign w21507 = w21504 ^ w21506 ;
  assign w21508 = ( ~w21376 & w21377 ) | ( ~w21376 & w21385 ) | ( w21377 & w21385 ) ;
  assign w21509 = w5710 | w18914 ;
  assign w21510 = w5494 & w16617 ;
  assign w21511 = ( ~w18914 & w21509 ) | ( ~w18914 & w21510 ) | ( w21509 & w21510 ) ;
  assign w21512 = ~w5948 & w18916 ;
  assign w21513 = w19366 & ~w21511 ;
  assign w21514 = ( w5497 & w21511 ) | ( w5497 & ~w21513 ) | ( w21511 & ~w21513 ) ;
  assign w21515 = ( w18916 & ~w21512 ) | ( w18916 & w21514 ) | ( ~w21512 & w21514 ) ;
  assign w21516 = \pi17 ^ w21515 ;
  assign w21517 = w21507 ^ w21508 ;
  assign w21518 = w21516 ^ w21517 ;
  assign w21519 = ~w6549 & w19529 ;
  assign w21520 = w6048 & ~w18912 ;
  assign w21521 = ( w19529 & ~w21519 ) | ( w19529 & w21520 ) | ( ~w21519 & w21520 ) ;
  assign w21522 = ~w6637 & w19713 ;
  assign w21523 = w19723 | w21521 ;
  assign w21524 = ( w6045 & w21521 ) | ( w6045 & w21523 ) | ( w21521 & w21523 ) ;
  assign w21525 = ( w19713 & ~w21522 ) | ( w19713 & w21524 ) | ( ~w21522 & w21524 ) ;
  assign w21526 = \pi14 ^ w21525 ;
  assign w21527 = ( ~w21387 & w21388 ) | ( ~w21387 & w21396 ) | ( w21388 & w21396 ) ;
  assign w21528 = w21518 ^ w21527 ;
  assign w21529 = w21526 ^ w21528 ;
  assign w21530 = ( ~w21398 & w21399 ) | ( ~w21398 & w21407 ) | ( w21399 & w21407 ) ;
  assign w21531 = w6949 | w20068 ;
  assign w21532 = w6748 & w19887 ;
  assign w21533 = ( ~w20068 & w21531 ) | ( ~w20068 & w21532 ) | ( w21531 & w21532 ) ;
  assign w21534 = ~w7154 & w20247 ;
  assign w21535 = w20257 & ~w21533 ;
  assign w21536 = ( w6751 & w21533 ) | ( w6751 & ~w21535 ) | ( w21533 & ~w21535 ) ;
  assign w21537 = ( w20247 & ~w21534 ) | ( w20247 & w21536 ) | ( ~w21534 & w21536 ) ;
  assign w21538 = \pi11 ^ w21537 ;
  assign w21539 = w21529 ^ w21530 ;
  assign w21540 = w21538 ^ w21539 ;
  assign w21541 = w21426 ^ w21430 ;
  assign w21542 = w21540 ^ w21541 ;
  assign w21543 = w21424 & ~w21542 ;
  assign w21544 = w21424 ^ w21542 ;
  assign w21545 = ( ~w21463 & w21471 ) | ( ~w21463 & w21472 ) | ( w21471 & w21472 ) ;
  assign w21546 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16646 ) | ( \pi31 & ~w16646 ) ;
  assign w21547 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21546 ) | ( ~\pi30 & w21546 ) ;
  assign w21548 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21546 ) | ( \pi30 & w21546 ) ;
  assign w21549 = ( \pi29 & w16648 ) | ( \pi29 & ~w21548 ) | ( w16648 & ~w21548 ) ;
  assign w21550 = ( ~w16644 & w21548 ) | ( ~w16644 & w21549 ) | ( w21548 & w21549 ) ;
  assign w21551 = ~\pi31 & w21550 ;
  assign w21552 = ( w21547 & ~w21549 ) | ( w21547 & w21551 ) | ( ~w21549 & w21551 ) ;
  assign w21553 = ( w37 & ~w17468 ) | ( w37 & w21552 ) | ( ~w17468 & w21552 ) ;
  assign w21554 = w21552 | w21553 ;
  assign w21555 = ( ~w21186 & w21441 ) | ( ~w21186 & w21459 ) | ( w21441 & w21459 ) ;
  assign w21556 = w980 | w1031 ;
  assign w21557 = w142 | w21556 ;
  assign w21558 = ( w74 & ~w142 ) | ( w74 & w388 ) | ( ~w142 & w388 ) ;
  assign w21559 = w21557 | w21558 ;
  assign w21560 = ( w361 & ~w505 ) | ( w361 & w21559 ) | ( ~w505 & w21559 ) ;
  assign w21561 = w4761 | w11473 ;
  assign w21562 = ( w505 & w1229 ) | ( w505 & ~w11473 ) | ( w1229 & ~w11473 ) ;
  assign w21563 = w21561 | w21562 ;
  assign w21564 = w21560 | w21563 ;
  assign w21565 = w3667 | w4784 ;
  assign w21566 = ( w1770 & w3667 ) | ( w1770 & ~w21564 ) | ( w3667 & ~w21564 ) ;
  assign w21567 = ~w21565 & w21566 ;
  assign w21568 = w220 | w2762 ;
  assign w21569 = ( ~w119 & w2762 ) | ( ~w119 & w21567 ) | ( w2762 & w21567 ) ;
  assign w21570 = ~w21568 & w21569 ;
  assign w21571 = ( w268 & w344 ) | ( w268 & ~w1001 ) | ( w344 & ~w1001 ) ;
  assign w21572 = ~w252 & w21570 ;
  assign w21573 = ( ~w252 & w1001 ) | ( ~w252 & w1030 ) | ( w1001 & w1030 ) ;
  assign w21574 = w21572 & ~w21573 ;
  assign w21575 = ~w21571 & w21574 ;
  assign w21576 = w21554 ^ w21555 ;
  assign w21577 = w21575 ^ w21576 ;
  assign w21578 = ( ~w21322 & w21439 ) | ( ~w21322 & w21461 ) | ( w21439 & w21461 ) ;
  assign w21579 = w3549 & ~w16638 ;
  assign w21580 = ( w3717 & w16640 ) | ( w3717 & w21579 ) | ( w16640 & w21579 ) ;
  assign w21581 = w3649 | w21580 ;
  assign w21582 = ( w16642 & w21580 ) | ( w16642 & w21581 ) | ( w21580 & w21581 ) ;
  assign w21583 = w21579 | w21582 ;
  assign w21584 = w3448 | w17783 ;
  assign w21585 = ( ~w17783 & w21583 ) | ( ~w17783 & w21584 ) | ( w21583 & w21584 ) ;
  assign w21586 = \pi29 ^ w21585 ;
  assign w21587 = w21577 ^ w21578 ;
  assign w21588 = w21586 ^ w21587 ;
  assign w21589 = w4143 | w16634 ;
  assign w21590 = w4052 & w16636 ;
  assign w21591 = ( ~w16634 & w21589 ) | ( ~w16634 & w21590 ) | ( w21589 & w21590 ) ;
  assign w21592 = w4147 | w18051 ;
  assign w21593 = w16632 | w21591 ;
  assign w21594 = ( w3964 & w21591 ) | ( w3964 & w21593 ) | ( w21591 & w21593 ) ;
  assign w21595 = ( ~w18051 & w21592 ) | ( ~w18051 & w21594 ) | ( w21592 & w21594 ) ;
  assign w21596 = \pi26 ^ w21595 ;
  assign w21597 = w21545 ^ w21588 ;
  assign w21598 = w21596 ^ w21597 ;
  assign w21599 = ( ~w21474 & w21482 ) | ( ~w21474 & w21483 ) | ( w21482 & w21483 ) ;
  assign w21600 = w4651 | w16628 ;
  assign w21601 = w4606 & ~w16630 ;
  assign w21602 = ( ~w16628 & w21600 ) | ( ~w16628 & w21601 ) | ( w21600 & w21601 ) ;
  assign w21603 = w4706 | w16626 ;
  assign w21604 = w18429 & ~w21602 ;
  assign w21605 = ( w4609 & w21602 ) | ( w4609 & ~w21604 ) | ( w21602 & ~w21604 ) ;
  assign w21606 = ( ~w16626 & w21603 ) | ( ~w16626 & w21605 ) | ( w21603 & w21605 ) ;
  assign w21607 = \pi23 ^ w21606 ;
  assign w21608 = w21598 ^ w21599 ;
  assign w21609 = w21607 ^ w21608 ;
  assign w21610 = ( ~w21485 & w21493 ) | ( ~w21485 & w21494 ) | ( w21493 & w21494 ) ;
  assign w21611 = ~w5343 & w16621 ;
  assign w21612 = w4905 & w16619 ;
  assign w21613 = ( w16621 & ~w21611 ) | ( w16621 & w21612 ) | ( ~w21611 & w21612 ) ;
  assign w21614 = ~w5395 & w16617 ;
  assign w21615 = w16732 | w21613 ;
  assign w21616 = ( w4908 & w21613 ) | ( w4908 & w21615 ) | ( w21613 & w21615 ) ;
  assign w21617 = ( w16617 & ~w21614 ) | ( w16617 & w21616 ) | ( ~w21614 & w21616 ) ;
  assign w21618 = \pi20 ^ w21617 ;
  assign w21619 = w21609 ^ w21610 ;
  assign w21620 = w21618 ^ w21619 ;
  assign w21621 = ( ~w21496 & w21504 ) | ( ~w21496 & w21505 ) | ( w21504 & w21505 ) ;
  assign w21622 = ~w5710 & w18916 ;
  assign w21623 = w5494 & ~w18914 ;
  assign w21624 = ( w18916 & ~w21622 ) | ( w18916 & w21623 ) | ( ~w21622 & w21623 ) ;
  assign w21625 = w5948 | w18912 ;
  assign w21626 = w18929 & ~w21624 ;
  assign w21627 = ( w5497 & w21624 ) | ( w5497 & ~w21626 ) | ( w21624 & ~w21626 ) ;
  assign w21628 = ( ~w18912 & w21625 ) | ( ~w18912 & w21627 ) | ( w21625 & w21627 ) ;
  assign w21629 = \pi17 ^ w21628 ;
  assign w21630 = w21620 ^ w21621 ;
  assign w21631 = w21629 ^ w21630 ;
  assign w21632 = ( ~w21507 & w21508 ) | ( ~w21507 & w21516 ) | ( w21508 & w21516 ) ;
  assign w21633 = ~w6549 & w19713 ;
  assign w21634 = w6048 & w19529 ;
  assign w21635 = ( w19713 & ~w21633 ) | ( w19713 & w21634 ) | ( ~w21633 & w21634 ) ;
  assign w21636 = ~w6637 & w19887 ;
  assign w21637 = w19898 | w21635 ;
  assign w21638 = ( w6045 & w21635 ) | ( w6045 & w21637 ) | ( w21635 & w21637 ) ;
  assign w21639 = ( w19887 & ~w21636 ) | ( w19887 & w21638 ) | ( ~w21636 & w21638 ) ;
  assign w21640 = \pi14 ^ w21639 ;
  assign w21641 = w21631 ^ w21632 ;
  assign w21642 = w21640 ^ w21641 ;
  assign w21643 = ( ~w21518 & w21526 ) | ( ~w21518 & w21527 ) | ( w21526 & w21527 ) ;
  assign w21644 = ~w6949 & w20247 ;
  assign w21645 = w6748 & ~w20068 ;
  assign w21646 = ( w20247 & ~w21644 ) | ( w20247 & w21645 ) | ( ~w21644 & w21645 ) ;
  assign w21647 = ~w7154 & w20404 ;
  assign w21648 = w20417 | w21646 ;
  assign w21649 = ( w6751 & w21646 ) | ( w6751 & w21648 ) | ( w21646 & w21648 ) ;
  assign w21650 = ( w20404 & ~w21647 ) | ( w20404 & w21649 ) | ( ~w21647 & w21649 ) ;
  assign w21651 = \pi11 ^ w21650 ;
  assign w21652 = w21642 ^ w21643 ;
  assign w21653 = w21651 ^ w21652 ;
  assign w21654 = ( ~w21529 & w21530 ) | ( ~w21529 & w21538 ) | ( w21530 & w21538 ) ;
  assign w21655 = ( w21426 & w21430 ) | ( w21426 & ~w21540 ) | ( w21430 & ~w21540 ) ;
  assign w21656 = w21653 ^ w21655 ;
  assign w21657 = w21654 ^ w21656 ;
  assign w21658 = w21543 ^ w21657 ;
  assign w21659 = ( ~w21577 & w21578 ) | ( ~w21577 & w21586 ) | ( w21578 & w21586 ) ;
  assign w21660 = ( w21554 & ~w21555 ) | ( w21554 & w21575 ) | ( ~w21555 & w21575 ) ;
  assign w21661 = w259 | w277 ;
  assign w21662 = w135 | w21661 ;
  assign w21663 = ( ~w135 & w147 ) | ( ~w135 & w2147 ) | ( w147 & w2147 ) ;
  assign w21664 = w21662 | w21663 ;
  assign w21665 = ( w390 & w491 ) | ( w390 & ~w534 ) | ( w491 & ~w534 ) ;
  assign w21666 = w890 | w21664 ;
  assign w21667 = ( w534 & w680 ) | ( w534 & ~w890 ) | ( w680 & ~w890 ) ;
  assign w21668 = w21666 | w21667 ;
  assign w21669 = w21665 | w21668 ;
  assign w21670 = ( ~w273 & w12166 ) | ( ~w273 & w21669 ) | ( w12166 & w21669 ) ;
  assign w21671 = w5255 | w10998 ;
  assign w21672 = ( w273 & w2782 ) | ( w273 & ~w10998 ) | ( w2782 & ~w10998 ) ;
  assign w21673 = w21671 | w21672 ;
  assign w21674 = w21670 | w21673 ;
  assign w21675 = w1275 | w1363 ;
  assign w21676 = w21163 | w21675 ;
  assign w21677 = ( w742 & ~w21163 ) | ( w742 & w21674 ) | ( ~w21163 & w21674 ) ;
  assign w21678 = w21676 | w21677 ;
  assign w21679 = ( w274 & w415 ) | ( w274 & ~w420 ) | ( w415 & ~w420 ) ;
  assign w21680 = w68 | w21678 ;
  assign w21681 = ( ~w68 & w420 ) | ( ~w68 & w530 ) | ( w420 & w530 ) ;
  assign w21682 = w21680 | w21681 ;
  assign w21683 = w21679 | w21682 ;
  assign w21684 = ( w21575 & w21660 ) | ( w21575 & w21683 ) | ( w21660 & w21683 ) ;
  assign w21685 = w21575 ^ w21660 ;
  assign w21686 = w21683 ^ w21685 ;
  assign w21687 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16644 ) | ( \pi31 & ~w16644 ) ;
  assign w21688 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21687 ) | ( ~\pi30 & w21687 ) ;
  assign w21689 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21687 ) | ( \pi30 & w21687 ) ;
  assign w21690 = ( \pi29 & w16646 ) | ( \pi29 & ~w21689 ) | ( w16646 & ~w21689 ) ;
  assign w21691 = ( w16642 & w21689 ) | ( w16642 & w21690 ) | ( w21689 & w21690 ) ;
  assign w21692 = ~\pi31 & w21691 ;
  assign w21693 = ( w21688 & ~w21690 ) | ( w21688 & w21692 ) | ( ~w21690 & w21692 ) ;
  assign w21694 = ( w37 & w17455 ) | ( w37 & w21693 ) | ( w17455 & w21693 ) ;
  assign w21695 = w21693 | w21694 ;
  assign w21696 = w3549 & w16636 ;
  assign w21697 = ( w3717 & ~w16638 ) | ( w3717 & w21696 ) | ( ~w16638 & w21696 ) ;
  assign w21698 = w3649 | w21697 ;
  assign w21699 = ( w16640 & w21697 ) | ( w16640 & w21698 ) | ( w21697 & w21698 ) ;
  assign w21700 = w21696 | w21699 ;
  assign w21701 = w3448 | w17770 ;
  assign w21702 = ( ~w17770 & w21700 ) | ( ~w17770 & w21701 ) | ( w21700 & w21701 ) ;
  assign w21703 = \pi29 ^ w21702 ;
  assign w21704 = w21686 ^ w21703 ;
  assign w21705 = w21695 ^ w21704 ;
  assign w21706 = ~w4143 & w16632 ;
  assign w21707 = w4052 & ~w16634 ;
  assign w21708 = ( w16632 & ~w21706 ) | ( w16632 & w21707 ) | ( ~w21706 & w21707 ) ;
  assign w21709 = w4147 | w18038 ;
  assign w21710 = w16630 & ~w21708 ;
  assign w21711 = ( w3964 & w21708 ) | ( w3964 & ~w21710 ) | ( w21708 & ~w21710 ) ;
  assign w21712 = ( ~w18038 & w21709 ) | ( ~w18038 & w21711 ) | ( w21709 & w21711 ) ;
  assign w21713 = \pi26 ^ w21712 ;
  assign w21714 = w21659 ^ w21705 ;
  assign w21715 = w21713 ^ w21714 ;
  assign w21716 = ( w21545 & ~w21588 ) | ( w21545 & w21596 ) | ( ~w21588 & w21596 ) ;
  assign w21717 = w4651 | w16626 ;
  assign w21718 = w4606 & ~w16628 ;
  assign w21719 = ( ~w16626 & w21717 ) | ( ~w16626 & w21718 ) | ( w21717 & w21718 ) ;
  assign w21720 = ~w4706 & w16619 ;
  assign w21721 = w18451 | w21719 ;
  assign w21722 = ( w4609 & w21719 ) | ( w4609 & w21721 ) | ( w21719 & w21721 ) ;
  assign w21723 = ( w16619 & ~w21720 ) | ( w16619 & w21722 ) | ( ~w21720 & w21722 ) ;
  assign w21724 = \pi23 ^ w21723 ;
  assign w21725 = w21715 ^ w21716 ;
  assign w21726 = w21724 ^ w21725 ;
  assign w21727 = ( ~w21598 & w21599 ) | ( ~w21598 & w21607 ) | ( w21599 & w21607 ) ;
  assign w21728 = ~w5343 & w16617 ;
  assign w21729 = w4905 & w16621 ;
  assign w21730 = ( w16617 & ~w21728 ) | ( w16617 & w21729 ) | ( ~w21728 & w21729 ) ;
  assign w21731 = w5395 | w18914 ;
  assign w21732 = w19350 & ~w21730 ;
  assign w21733 = ( w4908 & w21730 ) | ( w4908 & ~w21732 ) | ( w21730 & ~w21732 ) ;
  assign w21734 = ( ~w18914 & w21731 ) | ( ~w18914 & w21733 ) | ( w21731 & w21733 ) ;
  assign w21735 = \pi20 ^ w21734 ;
  assign w21736 = w21726 ^ w21727 ;
  assign w21737 = w21735 ^ w21736 ;
  assign w21738 = ( ~w21609 & w21610 ) | ( ~w21609 & w21618 ) | ( w21610 & w21618 ) ;
  assign w21739 = w5710 | w18912 ;
  assign w21740 = w5494 & w18916 ;
  assign w21741 = ( ~w18912 & w21739 ) | ( ~w18912 & w21740 ) | ( w21739 & w21740 ) ;
  assign w21742 = ~w5948 & w19529 ;
  assign w21743 = w19540 & ~w21741 ;
  assign w21744 = ( w5497 & w21741 ) | ( w5497 & ~w21743 ) | ( w21741 & ~w21743 ) ;
  assign w21745 = ( w19529 & ~w21742 ) | ( w19529 & w21744 ) | ( ~w21742 & w21744 ) ;
  assign w21746 = \pi17 ^ w21745 ;
  assign w21747 = w21737 ^ w21738 ;
  assign w21748 = w21746 ^ w21747 ;
  assign w21749 = ( ~w21620 & w21621 ) | ( ~w21620 & w21629 ) | ( w21621 & w21629 ) ;
  assign w21750 = ~w6549 & w19887 ;
  assign w21751 = w6048 & w19713 ;
  assign w21752 = ( w19887 & ~w21750 ) | ( w19887 & w21751 ) | ( ~w21750 & w21751 ) ;
  assign w21753 = w6637 | w20068 ;
  assign w21754 = w20081 & ~w21752 ;
  assign w21755 = ( w6045 & w21752 ) | ( w6045 & ~w21754 ) | ( w21752 & ~w21754 ) ;
  assign w21756 = ( ~w20068 & w21753 ) | ( ~w20068 & w21755 ) | ( w21753 & w21755 ) ;
  assign w21757 = \pi14 ^ w21756 ;
  assign w21758 = w21748 ^ w21749 ;
  assign w21759 = w21757 ^ w21758 ;
  assign w21760 = ( ~w21631 & w21632 ) | ( ~w21631 & w21640 ) | ( w21632 & w21640 ) ;
  assign w21761 = w7154 & w20404 ;
  assign w21762 = ( w6949 & w20404 ) | ( w6949 & w21761 ) | ( w20404 & w21761 ) ;
  assign w21763 = w6748 & w20247 ;
  assign w21764 = w21762 | w21763 ;
  assign w21765 = w6751 & ~w20414 ;
  assign w21766 = ( w6751 & w21764 ) | ( w6751 & ~w21765 ) | ( w21764 & ~w21765 ) ;
  assign w21767 = w21759 ^ w21766 ;
  assign w21768 = \pi11 ^ w21760 ;
  assign w21769 = w21767 ^ w21768 ;
  assign w21770 = ( ~w21642 & w21643 ) | ( ~w21642 & w21651 ) | ( w21643 & w21651 ) ;
  assign w21771 = ( ~w21653 & w21654 ) | ( ~w21653 & w21655 ) | ( w21654 & w21655 ) ;
  assign w21772 = w21769 ^ w21771 ;
  assign w21773 = w21770 ^ w21772 ;
  assign w21774 = w21543 & ~w21657 ;
  assign w21775 = w21773 & w21774 ;
  assign w21776 = w21773 ^ w21774 ;
  assign w21777 = ( w21769 & w21770 ) | ( w21769 & w21771 ) | ( w21770 & w21771 ) ;
  assign w21778 = w20414 | w21764 ;
  assign w21779 = ( w6751 & w21764 ) | ( w6751 & w21778 ) | ( w21764 & w21778 ) ;
  assign w21780 = \pi11 ^ w21779 ;
  assign w21781 = ( w21759 & w21760 ) | ( w21759 & w21780 ) | ( w21760 & w21780 ) ;
  assign w21782 = ( w21686 & w21695 ) | ( w21686 & w21703 ) | ( w21695 & w21703 ) ;
  assign w21783 = ( \pi29 & \pi31 ) | ( \pi29 & w16642 ) | ( \pi31 & w16642 ) ;
  assign w21784 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21783 ) | ( ~\pi30 & w21783 ) ;
  assign w21785 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21783 ) | ( \pi30 & w21783 ) ;
  assign w21786 = ( \pi29 & w16644 ) | ( \pi29 & ~w21785 ) | ( w16644 & ~w21785 ) ;
  assign w21787 = ( w16640 & w21785 ) | ( w16640 & w21786 ) | ( w21785 & w21786 ) ;
  assign w21788 = ~\pi31 & w21787 ;
  assign w21789 = ( w21784 & ~w21786 ) | ( w21784 & w21788 ) | ( ~w21786 & w21788 ) ;
  assign w21790 = ( w37 & ~w17760 ) | ( w37 & w21789 ) | ( ~w17760 & w21789 ) ;
  assign w21791 = w21789 | w21790 ;
  assign w21792 = w11496 ^ w20404 ;
  assign w21793 = ( \pi11 & w11496 ) | ( \pi11 & ~w21792 ) | ( w11496 & ~w21792 ) ;
  assign w21794 = ( w113 & w169 ) | ( w113 & ~w570 ) | ( w169 & ~w570 ) ;
  assign w21795 = w2257 | w4985 ;
  assign w21796 = ( w570 & w901 ) | ( w570 & ~w4985 ) | ( w901 & ~w4985 ) ;
  assign w21797 = w21795 | w21796 ;
  assign w21798 = w21794 | w21797 ;
  assign w21799 = ( ~w218 & w4964 ) | ( ~w218 & w21798 ) | ( w4964 & w21798 ) ;
  assign w21800 = w1443 & ~w3616 ;
  assign w21801 = ( w218 & w219 ) | ( w218 & w1443 ) | ( w219 & w1443 ) ;
  assign w21802 = w21800 & ~w21801 ;
  assign w21803 = ~w21799 & w21802 ;
  assign w21804 = ( w594 & w1281 ) | ( w594 & ~w1617 ) | ( w1281 & ~w1617 ) ;
  assign w21805 = ~w1472 & w21803 ;
  assign w21806 = ( ~w1472 & w1617 ) | ( ~w1472 & w3965 ) | ( w1617 & w3965 ) ;
  assign w21807 = w21805 & ~w21806 ;
  assign w21808 = ~w21804 & w21807 ;
  assign w21809 = w429 | w531 ;
  assign w21810 = w220 | w21809 ;
  assign w21811 = ( w220 & ~w350 ) | ( w220 & w21808 ) | ( ~w350 & w21808 ) ;
  assign w21812 = ~w21810 & w21811 ;
  assign w21813 = w21575 ^ w21793 ;
  assign w21814 = w21812 ^ w21813 ;
  assign w21815 = w21684 ^ w21814 ;
  assign w21816 = w21791 ^ w21815 ;
  assign w21817 = ~w3717 & w16636 ;
  assign w21818 = w3649 & ~w16638 ;
  assign w21819 = ( w16636 & ~w21817 ) | ( w16636 & w21818 ) | ( ~w21817 & w21818 ) ;
  assign w21820 = w3549 | w16634 ;
  assign w21821 = w16742 & ~w21819 ;
  assign w21822 = ( w3448 & w21819 ) | ( w3448 & ~w21821 ) | ( w21819 & ~w21821 ) ;
  assign w21823 = ( ~w16634 & w21820 ) | ( ~w16634 & w21822 ) | ( w21820 & w21822 ) ;
  assign w21824 = \pi29 ^ w21823 ;
  assign w21825 = w21782 ^ w21816 ;
  assign w21826 = w21824 ^ w21825 ;
  assign w21827 = w4143 | w16630 ;
  assign w21828 = w4052 & w16632 ;
  assign w21829 = ( ~w16630 & w21827 ) | ( ~w16630 & w21828 ) | ( w21827 & w21828 ) ;
  assign w21830 = ~w4147 & w18026 ;
  assign w21831 = w16628 & ~w21829 ;
  assign w21832 = ( w3964 & w21829 ) | ( w3964 & ~w21831 ) | ( w21829 & ~w21831 ) ;
  assign w21833 = ( w18026 & ~w21830 ) | ( w18026 & w21832 ) | ( ~w21830 & w21832 ) ;
  assign w21834 = \pi26 ^ w21833 ;
  assign w21835 = ( w21659 & w21705 ) | ( w21659 & w21713 ) | ( w21705 & w21713 ) ;
  assign w21836 = w21826 ^ w21835 ;
  assign w21837 = w21834 ^ w21836 ;
  assign w21838 = ~w4651 & w16619 ;
  assign w21839 = w4606 & ~w16626 ;
  assign w21840 = ( w16619 & ~w21838 ) | ( w16619 & w21839 ) | ( ~w21838 & w21839 ) ;
  assign w21841 = ~w4706 & w16621 ;
  assign w21842 = w18439 & ~w21840 ;
  assign w21843 = ( w4609 & w21840 ) | ( w4609 & ~w21842 ) | ( w21840 & ~w21842 ) ;
  assign w21844 = ( w16621 & ~w21841 ) | ( w16621 & w21843 ) | ( ~w21841 & w21843 ) ;
  assign w21845 = \pi23 ^ w21844 ;
  assign w21846 = ( w21715 & w21716 ) | ( w21715 & w21724 ) | ( w21716 & w21724 ) ;
  assign w21847 = w21837 ^ w21846 ;
  assign w21848 = w21845 ^ w21847 ;
  assign w21849 = ( w21726 & w21727 ) | ( w21726 & w21735 ) | ( w21727 & w21735 ) ;
  assign w21850 = w5343 | w18914 ;
  assign w21851 = w4905 & w16617 ;
  assign w21852 = ( ~w18914 & w21850 ) | ( ~w18914 & w21851 ) | ( w21850 & w21851 ) ;
  assign w21853 = ~w5395 & w18916 ;
  assign w21854 = w19366 & ~w21852 ;
  assign w21855 = ( w4908 & w21852 ) | ( w4908 & ~w21854 ) | ( w21852 & ~w21854 ) ;
  assign w21856 = ( w18916 & ~w21853 ) | ( w18916 & w21855 ) | ( ~w21853 & w21855 ) ;
  assign w21857 = \pi20 ^ w21856 ;
  assign w21858 = w21848 ^ w21849 ;
  assign w21859 = w21857 ^ w21858 ;
  assign w21860 = ~w5710 & w19529 ;
  assign w21861 = w5494 & ~w18912 ;
  assign w21862 = ( w19529 & ~w21860 ) | ( w19529 & w21861 ) | ( ~w21860 & w21861 ) ;
  assign w21863 = ~w5948 & w19713 ;
  assign w21864 = w19723 | w21862 ;
  assign w21865 = ( w5497 & w21862 ) | ( w5497 & w21864 ) | ( w21862 & w21864 ) ;
  assign w21866 = ( w19713 & ~w21863 ) | ( w19713 & w21865 ) | ( ~w21863 & w21865 ) ;
  assign w21867 = \pi17 ^ w21866 ;
  assign w21868 = ( w21737 & w21738 ) | ( w21737 & w21746 ) | ( w21738 & w21746 ) ;
  assign w21869 = w21859 ^ w21868 ;
  assign w21870 = w21867 ^ w21869 ;
  assign w21871 = ( w21748 & w21749 ) | ( w21748 & w21757 ) | ( w21749 & w21757 ) ;
  assign w21872 = w6549 | w20068 ;
  assign w21873 = w6048 & w19887 ;
  assign w21874 = ( ~w20068 & w21872 ) | ( ~w20068 & w21873 ) | ( w21872 & w21873 ) ;
  assign w21875 = ~w6637 & w20247 ;
  assign w21876 = w20257 & ~w21874 ;
  assign w21877 = ( w6045 & w21874 ) | ( w6045 & ~w21876 ) | ( w21874 & ~w21876 ) ;
  assign w21878 = ( w20247 & ~w21875 ) | ( w20247 & w21877 ) | ( ~w21875 & w21877 ) ;
  assign w21879 = \pi14 ^ w21878 ;
  assign w21880 = w21870 ^ w21871 ;
  assign w21881 = w21879 ^ w21880 ;
  assign w21882 = w21777 ^ w21781 ;
  assign w21883 = w21881 ^ w21882 ;
  assign w21884 = w21775 & ~w21883 ;
  assign w21885 = w21775 ^ w21883 ;
  assign w21886 = ( w21782 & ~w21816 ) | ( w21782 & w21824 ) | ( ~w21816 & w21824 ) ;
  assign w21887 = ( \pi29 & \pi31 ) | ( \pi29 & w16640 ) | ( \pi31 & w16640 ) ;
  assign w21888 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21887 ) | ( ~\pi30 & w21887 ) ;
  assign w21889 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21887 ) | ( \pi30 & w21887 ) ;
  assign w21890 = ( ~\pi29 & w16642 ) | ( ~\pi29 & w21889 ) | ( w16642 & w21889 ) ;
  assign w21891 = ( w16638 & ~w21889 ) | ( w16638 & w21890 ) | ( ~w21889 & w21890 ) ;
  assign w21892 = \pi31 | w21891 ;
  assign w21893 = ( w21888 & w21890 ) | ( w21888 & ~w21892 ) | ( w21890 & ~w21892 ) ;
  assign w21894 = ( w37 & ~w17783 ) | ( w37 & w21893 ) | ( ~w17783 & w21893 ) ;
  assign w21895 = w21893 | w21894 ;
  assign w21896 = ( w21575 & w21793 ) | ( w21575 & w21812 ) | ( w21793 & w21812 ) ;
  assign w21897 = w512 | w764 ;
  assign w21898 = w164 | w21897 ;
  assign w21899 = ( w122 & ~w164 ) | ( w122 & w419 ) | ( ~w164 & w419 ) ;
  assign w21900 = w21898 | w21899 ;
  assign w21901 = w3971 | w21900 ;
  assign w21902 = ( w320 & w624 ) | ( w320 & ~w21900 ) | ( w624 & ~w21900 ) ;
  assign w21903 = w21901 | w21902 ;
  assign w21904 = ( w20142 & w20470 ) | ( w20142 & ~w21903 ) | ( w20470 & ~w21903 ) ;
  assign w21905 = w10758 | w12181 ;
  assign w21906 = ( w10310 & ~w12181 ) | ( w10310 & w21903 ) | ( ~w12181 & w21903 ) ;
  assign w21907 = w21905 | w21906 ;
  assign w21908 = w21904 | w21907 ;
  assign w21909 = w466 | w822 ;
  assign w21910 = ( ~w822 & w1413 ) | ( ~w822 & w21908 ) | ( w1413 & w21908 ) ;
  assign w21911 = w21909 | w21910 ;
  assign w21912 = w758 | w1128 ;
  assign w21913 = w386 | w21912 ;
  assign w21914 = ( ~w386 & w467 ) | ( ~w386 & w21911 ) | ( w467 & w21911 ) ;
  assign w21915 = w21913 | w21914 ;
  assign w21916 = w21895 ^ w21896 ;
  assign w21917 = w21915 ^ w21916 ;
  assign w21918 = ( w21684 & w21791 ) | ( w21684 & ~w21814 ) | ( w21791 & ~w21814 ) ;
  assign w21919 = w3549 & w16632 ;
  assign w21920 = ( w3717 & ~w16634 ) | ( w3717 & w21919 ) | ( ~w16634 & w21919 ) ;
  assign w21921 = w3649 | w21920 ;
  assign w21922 = ( w16636 & w21920 ) | ( w16636 & w21921 ) | ( w21920 & w21921 ) ;
  assign w21923 = w21919 | w21922 ;
  assign w21924 = w3448 | w18051 ;
  assign w21925 = ( ~w18051 & w21923 ) | ( ~w18051 & w21924 ) | ( w21923 & w21924 ) ;
  assign w21926 = \pi29 ^ w21925 ;
  assign w21927 = w21917 ^ w21918 ;
  assign w21928 = w21926 ^ w21927 ;
  assign w21929 = w4143 | w16628 ;
  assign w21930 = w4052 & ~w16630 ;
  assign w21931 = ( ~w16628 & w21929 ) | ( ~w16628 & w21930 ) | ( w21929 & w21930 ) ;
  assign w21932 = w4147 | w18429 ;
  assign w21933 = w16626 & ~w21931 ;
  assign w21934 = ( w3964 & w21931 ) | ( w3964 & ~w21933 ) | ( w21931 & ~w21933 ) ;
  assign w21935 = ( ~w18429 & w21932 ) | ( ~w18429 & w21934 ) | ( w21932 & w21934 ) ;
  assign w21936 = \pi26 ^ w21935 ;
  assign w21937 = w21886 ^ w21928 ;
  assign w21938 = w21936 ^ w21937 ;
  assign w21939 = ( ~w21826 & w21834 ) | ( ~w21826 & w21835 ) | ( w21834 & w21835 ) ;
  assign w21940 = ~w4651 & w16621 ;
  assign w21941 = w4606 & w16619 ;
  assign w21942 = ( w16621 & ~w21940 ) | ( w16621 & w21941 ) | ( ~w21940 & w21941 ) ;
  assign w21943 = ~w4706 & w16617 ;
  assign w21944 = w16732 | w21942 ;
  assign w21945 = ( w4609 & w21942 ) | ( w4609 & w21944 ) | ( w21942 & w21944 ) ;
  assign w21946 = ( w16617 & ~w21943 ) | ( w16617 & w21945 ) | ( ~w21943 & w21945 ) ;
  assign w21947 = \pi23 ^ w21946 ;
  assign w21948 = w21938 ^ w21939 ;
  assign w21949 = w21947 ^ w21948 ;
  assign w21950 = ( ~w21837 & w21845 ) | ( ~w21837 & w21846 ) | ( w21845 & w21846 ) ;
  assign w21951 = ~w5343 & w18916 ;
  assign w21952 = w4905 & ~w18914 ;
  assign w21953 = ( w18916 & ~w21951 ) | ( w18916 & w21952 ) | ( ~w21951 & w21952 ) ;
  assign w21954 = w5395 | w18912 ;
  assign w21955 = w18929 & ~w21953 ;
  assign w21956 = ( w4908 & w21953 ) | ( w4908 & ~w21955 ) | ( w21953 & ~w21955 ) ;
  assign w21957 = ( ~w18912 & w21954 ) | ( ~w18912 & w21956 ) | ( w21954 & w21956 ) ;
  assign w21958 = \pi20 ^ w21957 ;
  assign w21959 = w21949 ^ w21950 ;
  assign w21960 = w21958 ^ w21959 ;
  assign w21961 = ( ~w21848 & w21849 ) | ( ~w21848 & w21857 ) | ( w21849 & w21857 ) ;
  assign w21962 = ~w5710 & w19713 ;
  assign w21963 = w5494 & w19529 ;
  assign w21964 = ( w19713 & ~w21962 ) | ( w19713 & w21963 ) | ( ~w21962 & w21963 ) ;
  assign w21965 = ~w5948 & w19887 ;
  assign w21966 = w19898 | w21964 ;
  assign w21967 = ( w5497 & w21964 ) | ( w5497 & w21966 ) | ( w21964 & w21966 ) ;
  assign w21968 = ( w19887 & ~w21965 ) | ( w19887 & w21967 ) | ( ~w21965 & w21967 ) ;
  assign w21969 = \pi17 ^ w21968 ;
  assign w21970 = w21960 ^ w21961 ;
  assign w21971 = w21969 ^ w21970 ;
  assign w21972 = ( ~w21859 & w21867 ) | ( ~w21859 & w21868 ) | ( w21867 & w21868 ) ;
  assign w21973 = ~w6549 & w20247 ;
  assign w21974 = w6048 & ~w20068 ;
  assign w21975 = ( w20247 & ~w21973 ) | ( w20247 & w21974 ) | ( ~w21973 & w21974 ) ;
  assign w21976 = ~w6637 & w20404 ;
  assign w21977 = w20417 | w21975 ;
  assign w21978 = ( w6045 & w21975 ) | ( w6045 & w21977 ) | ( w21975 & w21977 ) ;
  assign w21979 = ( w20404 & ~w21976 ) | ( w20404 & w21978 ) | ( ~w21976 & w21978 ) ;
  assign w21980 = \pi14 ^ w21979 ;
  assign w21981 = w21971 ^ w21972 ;
  assign w21982 = w21980 ^ w21981 ;
  assign w21983 = ( ~w21870 & w21871 ) | ( ~w21870 & w21879 ) | ( w21871 & w21879 ) ;
  assign w21984 = ( w21777 & w21781 ) | ( w21777 & ~w21881 ) | ( w21781 & ~w21881 ) ;
  assign w21985 = w21982 ^ w21984 ;
  assign w21986 = w21983 ^ w21985 ;
  assign w21987 = w21884 ^ w21986 ;
  assign w21988 = w21884 & w21986 ;
  assign w21989 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16638 ) | ( \pi31 & ~w16638 ) ;
  assign w21990 = ( \pi29 & ~\pi30 ) | ( \pi29 & w21989 ) | ( ~\pi30 & w21989 ) ;
  assign w21991 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w21989 ) | ( \pi30 & w21989 ) ;
  assign w21992 = ( ~\pi29 & w16640 ) | ( ~\pi29 & w21991 ) | ( w16640 & w21991 ) ;
  assign w21993 = ( w16636 & w21991 ) | ( w16636 & ~w21992 ) | ( w21991 & ~w21992 ) ;
  assign w21994 = ~\pi31 & w21993 ;
  assign w21995 = ( w21990 & w21992 ) | ( w21990 & w21994 ) | ( w21992 & w21994 ) ;
  assign w21996 = ( w37 & ~w17770 ) | ( w37 & w21995 ) | ( ~w17770 & w21995 ) ;
  assign w21997 = w21995 | w21996 ;
  assign w21998 = ( w114 & w230 ) | ( w114 & ~w277 ) | ( w230 & ~w277 ) ;
  assign w21999 = w2259 | w3190 ;
  assign w22000 = ( w277 & w385 ) | ( w277 & ~w2259 ) | ( w385 & ~w2259 ) ;
  assign w22001 = w21999 | w22000 ;
  assign w22002 = w21998 | w22001 ;
  assign w22003 = ( w3468 & w5161 ) | ( w3468 & w10473 ) | ( w5161 & w10473 ) ;
  assign w22004 = w2618 | w22002 ;
  assign w22005 = ( w2618 & w5161 ) | ( w2618 & ~w10076 ) | ( w5161 & ~w10076 ) ;
  assign w22006 = ~w22004 & w22005 ;
  assign w22007 = ~w22003 & w22006 ;
  assign w22008 = ( w317 & w561 ) | ( w317 & ~w663 ) | ( w561 & ~w663 ) ;
  assign w22009 = ~w125 & w22007 ;
  assign w22010 = ( ~w125 & w663 ) | ( ~w125 & w1128 ) | ( w663 & w1128 ) ;
  assign w22011 = w22009 & ~w22010 ;
  assign w22012 = ~w22008 & w22011 ;
  assign w22013 = ( w179 & w225 ) | ( w179 & ~w344 ) | ( w225 & ~w344 ) ;
  assign w22014 = ~w44 & w22012 ;
  assign w22015 = ( ~w44 & w344 ) | ( ~w44 & w430 ) | ( w344 & w430 ) ;
  assign w22016 = w22014 & ~w22015 ;
  assign w22017 = ~w22013 & w22016 ;
  assign w22018 = ( w21915 & ~w21997 ) | ( w21915 & w22017 ) | ( ~w21997 & w22017 ) ;
  assign w22019 = w21997 ^ w22017 ;
  assign w22020 = w21915 ^ w22019 ;
  assign w22021 = ( ~w21895 & w21896 ) | ( ~w21895 & w21915 ) | ( w21896 & w21915 ) ;
  assign w22022 = ( w21917 & w21918 ) | ( w21917 & w21926 ) | ( w21918 & w21926 ) ;
  assign w22023 = w22021 ^ w22022 ;
  assign w22024 = w22020 ^ w22023 ;
  assign w22025 = ~w3717 & w16632 ;
  assign w22026 = w3649 & ~w16634 ;
  assign w22027 = ( w16632 & ~w22025 ) | ( w16632 & w22026 ) | ( ~w22025 & w22026 ) ;
  assign w22028 = w3549 | w16630 ;
  assign w22029 = w18038 & ~w22027 ;
  assign w22030 = ( w3448 & w22027 ) | ( w3448 & ~w22029 ) | ( w22027 & ~w22029 ) ;
  assign w22031 = ( ~w16630 & w22028 ) | ( ~w16630 & w22030 ) | ( w22028 & w22030 ) ;
  assign w22032 = \pi29 ^ w22031 ;
  assign w22033 = w4143 | w16626 ;
  assign w22034 = w4052 & ~w16628 ;
  assign w22035 = ( ~w16626 & w22033 ) | ( ~w16626 & w22034 ) | ( w22033 & w22034 ) ;
  assign w22036 = ~w4147 & w18451 ;
  assign w22037 = w16619 | w22035 ;
  assign w22038 = ( w3964 & w22035 ) | ( w3964 & w22037 ) | ( w22035 & w22037 ) ;
  assign w22039 = ( w18451 & ~w22036 ) | ( w18451 & w22038 ) | ( ~w22036 & w22038 ) ;
  assign w22040 = \pi26 ^ w22039 ;
  assign w22041 = w22024 ^ w22040 ;
  assign w22042 = w22032 ^ w22041 ;
  assign w22043 = ( w21886 & w21928 ) | ( w21886 & w21936 ) | ( w21928 & w21936 ) ;
  assign w22044 = ~w4651 & w16617 ;
  assign w22045 = w4606 & w16621 ;
  assign w22046 = ( w16617 & ~w22044 ) | ( w16617 & w22045 ) | ( ~w22044 & w22045 ) ;
  assign w22047 = w4706 | w18914 ;
  assign w22048 = w19350 & ~w22046 ;
  assign w22049 = ( w4609 & w22046 ) | ( w4609 & ~w22048 ) | ( w22046 & ~w22048 ) ;
  assign w22050 = ( ~w18914 & w22047 ) | ( ~w18914 & w22049 ) | ( w22047 & w22049 ) ;
  assign w22051 = \pi23 ^ w22050 ;
  assign w22052 = w22042 ^ w22043 ;
  assign w22053 = w22051 ^ w22052 ;
  assign w22054 = ( w21938 & w21939 ) | ( w21938 & w21947 ) | ( w21939 & w21947 ) ;
  assign w22055 = w5343 | w18912 ;
  assign w22056 = w4905 & w18916 ;
  assign w22057 = ( ~w18912 & w22055 ) | ( ~w18912 & w22056 ) | ( w22055 & w22056 ) ;
  assign w22058 = ~w5395 & w19529 ;
  assign w22059 = w19540 & ~w22057 ;
  assign w22060 = ( w4908 & w22057 ) | ( w4908 & ~w22059 ) | ( w22057 & ~w22059 ) ;
  assign w22061 = ( w19529 & ~w22058 ) | ( w19529 & w22060 ) | ( ~w22058 & w22060 ) ;
  assign w22062 = \pi20 ^ w22061 ;
  assign w22063 = w22053 ^ w22054 ;
  assign w22064 = w22062 ^ w22063 ;
  assign w22065 = ( w21949 & w21950 ) | ( w21949 & w21958 ) | ( w21950 & w21958 ) ;
  assign w22066 = ~w5710 & w19887 ;
  assign w22067 = w5494 & w19713 ;
  assign w22068 = ( w19887 & ~w22066 ) | ( w19887 & w22067 ) | ( ~w22066 & w22067 ) ;
  assign w22069 = w5948 | w20068 ;
  assign w22070 = w20081 & ~w22068 ;
  assign w22071 = ( w5497 & w22068 ) | ( w5497 & ~w22070 ) | ( w22068 & ~w22070 ) ;
  assign w22072 = ( ~w20068 & w22069 ) | ( ~w20068 & w22071 ) | ( w22069 & w22071 ) ;
  assign w22073 = \pi17 ^ w22072 ;
  assign w22074 = w22064 ^ w22065 ;
  assign w22075 = w22073 ^ w22074 ;
  assign w22076 = ( w21960 & w21961 ) | ( w21960 & w21969 ) | ( w21961 & w21969 ) ;
  assign w22077 = w6637 & w20404 ;
  assign w22078 = ( w6549 & w20404 ) | ( w6549 & w22077 ) | ( w20404 & w22077 ) ;
  assign w22079 = w6048 & w20247 ;
  assign w22080 = w22078 | w22079 ;
  assign w22081 = w6045 & ~w20414 ;
  assign w22082 = ( w6045 & w22080 ) | ( w6045 & ~w22081 ) | ( w22080 & ~w22081 ) ;
  assign w22083 = w22075 ^ w22082 ;
  assign w22084 = \pi14 ^ w22076 ;
  assign w22085 = w22083 ^ w22084 ;
  assign w22086 = ( w21971 & w21972 ) | ( w21971 & w21980 ) | ( w21972 & w21980 ) ;
  assign w22087 = ( w21982 & w21983 ) | ( w21982 & w21984 ) | ( w21983 & w21984 ) ;
  assign w22088 = w22085 ^ w22087 ;
  assign w22089 = w22086 ^ w22088 ;
  assign w22090 = w21988 & ~w22089 ;
  assign w22091 = w21988 ^ w22089 ;
  assign w22092 = ( ~w22085 & w22086 ) | ( ~w22085 & w22087 ) | ( w22086 & w22087 ) ;
  assign w22093 = w20414 | w22080 ;
  assign w22094 = ( w6045 & w22080 ) | ( w6045 & w22093 ) | ( w22080 & w22093 ) ;
  assign w22095 = \pi14 ^ w22094 ;
  assign w22096 = ( ~w22075 & w22076 ) | ( ~w22075 & w22095 ) | ( w22076 & w22095 ) ;
  assign w22097 = ( \pi29 & \pi31 ) | ( \pi29 & w16636 ) | ( \pi31 & w16636 ) ;
  assign w22098 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22097 ) | ( ~\pi30 & w22097 ) ;
  assign w22099 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22097 ) | ( \pi30 & w22097 ) ;
  assign w22100 = ( \pi29 & w16638 ) | ( \pi29 & ~w22099 ) | ( w16638 & ~w22099 ) ;
  assign w22101 = ( ~w16634 & w22099 ) | ( ~w16634 & w22100 ) | ( w22099 & w22100 ) ;
  assign w22102 = ~\pi31 & w22101 ;
  assign w22103 = ( w22098 & ~w22100 ) | ( w22098 & w22102 ) | ( ~w22100 & w22102 ) ;
  assign w22104 = ( w37 & ~w16742 ) | ( w37 & w22103 ) | ( ~w16742 & w22103 ) ;
  assign w22105 = w22103 | w22104 ;
  assign w22106 = w11083 ^ w20404 ;
  assign w22107 = ( \pi14 & w11083 ) | ( \pi14 & ~w22106 ) | ( w11083 & ~w22106 ) ;
  assign w22108 = ( w165 & ~w390 ) | ( w165 & w2656 ) | ( ~w390 & w2656 ) ;
  assign w22109 = w1955 | w11540 ;
  assign w22110 = ( w390 & w723 ) | ( w390 & ~w1955 ) | ( w723 & ~w1955 ) ;
  assign w22111 = w22109 | w22110 ;
  assign w22112 = w22108 | w22111 ;
  assign w22113 = w11308 | w22112 ;
  assign w22114 = ( ~w1324 & w6362 ) | ( ~w1324 & w11308 ) | ( w6362 & w11308 ) ;
  assign w22115 = ~w22113 & w22114 ;
  assign w22116 = w996 | w2306 ;
  assign w22117 = ( w996 & ~w1165 ) | ( w996 & w22115 ) | ( ~w1165 & w22115 ) ;
  assign w22118 = ~w22116 & w22117 ;
  assign w22119 = w310 | w447 ;
  assign w22120 = ( w310 & ~w344 ) | ( w310 & w22118 ) | ( ~w344 & w22118 ) ;
  assign w22121 = ~w22119 & w22120 ;
  assign w22122 = w21915 ^ w22107 ;
  assign w22123 = w22121 ^ w22122 ;
  assign w22124 = w22018 ^ w22123 ;
  assign w22125 = w22105 ^ w22124 ;
  assign w22126 = w3717 | w16630 ;
  assign w22127 = w3649 & w16632 ;
  assign w22128 = ( ~w16630 & w22126 ) | ( ~w16630 & w22127 ) | ( w22126 & w22127 ) ;
  assign w22129 = w3549 | w16628 ;
  assign w22130 = w18026 | w22128 ;
  assign w22131 = ( w3448 & w22128 ) | ( w3448 & w22130 ) | ( w22128 & w22130 ) ;
  assign w22132 = ( ~w16628 & w22129 ) | ( ~w16628 & w22131 ) | ( w22129 & w22131 ) ;
  assign w22133 = \pi29 ^ w22132 ;
  assign w22134 = ( w22020 & ~w22021 ) | ( w22020 & w22022 ) | ( ~w22021 & w22022 ) ;
  assign w22135 = w22125 ^ w22134 ;
  assign w22136 = w22133 ^ w22135 ;
  assign w22137 = ~w4143 & w16619 ;
  assign w22138 = w4052 & ~w16626 ;
  assign w22139 = ( w16619 & ~w22137 ) | ( w16619 & w22138 ) | ( ~w22137 & w22138 ) ;
  assign w22140 = w4147 | w18439 ;
  assign w22141 = w16621 | w22139 ;
  assign w22142 = ( w3964 & w22139 ) | ( w3964 & w22141 ) | ( w22139 & w22141 ) ;
  assign w22143 = ( ~w18439 & w22140 ) | ( ~w18439 & w22142 ) | ( w22140 & w22142 ) ;
  assign w22144 = \pi26 ^ w22143 ;
  assign w22145 = ( ~w22024 & w22032 ) | ( ~w22024 & w22040 ) | ( w22032 & w22040 ) ;
  assign w22146 = w22136 ^ w22145 ;
  assign w22147 = w22144 ^ w22146 ;
  assign w22148 = ( ~w22042 & w22043 ) | ( ~w22042 & w22051 ) | ( w22043 & w22051 ) ;
  assign w22149 = w4651 | w18914 ;
  assign w22150 = w4606 & w16617 ;
  assign w22151 = ( ~w18914 & w22149 ) | ( ~w18914 & w22150 ) | ( w22149 & w22150 ) ;
  assign w22152 = ~w4706 & w18916 ;
  assign w22153 = w19366 & ~w22151 ;
  assign w22154 = ( w4609 & w22151 ) | ( w4609 & ~w22153 ) | ( w22151 & ~w22153 ) ;
  assign w22155 = ( w18916 & ~w22152 ) | ( w18916 & w22154 ) | ( ~w22152 & w22154 ) ;
  assign w22156 = \pi23 ^ w22155 ;
  assign w22157 = w22147 ^ w22148 ;
  assign w22158 = w22156 ^ w22157 ;
  assign w22159 = ~w5343 & w19529 ;
  assign w22160 = w4905 & ~w18912 ;
  assign w22161 = ( w19529 & ~w22159 ) | ( w19529 & w22160 ) | ( ~w22159 & w22160 ) ;
  assign w22162 = ~w5395 & w19713 ;
  assign w22163 = w19723 | w22161 ;
  assign w22164 = ( w4908 & w22161 ) | ( w4908 & w22163 ) | ( w22161 & w22163 ) ;
  assign w22165 = ( w19713 & ~w22162 ) | ( w19713 & w22164 ) | ( ~w22162 & w22164 ) ;
  assign w22166 = \pi20 ^ w22165 ;
  assign w22167 = ( ~w22053 & w22054 ) | ( ~w22053 & w22062 ) | ( w22054 & w22062 ) ;
  assign w22168 = w22158 ^ w22167 ;
  assign w22169 = w22166 ^ w22168 ;
  assign w22170 = ( ~w22064 & w22065 ) | ( ~w22064 & w22073 ) | ( w22065 & w22073 ) ;
  assign w22171 = w5710 | w20068 ;
  assign w22172 = w5494 & w19887 ;
  assign w22173 = ( ~w20068 & w22171 ) | ( ~w20068 & w22172 ) | ( w22171 & w22172 ) ;
  assign w22174 = ~w5948 & w20247 ;
  assign w22175 = w20257 & ~w22173 ;
  assign w22176 = ( w5497 & w22173 ) | ( w5497 & ~w22175 ) | ( w22173 & ~w22175 ) ;
  assign w22177 = ( w20247 & ~w22174 ) | ( w20247 & w22176 ) | ( ~w22174 & w22176 ) ;
  assign w22178 = \pi17 ^ w22177 ;
  assign w22179 = w22169 ^ w22170 ;
  assign w22180 = w22178 ^ w22179 ;
  assign w22181 = w22092 ^ w22096 ;
  assign w22182 = w22180 ^ w22181 ;
  assign w22183 = w22090 & ~w22182 ;
  assign w22184 = w22090 ^ w22182 ;
  assign w22185 = ( ~w22125 & w22133 ) | ( ~w22125 & w22134 ) | ( w22133 & w22134 ) ;
  assign w22186 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16634 ) | ( \pi31 & ~w16634 ) ;
  assign w22187 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22186 ) | ( ~\pi30 & w22186 ) ;
  assign w22188 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22186 ) | ( \pi30 & w22186 ) ;
  assign w22189 = ( ~\pi29 & w16636 ) | ( ~\pi29 & w22188 ) | ( w16636 & w22188 ) ;
  assign w22190 = ( w16632 & w22188 ) | ( w16632 & ~w22189 ) | ( w22188 & ~w22189 ) ;
  assign w22191 = ~\pi31 & w22190 ;
  assign w22192 = ( w22187 & w22189 ) | ( w22187 & w22191 ) | ( w22189 & w22191 ) ;
  assign w22193 = ( w37 & ~w18051 ) | ( w37 & w22192 ) | ( ~w18051 & w22192 ) ;
  assign w22194 = w22192 | w22193 ;
  assign w22195 = ( ~w21915 & w22107 ) | ( ~w21915 & w22121 ) | ( w22107 & w22121 ) ;
  assign w22196 = ( w165 & ~w254 ) | ( w165 & w2470 ) | ( ~w254 & w2470 ) ;
  assign w22197 = w3474 | w11589 ;
  assign w22198 = ( w254 & w339 ) | ( w254 & ~w3474 ) | ( w339 & ~w3474 ) ;
  assign w22199 = w22197 | w22198 ;
  assign w22200 = w22196 | w22199 ;
  assign w22201 = ( ~w488 & w997 ) | ( ~w488 & w5590 ) | ( w997 & w5590 ) ;
  assign w22202 = w4983 | w22200 ;
  assign w22203 = ( w488 & w490 ) | ( w488 & ~w22200 ) | ( w490 & ~w22200 ) ;
  assign w22204 = w22202 | w22203 ;
  assign w22205 = w22201 | w22204 ;
  assign w22206 = ( w468 & w1208 ) | ( w468 & ~w1836 ) | ( w1208 & ~w1836 ) ;
  assign w22207 = w2829 & ~w22205 ;
  assign w22208 = ( w1836 & w2452 ) | ( w1836 & w2829 ) | ( w2452 & w2829 ) ;
  assign w22209 = w22207 & ~w22208 ;
  assign w22210 = ~w22206 & w22209 ;
  assign w22211 = w201 | w345 ;
  assign w22212 = w115 | w22211 ;
  assign w22213 = ( w115 & ~w131 ) | ( w115 & w22210 ) | ( ~w131 & w22210 ) ;
  assign w22214 = ~w22212 & w22213 ;
  assign w22215 = w22194 ^ w22195 ;
  assign w22216 = w22214 ^ w22215 ;
  assign w22217 = ( ~w22018 & w22105 ) | ( ~w22018 & w22123 ) | ( w22105 & w22123 ) ;
  assign w22218 = w3549 & ~w16626 ;
  assign w22219 = ( w3717 & ~w16628 ) | ( w3717 & w22218 ) | ( ~w16628 & w22218 ) ;
  assign w22220 = w3649 | w22219 ;
  assign w22221 = ( ~w16630 & w22219 ) | ( ~w16630 & w22220 ) | ( w22219 & w22220 ) ;
  assign w22222 = w22218 | w22221 ;
  assign w22223 = w3448 | w18429 ;
  assign w22224 = ( ~w18429 & w22222 ) | ( ~w18429 & w22223 ) | ( w22222 & w22223 ) ;
  assign w22225 = \pi29 ^ w22224 ;
  assign w22226 = w22216 ^ w22217 ;
  assign w22227 = w22225 ^ w22226 ;
  assign w22228 = ~w4143 & w16621 ;
  assign w22229 = w4052 & w16619 ;
  assign w22230 = ( w16621 & ~w22228 ) | ( w16621 & w22229 ) | ( ~w22228 & w22229 ) ;
  assign w22231 = ~w4147 & w16732 ;
  assign w22232 = w16617 | w22230 ;
  assign w22233 = ( w3964 & w22230 ) | ( w3964 & w22232 ) | ( w22230 & w22232 ) ;
  assign w22234 = ( w16732 & ~w22231 ) | ( w16732 & w22233 ) | ( ~w22231 & w22233 ) ;
  assign w22235 = \pi26 ^ w22234 ;
  assign w22236 = w22185 ^ w22227 ;
  assign w22237 = w22235 ^ w22236 ;
  assign w22238 = ( ~w22136 & w22144 ) | ( ~w22136 & w22145 ) | ( w22144 & w22145 ) ;
  assign w22239 = ~w4651 & w18916 ;
  assign w22240 = w4606 & ~w18914 ;
  assign w22241 = ( w18916 & ~w22239 ) | ( w18916 & w22240 ) | ( ~w22239 & w22240 ) ;
  assign w22242 = w4706 | w18912 ;
  assign w22243 = w18929 & ~w22241 ;
  assign w22244 = ( w4609 & w22241 ) | ( w4609 & ~w22243 ) | ( w22241 & ~w22243 ) ;
  assign w22245 = ( ~w18912 & w22242 ) | ( ~w18912 & w22244 ) | ( w22242 & w22244 ) ;
  assign w22246 = \pi23 ^ w22245 ;
  assign w22247 = w22237 ^ w22238 ;
  assign w22248 = w22246 ^ w22247 ;
  assign w22249 = ( ~w22147 & w22148 ) | ( ~w22147 & w22156 ) | ( w22148 & w22156 ) ;
  assign w22250 = ~w5343 & w19713 ;
  assign w22251 = w4905 & w19529 ;
  assign w22252 = ( w19713 & ~w22250 ) | ( w19713 & w22251 ) | ( ~w22250 & w22251 ) ;
  assign w22253 = ~w5395 & w19887 ;
  assign w22254 = w19898 | w22252 ;
  assign w22255 = ( w4908 & w22252 ) | ( w4908 & w22254 ) | ( w22252 & w22254 ) ;
  assign w22256 = ( w19887 & ~w22253 ) | ( w19887 & w22255 ) | ( ~w22253 & w22255 ) ;
  assign w22257 = \pi20 ^ w22256 ;
  assign w22258 = w22248 ^ w22249 ;
  assign w22259 = w22257 ^ w22258 ;
  assign w22260 = ( ~w22158 & w22166 ) | ( ~w22158 & w22167 ) | ( w22166 & w22167 ) ;
  assign w22261 = ~w5710 & w20247 ;
  assign w22262 = w5494 & ~w20068 ;
  assign w22263 = ( w20247 & ~w22261 ) | ( w20247 & w22262 ) | ( ~w22261 & w22262 ) ;
  assign w22264 = ~w5948 & w20404 ;
  assign w22265 = w20417 | w22263 ;
  assign w22266 = ( w5497 & w22263 ) | ( w5497 & w22265 ) | ( w22263 & w22265 ) ;
  assign w22267 = ( w20404 & ~w22264 ) | ( w20404 & w22266 ) | ( ~w22264 & w22266 ) ;
  assign w22268 = \pi17 ^ w22267 ;
  assign w22269 = w22259 ^ w22260 ;
  assign w22270 = w22268 ^ w22269 ;
  assign w22271 = ( ~w22169 & w22170 ) | ( ~w22169 & w22178 ) | ( w22170 & w22178 ) ;
  assign w22272 = ( w22092 & w22096 ) | ( w22092 & ~w22180 ) | ( w22096 & ~w22180 ) ;
  assign w22273 = w22270 ^ w22272 ;
  assign w22274 = w22271 ^ w22273 ;
  assign w22275 = w22183 ^ w22274 ;
  assign w22276 = ( ~w22216 & w22217 ) | ( ~w22216 & w22225 ) | ( w22217 & w22225 ) ;
  assign w22277 = ( w22194 & ~w22195 ) | ( w22194 & w22214 ) | ( ~w22195 & w22214 ) ;
  assign w22278 = ( w103 & w220 ) | ( w103 & ~w361 ) | ( w220 & ~w361 ) ;
  assign w22279 = w1282 | w2096 ;
  assign w22280 = ( w361 & w362 ) | ( w361 & ~w2096 ) | ( w362 & ~w2096 ) ;
  assign w22281 = w22279 | w22280 ;
  assign w22282 = w22278 | w22281 ;
  assign w22283 = ( ~w758 & w10603 ) | ( ~w758 & w22282 ) | ( w10603 & w22282 ) ;
  assign w22284 = w1125 | w5137 ;
  assign w22285 = ( w758 & w821 ) | ( w758 & ~w5137 ) | ( w821 & ~w5137 ) ;
  assign w22286 = w22284 | w22285 ;
  assign w22287 = w22283 | w22286 ;
  assign w22288 = ( w1413 & ~w1835 ) | ( w1413 & w3832 ) | ( ~w1835 & w3832 ) ;
  assign w22289 = w2624 | w22287 ;
  assign w22290 = ( w1340 & w1835 ) | ( w1340 & ~w2624 ) | ( w1835 & ~w2624 ) ;
  assign w22291 = w22289 | w22290 ;
  assign w22292 = w22288 | w22291 ;
  assign w22293 = ( w219 & w274 ) | ( w219 & ~w488 ) | ( w274 & ~w488 ) ;
  assign w22294 = w202 | w22292 ;
  assign w22295 = ( ~w202 & w488 ) | ( ~w202 & w524 ) | ( w488 & w524 ) ;
  assign w22296 = w22294 | w22295 ;
  assign w22297 = w22293 | w22296 ;
  assign w22298 = ( w22214 & ~w22277 ) | ( w22214 & w22297 ) | ( ~w22277 & w22297 ) ;
  assign w22299 = w22277 ^ w22297 ;
  assign w22300 = w22214 ^ w22299 ;
  assign w22301 = ( \pi29 & \pi31 ) | ( \pi29 & w16632 ) | ( \pi31 & w16632 ) ;
  assign w22302 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22301 ) | ( ~\pi30 & w22301 ) ;
  assign w22303 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22301 ) | ( \pi30 & w22301 ) ;
  assign w22304 = ( \pi29 & w16634 ) | ( \pi29 & ~w22303 ) | ( w16634 & ~w22303 ) ;
  assign w22305 = ( ~w16630 & w22303 ) | ( ~w16630 & w22304 ) | ( w22303 & w22304 ) ;
  assign w22306 = ~\pi31 & w22305 ;
  assign w22307 = ( w22302 & ~w22304 ) | ( w22302 & w22306 ) | ( ~w22304 & w22306 ) ;
  assign w22308 = ( w37 & ~w18038 ) | ( w37 & w22307 ) | ( ~w18038 & w22307 ) ;
  assign w22309 = w22307 | w22308 ;
  assign w22310 = w3549 & w16619 ;
  assign w22311 = ( w3717 & ~w16626 ) | ( w3717 & w22310 ) | ( ~w16626 & w22310 ) ;
  assign w22312 = w3649 | w22311 ;
  assign w22313 = ( ~w16628 & w22311 ) | ( ~w16628 & w22312 ) | ( w22311 & w22312 ) ;
  assign w22314 = w22310 | w22313 ;
  assign w22315 = ~w3448 & w18451 ;
  assign w22316 = ( w18451 & w22314 ) | ( w18451 & ~w22315 ) | ( w22314 & ~w22315 ) ;
  assign w22317 = \pi29 ^ w22316 ;
  assign w22318 = w22300 ^ w22317 ;
  assign w22319 = w22309 ^ w22318 ;
  assign w22320 = ~w4143 & w16617 ;
  assign w22321 = w4052 & w16621 ;
  assign w22322 = ( w16617 & ~w22320 ) | ( w16617 & w22321 ) | ( ~w22320 & w22321 ) ;
  assign w22323 = w4147 | w19350 ;
  assign w22324 = w18914 & ~w22322 ;
  assign w22325 = ( w3964 & w22322 ) | ( w3964 & ~w22324 ) | ( w22322 & ~w22324 ) ;
  assign w22326 = ( ~w19350 & w22323 ) | ( ~w19350 & w22325 ) | ( w22323 & w22325 ) ;
  assign w22327 = \pi26 ^ w22326 ;
  assign w22328 = w22276 ^ w22319 ;
  assign w22329 = w22327 ^ w22328 ;
  assign w22330 = ( w22185 & ~w22227 ) | ( w22185 & w22235 ) | ( ~w22227 & w22235 ) ;
  assign w22331 = w4651 | w18912 ;
  assign w22332 = w4606 & w18916 ;
  assign w22333 = ( ~w18912 & w22331 ) | ( ~w18912 & w22332 ) | ( w22331 & w22332 ) ;
  assign w22334 = ~w4706 & w19529 ;
  assign w22335 = w19540 & ~w22333 ;
  assign w22336 = ( w4609 & w22333 ) | ( w4609 & ~w22335 ) | ( w22333 & ~w22335 ) ;
  assign w22337 = ( w19529 & ~w22334 ) | ( w19529 & w22336 ) | ( ~w22334 & w22336 ) ;
  assign w22338 = \pi23 ^ w22337 ;
  assign w22339 = w22329 ^ w22330 ;
  assign w22340 = w22338 ^ w22339 ;
  assign w22341 = ( ~w22237 & w22238 ) | ( ~w22237 & w22246 ) | ( w22238 & w22246 ) ;
  assign w22342 = ~w5343 & w19887 ;
  assign w22343 = w4905 & w19713 ;
  assign w22344 = ( w19887 & ~w22342 ) | ( w19887 & w22343 ) | ( ~w22342 & w22343 ) ;
  assign w22345 = w5395 | w20068 ;
  assign w22346 = w20081 & ~w22344 ;
  assign w22347 = ( w4908 & w22344 ) | ( w4908 & ~w22346 ) | ( w22344 & ~w22346 ) ;
  assign w22348 = ( ~w20068 & w22345 ) | ( ~w20068 & w22347 ) | ( w22345 & w22347 ) ;
  assign w22349 = \pi20 ^ w22348 ;
  assign w22350 = w22340 ^ w22341 ;
  assign w22351 = w22349 ^ w22350 ;
  assign w22352 = ( ~w22248 & w22249 ) | ( ~w22248 & w22257 ) | ( w22249 & w22257 ) ;
  assign w22353 = w5948 & w20404 ;
  assign w22354 = ( w5710 & w20404 ) | ( w5710 & w22353 ) | ( w20404 & w22353 ) ;
  assign w22355 = w5494 & w20247 ;
  assign w22356 = w22354 | w22355 ;
  assign w22357 = w5497 & ~w20414 ;
  assign w22358 = ( w5497 & w22356 ) | ( w5497 & ~w22357 ) | ( w22356 & ~w22357 ) ;
  assign w22359 = w22351 ^ w22358 ;
  assign w22360 = \pi17 ^ w22352 ;
  assign w22361 = w22359 ^ w22360 ;
  assign w22362 = ( ~w22259 & w22260 ) | ( ~w22259 & w22268 ) | ( w22260 & w22268 ) ;
  assign w22363 = ( ~w22270 & w22271 ) | ( ~w22270 & w22272 ) | ( w22271 & w22272 ) ;
  assign w22364 = w22362 ^ w22363 ;
  assign w22365 = w22361 ^ w22364 ;
  assign w22366 = w22183 & ~w22274 ;
  assign w22367 = w22365 & w22366 ;
  assign w22368 = w22365 ^ w22366 ;
  assign w22369 = ( w22361 & w22362 ) | ( w22361 & w22363 ) | ( w22362 & w22363 ) ;
  assign w22370 = w20414 | w22356 ;
  assign w22371 = ( w5497 & w22356 ) | ( w5497 & w22370 ) | ( w22356 & w22370 ) ;
  assign w22372 = \pi17 ^ w22371 ;
  assign w22373 = ( w22351 & w22352 ) | ( w22351 & w22372 ) | ( w22352 & w22372 ) ;
  assign w22374 = ( w22329 & w22330 ) | ( w22329 & w22338 ) | ( w22330 & w22338 ) ;
  assign w22375 = ( w22276 & w22319 ) | ( w22276 & w22327 ) | ( w22319 & w22327 ) ;
  assign w22376 = w4143 | w18914 ;
  assign w22377 = w4052 & w16617 ;
  assign w22378 = ( ~w18914 & w22376 ) | ( ~w18914 & w22377 ) | ( w22376 & w22377 ) ;
  assign w22379 = w4147 | w19366 ;
  assign w22380 = w18916 | w22378 ;
  assign w22381 = ( w3964 & w22378 ) | ( w3964 & w22380 ) | ( w22378 & w22380 ) ;
  assign w22382 = ( ~w19366 & w22379 ) | ( ~w19366 & w22381 ) | ( w22379 & w22381 ) ;
  assign w22383 = \pi26 ^ w22382 ;
  assign w22384 = ( w22300 & w22309 ) | ( w22300 & w22317 ) | ( w22309 & w22317 ) ;
  assign w22385 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16630 ) | ( \pi31 & ~w16630 ) ;
  assign w22386 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22385 ) | ( ~\pi30 & w22385 ) ;
  assign w22387 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22385 ) | ( \pi30 & w22385 ) ;
  assign w22388 = ( ~\pi29 & w16632 ) | ( ~\pi29 & w22387 ) | ( w16632 & w22387 ) ;
  assign w22389 = ( w16628 & ~w22387 ) | ( w16628 & w22388 ) | ( ~w22387 & w22388 ) ;
  assign w22390 = \pi31 | w22389 ;
  assign w22391 = ( w22386 & w22388 ) | ( w22386 & ~w22390 ) | ( w22388 & ~w22390 ) ;
  assign w22392 = ( w37 & w18026 ) | ( w37 & w22391 ) | ( w18026 & w22391 ) ;
  assign w22393 = w22391 | w22392 ;
  assign w22394 = w10960 ^ w20404 ;
  assign w22395 = ( \pi17 & w10960 ) | ( \pi17 & ~w22394 ) | ( w10960 & ~w22394 ) ;
  assign w22396 = ( w133 & w257 ) | ( w133 & ~w511 ) | ( w257 & ~w511 ) ;
  assign w22397 = w82 | w1166 ;
  assign w22398 = ( w511 & w513 ) | ( w511 & ~w1166 ) | ( w513 & ~w1166 ) ;
  assign w22399 = w22397 | w22398 ;
  assign w22400 = w22396 | w22399 ;
  assign w22401 = ( w226 & ~w1836 ) | ( w226 & w22400 ) | ( ~w1836 & w22400 ) ;
  assign w22402 = w2856 | w22401 ;
  assign w22403 = ( w442 & w896 ) | ( w442 & ~w22402 ) | ( w896 & ~w22402 ) ;
  assign w22404 = w3371 | w4783 ;
  assign w22405 = ( ~w4783 & w10249 ) | ( ~w4783 & w22402 ) | ( w10249 & w22402 ) ;
  assign w22406 = w22404 | w22405 ;
  assign w22407 = w22403 | w22406 ;
  assign w22408 = ( w259 & w260 ) | ( w259 & ~w281 ) | ( w260 & ~w281 ) ;
  assign w22409 = w206 | w22407 ;
  assign w22410 = ( ~w206 & w281 ) | ( ~w206 & w318 ) | ( w281 & w318 ) ;
  assign w22411 = w22409 | w22410 ;
  assign w22412 = w22408 | w22411 ;
  assign w22413 = ( ~w524 & w783 ) | ( ~w524 & w22412 ) | ( w783 & w22412 ) ;
  assign w22414 = w524 | w22413 ;
  assign w22415 = w22297 ^ w22395 ;
  assign w22416 = w22414 ^ w22415 ;
  assign w22417 = w22298 ^ w22416 ;
  assign w22418 = w22393 ^ w22417 ;
  assign w22419 = ~w3717 & w16619 ;
  assign w22420 = w3649 & ~w16626 ;
  assign w22421 = ( w16619 & ~w22419 ) | ( w16619 & w22420 ) | ( ~w22419 & w22420 ) ;
  assign w22422 = ~w3549 & w16621 ;
  assign w22423 = w18439 & ~w22421 ;
  assign w22424 = ( w3448 & w22421 ) | ( w3448 & ~w22423 ) | ( w22421 & ~w22423 ) ;
  assign w22425 = ( w16621 & ~w22422 ) | ( w16621 & w22424 ) | ( ~w22422 & w22424 ) ;
  assign w22426 = \pi29 ^ w22425 ;
  assign w22427 = w22384 ^ w22418 ;
  assign w22428 = w22426 ^ w22427 ;
  assign w22429 = w22375 ^ w22428 ;
  assign w22430 = w22383 ^ w22429 ;
  assign w22431 = ~w4651 & w19529 ;
  assign w22432 = w4606 & ~w18912 ;
  assign w22433 = ( w19529 & ~w22431 ) | ( w19529 & w22432 ) | ( ~w22431 & w22432 ) ;
  assign w22434 = ~w4706 & w19713 ;
  assign w22435 = w19723 | w22433 ;
  assign w22436 = ( w4609 & w22433 ) | ( w4609 & w22435 ) | ( w22433 & w22435 ) ;
  assign w22437 = ( w19713 & ~w22434 ) | ( w19713 & w22436 ) | ( ~w22434 & w22436 ) ;
  assign w22438 = \pi23 ^ w22437 ;
  assign w22439 = w22374 ^ w22430 ;
  assign w22440 = w22438 ^ w22439 ;
  assign w22441 = ( w22340 & w22341 ) | ( w22340 & w22349 ) | ( w22341 & w22349 ) ;
  assign w22442 = w5343 | w20068 ;
  assign w22443 = w4905 & w19887 ;
  assign w22444 = ( ~w20068 & w22442 ) | ( ~w20068 & w22443 ) | ( w22442 & w22443 ) ;
  assign w22445 = ~w5395 & w20247 ;
  assign w22446 = w20257 & ~w22444 ;
  assign w22447 = ( w4908 & w22444 ) | ( w4908 & ~w22446 ) | ( w22444 & ~w22446 ) ;
  assign w22448 = ( w20247 & ~w22445 ) | ( w20247 & w22447 ) | ( ~w22445 & w22447 ) ;
  assign w22449 = \pi20 ^ w22448 ;
  assign w22450 = w22440 ^ w22441 ;
  assign w22451 = w22449 ^ w22450 ;
  assign w22452 = w22369 ^ w22373 ;
  assign w22453 = w22451 ^ w22452 ;
  assign w22454 = w22367 & w22453 ;
  assign w22455 = w22367 ^ w22453 ;
  assign w22456 = ( w22384 & w22418 ) | ( w22384 & w22426 ) | ( w22418 & w22426 ) ;
  assign w22457 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16628 ) | ( \pi31 & ~w16628 ) ;
  assign w22458 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22457 ) | ( ~\pi30 & w22457 ) ;
  assign w22459 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22457 ) | ( \pi30 & w22457 ) ;
  assign w22460 = ( \pi29 & w16630 ) | ( \pi29 & ~w22459 ) | ( w16630 & ~w22459 ) ;
  assign w22461 = ( ~w16626 & w22459 ) | ( ~w16626 & w22460 ) | ( w22459 & w22460 ) ;
  assign w22462 = ~\pi31 & w22461 ;
  assign w22463 = ( w22458 & ~w22460 ) | ( w22458 & w22462 ) | ( ~w22460 & w22462 ) ;
  assign w22464 = ( w37 & ~w18429 ) | ( w37 & w22463 ) | ( ~w18429 & w22463 ) ;
  assign w22465 = w22463 | w22464 ;
  assign w22466 = ( w22297 & ~w22395 ) | ( w22297 & w22414 ) | ( ~w22395 & w22414 ) ;
  assign w22467 = w340 | w860 ;
  assign w22468 = w220 | w22467 ;
  assign w22469 = ( w68 & ~w220 ) | ( w68 & w310 ) | ( ~w220 & w310 ) ;
  assign w22470 = w22468 | w22469 ;
  assign w22471 = w492 | w606 ;
  assign w22472 = w144 | w22471 ;
  assign w22473 = ( ~w144 & w413 ) | ( ~w144 & w22470 ) | ( w413 & w22470 ) ;
  assign w22474 = w22472 | w22473 ;
  assign w22475 = ( w2663 & w3599 ) | ( w2663 & ~w22474 ) | ( w3599 & ~w22474 ) ;
  assign w22476 = ~w6135 & w21307 ;
  assign w22477 = ( w416 & w21307 ) | ( w416 & w22474 ) | ( w21307 & w22474 ) ;
  assign w22478 = w22476 & ~w22477 ;
  assign w22479 = ~w22475 & w22478 ;
  assign w22480 = w313 | w314 ;
  assign w22481 = w410 | w22480 ;
  assign w22482 = ( w410 & ~w4174 ) | ( w410 & w22479 ) | ( ~w4174 & w22479 ) ;
  assign w22483 = ~w22481 & w22482 ;
  assign w22484 = w533 | w625 ;
  assign w22485 = w178 | w22484 ;
  assign w22486 = ( w178 & ~w262 ) | ( w178 & w22483 ) | ( ~w262 & w22483 ) ;
  assign w22487 = ~w22485 & w22486 ;
  assign w22488 = w22465 ^ w22466 ;
  assign w22489 = w22487 ^ w22488 ;
  assign w22490 = ( w22298 & ~w22393 ) | ( w22298 & w22416 ) | ( ~w22393 & w22416 ) ;
  assign w22491 = ~w3717 & w16621 ;
  assign w22492 = w3649 & w16619 ;
  assign w22493 = ( w16621 & ~w22491 ) | ( w16621 & w22492 ) | ( ~w22491 & w22492 ) ;
  assign w22494 = ~w3549 & w16617 ;
  assign w22495 = w16732 | w22493 ;
  assign w22496 = ( w3448 & w22493 ) | ( w3448 & w22495 ) | ( w22493 & w22495 ) ;
  assign w22497 = ( w16617 & ~w22494 ) | ( w16617 & w22496 ) | ( ~w22494 & w22496 ) ;
  assign w22498 = \pi29 ^ w22497 ;
  assign w22499 = w22489 ^ w22490 ;
  assign w22500 = w22498 ^ w22499 ;
  assign w22501 = ~w4143 & w18916 ;
  assign w22502 = w4052 & ~w18914 ;
  assign w22503 = ( w18916 & ~w22501 ) | ( w18916 & w22502 ) | ( ~w22501 & w22502 ) ;
  assign w22504 = w4147 | w18929 ;
  assign w22505 = w18912 & ~w22503 ;
  assign w22506 = ( w3964 & w22503 ) | ( w3964 & ~w22505 ) | ( w22503 & ~w22505 ) ;
  assign w22507 = ( ~w18929 & w22504 ) | ( ~w18929 & w22506 ) | ( w22504 & w22506 ) ;
  assign w22508 = \pi26 ^ w22507 ;
  assign w22509 = w22456 ^ w22500 ;
  assign w22510 = w22508 ^ w22509 ;
  assign w22511 = ( w22375 & w22383 ) | ( w22375 & w22428 ) | ( w22383 & w22428 ) ;
  assign w22512 = ~w4651 & w19713 ;
  assign w22513 = w4606 & w19529 ;
  assign w22514 = ( w19713 & ~w22512 ) | ( w19713 & w22513 ) | ( ~w22512 & w22513 ) ;
  assign w22515 = ~w4706 & w19887 ;
  assign w22516 = w19898 | w22514 ;
  assign w22517 = ( w4609 & w22514 ) | ( w4609 & w22516 ) | ( w22514 & w22516 ) ;
  assign w22518 = ( w19887 & ~w22515 ) | ( w19887 & w22517 ) | ( ~w22515 & w22517 ) ;
  assign w22519 = \pi23 ^ w22518 ;
  assign w22520 = w22510 ^ w22511 ;
  assign w22521 = w22519 ^ w22520 ;
  assign w22522 = ( w22374 & w22430 ) | ( w22374 & w22438 ) | ( w22430 & w22438 ) ;
  assign w22523 = ~w5343 & w20247 ;
  assign w22524 = w4905 & ~w20068 ;
  assign w22525 = ( w20247 & ~w22523 ) | ( w20247 & w22524 ) | ( ~w22523 & w22524 ) ;
  assign w22526 = ~w5395 & w20404 ;
  assign w22527 = w20417 | w22525 ;
  assign w22528 = ( w4908 & w22525 ) | ( w4908 & w22527 ) | ( w22525 & w22527 ) ;
  assign w22529 = ( w20404 & ~w22526 ) | ( w20404 & w22528 ) | ( ~w22526 & w22528 ) ;
  assign w22530 = \pi20 ^ w22529 ;
  assign w22531 = w22521 ^ w22522 ;
  assign w22532 = w22530 ^ w22531 ;
  assign w22533 = ( w22440 & w22441 ) | ( w22440 & w22449 ) | ( w22441 & w22449 ) ;
  assign w22534 = ( w22369 & w22373 ) | ( w22369 & w22451 ) | ( w22373 & w22451 ) ;
  assign w22535 = w22532 ^ w22534 ;
  assign w22536 = w22533 ^ w22535 ;
  assign w22537 = w22454 ^ w22536 ;
  assign w22538 = w22454 & ~w22536 ;
  assign w22539 = ( \pi29 & \pi31 ) | ( \pi29 & ~w16626 ) | ( \pi31 & ~w16626 ) ;
  assign w22540 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22539 ) | ( ~\pi30 & w22539 ) ;
  assign w22541 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22539 ) | ( \pi30 & w22539 ) ;
  assign w22542 = ( \pi29 & w16628 ) | ( \pi29 & ~w22541 ) | ( w16628 & ~w22541 ) ;
  assign w22543 = ( w16619 & w22541 ) | ( w16619 & w22542 ) | ( w22541 & w22542 ) ;
  assign w22544 = ~\pi31 & w22543 ;
  assign w22545 = ( w22540 & ~w22542 ) | ( w22540 & w22544 ) | ( ~w22542 & w22544 ) ;
  assign w22546 = ( w37 & w18451 ) | ( w37 & w22545 ) | ( w18451 & w22545 ) ;
  assign w22547 = w22545 | w22546 ;
  assign w22548 = ( w143 & w220 ) | ( w143 & ~w342 ) | ( w220 & ~w342 ) ;
  assign w22549 = w103 | w1282 ;
  assign w22550 = ( ~w103 & w342 ) | ( ~w103 & w1031 ) | ( w342 & w1031 ) ;
  assign w22551 = w22549 | w22550 ;
  assign w22552 = w22548 | w22551 ;
  assign w22553 = w2782 | w22552 ;
  assign w22554 = w4463 & ~w22553 ;
  assign w22555 = ( w3347 & w4463 ) | ( w3347 & w6190 ) | ( w4463 & w6190 ) ;
  assign w22556 = w22554 & ~w22555 ;
  assign w22557 = ( w198 & w205 ) | ( w198 & ~w206 ) | ( w205 & ~w206 ) ;
  assign w22558 = ~w487 & w22556 ;
  assign w22559 = ( w206 & w269 ) | ( w206 & ~w487 ) | ( w269 & ~w487 ) ;
  assign w22560 = w22558 & ~w22559 ;
  assign w22561 = ~w22557 & w22560 ;
  assign w22562 = ( w92 & w111 ) | ( w92 & ~w606 ) | ( w111 & ~w606 ) ;
  assign w22563 = ~w20728 & w22561 ;
  assign w22564 = ( w606 & w1126 ) | ( w606 & ~w20728 ) | ( w1126 & ~w20728 ) ;
  assign w22565 = w22563 & ~w22564 ;
  assign w22566 = ~w22562 & w22565 ;
  assign w22567 = ( w22487 & w22547 ) | ( w22487 & ~w22566 ) | ( w22547 & ~w22566 ) ;
  assign w22568 = w22487 ^ w22547 ;
  assign w22569 = w22566 ^ w22568 ;
  assign w22570 = ( w22465 & w22466 ) | ( w22465 & w22487 ) | ( w22466 & w22487 ) ;
  assign w22571 = ( w22489 & ~w22490 ) | ( w22489 & w22498 ) | ( ~w22490 & w22498 ) ;
  assign w22572 = w22570 ^ w22571 ;
  assign w22573 = w22569 ^ w22572 ;
  assign w22574 = ~w3717 & w16617 ;
  assign w22575 = w3649 & w16621 ;
  assign w22576 = ( w16617 & ~w22574 ) | ( w16617 & w22575 ) | ( ~w22574 & w22575 ) ;
  assign w22577 = w3549 | w18914 ;
  assign w22578 = w19350 & ~w22576 ;
  assign w22579 = ( w3448 & w22576 ) | ( w3448 & ~w22578 ) | ( w22576 & ~w22578 ) ;
  assign w22580 = ( ~w18914 & w22577 ) | ( ~w18914 & w22579 ) | ( w22577 & w22579 ) ;
  assign w22581 = \pi29 ^ w22580 ;
  assign w22582 = w4143 | w18912 ;
  assign w22583 = w4052 & w18916 ;
  assign w22584 = ( ~w18912 & w22582 ) | ( ~w18912 & w22583 ) | ( w22582 & w22583 ) ;
  assign w22585 = w4147 | w19540 ;
  assign w22586 = w19529 | w22584 ;
  assign w22587 = ( w3964 & w22584 ) | ( w3964 & w22586 ) | ( w22584 & w22586 ) ;
  assign w22588 = ( ~w19540 & w22585 ) | ( ~w19540 & w22587 ) | ( w22585 & w22587 ) ;
  assign w22589 = \pi26 ^ w22588 ;
  assign w22590 = w22573 ^ w22589 ;
  assign w22591 = w22581 ^ w22590 ;
  assign w22592 = ( w22456 & ~w22500 ) | ( w22456 & w22508 ) | ( ~w22500 & w22508 ) ;
  assign w22593 = ~w4651 & w19887 ;
  assign w22594 = w4606 & w19713 ;
  assign w22595 = ( w19887 & ~w22593 ) | ( w19887 & w22594 ) | ( ~w22593 & w22594 ) ;
  assign w22596 = w4706 | w20068 ;
  assign w22597 = w20081 & ~w22595 ;
  assign w22598 = ( w4609 & w22595 ) | ( w4609 & ~w22597 ) | ( w22595 & ~w22597 ) ;
  assign w22599 = ( ~w20068 & w22596 ) | ( ~w20068 & w22598 ) | ( w22596 & w22598 ) ;
  assign w22600 = \pi23 ^ w22599 ;
  assign w22601 = w22591 ^ w22592 ;
  assign w22602 = w22600 ^ w22601 ;
  assign w22603 = ( ~w22510 & w22511 ) | ( ~w22510 & w22519 ) | ( w22511 & w22519 ) ;
  assign w22604 = w5395 & w20404 ;
  assign w22605 = ( w5343 & w20404 ) | ( w5343 & w22604 ) | ( w20404 & w22604 ) ;
  assign w22606 = w4905 & w20247 ;
  assign w22607 = w22605 | w22606 ;
  assign w22608 = w4908 & ~w20414 ;
  assign w22609 = ( w4908 & w22607 ) | ( w4908 & ~w22608 ) | ( w22607 & ~w22608 ) ;
  assign w22610 = w22602 ^ w22609 ;
  assign w22611 = \pi20 ^ w22603 ;
  assign w22612 = w22610 ^ w22611 ;
  assign w22613 = ( ~w22521 & w22522 ) | ( ~w22521 & w22530 ) | ( w22522 & w22530 ) ;
  assign w22614 = ( ~w22532 & w22533 ) | ( ~w22532 & w22534 ) | ( w22533 & w22534 ) ;
  assign w22615 = w22613 ^ w22614 ;
  assign w22616 = w22612 ^ w22615 ;
  assign w22617 = w22538 & ~w22616 ;
  assign w22618 = w22538 ^ w22616 ;
  assign w22619 = ( ~w22612 & w22613 ) | ( ~w22612 & w22614 ) | ( w22613 & w22614 ) ;
  assign w22620 = w20414 | w22607 ;
  assign w22621 = ( w4908 & w22607 ) | ( w4908 & w22620 ) | ( w22607 & w22620 ) ;
  assign w22622 = \pi20 ^ w22621 ;
  assign w22623 = ( ~w22602 & w22603 ) | ( ~w22602 & w22622 ) | ( w22603 & w22622 ) ;
  assign w22624 = ( \pi29 & \pi31 ) | ( \pi29 & w16619 ) | ( \pi31 & w16619 ) ;
  assign w22625 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22624 ) | ( ~\pi30 & w22624 ) ;
  assign w22626 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22624 ) | ( \pi30 & w22624 ) ;
  assign w22627 = ( \pi29 & w16626 ) | ( \pi29 & ~w22626 ) | ( w16626 & ~w22626 ) ;
  assign w22628 = ( w16621 & w22626 ) | ( w16621 & w22627 ) | ( w22626 & w22627 ) ;
  assign w22629 = ~\pi31 & w22628 ;
  assign w22630 = ( w22625 & ~w22627 ) | ( w22625 & w22629 ) | ( ~w22627 & w22629 ) ;
  assign w22631 = ( w37 & ~w18439 ) | ( w37 & w22630 ) | ( ~w18439 & w22630 ) ;
  assign w22632 = w22630 | w22631 ;
  assign w22633 = w10740 ^ w20404 ;
  assign w22634 = ( \pi20 & w10740 ) | ( \pi20 & ~w22633 ) | ( w10740 & ~w22633 ) ;
  assign w22635 = ( w390 & w466 ) | ( w390 & ~w663 ) | ( w466 & ~w663 ) ;
  assign w22636 = w517 | w528 ;
  assign w22637 = ( ~w528 & w663 ) | ( ~w528 & w1030 ) | ( w663 & w1030 ) ;
  assign w22638 = w22636 | w22637 ;
  assign w22639 = w22635 | w22638 ;
  assign w22640 = ( w11968 & w12706 ) | ( w11968 & w22639 ) | ( w12706 & w22639 ) ;
  assign w22641 = w12706 & ~w22640 ;
  assign w22642 = ( w495 & ~w536 ) | ( w495 & w22641 ) | ( ~w536 & w22641 ) ;
  assign w22643 = w1029 | w4379 ;
  assign w22644 = ( w495 & w513 ) | ( w495 & ~w4379 ) | ( w513 & ~w4379 ) ;
  assign w22645 = w22643 | w22644 ;
  assign w22646 = w22642 & ~w22645 ;
  assign w22647 = ( w120 & ~w311 ) | ( w120 & w1615 ) | ( ~w311 & w1615 ) ;
  assign w22648 = ~w2624 & w22646 ;
  assign w22649 = ( w311 & w561 ) | ( w311 & ~w2624 ) | ( w561 & ~w2624 ) ;
  assign w22650 = w22648 & ~w22649 ;
  assign w22651 = ~w22647 & w22650 ;
  assign w22652 = ( w176 & w413 ) | ( w176 & ~w447 ) | ( w413 & ~w447 ) ;
  assign w22653 = ~w163 & w22651 ;
  assign w22654 = ( ~w163 & w447 ) | ( ~w163 & w726 ) | ( w447 & w726 ) ;
  assign w22655 = w22653 & ~w22654 ;
  assign w22656 = ~w22652 & w22655 ;
  assign w22657 = w22487 ^ w22634 ;
  assign w22658 = w22656 ^ w22657 ;
  assign w22659 = w22567 ^ w22658 ;
  assign w22660 = w22632 ^ w22659 ;
  assign w22661 = ( ~w22569 & w22570 ) | ( ~w22569 & w22571 ) | ( w22570 & w22571 ) ;
  assign w22662 = w3717 | w18914 ;
  assign w22663 = w3649 & w16617 ;
  assign w22664 = ( ~w18914 & w22662 ) | ( ~w18914 & w22663 ) | ( w22662 & w22663 ) ;
  assign w22665 = ~w3549 & w18916 ;
  assign w22666 = w19366 & ~w22664 ;
  assign w22667 = ( w3448 & w22664 ) | ( w3448 & ~w22666 ) | ( w22664 & ~w22666 ) ;
  assign w22668 = ( w18916 & ~w22665 ) | ( w18916 & w22667 ) | ( ~w22665 & w22667 ) ;
  assign w22669 = \pi29 ^ w22668 ;
  assign w22670 = w22660 ^ w22661 ;
  assign w22671 = w22669 ^ w22670 ;
  assign w22672 = ~w4143 & w19529 ;
  assign w22673 = w4052 & ~w18912 ;
  assign w22674 = ( w19529 & ~w22672 ) | ( w19529 & w22673 ) | ( ~w22672 & w22673 ) ;
  assign w22675 = ~w4147 & w19723 ;
  assign w22676 = w19713 | w22674 ;
  assign w22677 = ( w3964 & w22674 ) | ( w3964 & w22676 ) | ( w22674 & w22676 ) ;
  assign w22678 = ( w19723 & ~w22675 ) | ( w19723 & w22677 ) | ( ~w22675 & w22677 ) ;
  assign w22679 = \pi26 ^ w22678 ;
  assign w22680 = ( ~w22573 & w22581 ) | ( ~w22573 & w22589 ) | ( w22581 & w22589 ) ;
  assign w22681 = w22671 ^ w22680 ;
  assign w22682 = w22679 ^ w22681 ;
  assign w22683 = ( ~w22591 & w22592 ) | ( ~w22591 & w22600 ) | ( w22592 & w22600 ) ;
  assign w22684 = w4651 | w20068 ;
  assign w22685 = w4606 & w19887 ;
  assign w22686 = ( ~w20068 & w22684 ) | ( ~w20068 & w22685 ) | ( w22684 & w22685 ) ;
  assign w22687 = ~w4706 & w20247 ;
  assign w22688 = w20257 & ~w22686 ;
  assign w22689 = ( w4609 & w22686 ) | ( w4609 & ~w22688 ) | ( w22686 & ~w22688 ) ;
  assign w22690 = ( w20247 & ~w22687 ) | ( w20247 & w22689 ) | ( ~w22687 & w22689 ) ;
  assign w22691 = \pi23 ^ w22690 ;
  assign w22692 = w22682 ^ w22683 ;
  assign w22693 = w22691 ^ w22692 ;
  assign w22694 = w22619 ^ w22623 ;
  assign w22695 = w22693 ^ w22694 ;
  assign w22696 = w22617 & ~w22695 ;
  assign w22697 = w22617 ^ w22695 ;
  assign w22698 = ( ~w22660 & w22661 ) | ( ~w22660 & w22669 ) | ( w22661 & w22669 ) ;
  assign w22699 = ( \pi29 & \pi31 ) | ( \pi29 & w16621 ) | ( \pi31 & w16621 ) ;
  assign w22700 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22699 ) | ( ~\pi30 & w22699 ) ;
  assign w22701 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22699 ) | ( \pi30 & w22699 ) ;
  assign w22702 = ( ~\pi29 & w16619 ) | ( ~\pi29 & w22701 ) | ( w16619 & w22701 ) ;
  assign w22703 = ( w16617 & w22701 ) | ( w16617 & ~w22702 ) | ( w22701 & ~w22702 ) ;
  assign w22704 = ~\pi31 & w22703 ;
  assign w22705 = ( w22700 & w22702 ) | ( w22700 & w22704 ) | ( w22702 & w22704 ) ;
  assign w22706 = ( w37 & w16732 ) | ( w37 & w22705 ) | ( w16732 & w22705 ) ;
  assign w22707 = w22705 | w22706 ;
  assign w22708 = ( w22487 & w22634 ) | ( w22487 & w22656 ) | ( w22634 & w22656 ) ;
  assign w22709 = ( w496 & w608 ) | ( w496 & ~w899 ) | ( w608 & ~w899 ) ;
  assign w22710 = w86 | w495 ;
  assign w22711 = ( ~w495 & w899 ) | ( ~w495 & w1031 ) | ( w899 & w1031 ) ;
  assign w22712 = w22710 | w22711 ;
  assign w22713 = w22709 | w22712 ;
  assign w22714 = w1051 | w22713 ;
  assign w22715 = ( ~w1051 & w1684 ) | ( ~w1051 & w11601 ) | ( w1684 & w11601 ) ;
  assign w22716 = w22714 | w22715 ;
  assign w22717 = ( w1727 & w3114 ) | ( w1727 & ~w12830 ) | ( w3114 & ~w12830 ) ;
  assign w22718 = w3371 | w22716 ;
  assign w22719 = ( w1281 & w12830 ) | ( w1281 & ~w22716 ) | ( w12830 & ~w22716 ) ;
  assign w22720 = w22718 | w22719 ;
  assign w22721 = w22717 | w22720 ;
  assign w22722 = ( w198 & w280 ) | ( w198 & ~w606 ) | ( w280 & ~w606 ) ;
  assign w22723 = w114 | w22721 ;
  assign w22724 = ( ~w114 & w606 ) | ( ~w114 & w1274 ) | ( w606 & w1274 ) ;
  assign w22725 = w22723 | w22724 ;
  assign w22726 = w22722 | w22725 ;
  assign w22727 = w22707 ^ w22708 ;
  assign w22728 = w22726 ^ w22727 ;
  assign w22729 = ( w22567 & w22632 ) | ( w22567 & ~w22658 ) | ( w22632 & ~w22658 ) ;
  assign w22730 = ~w3717 & w18916 ;
  assign w22731 = w3649 & ~w18914 ;
  assign w22732 = ( w18916 & ~w22730 ) | ( w18916 & w22731 ) | ( ~w22730 & w22731 ) ;
  assign w22733 = w3549 | w18912 ;
  assign w22734 = w18929 & ~w22732 ;
  assign w22735 = ( w3448 & w22732 ) | ( w3448 & ~w22734 ) | ( w22732 & ~w22734 ) ;
  assign w22736 = ( ~w18912 & w22733 ) | ( ~w18912 & w22735 ) | ( w22733 & w22735 ) ;
  assign w22737 = \pi29 ^ w22736 ;
  assign w22738 = w22728 ^ w22729 ;
  assign w22739 = w22737 ^ w22738 ;
  assign w22740 = ~w4143 & w19713 ;
  assign w22741 = w4052 & w19529 ;
  assign w22742 = ( w19713 & ~w22740 ) | ( w19713 & w22741 ) | ( ~w22740 & w22741 ) ;
  assign w22743 = ~w4147 & w19898 ;
  assign w22744 = w19887 | w22742 ;
  assign w22745 = ( w3964 & w22742 ) | ( w3964 & w22744 ) | ( w22742 & w22744 ) ;
  assign w22746 = ( w19898 & ~w22743 ) | ( w19898 & w22745 ) | ( ~w22743 & w22745 ) ;
  assign w22747 = \pi26 ^ w22746 ;
  assign w22748 = w22698 ^ w22739 ;
  assign w22749 = w22747 ^ w22748 ;
  assign w22750 = ( ~w22671 & w22679 ) | ( ~w22671 & w22680 ) | ( w22679 & w22680 ) ;
  assign w22751 = ~w4651 & w20247 ;
  assign w22752 = w4606 & ~w20068 ;
  assign w22753 = ( w20247 & ~w22751 ) | ( w20247 & w22752 ) | ( ~w22751 & w22752 ) ;
  assign w22754 = ~w4706 & w20404 ;
  assign w22755 = w20417 | w22753 ;
  assign w22756 = ( w4609 & w22753 ) | ( w4609 & w22755 ) | ( w22753 & w22755 ) ;
  assign w22757 = ( w20404 & ~w22754 ) | ( w20404 & w22756 ) | ( ~w22754 & w22756 ) ;
  assign w22758 = \pi23 ^ w22757 ;
  assign w22759 = w22749 ^ w22750 ;
  assign w22760 = w22758 ^ w22759 ;
  assign w22761 = ( ~w22682 & w22683 ) | ( ~w22682 & w22691 ) | ( w22683 & w22691 ) ;
  assign w22762 = ( w22619 & w22623 ) | ( w22619 & ~w22693 ) | ( w22623 & ~w22693 ) ;
  assign w22763 = w22760 ^ w22762 ;
  assign w22764 = w22761 ^ w22763 ;
  assign w22765 = w22696 ^ w22764 ;
  assign w22766 = ( ~w22707 & w22708 ) | ( ~w22707 & w22726 ) | ( w22708 & w22726 ) ;
  assign w22767 = w492 | w697 ;
  assign w22768 = w253 | w22767 ;
  assign w22769 = ( w86 & ~w253 ) | ( w86 & w411 ) | ( ~w253 & w411 ) ;
  assign w22770 = w22768 | w22769 ;
  assign w22771 = ( ~w229 & w12620 ) | ( ~w229 & w22770 ) | ( w12620 & w22770 ) ;
  assign w22772 = w4311 | w18776 ;
  assign w22773 = ( w229 & w509 ) | ( w229 & ~w18776 ) | ( w509 & ~w18776 ) ;
  assign w22774 = w22772 | w22773 ;
  assign w22775 = w22771 | w22774 ;
  assign w22776 = ( w267 & w731 ) | ( w267 & ~w1281 ) | ( w731 & ~w1281 ) ;
  assign w22777 = w21292 | w22775 ;
  assign w22778 = ( w1281 & w2782 ) | ( w1281 & ~w21292 ) | ( w2782 & ~w21292 ) ;
  assign w22779 = w22777 | w22778 ;
  assign w22780 = w22776 | w22779 ;
  assign w22781 = ( w210 & w284 ) | ( w210 & ~w317 ) | ( w284 & ~w317 ) ;
  assign w22782 = w16910 & ~w22780 ;
  assign w22783 = ( w317 & w724 ) | ( w317 & w16910 ) | ( w724 & w16910 ) ;
  assign w22784 = w22782 & ~w22783 ;
  assign w22785 = ~w22781 & w22784 ;
  assign w22786 = ( w22726 & ~w22766 ) | ( w22726 & w22785 ) | ( ~w22766 & w22785 ) ;
  assign w22787 = w22766 ^ w22785 ;
  assign w22788 = w22726 ^ w22787 ;
  assign w22789 = ( \pi29 & \pi31 ) | ( \pi29 & w16617 ) | ( \pi31 & w16617 ) ;
  assign w22790 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22789 ) | ( ~\pi30 & w22789 ) ;
  assign w22791 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22789 ) | ( \pi30 & w22789 ) ;
  assign w22792 = ( ~\pi29 & w16621 ) | ( ~\pi29 & w22791 ) | ( w16621 & w22791 ) ;
  assign w22793 = ( w18914 & ~w22791 ) | ( w18914 & w22792 ) | ( ~w22791 & w22792 ) ;
  assign w22794 = \pi31 | w22793 ;
  assign w22795 = ( w22790 & w22792 ) | ( w22790 & ~w22794 ) | ( w22792 & ~w22794 ) ;
  assign w22796 = ( w37 & ~w19350 ) | ( w37 & w22795 ) | ( ~w19350 & w22795 ) ;
  assign w22797 = w22795 | w22796 ;
  assign w22798 = ( w22728 & w22729 ) | ( w22728 & w22737 ) | ( w22729 & w22737 ) ;
  assign w22799 = w22788 ^ w22798 ;
  assign w22800 = w22797 ^ w22799 ;
  assign w22801 = w3717 | w18912 ;
  assign w22802 = w3649 & w18916 ;
  assign w22803 = ( ~w18912 & w22801 ) | ( ~w18912 & w22802 ) | ( w22801 & w22802 ) ;
  assign w22804 = ~w3549 & w19529 ;
  assign w22805 = w19540 & ~w22803 ;
  assign w22806 = ( w3448 & w22803 ) | ( w3448 & ~w22805 ) | ( w22803 & ~w22805 ) ;
  assign w22807 = ( w19529 & ~w22804 ) | ( w19529 & w22806 ) | ( ~w22804 & w22806 ) ;
  assign w22808 = \pi29 ^ w22807 ;
  assign w22809 = ~w4143 & w19887 ;
  assign w22810 = w4052 & w19713 ;
  assign w22811 = ( w19887 & ~w22809 ) | ( w19887 & w22810 ) | ( ~w22809 & w22810 ) ;
  assign w22812 = w4147 | w20081 ;
  assign w22813 = w20068 & ~w22811 ;
  assign w22814 = ( w3964 & w22811 ) | ( w3964 & ~w22813 ) | ( w22811 & ~w22813 ) ;
  assign w22815 = ( ~w20081 & w22812 ) | ( ~w20081 & w22814 ) | ( w22812 & w22814 ) ;
  assign w22816 = \pi26 ^ w22815 ;
  assign w22817 = w22800 ^ w22816 ;
  assign w22818 = w22808 ^ w22817 ;
  assign w22819 = ( w22698 & w22739 ) | ( w22698 & w22747 ) | ( w22739 & w22747 ) ;
  assign w22820 = w4706 & w20404 ;
  assign w22821 = ( w4651 & w20404 ) | ( w4651 & w22820 ) | ( w20404 & w22820 ) ;
  assign w22822 = w4606 & w20247 ;
  assign w22823 = w22821 | w22822 ;
  assign w22824 = w4609 & ~w20414 ;
  assign w22825 = ( w4609 & w22823 ) | ( w4609 & ~w22824 ) | ( w22823 & ~w22824 ) ;
  assign w22826 = w22819 ^ w22825 ;
  assign w22827 = \pi23 ^ w22818 ;
  assign w22828 = w22826 ^ w22827 ;
  assign w22829 = ( w22749 & w22750 ) | ( w22749 & w22758 ) | ( w22750 & w22758 ) ;
  assign w22830 = ( w22760 & w22761 ) | ( w22760 & w22762 ) | ( w22761 & w22762 ) ;
  assign w22831 = w22828 ^ w22830 ;
  assign w22832 = w22829 ^ w22831 ;
  assign w22833 = w22696 & w22764 ;
  assign w22834 = ~w22832 & w22833 ;
  assign w22835 = w22832 ^ w22833 ;
  assign w22836 = ( ~w22828 & w22829 ) | ( ~w22828 & w22830 ) | ( w22829 & w22830 ) ;
  assign w22837 = w20414 | w22823 ;
  assign w22838 = ( w4609 & w22823 ) | ( w4609 & w22837 ) | ( w22823 & w22837 ) ;
  assign w22839 = \pi23 ^ w22838 ;
  assign w22840 = ( ~w22818 & w22819 ) | ( ~w22818 & w22839 ) | ( w22819 & w22839 ) ;
  assign w22841 = ( ~w22800 & w22808 ) | ( ~w22800 & w22816 ) | ( w22808 & w22816 ) ;
  assign w22842 = w4143 | w20068 ;
  assign w22843 = w4052 & w19887 ;
  assign w22844 = ( ~w20068 & w22842 ) | ( ~w20068 & w22843 ) | ( w22842 & w22843 ) ;
  assign w22845 = w4147 | w20257 ;
  assign w22846 = w20247 | w22844 ;
  assign w22847 = ( w3964 & w22844 ) | ( w3964 & w22846 ) | ( w22844 & w22846 ) ;
  assign w22848 = ( ~w20257 & w22845 ) | ( ~w20257 & w22847 ) | ( w22845 & w22847 ) ;
  assign w22849 = \pi26 ^ w22848 ;
  assign w22850 = ( \pi29 & \pi31 ) | ( \pi29 & ~w18914 ) | ( \pi31 & ~w18914 ) ;
  assign w22851 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22850 ) | ( ~\pi30 & w22850 ) ;
  assign w22852 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22850 ) | ( \pi30 & w22850 ) ;
  assign w22853 = ( ~\pi29 & w16617 ) | ( ~\pi29 & w22852 ) | ( w16617 & w22852 ) ;
  assign w22854 = ( w18916 & w22852 ) | ( w18916 & ~w22853 ) | ( w22852 & ~w22853 ) ;
  assign w22855 = ~\pi31 & w22854 ;
  assign w22856 = ( w22851 & w22853 ) | ( w22851 & w22855 ) | ( w22853 & w22855 ) ;
  assign w22857 = ( w37 & ~w19366 ) | ( w37 & w22856 ) | ( ~w19366 & w22856 ) ;
  assign w22858 = w22856 | w22857 ;
  assign w22859 = w16576 ^ w20404 ;
  assign w22860 = ( \pi23 & w16576 ) | ( \pi23 & ~w22859 ) | ( w16576 & ~w22859 ) ;
  assign w22861 = w1181 | w4797 ;
  assign w22862 = ( ~w1181 & w1814 ) | ( ~w1181 & w10517 ) | ( w1814 & w10517 ) ;
  assign w22863 = w22861 | w22862 ;
  assign w22864 = w956 | w3949 ;
  assign w22865 = w4099 & ~w22864 ;
  assign w22866 = ( w270 & w4099 ) | ( w270 & w22863 ) | ( w4099 & w22863 ) ;
  assign w22867 = w22865 & ~w22866 ;
  assign w22868 = ~w168 & w22867 ;
  assign w22869 = ( ~w168 & w408 ) | ( ~w168 & w509 ) | ( w408 & w509 ) ;
  assign w22870 = w22868 & ~w22869 ;
  assign w22871 = ~w1540 & w22870 ;
  assign w22872 = ( w516 & w570 ) | ( w516 & ~w837 ) | ( w570 & ~w837 ) ;
  assign w22873 = ~w205 & w22871 ;
  assign w22874 = ( ~w205 & w837 ) | ( ~w205 & w1031 ) | ( w837 & w1031 ) ;
  assign w22875 = w22873 & ~w22874 ;
  assign w22876 = ~w22872 & w22875 ;
  assign w22877 = w22860 ^ w22876 ;
  assign w22878 = w22785 ^ w22877 ;
  assign w22879 = w22786 ^ w22878 ;
  assign w22880 = w22858 ^ w22879 ;
  assign w22881 = ( ~w22788 & w22797 ) | ( ~w22788 & w22798 ) | ( w22797 & w22798 ) ;
  assign w22882 = ~w3717 & w19529 ;
  assign w22883 = w3649 & ~w18912 ;
  assign w22884 = ( w19529 & ~w22882 ) | ( w19529 & w22883 ) | ( ~w22882 & w22883 ) ;
  assign w22885 = ~w3549 & w19713 ;
  assign w22886 = w19723 | w22884 ;
  assign w22887 = ( w3448 & w22884 ) | ( w3448 & w22886 ) | ( w22884 & w22886 ) ;
  assign w22888 = ( w19713 & ~w22885 ) | ( w19713 & w22887 ) | ( ~w22885 & w22887 ) ;
  assign w22889 = \pi29 ^ w22888 ;
  assign w22890 = w22880 ^ w22881 ;
  assign w22891 = w22889 ^ w22890 ;
  assign w22892 = w22841 ^ w22891 ;
  assign w22893 = w22849 ^ w22892 ;
  assign w22894 = w22836 ^ w22840 ;
  assign w22895 = w22893 ^ w22894 ;
  assign w22896 = w22834 & ~w22895 ;
  assign w22897 = w22834 ^ w22895 ;
  assign w22898 = ( ~w22880 & w22881 ) | ( ~w22880 & w22889 ) | ( w22881 & w22889 ) ;
  assign w22899 = ( \pi29 & \pi31 ) | ( \pi29 & w18916 ) | ( \pi31 & w18916 ) ;
  assign w22900 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22899 ) | ( ~\pi30 & w22899 ) ;
  assign w22901 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22899 ) | ( \pi30 & w22899 ) ;
  assign w22902 = ( \pi29 & w18914 ) | ( \pi29 & ~w22901 ) | ( w18914 & ~w22901 ) ;
  assign w22903 = ( ~w18912 & w22901 ) | ( ~w18912 & w22902 ) | ( w22901 & w22902 ) ;
  assign w22904 = ~\pi31 & w22903 ;
  assign w22905 = ( w22900 & ~w22902 ) | ( w22900 & w22904 ) | ( ~w22902 & w22904 ) ;
  assign w22906 = ( w37 & ~w18929 ) | ( w37 & w22905 ) | ( ~w18929 & w22905 ) ;
  assign w22907 = w22905 | w22906 ;
  assign w22908 = ( w22785 & w22860 ) | ( w22785 & w22876 ) | ( w22860 & w22876 ) ;
  assign w22909 = w674 | w901 ;
  assign w22910 = w221 | w22909 ;
  assign w22911 = ( ~w221 & w640 ) | ( ~w221 & w1165 ) | ( w640 & w1165 ) ;
  assign w22912 = w22910 | w22911 ;
  assign w22913 = ( ~w51 & w18888 ) | ( ~w51 & w22912 ) | ( w18888 & w22912 ) ;
  assign w22914 = w6244 | w12617 ;
  assign w22915 = ( w51 & w219 ) | ( w51 & ~w6244 ) | ( w219 & ~w6244 ) ;
  assign w22916 = w22914 | w22915 ;
  assign w22917 = w22913 | w22916 ;
  assign w22918 = ( w1208 & w1400 ) | ( w1208 & ~w1566 ) | ( w1400 & ~w1566 ) ;
  assign w22919 = w4026 | w22917 ;
  assign w22920 = ( w1566 & ~w4026 ) | ( w1566 & w4092 ) | ( ~w4026 & w4092 ) ;
  assign w22921 = w22919 | w22920 ;
  assign w22922 = w22918 | w22921 ;
  assign w22923 = w64 | w413 ;
  assign w22924 = ( ~w64 & w1837 ) | ( ~w64 & w22922 ) | ( w1837 & w22922 ) ;
  assign w22925 = w22923 | w22924 ;
  assign w22926 = w227 | w463 ;
  assign w22927 = ( ~w227 & w280 ) | ( ~w227 & w22925 ) | ( w280 & w22925 ) ;
  assign w22928 = w22926 | w22927 ;
  assign w22929 = w22907 ^ w22908 ;
  assign w22930 = w22928 ^ w22929 ;
  assign w22931 = ( w22786 & w22858 ) | ( w22786 & ~w22878 ) | ( w22858 & ~w22878 ) ;
  assign w22932 = ~w3717 & w19713 ;
  assign w22933 = w3649 & w19529 ;
  assign w22934 = ( w19713 & ~w22932 ) | ( w19713 & w22933 ) | ( ~w22932 & w22933 ) ;
  assign w22935 = ~w3549 & w19887 ;
  assign w22936 = w19898 | w22934 ;
  assign w22937 = ( w3448 & w22934 ) | ( w3448 & w22936 ) | ( w22934 & w22936 ) ;
  assign w22938 = ( w19887 & ~w22935 ) | ( w19887 & w22937 ) | ( ~w22935 & w22937 ) ;
  assign w22939 = \pi29 ^ w22938 ;
  assign w22940 = w22930 ^ w22931 ;
  assign w22941 = w22939 ^ w22940 ;
  assign w22942 = ~w4143 & w20247 ;
  assign w22943 = w4052 & ~w20068 ;
  assign w22944 = ( w20247 & ~w22942 ) | ( w20247 & w22943 ) | ( ~w22942 & w22943 ) ;
  assign w22945 = ~w4147 & w20417 ;
  assign w22946 = w20404 | w22944 ;
  assign w22947 = ( w3964 & w22944 ) | ( w3964 & w22946 ) | ( w22944 & w22946 ) ;
  assign w22948 = ( w20417 & ~w22945 ) | ( w20417 & w22947 ) | ( ~w22945 & w22947 ) ;
  assign w22949 = \pi26 ^ w22948 ;
  assign w22950 = w22898 ^ w22941 ;
  assign w22951 = w22949 ^ w22950 ;
  assign w22952 = ( w22841 & w22849 ) | ( w22841 & ~w22891 ) | ( w22849 & ~w22891 ) ;
  assign w22953 = ( w22836 & w22840 ) | ( w22836 & ~w22893 ) | ( w22840 & ~w22893 ) ;
  assign w22954 = w22951 ^ w22953 ;
  assign w22955 = w22952 ^ w22954 ;
  assign w22956 = w22896 ^ w22955 ;
  assign w22957 = w22896 & w22955 ;
  assign w22958 = ( w22951 & w22952 ) | ( w22951 & w22953 ) | ( w22952 & w22953 ) ;
  assign w22959 = ( w22898 & w22941 ) | ( w22898 & w22949 ) | ( w22941 & w22949 ) ;
  assign w22960 = ( ~w22907 & w22908 ) | ( ~w22907 & w22928 ) | ( w22908 & w22928 ) ;
  assign w22961 = ( w2371 & w3927 ) | ( w2371 & w18888 ) | ( w3927 & w18888 ) ;
  assign w22962 = w3937 | w10423 ;
  assign w22963 = ( w3927 & ~w4101 ) | ( w3927 & w10423 ) | ( ~w4101 & w10423 ) ;
  assign w22964 = ~w22962 & w22963 ;
  assign w22965 = ~w22961 & w22964 ;
  assign w22966 = ( w837 & ~w4073 ) | ( w837 & w22965 ) | ( ~w4073 & w22965 ) ;
  assign w22967 = ~w837 & w22966 ;
  assign w22968 = w22928 ^ w22960 ;
  assign w22969 = w22967 ^ w22968 ;
  assign w22970 = ( \pi29 & \pi31 ) | ( \pi29 & ~w18912 ) | ( \pi31 & ~w18912 ) ;
  assign w22971 = ( \pi29 & ~\pi30 ) | ( \pi29 & w22970 ) | ( ~\pi30 & w22970 ) ;
  assign w22972 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w22970 ) | ( \pi30 & w22970 ) ;
  assign w22973 = ( ~\pi29 & w18916 ) | ( ~\pi29 & w22972 ) | ( w18916 & w22972 ) ;
  assign w22974 = ( w19529 & w22972 ) | ( w19529 & ~w22973 ) | ( w22972 & ~w22973 ) ;
  assign w22975 = ~\pi31 & w22974 ;
  assign w22976 = ( w22971 & w22973 ) | ( w22971 & w22975 ) | ( w22973 & w22975 ) ;
  assign w22977 = ( w37 & ~w19540 ) | ( w37 & w22976 ) | ( ~w19540 & w22976 ) ;
  assign w22978 = w22976 | w22977 ;
  assign w22979 = ( w22930 & w22931 ) | ( w22930 & w22939 ) | ( w22931 & w22939 ) ;
  assign w22980 = w22969 ^ w22979 ;
  assign w22981 = w22978 ^ w22980 ;
  assign w22982 = ~w4052 & w20247 ;
  assign w22983 = w18851 & w20404 ;
  assign w22984 = ( w20247 & ~w22982 ) | ( w20247 & w22983 ) | ( ~w22982 & w22983 ) ;
  assign w22985 = ~w4147 & w20414 ;
  assign w22986 = ( w20414 & w22984 ) | ( w20414 & ~w22985 ) | ( w22984 & ~w22985 ) ;
  assign w22987 = \pi26 ^ w22986 ;
  assign w22988 = ~w3717 & w19887 ;
  assign w22989 = w3649 & w19713 ;
  assign w22990 = ( w19887 & ~w22988 ) | ( w19887 & w22989 ) | ( ~w22988 & w22989 ) ;
  assign w22991 = w3549 | w20068 ;
  assign w22992 = w20081 & ~w22990 ;
  assign w22993 = ( w3448 & w22990 ) | ( w3448 & ~w22992 ) | ( w22990 & ~w22992 ) ;
  assign w22994 = ( ~w20068 & w22991 ) | ( ~w20068 & w22993 ) | ( w22991 & w22993 ) ;
  assign w22995 = \pi29 ^ w22994 ;
  assign w22996 = w22981 ^ w22987 ;
  assign w22997 = w22995 ^ w22996 ;
  assign w22998 = w22959 ^ w22997 ;
  assign w22999 = w22957 ^ w22998 ;
  assign w23000 = w22958 ^ w22999 ;
  assign w23001 = w3717 | w20068 ;
  assign w23002 = w3649 & w19887 ;
  assign w23003 = ( ~w20068 & w23001 ) | ( ~w20068 & w23002 ) | ( w23001 & w23002 ) ;
  assign w23004 = ~w3549 & w20247 ;
  assign w23005 = w3448 | w20257 ;
  assign w23006 = ( ~w20257 & w23003 ) | ( ~w20257 & w23005 ) | ( w23003 & w23005 ) ;
  assign w23007 = ( w20247 & ~w23004 ) | ( w20247 & w23006 ) | ( ~w23004 & w23006 ) ;
  assign w23008 = ( \pi29 & \pi31 ) | ( \pi29 & w19529 ) | ( \pi31 & w19529 ) ;
  assign w23009 = ( \pi29 & ~\pi30 ) | ( \pi29 & w23008 ) | ( ~\pi30 & w23008 ) ;
  assign w23010 = ( ~\pi29 & \pi30 ) | ( ~\pi29 & w23008 ) | ( \pi30 & w23008 ) ;
  assign w23011 = ( \pi29 & w18912 ) | ( \pi29 & ~w23010 ) | ( w18912 & ~w23010 ) ;
  assign w23012 = ( w19713 & w23010 ) | ( w19713 & w23011 ) | ( w23010 & w23011 ) ;
  assign w23013 = ~\pi31 & w23012 ;
  assign w23014 = ( w23009 & ~w23011 ) | ( w23009 & w23013 ) | ( ~w23011 & w23013 ) ;
  assign w23015 = w19723 | w23014 ;
  assign w23016 = ( w37 & w23014 ) | ( w37 & w23015 ) | ( w23014 & w23015 ) ;
  assign w23017 = ( w22928 & w22960 ) | ( w22928 & w22967 ) | ( w22960 & w22967 ) ;
  assign w23018 = w23016 ^ w23017 ;
  assign w23019 = w23007 ^ w23018 ;
  assign w23020 = ( ~w22969 & w22978 ) | ( ~w22969 & w22979 ) | ( w22978 & w22979 ) ;
  assign w23021 = w23019 ^ w23020 ;
  assign w23022 = \pi29 ^ w23021 ;
  assign w23023 = ~w4052 & w18851 ;
  assign w23024 = ( w4052 & ~w4147 ) | ( w4052 & w23023 ) | ( ~w4147 & w23023 ) ;
  assign w23025 = ( w4147 & w20404 ) | ( w4147 & w23024 ) | ( w20404 & w23024 ) ;
  assign w23026 = w22928 ^ w23025 ;
  assign w23027 = \pi26 ^ w23026 ;
  assign w23028 = w605 | w3959 ;
  assign w23029 = w4596 | w23028 ;
  assign w23030 = w23027 ^ w23029 ;
  assign w23031 = ( ~w22981 & w22987 ) | ( ~w22981 & w22995 ) | ( w22987 & w22995 ) ;
  assign w23032 = w23022 ^ w23030 ;
  assign w23033 = w23031 ^ w23032 ;
  assign w23034 = w22957 ^ w22958 ;
  assign w23035 = ( w22957 & w22958 ) | ( w22957 & ~w23034 ) | ( w22958 & ~w23034 ) ;
  assign w23036 = w23033 ^ w23035 ;
  assign w23037 = ( w22959 & ~w22997 ) | ( w22959 & w23034 ) | ( ~w22997 & w23034 ) ;
  assign w23038 = w23036 ^ w23037 ;
  assign \po00 = w19548 ;
  assign \po01 = w19730 ;
  assign \po02 = ~w19905 ;
  assign \po03 = ~w20088 ;
  assign \po04 = ~w20264 ;
  assign \po05 = ~w20424 ;
  assign \po06 = ~w20579 ;
  assign \po07 = ~w20722 ;
  assign \po08 = w20868 ;
  assign \po09 = w21001 ;
  assign \po10 = w21136 ;
  assign \po11 = w21282 ;
  assign \po12 = ~w21425 ;
  assign \po13 = ~w21544 ;
  assign \po14 = ~w21658 ;
  assign \po15 = w21776 ;
  assign \po16 = ~w21885 ;
  assign \po17 = w21987 ;
  assign \po18 = ~w22091 ;
  assign \po19 = ~w22184 ;
  assign \po20 = ~w22275 ;
  assign \po21 = w22368 ;
  assign \po22 = w22455 ;
  assign \po23 = ~w22537 ;
  assign \po24 = ~w22618 ;
  assign \po25 = ~w22697 ;
  assign \po26 = w22765 ;
  assign \po27 = ~w22835 ;
  assign \po28 = ~w22897 ;
  assign \po29 = w22956 ;
  assign \po30 = ~w23000 ;
  assign \po31 = w23038 ;
endmodule
