module multiplier( \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 , \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 );
  input \pi000 , \pi001 , \pi002 , \pi003 , \pi004 , \pi005 , \pi006 , \pi007 , \pi008 , \pi009 , \pi010 , \pi011 , \pi012 , \pi013 , \pi014 , \pi015 , \pi016 , \pi017 , \pi018 , \pi019 , \pi020 , \pi021 , \pi022 , \pi023 , \pi024 , \pi025 , \pi026 , \pi027 , \pi028 , \pi029 , \pi030 , \pi031 , \pi032 , \pi033 , \pi034 , \pi035 , \pi036 , \pi037 , \pi038 , \pi039 , \pi040 , \pi041 , \pi042 , \pi043 , \pi044 , \pi045 , \pi046 , \pi047 , \pi048 , \pi049 , \pi050 , \pi051 , \pi052 , \pi053 , \pi054 , \pi055 , \pi056 , \pi057 , \pi058 , \pi059 , \pi060 , \pi061 , \pi062 , \pi063 , \pi064 , \pi065 , \pi066 , \pi067 , \pi068 , \pi069 , \pi070 , \pi071 , \pi072 , \pi073 , \pi074 , \pi075 , \pi076 , \pi077 , \pi078 , \pi079 , \pi080 , \pi081 , \pi082 , \pi083 , \pi084 , \pi085 , \pi086 , \pi087 , \pi088 , \pi089 , \pi090 , \pi091 , \pi092 , \pi093 , \pi094 , \pi095 , \pi096 , \pi097 , \pi098 , \pi099 , \pi100 , \pi101 , \pi102 , \pi103 , \pi104 , \pi105 , \pi106 , \pi107 , \pi108 , \pi109 , \pi110 , \pi111 , \pi112 , \pi113 , \pi114 , \pi115 , \pi116 , \pi117 , \pi118 , \pi119 , \pi120 , \pi121 , \pi122 , \pi123 , \pi124 , \pi125 , \pi126 , \pi127 ;
  output \po000 , \po001 , \po002 , \po003 , \po004 , \po005 , \po006 , \po007 , \po008 , \po009 , \po010 , \po011 , \po012 , \po013 , \po014 , \po015 , \po016 , \po017 , \po018 , \po019 , \po020 , \po021 , \po022 , \po023 , \po024 , \po025 , \po026 , \po027 , \po028 , \po029 , \po030 , \po031 , \po032 , \po033 , \po034 , \po035 , \po036 , \po037 , \po038 , \po039 , \po040 , \po041 , \po042 , \po043 , \po044 , \po045 , \po046 , \po047 , \po048 , \po049 , \po050 , \po051 , \po052 , \po053 , \po054 , \po055 , \po056 , \po057 , \po058 , \po059 , \po060 , \po061 , \po062 , \po063 , \po064 , \po065 , \po066 , \po067 , \po068 , \po069 , \po070 , \po071 , \po072 , \po073 , \po074 , \po075 , \po076 , \po077 , \po078 , \po079 , \po080 , \po081 , \po082 , \po083 , \po084 , \po085 , \po086 , \po087 , \po088 , \po089 , \po090 , \po091 , \po092 , \po093 , \po094 , \po095 , \po096 , \po097 , \po098 , \po099 , \po100 , \po101 , \po102 , \po103 , \po104 , \po105 , \po106 , \po107 , \po108 , \po109 , \po110 , \po111 , \po112 , \po113 , \po114 , \po115 , \po116 , \po117 , \po118 , \po119 , \po120 , \po121 , \po122 , \po123 , \po124 , \po125 , \po126 , \po127 ;
  wire zero , w129 , w130 , w131 , w132 , w133 , w134 , w135 , w136 , w137 , w138 , w139 , w140 , w141 , w142 , w143 , w144 , w145 , w146 , w147 , w148 , w149 , w150 , w151 , w152 , w153 , w154 , w155 , w156 , w157 , w158 , w159 , w160 , w161 , w162 , w163 , w164 , w165 , w166 , w167 , w168 , w169 , w170 , w171 , w172 , w173 , w174 , w175 , w176 , w177 , w178 , w179 , w180 , w181 , w182 , w183 , w184 , w185 , w186 , w187 , w188 , w189 , w190 , w191 , w192 , w193 , w194 , w195 , w196 , w197 , w198 , w199 , w200 , w201 , w202 , w203 , w204 , w205 , w206 , w207 , w208 , w209 , w210 , w211 , w212 , w213 , w214 , w215 , w216 , w217 , w218 , w219 , w220 , w221 , w222 , w223 , w224 , w225 , w226 , w227 , w228 , w229 , w230 , w231 , w232 , w233 , w234 , w235 , w236 , w237 , w238 , w239 , w240 , w241 , w242 , w243 , w244 , w245 , w246 , w247 , w248 , w249 , w250 , w251 , w252 , w253 , w254 , w255 , w256 , w257 , w258 , w259 , w260 , w261 , w262 , w263 , w264 , w265 , w266 , w267 , w268 , w269 , w270 , w271 , w272 , w273 , w274 , w275 , w276 , w277 , w278 , w279 , w280 , w281 , w282 , w283 , w284 , w285 , w286 , w287 , w288 , w289 , w290 , w291 , w292 , w293 , w294 , w295 , w296 , w297 , w298 , w299 , w300 , w301 , w302 , w303 , w304 , w305 , w306 , w307 , w308 , w309 , w310 , w311 , w312 , w313 , w314 , w315 , w316 , w317 , w318 , w319 , w320 , w321 , w322 , w323 , w324 , w325 , w326 , w327 , w328 , w329 , w330 , w331 , w332 , w333 , w334 , w335 , w336 , w337 , w338 , w339 , w340 , w341 , w342 , w343 , w344 , w345 , w346 , w347 , w348 , w349 , w350 , w351 , w352 , w353 , w354 , w355 , w356 , w357 , w358 , w359 , w360 , w361 , w362 , w363 , w364 , w365 , w366 , w367 , w368 , w369 , w370 , w371 , w372 , w373 , w374 , w375 , w376 , w377 , w378 , w379 , w380 , w381 , w382 , w383 , w384 , w385 , w386 , w387 , w388 , w389 , w390 , w391 , w392 , w393 , w394 , w395 , w396 , w397 , w398 , w399 , w400 , w401 , w402 , w403 , w404 , w405 , w406 , w407 , w408 , w409 , w410 , w411 , w412 , w413 , w414 , w415 , w416 , w417 , w418 , w419 , w420 , w421 , w422 , w423 , w424 , w425 , w426 , w427 , w428 , w429 , w430 , w431 , w432 , w433 , w434 , w435 , w436 , w437 , w438 , w439 , w440 , w441 , w442 , w443 , w444 , w445 , w446 , w447 , w448 , w449 , w450 , w451 , w452 , w453 , w454 , w455 , w456 , w457 , w458 , w459 , w460 , w461 , w462 , w463 , w464 , w465 , w466 , w467 , w468 , w469 , w470 , w471 , w472 , w473 , w474 , w475 , w476 , w477 , w478 , w479 , w480 , w481 , w482 , w483 , w484 , w485 , w486 , w487 , w488 , w489 , w490 , w491 , w492 , w493 , w494 , w495 , w496 , w497 , w498 , w499 , w500 , w501 , w502 , w503 , w504 , w505 , w506 , w507 , w508 , w509 , w510 , w511 , w512 , w513 , w514 , w515 , w516 , w517 , w518 , w519 , w520 , w521 , w522 , w523 , w524 , w525 , w526 , w527 , w528 , w529 , w530 , w531 , w532 , w533 , w534 , w535 , w536 , w537 , w538 , w539 , w540 , w541 , w542 , w543 , w544 , w545 , w546 , w547 , w548 , w549 , w550 , w551 , w552 , w553 , w554 , w555 , w556 , w557 , w558 , w559 , w560 , w561 , w562 , w563 , w564 , w565 , w566 , w567 , w568 , w569 , w570 , w571 , w572 , w573 , w574 , w575 , w576 , w577 , w578 , w579 , w580 , w581 , w582 , w583 , w584 , w585 , w586 , w587 , w588 , w589 , w590 , w591 , w592 , w593 , w594 , w595 , w596 , w597 , w598 , w599 , w600 , w601 , w602 , w603 , w604 , w605 , w606 , w607 , w608 , w609 , w610 , w611 , w612 , w613 , w614 , w615 , w616 , w617 , w618 , w619 , w620 , w621 , w622 , w623 , w624 , w625 , w626 , w627 , w628 , w629 , w630 , w631 , w632 , w633 , w634 , w635 , w636 , w637 , w638 , w639 , w640 , w641 , w642 , w643 , w644 , w645 , w646 , w647 , w648 , w649 , w650 , w651 , w652 , w653 , w654 , w655 , w656 , w657 , w658 , w659 , w660 , w661 , w662 , w663 , w664 , w665 , w666 , w667 , w668 , w669 , w670 , w671 , w672 , w673 , w674 , w675 , w676 , w677 , w678 , w679 , w680 , w681 , w682 , w683 , w684 , w685 , w686 , w687 , w688 , w689 , w690 , w691 , w692 , w693 , w694 , w695 , w696 , w697 , w698 , w699 , w700 , w701 , w702 , w703 , w704 , w705 , w706 , w707 , w708 , w709 , w710 , w711 , w712 , w713 , w714 , w715 , w716 , w717 , w718 , w719 , w720 , w721 , w722 , w723 , w724 , w725 , w726 , w727 , w728 , w729 , w730 , w731 , w732 , w733 , w734 , w735 , w736 , w737 , w738 , w739 , w740 , w741 , w742 , w743 , w744 , w745 , w746 , w747 , w748 , w749 , w750 , w751 , w752 , w753 , w754 , w755 , w756 , w757 , w758 , w759 , w760 , w761 , w762 , w763 , w764 , w765 , w766 , w767 , w768 , w769 , w770 , w771 , w772 , w773 , w774 , w775 , w776 , w777 , w778 , w779 , w780 , w781 , w782 , w783 , w784 , w785 , w786 , w787 , w788 , w789 , w790 , w791 , w792 , w793 , w794 , w795 , w796 , w797 , w798 , w799 , w800 , w801 , w802 , w803 , w804 , w805 , w806 , w807 , w808 , w809 , w810 , w811 , w812 , w813 , w814 , w815 , w816 , w817 , w818 , w819 , w820 , w821 , w822 , w823 , w824 , w825 , w826 , w827 , w828 , w829 , w830 , w831 , w832 , w833 , w834 , w835 , w836 , w837 , w838 , w839 , w840 , w841 , w842 , w843 , w844 , w845 , w846 , w847 , w848 , w849 , w850 , w851 , w852 , w853 , w854 , w855 , w856 , w857 , w858 , w859 , w860 , w861 , w862 , w863 , w864 , w865 , w866 , w867 , w868 , w869 , w870 , w871 , w872 , w873 , w874 , w875 , w876 , w877 , w878 , w879 , w880 , w881 , w882 , w883 , w884 , w885 , w886 , w887 , w888 , w889 , w890 , w891 , w892 , w893 , w894 , w895 , w896 , w897 , w898 , w899 , w900 , w901 , w902 , w903 , w904 , w905 , w906 , w907 , w908 , w909 , w910 , w911 , w912 , w913 , w914 , w915 , w916 , w917 , w918 , w919 , w920 , w921 , w922 , w923 , w924 , w925 , w926 , w927 , w928 , w929 , w930 , w931 , w932 , w933 , w934 , w935 , w936 , w937 , w938 , w939 , w940 , w941 , w942 , w943 , w944 , w945 , w946 , w947 , w948 , w949 , w950 , w951 , w952 , w953 , w954 , w955 , w956 , w957 , w958 , w959 , w960 , w961 , w962 , w963 , w964 , w965 , w966 , w967 , w968 , w969 , w970 , w971 , w972 , w973 , w974 , w975 , w976 , w977 , w978 , w979 , w980 , w981 , w982 , w983 , w984 , w985 , w986 , w987 , w988 , w989 , w990 , w991 , w992 , w993 , w994 , w995 , w996 , w997 , w998 , w999 , w1000 , w1001 , w1002 , w1003 , w1004 , w1005 , w1006 , w1007 , w1008 , w1009 , w1010 , w1011 , w1012 , w1013 , w1014 , w1015 , w1016 , w1017 , w1018 , w1019 , w1020 , w1021 , w1022 , w1023 , w1024 , w1025 , w1026 , w1027 , w1028 , w1029 , w1030 , w1031 , w1032 , w1033 , w1034 , w1035 , w1036 , w1037 , w1038 , w1039 , w1040 , w1041 , w1042 , w1043 , w1044 , w1045 , w1046 , w1047 , w1048 , w1049 , w1050 , w1051 , w1052 , w1053 , w1054 , w1055 , w1056 , w1057 , w1058 , w1059 , w1060 , w1061 , w1062 , w1063 , w1064 , w1065 , w1066 , w1067 , w1068 , w1069 , w1070 , w1071 , w1072 , w1073 , w1074 , w1075 , w1076 , w1077 , w1078 , w1079 , w1080 , w1081 , w1082 , w1083 , w1084 , w1085 , w1086 , w1087 , w1088 , w1089 , w1090 , w1091 , w1092 , w1093 , w1094 , w1095 , w1096 , w1097 , w1098 , w1099 , w1100 , w1101 , w1102 , w1103 , w1104 , w1105 , w1106 , w1107 , w1108 , w1109 , w1110 , w1111 , w1112 , w1113 , w1114 , w1115 , w1116 , w1117 , w1118 , w1119 , w1120 , w1121 , w1122 , w1123 , w1124 , w1125 , w1126 , w1127 , w1128 , w1129 , w1130 , w1131 , w1132 , w1133 , w1134 , w1135 , w1136 , w1137 , w1138 , w1139 , w1140 , w1141 , w1142 , w1143 , w1144 , w1145 , w1146 , w1147 , w1148 , w1149 , w1150 , w1151 , w1152 , w1153 , w1154 , w1155 , w1156 , w1157 , w1158 , w1159 , w1160 , w1161 , w1162 , w1163 , w1164 , w1165 , w1166 , w1167 , w1168 , w1169 , w1170 , w1171 , w1172 , w1173 , w1174 , w1175 , w1176 , w1177 , w1178 , w1179 , w1180 , w1181 , w1182 , w1183 , w1184 , w1185 , w1186 , w1187 , w1188 , w1189 , w1190 , w1191 , w1192 , w1193 , w1194 , w1195 , w1196 , w1197 , w1198 , w1199 , w1200 , w1201 , w1202 , w1203 , w1204 , w1205 , w1206 , w1207 , w1208 , w1209 , w1210 , w1211 , w1212 , w1213 , w1214 , w1215 , w1216 , w1217 , w1218 , w1219 , w1220 , w1221 , w1222 , w1223 , w1224 , w1225 , w1226 , w1227 , w1228 , w1229 , w1230 , w1231 , w1232 , w1233 , w1234 , w1235 , w1236 , w1237 , w1238 , w1239 , w1240 , w1241 , w1242 , w1243 , w1244 , w1245 , w1246 , w1247 , w1248 , w1249 , w1250 , w1251 , w1252 , w1253 , w1254 , w1255 , w1256 , w1257 , w1258 , w1259 , w1260 , w1261 , w1262 , w1263 , w1264 , w1265 , w1266 , w1267 , w1268 , w1269 , w1270 , w1271 , w1272 , w1273 , w1274 , w1275 , w1276 , w1277 , w1278 , w1279 , w1280 , w1281 , w1282 , w1283 , w1284 , w1285 , w1286 , w1287 , w1288 , w1289 , w1290 , w1291 , w1292 , w1293 , w1294 , w1295 , w1296 , w1297 , w1298 , w1299 , w1300 , w1301 , w1302 , w1303 , w1304 , w1305 , w1306 , w1307 , w1308 , w1309 , w1310 , w1311 , w1312 , w1313 , w1314 , w1315 , w1316 , w1317 , w1318 , w1319 , w1320 , w1321 , w1322 , w1323 , w1324 , w1325 , w1326 , w1327 , w1328 , w1329 , w1330 , w1331 , w1332 , w1333 , w1334 , w1335 , w1336 , w1337 , w1338 , w1339 , w1340 , w1341 , w1342 , w1343 , w1344 , w1345 , w1346 , w1347 , w1348 , w1349 , w1350 , w1351 , w1352 , w1353 , w1354 , w1355 , w1356 , w1357 , w1358 , w1359 , w1360 , w1361 , w1362 , w1363 , w1364 , w1365 , w1366 , w1367 , w1368 , w1369 , w1370 , w1371 , w1372 , w1373 , w1374 , w1375 , w1376 , w1377 , w1378 , w1379 , w1380 , w1381 , w1382 , w1383 , w1384 , w1385 , w1386 , w1387 , w1388 , w1389 , w1390 , w1391 , w1392 , w1393 , w1394 , w1395 , w1396 , w1397 , w1398 , w1399 , w1400 , w1401 , w1402 , w1403 , w1404 , w1405 , w1406 , w1407 , w1408 , w1409 , w1410 , w1411 , w1412 , w1413 , w1414 , w1415 , w1416 , w1417 , w1418 , w1419 , w1420 , w1421 , w1422 , w1423 , w1424 , w1425 , w1426 , w1427 , w1428 , w1429 , w1430 , w1431 , w1432 , w1433 , w1434 , w1435 , w1436 , w1437 , w1438 , w1439 , w1440 , w1441 , w1442 , w1443 , w1444 , w1445 , w1446 , w1447 , w1448 , w1449 , w1450 , w1451 , w1452 , w1453 , w1454 , w1455 , w1456 , w1457 , w1458 , w1459 , w1460 , w1461 , w1462 , w1463 , w1464 , w1465 , w1466 , w1467 , w1468 , w1469 , w1470 , w1471 , w1472 , w1473 , w1474 , w1475 , w1476 , w1477 , w1478 , w1479 , w1480 , w1481 , w1482 , w1483 , w1484 , w1485 , w1486 , w1487 , w1488 , w1489 , w1490 , w1491 , w1492 , w1493 , w1494 , w1495 , w1496 , w1497 , w1498 , w1499 , w1500 , w1501 , w1502 , w1503 , w1504 , w1505 , w1506 , w1507 , w1508 , w1509 , w1510 , w1511 , w1512 , w1513 , w1514 , w1515 , w1516 , w1517 , w1518 , w1519 , w1520 , w1521 , w1522 , w1523 , w1524 , w1525 , w1526 , w1527 , w1528 , w1529 , w1530 , w1531 , w1532 , w1533 , w1534 , w1535 , w1536 , w1537 , w1538 , w1539 , w1540 , w1541 , w1542 , w1543 , w1544 , w1545 , w1546 , w1547 , w1548 , w1549 , w1550 , w1551 , w1552 , w1553 , w1554 , w1555 , w1556 , w1557 , w1558 , w1559 , w1560 , w1561 , w1562 , w1563 , w1564 , w1565 , w1566 , w1567 , w1568 , w1569 , w1570 , w1571 , w1572 , w1573 , w1574 , w1575 , w1576 , w1577 , w1578 , w1579 , w1580 , w1581 , w1582 , w1583 , w1584 , w1585 , w1586 , w1587 , w1588 , w1589 , w1590 , w1591 , w1592 , w1593 , w1594 , w1595 , w1596 , w1597 , w1598 , w1599 , w1600 , w1601 , w1602 , w1603 , w1604 , w1605 , w1606 , w1607 , w1608 , w1609 , w1610 , w1611 , w1612 , w1613 , w1614 , w1615 , w1616 , w1617 , w1618 , w1619 , w1620 , w1621 , w1622 , w1623 , w1624 , w1625 , w1626 , w1627 , w1628 , w1629 , w1630 , w1631 , w1632 , w1633 , w1634 , w1635 , w1636 , w1637 , w1638 , w1639 , w1640 , w1641 , w1642 , w1643 , w1644 , w1645 , w1646 , w1647 , w1648 , w1649 , w1650 , w1651 , w1652 , w1653 , w1654 , w1655 , w1656 , w1657 , w1658 , w1659 , w1660 , w1661 , w1662 , w1663 , w1664 , w1665 , w1666 , w1667 , w1668 , w1669 , w1670 , w1671 , w1672 , w1673 , w1674 , w1675 , w1676 , w1677 , w1678 , w1679 , w1680 , w1681 , w1682 , w1683 , w1684 , w1685 , w1686 , w1687 , w1688 , w1689 , w1690 , w1691 , w1692 , w1693 , w1694 , w1695 , w1696 , w1697 , w1698 , w1699 , w1700 , w1701 , w1702 , w1703 , w1704 , w1705 , w1706 , w1707 , w1708 , w1709 , w1710 , w1711 , w1712 , w1713 , w1714 , w1715 , w1716 , w1717 , w1718 , w1719 , w1720 , w1721 , w1722 , w1723 , w1724 , w1725 , w1726 , w1727 , w1728 , w1729 , w1730 , w1731 , w1732 , w1733 , w1734 , w1735 , w1736 , w1737 , w1738 , w1739 , w1740 , w1741 , w1742 , w1743 , w1744 , w1745 , w1746 , w1747 , w1748 , w1749 , w1750 , w1751 , w1752 , w1753 , w1754 , w1755 , w1756 , w1757 , w1758 , w1759 , w1760 , w1761 , w1762 , w1763 , w1764 , w1765 , w1766 , w1767 , w1768 , w1769 , w1770 , w1771 , w1772 , w1773 , w1774 , w1775 , w1776 , w1777 , w1778 , w1779 , w1780 , w1781 , w1782 , w1783 , w1784 , w1785 , w1786 , w1787 , w1788 , w1789 , w1790 , w1791 , w1792 , w1793 , w1794 , w1795 , w1796 , w1797 , w1798 , w1799 , w1800 , w1801 , w1802 , w1803 , w1804 , w1805 , w1806 , w1807 , w1808 , w1809 , w1810 , w1811 , w1812 , w1813 , w1814 , w1815 , w1816 , w1817 , w1818 , w1819 , w1820 , w1821 , w1822 , w1823 , w1824 , w1825 , w1826 , w1827 , w1828 , w1829 , w1830 , w1831 , w1832 , w1833 , w1834 , w1835 , w1836 , w1837 , w1838 , w1839 , w1840 , w1841 , w1842 , w1843 , w1844 , w1845 , w1846 , w1847 , w1848 , w1849 , w1850 , w1851 , w1852 , w1853 , w1854 , w1855 , w1856 , w1857 , w1858 , w1859 , w1860 , w1861 , w1862 , w1863 , w1864 , w1865 , w1866 , w1867 , w1868 , w1869 , w1870 , w1871 , w1872 , w1873 , w1874 , w1875 , w1876 , w1877 , w1878 , w1879 , w1880 , w1881 , w1882 , w1883 , w1884 , w1885 , w1886 , w1887 , w1888 , w1889 , w1890 , w1891 , w1892 , w1893 , w1894 , w1895 , w1896 , w1897 , w1898 , w1899 , w1900 , w1901 , w1902 , w1903 , w1904 , w1905 , w1906 , w1907 , w1908 , w1909 , w1910 , w1911 , w1912 , w1913 , w1914 , w1915 , w1916 , w1917 , w1918 , w1919 , w1920 , w1921 , w1922 , w1923 , w1924 , w1925 , w1926 , w1927 , w1928 , w1929 , w1930 , w1931 , w1932 , w1933 , w1934 , w1935 , w1936 , w1937 , w1938 , w1939 , w1940 , w1941 , w1942 , w1943 , w1944 , w1945 , w1946 , w1947 , w1948 , w1949 , w1950 , w1951 , w1952 , w1953 , w1954 , w1955 , w1956 , w1957 , w1958 , w1959 , w1960 , w1961 , w1962 , w1963 , w1964 , w1965 , w1966 , w1967 , w1968 , w1969 , w1970 , w1971 , w1972 , w1973 , w1974 , w1975 , w1976 , w1977 , w1978 , w1979 , w1980 , w1981 , w1982 , w1983 , w1984 , w1985 , w1986 , w1987 , w1988 , w1989 , w1990 , w1991 , w1992 , w1993 , w1994 , w1995 , w1996 , w1997 , w1998 , w1999 , w2000 , w2001 , w2002 , w2003 , w2004 , w2005 , w2006 , w2007 , w2008 , w2009 , w2010 , w2011 , w2012 , w2013 , w2014 , w2015 , w2016 , w2017 , w2018 , w2019 , w2020 , w2021 , w2022 , w2023 , w2024 , w2025 , w2026 , w2027 , w2028 , w2029 , w2030 , w2031 , w2032 , w2033 , w2034 , w2035 , w2036 , w2037 , w2038 , w2039 , w2040 , w2041 , w2042 , w2043 , w2044 , w2045 , w2046 , w2047 , w2048 , w2049 , w2050 , w2051 , w2052 , w2053 , w2054 , w2055 , w2056 , w2057 , w2058 , w2059 , w2060 , w2061 , w2062 , w2063 , w2064 , w2065 , w2066 , w2067 , w2068 , w2069 , w2070 , w2071 , w2072 , w2073 , w2074 , w2075 , w2076 , w2077 , w2078 , w2079 , w2080 , w2081 , w2082 , w2083 , w2084 , w2085 , w2086 , w2087 , w2088 , w2089 , w2090 , w2091 , w2092 , w2093 , w2094 , w2095 , w2096 , w2097 , w2098 , w2099 , w2100 , w2101 , w2102 , w2103 , w2104 , w2105 , w2106 , w2107 , w2108 , w2109 , w2110 , w2111 , w2112 , w2113 , w2114 , w2115 , w2116 , w2117 , w2118 , w2119 , w2120 , w2121 , w2122 , w2123 , w2124 , w2125 , w2126 , w2127 , w2128 , w2129 , w2130 , w2131 , w2132 , w2133 , w2134 , w2135 , w2136 , w2137 , w2138 , w2139 , w2140 , w2141 , w2142 , w2143 , w2144 , w2145 , w2146 , w2147 , w2148 , w2149 , w2150 , w2151 , w2152 , w2153 , w2154 , w2155 , w2156 , w2157 , w2158 , w2159 , w2160 , w2161 , w2162 , w2163 , w2164 , w2165 , w2166 , w2167 , w2168 , w2169 , w2170 , w2171 , w2172 , w2173 , w2174 , w2175 , w2176 , w2177 , w2178 , w2179 , w2180 , w2181 , w2182 , w2183 , w2184 , w2185 , w2186 , w2187 , w2188 , w2189 , w2190 , w2191 , w2192 , w2193 , w2194 , w2195 , w2196 , w2197 , w2198 , w2199 , w2200 , w2201 , w2202 , w2203 , w2204 , w2205 , w2206 , w2207 , w2208 , w2209 , w2210 , w2211 , w2212 , w2213 , w2214 , w2215 , w2216 , w2217 , w2218 , w2219 , w2220 , w2221 , w2222 , w2223 , w2224 , w2225 , w2226 , w2227 , w2228 , w2229 , w2230 , w2231 , w2232 , w2233 , w2234 , w2235 , w2236 , w2237 , w2238 , w2239 , w2240 , w2241 , w2242 , w2243 , w2244 , w2245 , w2246 , w2247 , w2248 , w2249 , w2250 , w2251 , w2252 , w2253 , w2254 , w2255 , w2256 , w2257 , w2258 , w2259 , w2260 , w2261 , w2262 , w2263 , w2264 , w2265 , w2266 , w2267 , w2268 , w2269 , w2270 , w2271 , w2272 , w2273 , w2274 , w2275 , w2276 , w2277 , w2278 , w2279 , w2280 , w2281 , w2282 , w2283 , w2284 , w2285 , w2286 , w2287 , w2288 , w2289 , w2290 , w2291 , w2292 , w2293 , w2294 , w2295 , w2296 , w2297 , w2298 , w2299 , w2300 , w2301 , w2302 , w2303 , w2304 , w2305 , w2306 , w2307 , w2308 , w2309 , w2310 , w2311 , w2312 , w2313 , w2314 , w2315 , w2316 , w2317 , w2318 , w2319 , w2320 , w2321 , w2322 , w2323 , w2324 , w2325 , w2326 , w2327 , w2328 , w2329 , w2330 , w2331 , w2332 , w2333 , w2334 , w2335 , w2336 , w2337 , w2338 , w2339 , w2340 , w2341 , w2342 , w2343 , w2344 , w2345 , w2346 , w2347 , w2348 , w2349 , w2350 , w2351 , w2352 , w2353 , w2354 , w2355 , w2356 , w2357 , w2358 , w2359 , w2360 , w2361 , w2362 , w2363 , w2364 , w2365 , w2366 , w2367 , w2368 , w2369 , w2370 , w2371 , w2372 , w2373 , w2374 , w2375 , w2376 , w2377 , w2378 , w2379 , w2380 , w2381 , w2382 , w2383 , w2384 , w2385 , w2386 , w2387 , w2388 , w2389 , w2390 , w2391 , w2392 , w2393 , w2394 , w2395 , w2396 , w2397 , w2398 , w2399 , w2400 , w2401 , w2402 , w2403 , w2404 , w2405 , w2406 , w2407 , w2408 , w2409 , w2410 , w2411 , w2412 , w2413 , w2414 , w2415 , w2416 , w2417 , w2418 , w2419 , w2420 , w2421 , w2422 , w2423 , w2424 , w2425 , w2426 , w2427 , w2428 , w2429 , w2430 , w2431 , w2432 , w2433 , w2434 , w2435 , w2436 , w2437 , w2438 , w2439 , w2440 , w2441 , w2442 , w2443 , w2444 , w2445 , w2446 , w2447 , w2448 , w2449 , w2450 , w2451 , w2452 , w2453 , w2454 , w2455 , w2456 , w2457 , w2458 , w2459 , w2460 , w2461 , w2462 , w2463 , w2464 , w2465 , w2466 , w2467 , w2468 , w2469 , w2470 , w2471 , w2472 , w2473 , w2474 , w2475 , w2476 , w2477 , w2478 , w2479 , w2480 , w2481 , w2482 , w2483 , w2484 , w2485 , w2486 , w2487 , w2488 , w2489 , w2490 , w2491 , w2492 , w2493 , w2494 , w2495 , w2496 , w2497 , w2498 , w2499 , w2500 , w2501 , w2502 , w2503 , w2504 , w2505 , w2506 , w2507 , w2508 , w2509 , w2510 , w2511 , w2512 , w2513 , w2514 , w2515 , w2516 , w2517 , w2518 , w2519 , w2520 , w2521 , w2522 , w2523 , w2524 , w2525 , w2526 , w2527 , w2528 , w2529 , w2530 , w2531 , w2532 , w2533 , w2534 , w2535 , w2536 , w2537 , w2538 , w2539 , w2540 , w2541 , w2542 , w2543 , w2544 , w2545 , w2546 , w2547 , w2548 , w2549 , w2550 , w2551 , w2552 , w2553 , w2554 , w2555 , w2556 , w2557 , w2558 , w2559 , w2560 , w2561 , w2562 , w2563 , w2564 , w2565 , w2566 , w2567 , w2568 , w2569 , w2570 , w2571 , w2572 , w2573 , w2574 , w2575 , w2576 , w2577 , w2578 , w2579 , w2580 , w2581 , w2582 , w2583 , w2584 , w2585 , w2586 , w2587 , w2588 , w2589 , w2590 , w2591 , w2592 , w2593 , w2594 , w2595 , w2596 , w2597 , w2598 , w2599 , w2600 , w2601 , w2602 , w2603 , w2604 , w2605 , w2606 , w2607 , w2608 , w2609 , w2610 , w2611 , w2612 , w2613 , w2614 , w2615 , w2616 , w2617 , w2618 , w2619 , w2620 , w2621 , w2622 , w2623 , w2624 , w2625 , w2626 , w2627 , w2628 , w2629 , w2630 , w2631 , w2632 , w2633 , w2634 , w2635 , w2636 , w2637 , w2638 , w2639 , w2640 , w2641 , w2642 , w2643 , w2644 , w2645 , w2646 , w2647 , w2648 , w2649 , w2650 , w2651 , w2652 , w2653 , w2654 , w2655 , w2656 , w2657 , w2658 , w2659 , w2660 , w2661 , w2662 , w2663 , w2664 , w2665 , w2666 , w2667 , w2668 , w2669 , w2670 , w2671 , w2672 , w2673 , w2674 , w2675 , w2676 , w2677 , w2678 , w2679 , w2680 , w2681 , w2682 , w2683 , w2684 , w2685 , w2686 , w2687 , w2688 , w2689 , w2690 , w2691 , w2692 , w2693 , w2694 , w2695 , w2696 , w2697 , w2698 , w2699 , w2700 , w2701 , w2702 , w2703 , w2704 , w2705 , w2706 , w2707 , w2708 , w2709 , w2710 , w2711 , w2712 , w2713 , w2714 , w2715 , w2716 , w2717 , w2718 , w2719 , w2720 , w2721 , w2722 , w2723 , w2724 , w2725 , w2726 , w2727 , w2728 , w2729 , w2730 , w2731 , w2732 , w2733 , w2734 , w2735 , w2736 , w2737 , w2738 , w2739 , w2740 , w2741 , w2742 , w2743 , w2744 , w2745 , w2746 , w2747 , w2748 , w2749 , w2750 , w2751 , w2752 , w2753 , w2754 , w2755 , w2756 , w2757 , w2758 , w2759 , w2760 , w2761 , w2762 , w2763 , w2764 , w2765 , w2766 , w2767 , w2768 , w2769 , w2770 , w2771 , w2772 , w2773 , w2774 , w2775 , w2776 , w2777 , w2778 , w2779 , w2780 , w2781 , w2782 , w2783 , w2784 , w2785 , w2786 , w2787 , w2788 , w2789 , w2790 , w2791 , w2792 , w2793 , w2794 , w2795 , w2796 , w2797 , w2798 , w2799 , w2800 , w2801 , w2802 , w2803 , w2804 , w2805 , w2806 , w2807 , w2808 , w2809 , w2810 , w2811 , w2812 , w2813 , w2814 , w2815 , w2816 , w2817 , w2818 , w2819 , w2820 , w2821 , w2822 , w2823 , w2824 , w2825 , w2826 , w2827 , w2828 , w2829 , w2830 , w2831 , w2832 , w2833 , w2834 , w2835 , w2836 , w2837 , w2838 , w2839 , w2840 , w2841 , w2842 , w2843 , w2844 , w2845 , w2846 , w2847 , w2848 , w2849 , w2850 , w2851 , w2852 , w2853 , w2854 , w2855 , w2856 , w2857 , w2858 , w2859 , w2860 , w2861 , w2862 , w2863 , w2864 , w2865 , w2866 , w2867 , w2868 , w2869 , w2870 , w2871 , w2872 , w2873 , w2874 , w2875 , w2876 , w2877 , w2878 , w2879 , w2880 , w2881 , w2882 , w2883 , w2884 , w2885 , w2886 , w2887 , w2888 , w2889 , w2890 , w2891 , w2892 , w2893 , w2894 , w2895 , w2896 , w2897 , w2898 , w2899 , w2900 , w2901 , w2902 , w2903 , w2904 , w2905 , w2906 , w2907 , w2908 , w2909 , w2910 , w2911 , w2912 , w2913 , w2914 , w2915 , w2916 , w2917 , w2918 , w2919 , w2920 , w2921 , w2922 , w2923 , w2924 , w2925 , w2926 , w2927 , w2928 , w2929 , w2930 , w2931 , w2932 , w2933 , w2934 , w2935 , w2936 , w2937 , w2938 , w2939 , w2940 , w2941 , w2942 , w2943 , w2944 , w2945 , w2946 , w2947 , w2948 , w2949 , w2950 , w2951 , w2952 , w2953 , w2954 , w2955 , w2956 , w2957 , w2958 , w2959 , w2960 , w2961 , w2962 , w2963 , w2964 , w2965 , w2966 , w2967 , w2968 , w2969 , w2970 , w2971 , w2972 , w2973 , w2974 , w2975 , w2976 , w2977 , w2978 , w2979 , w2980 , w2981 , w2982 , w2983 , w2984 , w2985 , w2986 , w2987 , w2988 , w2989 , w2990 , w2991 , w2992 , w2993 , w2994 , w2995 , w2996 , w2997 , w2998 , w2999 , w3000 , w3001 , w3002 , w3003 , w3004 , w3005 , w3006 , w3007 , w3008 , w3009 , w3010 , w3011 , w3012 , w3013 , w3014 , w3015 , w3016 , w3017 , w3018 , w3019 , w3020 , w3021 , w3022 , w3023 , w3024 , w3025 , w3026 , w3027 , w3028 , w3029 , w3030 , w3031 , w3032 , w3033 , w3034 , w3035 , w3036 , w3037 , w3038 , w3039 , w3040 , w3041 , w3042 , w3043 , w3044 , w3045 , w3046 , w3047 , w3048 , w3049 , w3050 , w3051 , w3052 , w3053 , w3054 , w3055 , w3056 , w3057 , w3058 , w3059 , w3060 , w3061 , w3062 , w3063 , w3064 , w3065 , w3066 , w3067 , w3068 , w3069 , w3070 , w3071 , w3072 , w3073 , w3074 , w3075 , w3076 , w3077 , w3078 , w3079 , w3080 , w3081 , w3082 , w3083 , w3084 , w3085 , w3086 , w3087 , w3088 , w3089 , w3090 , w3091 , w3092 , w3093 , w3094 , w3095 , w3096 , w3097 , w3098 , w3099 , w3100 , w3101 , w3102 , w3103 , w3104 , w3105 , w3106 , w3107 , w3108 , w3109 , w3110 , w3111 , w3112 , w3113 , w3114 , w3115 , w3116 , w3117 , w3118 , w3119 , w3120 , w3121 , w3122 , w3123 , w3124 , w3125 , w3126 , w3127 , w3128 , w3129 , w3130 , w3131 , w3132 , w3133 , w3134 , w3135 , w3136 , w3137 , w3138 , w3139 , w3140 , w3141 , w3142 , w3143 , w3144 , w3145 , w3146 , w3147 , w3148 , w3149 , w3150 , w3151 , w3152 , w3153 , w3154 , w3155 , w3156 , w3157 , w3158 , w3159 , w3160 , w3161 , w3162 , w3163 , w3164 , w3165 , w3166 , w3167 , w3168 , w3169 , w3170 , w3171 , w3172 , w3173 , w3174 , w3175 , w3176 , w3177 , w3178 , w3179 , w3180 , w3181 , w3182 , w3183 , w3184 , w3185 , w3186 , w3187 , w3188 , w3189 , w3190 , w3191 , w3192 , w3193 , w3194 , w3195 , w3196 , w3197 , w3198 , w3199 , w3200 , w3201 , w3202 , w3203 , w3204 , w3205 , w3206 , w3207 , w3208 , w3209 , w3210 , w3211 , w3212 , w3213 , w3214 , w3215 , w3216 , w3217 , w3218 , w3219 , w3220 , w3221 , w3222 , w3223 , w3224 , w3225 , w3226 , w3227 , w3228 , w3229 , w3230 , w3231 , w3232 , w3233 , w3234 , w3235 , w3236 , w3237 , w3238 , w3239 , w3240 , w3241 , w3242 , w3243 , w3244 , w3245 , w3246 , w3247 , w3248 , w3249 , w3250 , w3251 , w3252 , w3253 , w3254 , w3255 , w3256 , w3257 , w3258 , w3259 , w3260 , w3261 , w3262 , w3263 , w3264 , w3265 , w3266 , w3267 , w3268 , w3269 , w3270 , w3271 , w3272 , w3273 , w3274 , w3275 , w3276 , w3277 , w3278 , w3279 , w3280 , w3281 , w3282 , w3283 , w3284 , w3285 , w3286 , w3287 , w3288 , w3289 , w3290 , w3291 , w3292 , w3293 , w3294 , w3295 , w3296 , w3297 , w3298 , w3299 , w3300 , w3301 , w3302 , w3303 , w3304 , w3305 , w3306 , w3307 , w3308 , w3309 , w3310 , w3311 , w3312 , w3313 , w3314 , w3315 , w3316 , w3317 , w3318 , w3319 , w3320 , w3321 , w3322 , w3323 , w3324 , w3325 , w3326 , w3327 , w3328 , w3329 , w3330 , w3331 , w3332 , w3333 , w3334 , w3335 , w3336 , w3337 , w3338 , w3339 , w3340 , w3341 , w3342 , w3343 , w3344 , w3345 , w3346 , w3347 , w3348 , w3349 , w3350 , w3351 , w3352 , w3353 , w3354 , w3355 , w3356 , w3357 , w3358 , w3359 , w3360 , w3361 , w3362 , w3363 , w3364 , w3365 , w3366 , w3367 , w3368 , w3369 , w3370 , w3371 , w3372 , w3373 , w3374 , w3375 , w3376 , w3377 , w3378 , w3379 , w3380 , w3381 , w3382 , w3383 , w3384 , w3385 , w3386 , w3387 , w3388 , w3389 , w3390 , w3391 , w3392 , w3393 , w3394 , w3395 , w3396 , w3397 , w3398 , w3399 , w3400 , w3401 , w3402 , w3403 , w3404 , w3405 , w3406 , w3407 , w3408 , w3409 , w3410 , w3411 , w3412 , w3413 , w3414 , w3415 , w3416 , w3417 , w3418 , w3419 , w3420 , w3421 , w3422 , w3423 , w3424 , w3425 , w3426 , w3427 , w3428 , w3429 , w3430 , w3431 , w3432 , w3433 , w3434 , w3435 , w3436 , w3437 , w3438 , w3439 , w3440 , w3441 , w3442 , w3443 , w3444 , w3445 , w3446 , w3447 , w3448 , w3449 , w3450 , w3451 , w3452 , w3453 , w3454 , w3455 , w3456 , w3457 , w3458 , w3459 , w3460 , w3461 , w3462 , w3463 , w3464 , w3465 , w3466 , w3467 , w3468 , w3469 , w3470 , w3471 , w3472 , w3473 , w3474 , w3475 , w3476 , w3477 , w3478 , w3479 , w3480 , w3481 , w3482 , w3483 , w3484 , w3485 , w3486 , w3487 , w3488 , w3489 , w3490 , w3491 , w3492 , w3493 , w3494 , w3495 , w3496 , w3497 , w3498 , w3499 , w3500 , w3501 , w3502 , w3503 , w3504 , w3505 , w3506 , w3507 , w3508 , w3509 , w3510 , w3511 , w3512 , w3513 , w3514 , w3515 , w3516 , w3517 , w3518 , w3519 , w3520 , w3521 , w3522 , w3523 , w3524 , w3525 , w3526 , w3527 , w3528 , w3529 , w3530 , w3531 , w3532 , w3533 , w3534 , w3535 , w3536 , w3537 , w3538 , w3539 , w3540 , w3541 , w3542 , w3543 , w3544 , w3545 , w3546 , w3547 , w3548 , w3549 , w3550 , w3551 , w3552 , w3553 , w3554 , w3555 , w3556 , w3557 , w3558 , w3559 , w3560 , w3561 , w3562 , w3563 , w3564 , w3565 , w3566 , w3567 , w3568 , w3569 , w3570 , w3571 , w3572 , w3573 , w3574 , w3575 , w3576 , w3577 , w3578 , w3579 , w3580 , w3581 , w3582 , w3583 , w3584 , w3585 , w3586 , w3587 , w3588 , w3589 , w3590 , w3591 , w3592 , w3593 , w3594 , w3595 , w3596 , w3597 , w3598 , w3599 , w3600 , w3601 , w3602 , w3603 , w3604 , w3605 , w3606 , w3607 , w3608 , w3609 , w3610 , w3611 , w3612 , w3613 , w3614 , w3615 , w3616 , w3617 , w3618 , w3619 , w3620 , w3621 , w3622 , w3623 , w3624 , w3625 , w3626 , w3627 , w3628 , w3629 , w3630 , w3631 , w3632 , w3633 , w3634 , w3635 , w3636 , w3637 , w3638 , w3639 , w3640 , w3641 , w3642 , w3643 , w3644 , w3645 , w3646 , w3647 , w3648 , w3649 , w3650 , w3651 , w3652 , w3653 , w3654 , w3655 , w3656 , w3657 , w3658 , w3659 , w3660 , w3661 , w3662 , w3663 , w3664 , w3665 , w3666 , w3667 , w3668 , w3669 , w3670 , w3671 , w3672 , w3673 , w3674 , w3675 , w3676 , w3677 , w3678 , w3679 , w3680 , w3681 , w3682 , w3683 , w3684 , w3685 , w3686 , w3687 , w3688 , w3689 , w3690 , w3691 , w3692 , w3693 , w3694 , w3695 , w3696 , w3697 , w3698 , w3699 , w3700 , w3701 , w3702 , w3703 , w3704 , w3705 , w3706 , w3707 , w3708 , w3709 , w3710 , w3711 , w3712 , w3713 , w3714 , w3715 , w3716 , w3717 , w3718 , w3719 , w3720 , w3721 , w3722 , w3723 , w3724 , w3725 , w3726 , w3727 , w3728 , w3729 , w3730 , w3731 , w3732 , w3733 , w3734 , w3735 , w3736 , w3737 , w3738 , w3739 , w3740 , w3741 , w3742 , w3743 , w3744 , w3745 , w3746 , w3747 , w3748 , w3749 , w3750 , w3751 , w3752 , w3753 , w3754 , w3755 , w3756 , w3757 , w3758 , w3759 , w3760 , w3761 , w3762 , w3763 , w3764 , w3765 , w3766 , w3767 , w3768 , w3769 , w3770 , w3771 , w3772 , w3773 , w3774 , w3775 , w3776 , w3777 , w3778 , w3779 , w3780 , w3781 , w3782 , w3783 , w3784 , w3785 , w3786 , w3787 , w3788 , w3789 , w3790 , w3791 , w3792 , w3793 , w3794 , w3795 , w3796 , w3797 , w3798 , w3799 , w3800 , w3801 , w3802 , w3803 , w3804 , w3805 , w3806 , w3807 , w3808 , w3809 , w3810 , w3811 , w3812 , w3813 , w3814 , w3815 , w3816 , w3817 , w3818 , w3819 , w3820 , w3821 , w3822 , w3823 , w3824 , w3825 , w3826 , w3827 , w3828 , w3829 , w3830 , w3831 , w3832 , w3833 , w3834 , w3835 , w3836 , w3837 , w3838 , w3839 , w3840 , w3841 , w3842 , w3843 , w3844 , w3845 , w3846 , w3847 , w3848 , w3849 , w3850 , w3851 , w3852 , w3853 , w3854 , w3855 , w3856 , w3857 , w3858 , w3859 , w3860 , w3861 , w3862 , w3863 , w3864 , w3865 , w3866 , w3867 , w3868 , w3869 , w3870 , w3871 , w3872 , w3873 , w3874 , w3875 , w3876 , w3877 , w3878 , w3879 , w3880 , w3881 , w3882 , w3883 , w3884 , w3885 , w3886 , w3887 , w3888 , w3889 , w3890 , w3891 , w3892 , w3893 , w3894 , w3895 , w3896 , w3897 , w3898 , w3899 , w3900 , w3901 , w3902 , w3903 , w3904 , w3905 , w3906 , w3907 , w3908 , w3909 , w3910 , w3911 , w3912 , w3913 , w3914 , w3915 , w3916 , w3917 , w3918 , w3919 , w3920 , w3921 , w3922 , w3923 , w3924 , w3925 , w3926 , w3927 , w3928 , w3929 , w3930 , w3931 , w3932 , w3933 , w3934 , w3935 , w3936 , w3937 , w3938 , w3939 , w3940 , w3941 , w3942 , w3943 , w3944 , w3945 , w3946 , w3947 , w3948 , w3949 , w3950 , w3951 , w3952 , w3953 , w3954 , w3955 , w3956 , w3957 , w3958 , w3959 , w3960 , w3961 , w3962 , w3963 , w3964 , w3965 , w3966 , w3967 , w3968 , w3969 , w3970 , w3971 , w3972 , w3973 , w3974 , w3975 , w3976 , w3977 , w3978 , w3979 , w3980 , w3981 , w3982 , w3983 , w3984 , w3985 , w3986 , w3987 , w3988 , w3989 , w3990 , w3991 , w3992 , w3993 , w3994 , w3995 , w3996 , w3997 , w3998 , w3999 , w4000 , w4001 , w4002 , w4003 , w4004 , w4005 , w4006 , w4007 , w4008 , w4009 , w4010 , w4011 , w4012 , w4013 , w4014 , w4015 , w4016 , w4017 , w4018 , w4019 , w4020 , w4021 , w4022 , w4023 , w4024 , w4025 , w4026 , w4027 , w4028 , w4029 , w4030 , w4031 , w4032 , w4033 , w4034 , w4035 , w4036 , w4037 , w4038 , w4039 , w4040 , w4041 , w4042 , w4043 , w4044 , w4045 , w4046 , w4047 , w4048 , w4049 , w4050 , w4051 , w4052 , w4053 , w4054 , w4055 , w4056 , w4057 , w4058 , w4059 , w4060 , w4061 , w4062 , w4063 , w4064 , w4065 , w4066 , w4067 , w4068 , w4069 , w4070 , w4071 , w4072 , w4073 , w4074 , w4075 , w4076 , w4077 , w4078 , w4079 , w4080 , w4081 , w4082 , w4083 , w4084 , w4085 , w4086 , w4087 , w4088 , w4089 , w4090 , w4091 , w4092 , w4093 , w4094 , w4095 , w4096 , w4097 , w4098 , w4099 , w4100 , w4101 , w4102 , w4103 , w4104 , w4105 , w4106 , w4107 , w4108 , w4109 , w4110 , w4111 , w4112 , w4113 , w4114 , w4115 , w4116 , w4117 , w4118 , w4119 , w4120 , w4121 , w4122 , w4123 , w4124 , w4125 , w4126 , w4127 , w4128 , w4129 , w4130 , w4131 , w4132 , w4133 , w4134 , w4135 , w4136 , w4137 , w4138 , w4139 , w4140 , w4141 , w4142 , w4143 , w4144 , w4145 , w4146 , w4147 , w4148 , w4149 , w4150 , w4151 , w4152 , w4153 , w4154 , w4155 , w4156 , w4157 , w4158 , w4159 , w4160 , w4161 , w4162 , w4163 , w4164 , w4165 , w4166 , w4167 , w4168 , w4169 , w4170 , w4171 , w4172 , w4173 , w4174 , w4175 , w4176 , w4177 , w4178 , w4179 , w4180 , w4181 , w4182 , w4183 , w4184 , w4185 , w4186 , w4187 , w4188 , w4189 , w4190 , w4191 , w4192 , w4193 , w4194 , w4195 , w4196 , w4197 , w4198 , w4199 , w4200 , w4201 , w4202 , w4203 , w4204 , w4205 , w4206 , w4207 , w4208 , w4209 , w4210 , w4211 , w4212 , w4213 , w4214 , w4215 , w4216 , w4217 , w4218 , w4219 , w4220 , w4221 , w4222 , w4223 , w4224 , w4225 , w4226 , w4227 , w4228 , w4229 , w4230 , w4231 , w4232 , w4233 , w4234 , w4235 , w4236 , w4237 , w4238 , w4239 , w4240 , w4241 , w4242 , w4243 , w4244 , w4245 , w4246 , w4247 , w4248 , w4249 , w4250 , w4251 , w4252 , w4253 , w4254 , w4255 , w4256 , w4257 , w4258 , w4259 , w4260 , w4261 , w4262 , w4263 , w4264 , w4265 , w4266 , w4267 , w4268 , w4269 , w4270 , w4271 , w4272 , w4273 , w4274 , w4275 , w4276 , w4277 , w4278 , w4279 , w4280 , w4281 , w4282 , w4283 , w4284 , w4285 , w4286 , w4287 , w4288 , w4289 , w4290 , w4291 , w4292 , w4293 , w4294 , w4295 , w4296 , w4297 , w4298 , w4299 , w4300 , w4301 , w4302 , w4303 , w4304 , w4305 , w4306 , w4307 , w4308 , w4309 , w4310 , w4311 , w4312 , w4313 , w4314 , w4315 , w4316 , w4317 , w4318 , w4319 , w4320 , w4321 , w4322 , w4323 , w4324 , w4325 , w4326 , w4327 , w4328 , w4329 , w4330 , w4331 , w4332 , w4333 , w4334 , w4335 , w4336 , w4337 , w4338 , w4339 , w4340 , w4341 , w4342 , w4343 , w4344 , w4345 , w4346 , w4347 , w4348 , w4349 , w4350 , w4351 , w4352 , w4353 , w4354 , w4355 , w4356 , w4357 , w4358 , w4359 , w4360 , w4361 , w4362 , w4363 , w4364 , w4365 , w4366 , w4367 , w4368 , w4369 , w4370 , w4371 , w4372 , w4373 , w4374 , w4375 , w4376 , w4377 , w4378 , w4379 , w4380 , w4381 , w4382 , w4383 , w4384 , w4385 , w4386 , w4387 , w4388 , w4389 , w4390 , w4391 , w4392 , w4393 , w4394 , w4395 , w4396 , w4397 , w4398 , w4399 , w4400 , w4401 , w4402 , w4403 , w4404 , w4405 , w4406 , w4407 , w4408 , w4409 , w4410 , w4411 , w4412 , w4413 , w4414 , w4415 , w4416 , w4417 , w4418 , w4419 , w4420 , w4421 , w4422 , w4423 , w4424 , w4425 , w4426 , w4427 , w4428 , w4429 , w4430 , w4431 , w4432 , w4433 , w4434 , w4435 , w4436 , w4437 , w4438 , w4439 , w4440 , w4441 , w4442 , w4443 , w4444 , w4445 , w4446 , w4447 , w4448 , w4449 , w4450 , w4451 , w4452 , w4453 , w4454 , w4455 , w4456 , w4457 , w4458 , w4459 , w4460 , w4461 , w4462 , w4463 , w4464 , w4465 , w4466 , w4467 , w4468 , w4469 , w4470 , w4471 , w4472 , w4473 , w4474 , w4475 , w4476 , w4477 , w4478 , w4479 , w4480 , w4481 , w4482 , w4483 , w4484 , w4485 , w4486 , w4487 , w4488 , w4489 , w4490 , w4491 , w4492 , w4493 , w4494 , w4495 , w4496 , w4497 , w4498 , w4499 , w4500 , w4501 , w4502 , w4503 , w4504 , w4505 , w4506 , w4507 , w4508 , w4509 , w4510 , w4511 , w4512 , w4513 , w4514 , w4515 , w4516 , w4517 , w4518 , w4519 , w4520 , w4521 , w4522 , w4523 , w4524 , w4525 , w4526 , w4527 , w4528 , w4529 , w4530 , w4531 , w4532 , w4533 , w4534 , w4535 , w4536 , w4537 , w4538 , w4539 , w4540 , w4541 , w4542 , w4543 , w4544 , w4545 , w4546 , w4547 , w4548 , w4549 , w4550 , w4551 , w4552 , w4553 , w4554 , w4555 , w4556 , w4557 , w4558 , w4559 , w4560 , w4561 , w4562 , w4563 , w4564 , w4565 , w4566 , w4567 , w4568 , w4569 , w4570 , w4571 , w4572 , w4573 , w4574 , w4575 , w4576 , w4577 , w4578 , w4579 , w4580 , w4581 , w4582 , w4583 , w4584 , w4585 , w4586 , w4587 , w4588 , w4589 , w4590 , w4591 , w4592 , w4593 , w4594 , w4595 , w4596 , w4597 , w4598 , w4599 , w4600 , w4601 , w4602 , w4603 , w4604 , w4605 , w4606 , w4607 , w4608 , w4609 , w4610 , w4611 , w4612 , w4613 , w4614 , w4615 , w4616 , w4617 , w4618 , w4619 , w4620 , w4621 , w4622 , w4623 , w4624 , w4625 , w4626 , w4627 , w4628 , w4629 , w4630 , w4631 , w4632 , w4633 , w4634 , w4635 , w4636 , w4637 , w4638 , w4639 , w4640 , w4641 , w4642 , w4643 , w4644 , w4645 , w4646 , w4647 , w4648 , w4649 , w4650 , w4651 , w4652 , w4653 , w4654 , w4655 , w4656 , w4657 , w4658 , w4659 , w4660 , w4661 , w4662 , w4663 , w4664 , w4665 , w4666 , w4667 , w4668 , w4669 , w4670 , w4671 , w4672 , w4673 , w4674 , w4675 , w4676 , w4677 , w4678 , w4679 , w4680 , w4681 , w4682 , w4683 , w4684 , w4685 , w4686 , w4687 , w4688 , w4689 , w4690 , w4691 , w4692 , w4693 , w4694 , w4695 , w4696 , w4697 , w4698 , w4699 , w4700 , w4701 , w4702 , w4703 , w4704 , w4705 , w4706 , w4707 , w4708 , w4709 , w4710 , w4711 , w4712 , w4713 , w4714 , w4715 , w4716 , w4717 , w4718 , w4719 , w4720 , w4721 , w4722 , w4723 , w4724 , w4725 , w4726 , w4727 , w4728 , w4729 , w4730 , w4731 , w4732 , w4733 , w4734 , w4735 , w4736 , w4737 , w4738 , w4739 , w4740 , w4741 , w4742 , w4743 , w4744 , w4745 , w4746 , w4747 , w4748 , w4749 , w4750 , w4751 , w4752 , w4753 , w4754 , w4755 , w4756 , w4757 , w4758 , w4759 , w4760 , w4761 , w4762 , w4763 , w4764 , w4765 , w4766 , w4767 , w4768 , w4769 , w4770 , w4771 , w4772 , w4773 , w4774 , w4775 , w4776 , w4777 , w4778 , w4779 , w4780 , w4781 , w4782 , w4783 , w4784 , w4785 , w4786 , w4787 , w4788 , w4789 , w4790 , w4791 , w4792 , w4793 , w4794 , w4795 , w4796 , w4797 , w4798 , w4799 , w4800 , w4801 , w4802 , w4803 , w4804 , w4805 , w4806 , w4807 , w4808 , w4809 , w4810 , w4811 , w4812 , w4813 , w4814 , w4815 , w4816 , w4817 , w4818 , w4819 , w4820 , w4821 , w4822 , w4823 , w4824 , w4825 , w4826 , w4827 , w4828 , w4829 , w4830 , w4831 , w4832 , w4833 , w4834 , w4835 , w4836 , w4837 , w4838 , w4839 , w4840 , w4841 , w4842 , w4843 , w4844 , w4845 , w4846 , w4847 , w4848 , w4849 , w4850 , w4851 , w4852 , w4853 , w4854 , w4855 , w4856 , w4857 , w4858 , w4859 , w4860 , w4861 , w4862 , w4863 , w4864 , w4865 , w4866 , w4867 , w4868 , w4869 , w4870 , w4871 , w4872 , w4873 , w4874 , w4875 , w4876 , w4877 , w4878 , w4879 , w4880 , w4881 , w4882 , w4883 , w4884 , w4885 , w4886 , w4887 , w4888 , w4889 , w4890 , w4891 , w4892 , w4893 , w4894 , w4895 , w4896 , w4897 , w4898 , w4899 , w4900 , w4901 , w4902 , w4903 , w4904 , w4905 , w4906 , w4907 , w4908 , w4909 , w4910 , w4911 , w4912 , w4913 , w4914 , w4915 , w4916 , w4917 , w4918 , w4919 , w4920 , w4921 , w4922 , w4923 , w4924 , w4925 , w4926 , w4927 , w4928 , w4929 , w4930 , w4931 , w4932 , w4933 , w4934 , w4935 , w4936 , w4937 , w4938 , w4939 , w4940 , w4941 , w4942 , w4943 , w4944 , w4945 , w4946 , w4947 , w4948 , w4949 , w4950 , w4951 , w4952 , w4953 , w4954 , w4955 , w4956 , w4957 , w4958 , w4959 , w4960 , w4961 , w4962 , w4963 , w4964 , w4965 , w4966 , w4967 , w4968 , w4969 , w4970 , w4971 , w4972 , w4973 , w4974 , w4975 , w4976 , w4977 , w4978 , w4979 , w4980 , w4981 , w4982 , w4983 , w4984 , w4985 , w4986 , w4987 , w4988 , w4989 , w4990 , w4991 , w4992 , w4993 , w4994 , w4995 , w4996 , w4997 , w4998 , w4999 , w5000 , w5001 , w5002 , w5003 , w5004 , w5005 , w5006 , w5007 , w5008 , w5009 , w5010 , w5011 , w5012 , w5013 , w5014 , w5015 , w5016 , w5017 , w5018 , w5019 , w5020 , w5021 , w5022 , w5023 , w5024 , w5025 , w5026 , w5027 , w5028 , w5029 , w5030 , w5031 , w5032 , w5033 , w5034 , w5035 , w5036 , w5037 , w5038 , w5039 , w5040 , w5041 , w5042 , w5043 , w5044 , w5045 , w5046 , w5047 , w5048 , w5049 , w5050 , w5051 , w5052 , w5053 , w5054 , w5055 , w5056 , w5057 , w5058 , w5059 , w5060 , w5061 , w5062 , w5063 , w5064 , w5065 , w5066 , w5067 , w5068 , w5069 , w5070 , w5071 , w5072 , w5073 , w5074 , w5075 , w5076 , w5077 , w5078 , w5079 , w5080 , w5081 , w5082 , w5083 , w5084 , w5085 , w5086 , w5087 , w5088 , w5089 , w5090 , w5091 , w5092 , w5093 , w5094 , w5095 , w5096 , w5097 , w5098 , w5099 , w5100 , w5101 , w5102 , w5103 , w5104 , w5105 , w5106 , w5107 , w5108 , w5109 , w5110 , w5111 , w5112 , w5113 , w5114 , w5115 , w5116 , w5117 , w5118 , w5119 , w5120 , w5121 , w5122 , w5123 , w5124 , w5125 , w5126 , w5127 , w5128 , w5129 , w5130 , w5131 , w5132 , w5133 , w5134 , w5135 , w5136 , w5137 , w5138 , w5139 , w5140 , w5141 , w5142 , w5143 , w5144 , w5145 , w5146 , w5147 , w5148 , w5149 , w5150 , w5151 , w5152 , w5153 , w5154 , w5155 , w5156 , w5157 , w5158 , w5159 , w5160 , w5161 , w5162 , w5163 , w5164 , w5165 , w5166 , w5167 , w5168 , w5169 , w5170 , w5171 , w5172 , w5173 , w5174 , w5175 , w5176 , w5177 , w5178 , w5179 , w5180 , w5181 , w5182 , w5183 , w5184 , w5185 , w5186 , w5187 , w5188 , w5189 , w5190 , w5191 , w5192 , w5193 , w5194 , w5195 , w5196 , w5197 , w5198 , w5199 , w5200 , w5201 , w5202 , w5203 , w5204 , w5205 , w5206 , w5207 , w5208 , w5209 , w5210 , w5211 , w5212 , w5213 , w5214 , w5215 , w5216 , w5217 , w5218 , w5219 , w5220 , w5221 , w5222 , w5223 , w5224 , w5225 , w5226 , w5227 , w5228 , w5229 , w5230 , w5231 , w5232 , w5233 , w5234 , w5235 , w5236 , w5237 , w5238 , w5239 , w5240 , w5241 , w5242 , w5243 , w5244 , w5245 , w5246 , w5247 , w5248 , w5249 , w5250 , w5251 , w5252 , w5253 , w5254 , w5255 , w5256 , w5257 , w5258 , w5259 , w5260 , w5261 , w5262 , w5263 , w5264 , w5265 , w5266 , w5267 , w5268 , w5269 , w5270 , w5271 , w5272 , w5273 , w5274 , w5275 , w5276 , w5277 , w5278 , w5279 , w5280 , w5281 , w5282 , w5283 , w5284 , w5285 , w5286 , w5287 , w5288 , w5289 , w5290 , w5291 , w5292 , w5293 , w5294 , w5295 , w5296 , w5297 , w5298 , w5299 , w5300 , w5301 , w5302 , w5303 , w5304 , w5305 , w5306 , w5307 , w5308 , w5309 , w5310 , w5311 , w5312 , w5313 , w5314 , w5315 , w5316 , w5317 , w5318 , w5319 , w5320 , w5321 , w5322 , w5323 , w5324 , w5325 , w5326 , w5327 , w5328 , w5329 , w5330 , w5331 , w5332 , w5333 , w5334 , w5335 , w5336 , w5337 , w5338 , w5339 , w5340 , w5341 , w5342 , w5343 , w5344 , w5345 , w5346 , w5347 , w5348 , w5349 , w5350 , w5351 , w5352 , w5353 , w5354 , w5355 , w5356 , w5357 , w5358 , w5359 , w5360 , w5361 , w5362 , w5363 , w5364 , w5365 , w5366 , w5367 , w5368 , w5369 , w5370 , w5371 , w5372 , w5373 , w5374 , w5375 , w5376 , w5377 , w5378 , w5379 , w5380 , w5381 , w5382 , w5383 , w5384 , w5385 , w5386 , w5387 , w5388 , w5389 , w5390 , w5391 , w5392 , w5393 , w5394 , w5395 , w5396 , w5397 , w5398 , w5399 , w5400 , w5401 , w5402 , w5403 , w5404 , w5405 , w5406 , w5407 , w5408 , w5409 , w5410 , w5411 , w5412 , w5413 , w5414 , w5415 , w5416 , w5417 , w5418 , w5419 , w5420 , w5421 , w5422 , w5423 , w5424 , w5425 , w5426 , w5427 , w5428 , w5429 , w5430 , w5431 , w5432 , w5433 , w5434 , w5435 , w5436 , w5437 , w5438 , w5439 , w5440 , w5441 , w5442 , w5443 , w5444 , w5445 , w5446 , w5447 , w5448 , w5449 , w5450 , w5451 , w5452 , w5453 , w5454 , w5455 , w5456 , w5457 , w5458 , w5459 , w5460 , w5461 , w5462 , w5463 , w5464 , w5465 , w5466 , w5467 , w5468 , w5469 , w5470 , w5471 , w5472 , w5473 , w5474 , w5475 , w5476 , w5477 , w5478 , w5479 , w5480 , w5481 , w5482 , w5483 , w5484 , w5485 , w5486 , w5487 , w5488 , w5489 , w5490 , w5491 , w5492 , w5493 , w5494 , w5495 , w5496 , w5497 , w5498 , w5499 , w5500 , w5501 , w5502 , w5503 , w5504 , w5505 , w5506 , w5507 , w5508 , w5509 , w5510 , w5511 , w5512 , w5513 , w5514 , w5515 , w5516 , w5517 , w5518 , w5519 , w5520 , w5521 , w5522 , w5523 , w5524 , w5525 , w5526 , w5527 , w5528 , w5529 , w5530 , w5531 , w5532 , w5533 , w5534 , w5535 , w5536 , w5537 , w5538 , w5539 , w5540 , w5541 , w5542 , w5543 , w5544 , w5545 , w5546 , w5547 , w5548 , w5549 , w5550 , w5551 , w5552 , w5553 , w5554 , w5555 , w5556 , w5557 , w5558 , w5559 , w5560 , w5561 , w5562 , w5563 , w5564 , w5565 , w5566 , w5567 , w5568 , w5569 , w5570 , w5571 , w5572 , w5573 , w5574 , w5575 , w5576 , w5577 , w5578 , w5579 , w5580 , w5581 , w5582 , w5583 , w5584 , w5585 , w5586 , w5587 , w5588 , w5589 , w5590 , w5591 , w5592 , w5593 , w5594 , w5595 , w5596 , w5597 , w5598 , w5599 , w5600 , w5601 , w5602 , w5603 , w5604 , w5605 , w5606 , w5607 , w5608 , w5609 , w5610 , w5611 , w5612 , w5613 , w5614 , w5615 , w5616 , w5617 , w5618 , w5619 , w5620 , w5621 , w5622 , w5623 , w5624 , w5625 , w5626 , w5627 , w5628 , w5629 , w5630 , w5631 , w5632 , w5633 , w5634 , w5635 , w5636 , w5637 , w5638 , w5639 , w5640 , w5641 , w5642 , w5643 , w5644 , w5645 , w5646 , w5647 , w5648 , w5649 , w5650 , w5651 , w5652 , w5653 , w5654 , w5655 , w5656 , w5657 , w5658 , w5659 , w5660 , w5661 , w5662 , w5663 , w5664 , w5665 , w5666 , w5667 , w5668 , w5669 , w5670 , w5671 , w5672 , w5673 , w5674 , w5675 , w5676 , w5677 , w5678 , w5679 , w5680 , w5681 , w5682 , w5683 , w5684 , w5685 , w5686 , w5687 , w5688 , w5689 , w5690 , w5691 , w5692 , w5693 , w5694 , w5695 , w5696 , w5697 , w5698 , w5699 , w5700 , w5701 , w5702 , w5703 , w5704 , w5705 , w5706 , w5707 , w5708 , w5709 , w5710 , w5711 , w5712 , w5713 , w5714 , w5715 , w5716 , w5717 , w5718 , w5719 , w5720 , w5721 , w5722 , w5723 , w5724 , w5725 , w5726 , w5727 , w5728 , w5729 , w5730 , w5731 , w5732 , w5733 , w5734 , w5735 , w5736 , w5737 , w5738 , w5739 , w5740 , w5741 , w5742 , w5743 , w5744 , w5745 , w5746 , w5747 , w5748 , w5749 , w5750 , w5751 , w5752 , w5753 , w5754 , w5755 , w5756 , w5757 , w5758 , w5759 , w5760 , w5761 , w5762 , w5763 , w5764 , w5765 , w5766 , w5767 , w5768 , w5769 , w5770 , w5771 , w5772 , w5773 , w5774 , w5775 , w5776 , w5777 , w5778 , w5779 , w5780 , w5781 , w5782 , w5783 , w5784 , w5785 , w5786 , w5787 , w5788 , w5789 , w5790 , w5791 , w5792 , w5793 , w5794 , w5795 , w5796 , w5797 , w5798 , w5799 , w5800 , w5801 , w5802 , w5803 , w5804 , w5805 , w5806 , w5807 , w5808 , w5809 , w5810 , w5811 , w5812 , w5813 , w5814 , w5815 , w5816 , w5817 , w5818 , w5819 , w5820 , w5821 , w5822 , w5823 , w5824 , w5825 , w5826 , w5827 , w5828 , w5829 , w5830 , w5831 , w5832 , w5833 , w5834 , w5835 , w5836 , w5837 , w5838 , w5839 , w5840 , w5841 , w5842 , w5843 , w5844 , w5845 , w5846 , w5847 , w5848 , w5849 , w5850 , w5851 , w5852 , w5853 , w5854 , w5855 , w5856 , w5857 , w5858 , w5859 , w5860 , w5861 , w5862 , w5863 , w5864 , w5865 , w5866 , w5867 , w5868 , w5869 , w5870 , w5871 , w5872 , w5873 , w5874 , w5875 , w5876 , w5877 , w5878 , w5879 , w5880 , w5881 , w5882 , w5883 , w5884 , w5885 , w5886 , w5887 , w5888 , w5889 , w5890 , w5891 , w5892 , w5893 , w5894 , w5895 , w5896 , w5897 , w5898 , w5899 , w5900 , w5901 , w5902 , w5903 , w5904 , w5905 , w5906 , w5907 , w5908 , w5909 , w5910 , w5911 , w5912 , w5913 , w5914 , w5915 , w5916 , w5917 , w5918 , w5919 , w5920 , w5921 , w5922 , w5923 , w5924 , w5925 , w5926 , w5927 , w5928 , w5929 , w5930 , w5931 , w5932 , w5933 , w5934 , w5935 , w5936 , w5937 , w5938 , w5939 , w5940 , w5941 , w5942 , w5943 , w5944 , w5945 , w5946 , w5947 , w5948 , w5949 , w5950 , w5951 , w5952 , w5953 , w5954 , w5955 , w5956 , w5957 , w5958 , w5959 , w5960 , w5961 , w5962 , w5963 , w5964 , w5965 , w5966 , w5967 , w5968 , w5969 , w5970 , w5971 , w5972 , w5973 , w5974 , w5975 , w5976 , w5977 , w5978 , w5979 , w5980 , w5981 , w5982 , w5983 , w5984 , w5985 , w5986 , w5987 , w5988 , w5989 , w5990 , w5991 , w5992 , w5993 , w5994 , w5995 , w5996 , w5997 , w5998 , w5999 , w6000 , w6001 , w6002 , w6003 , w6004 , w6005 , w6006 , w6007 , w6008 , w6009 , w6010 , w6011 , w6012 , w6013 , w6014 , w6015 , w6016 , w6017 , w6018 , w6019 , w6020 , w6021 , w6022 , w6023 , w6024 , w6025 , w6026 , w6027 , w6028 , w6029 , w6030 , w6031 , w6032 , w6033 , w6034 , w6035 , w6036 , w6037 , w6038 , w6039 , w6040 , w6041 , w6042 , w6043 , w6044 , w6045 , w6046 , w6047 , w6048 , w6049 , w6050 , w6051 , w6052 , w6053 , w6054 , w6055 , w6056 , w6057 , w6058 , w6059 , w6060 , w6061 , w6062 , w6063 , w6064 , w6065 , w6066 , w6067 , w6068 , w6069 , w6070 , w6071 , w6072 , w6073 , w6074 , w6075 , w6076 , w6077 , w6078 , w6079 , w6080 , w6081 , w6082 , w6083 , w6084 , w6085 , w6086 , w6087 , w6088 , w6089 , w6090 , w6091 , w6092 , w6093 , w6094 , w6095 , w6096 , w6097 , w6098 , w6099 , w6100 , w6101 , w6102 , w6103 , w6104 , w6105 , w6106 , w6107 , w6108 , w6109 , w6110 , w6111 , w6112 , w6113 , w6114 , w6115 , w6116 , w6117 , w6118 , w6119 , w6120 , w6121 , w6122 , w6123 , w6124 , w6125 , w6126 , w6127 , w6128 , w6129 , w6130 , w6131 , w6132 , w6133 , w6134 , w6135 , w6136 , w6137 , w6138 , w6139 , w6140 , w6141 , w6142 , w6143 , w6144 , w6145 , w6146 , w6147 , w6148 , w6149 , w6150 , w6151 , w6152 , w6153 , w6154 , w6155 , w6156 , w6157 , w6158 , w6159 , w6160 , w6161 , w6162 , w6163 , w6164 , w6165 , w6166 , w6167 , w6168 , w6169 , w6170 , w6171 , w6172 , w6173 , w6174 , w6175 , w6176 , w6177 , w6178 , w6179 , w6180 , w6181 , w6182 , w6183 , w6184 , w6185 , w6186 , w6187 , w6188 , w6189 , w6190 , w6191 , w6192 , w6193 , w6194 , w6195 , w6196 , w6197 , w6198 , w6199 , w6200 , w6201 , w6202 , w6203 , w6204 , w6205 , w6206 , w6207 , w6208 , w6209 , w6210 , w6211 , w6212 , w6213 , w6214 , w6215 , w6216 , w6217 , w6218 , w6219 , w6220 , w6221 , w6222 , w6223 , w6224 , w6225 , w6226 , w6227 , w6228 , w6229 , w6230 , w6231 , w6232 , w6233 , w6234 , w6235 , w6236 , w6237 , w6238 , w6239 , w6240 , w6241 , w6242 , w6243 , w6244 , w6245 , w6246 , w6247 , w6248 , w6249 , w6250 , w6251 , w6252 , w6253 , w6254 , w6255 , w6256 , w6257 , w6258 , w6259 , w6260 , w6261 , w6262 , w6263 , w6264 , w6265 , w6266 , w6267 , w6268 , w6269 , w6270 , w6271 , w6272 , w6273 , w6274 , w6275 , w6276 , w6277 , w6278 , w6279 , w6280 , w6281 , w6282 , w6283 , w6284 , w6285 , w6286 , w6287 , w6288 , w6289 , w6290 , w6291 , w6292 , w6293 , w6294 , w6295 , w6296 , w6297 , w6298 , w6299 , w6300 , w6301 , w6302 , w6303 , w6304 , w6305 , w6306 , w6307 , w6308 , w6309 , w6310 , w6311 , w6312 , w6313 , w6314 , w6315 , w6316 , w6317 , w6318 , w6319 , w6320 , w6321 , w6322 , w6323 , w6324 , w6325 , w6326 , w6327 , w6328 , w6329 , w6330 , w6331 , w6332 , w6333 , w6334 , w6335 , w6336 , w6337 , w6338 , w6339 , w6340 , w6341 , w6342 , w6343 , w6344 , w6345 , w6346 , w6347 , w6348 , w6349 , w6350 , w6351 , w6352 , w6353 , w6354 , w6355 , w6356 , w6357 , w6358 , w6359 , w6360 , w6361 , w6362 , w6363 , w6364 , w6365 , w6366 , w6367 , w6368 , w6369 , w6370 , w6371 , w6372 , w6373 , w6374 , w6375 , w6376 , w6377 , w6378 , w6379 , w6380 , w6381 , w6382 , w6383 , w6384 , w6385 , w6386 , w6387 , w6388 , w6389 , w6390 , w6391 , w6392 , w6393 , w6394 , w6395 , w6396 , w6397 , w6398 , w6399 , w6400 , w6401 , w6402 , w6403 , w6404 , w6405 , w6406 , w6407 , w6408 , w6409 , w6410 , w6411 , w6412 , w6413 , w6414 , w6415 , w6416 , w6417 , w6418 , w6419 , w6420 , w6421 , w6422 , w6423 , w6424 , w6425 , w6426 , w6427 , w6428 , w6429 , w6430 , w6431 , w6432 , w6433 , w6434 , w6435 , w6436 , w6437 , w6438 , w6439 , w6440 , w6441 , w6442 , w6443 , w6444 , w6445 , w6446 , w6447 , w6448 , w6449 , w6450 , w6451 , w6452 , w6453 , w6454 , w6455 , w6456 , w6457 , w6458 , w6459 , w6460 , w6461 , w6462 , w6463 , w6464 , w6465 , w6466 , w6467 , w6468 , w6469 , w6470 , w6471 , w6472 , w6473 , w6474 , w6475 , w6476 , w6477 , w6478 , w6479 , w6480 , w6481 , w6482 , w6483 , w6484 , w6485 , w6486 , w6487 , w6488 , w6489 , w6490 , w6491 , w6492 , w6493 , w6494 , w6495 , w6496 , w6497 , w6498 , w6499 , w6500 , w6501 , w6502 , w6503 , w6504 , w6505 , w6506 , w6507 , w6508 , w6509 , w6510 , w6511 , w6512 , w6513 , w6514 , w6515 , w6516 , w6517 , w6518 , w6519 , w6520 , w6521 , w6522 , w6523 , w6524 , w6525 , w6526 , w6527 , w6528 , w6529 , w6530 , w6531 , w6532 , w6533 , w6534 , w6535 , w6536 , w6537 , w6538 , w6539 , w6540 , w6541 , w6542 , w6543 , w6544 , w6545 , w6546 , w6547 , w6548 , w6549 , w6550 , w6551 , w6552 , w6553 , w6554 , w6555 , w6556 , w6557 , w6558 , w6559 , w6560 , w6561 , w6562 , w6563 , w6564 , w6565 , w6566 , w6567 , w6568 , w6569 , w6570 , w6571 , w6572 , w6573 , w6574 , w6575 , w6576 , w6577 , w6578 , w6579 , w6580 , w6581 , w6582 , w6583 , w6584 , w6585 , w6586 , w6587 , w6588 , w6589 , w6590 , w6591 , w6592 , w6593 , w6594 , w6595 , w6596 , w6597 , w6598 , w6599 , w6600 , w6601 , w6602 , w6603 , w6604 , w6605 , w6606 , w6607 , w6608 , w6609 , w6610 , w6611 , w6612 , w6613 , w6614 , w6615 , w6616 , w6617 , w6618 , w6619 , w6620 , w6621 , w6622 , w6623 , w6624 , w6625 , w6626 , w6627 , w6628 , w6629 , w6630 , w6631 , w6632 , w6633 , w6634 , w6635 , w6636 , w6637 , w6638 , w6639 , w6640 , w6641 , w6642 , w6643 , w6644 , w6645 , w6646 , w6647 , w6648 , w6649 , w6650 , w6651 , w6652 , w6653 , w6654 , w6655 , w6656 , w6657 , w6658 , w6659 , w6660 , w6661 , w6662 , w6663 , w6664 , w6665 , w6666 , w6667 , w6668 , w6669 , w6670 , w6671 , w6672 , w6673 , w6674 , w6675 , w6676 , w6677 , w6678 , w6679 , w6680 , w6681 , w6682 , w6683 , w6684 , w6685 , w6686 , w6687 , w6688 , w6689 , w6690 , w6691 , w6692 , w6693 , w6694 , w6695 , w6696 , w6697 , w6698 , w6699 , w6700 , w6701 , w6702 , w6703 , w6704 , w6705 , w6706 , w6707 , w6708 , w6709 , w6710 , w6711 , w6712 , w6713 , w6714 , w6715 , w6716 , w6717 , w6718 , w6719 , w6720 , w6721 , w6722 , w6723 , w6724 , w6725 , w6726 , w6727 , w6728 , w6729 , w6730 , w6731 , w6732 , w6733 , w6734 , w6735 , w6736 , w6737 , w6738 , w6739 , w6740 , w6741 , w6742 , w6743 , w6744 , w6745 , w6746 , w6747 , w6748 , w6749 , w6750 , w6751 , w6752 , w6753 , w6754 , w6755 , w6756 , w6757 , w6758 , w6759 , w6760 , w6761 , w6762 , w6763 , w6764 , w6765 , w6766 , w6767 , w6768 , w6769 , w6770 , w6771 , w6772 , w6773 , w6774 , w6775 , w6776 , w6777 , w6778 , w6779 , w6780 , w6781 , w6782 , w6783 , w6784 , w6785 , w6786 , w6787 , w6788 , w6789 , w6790 , w6791 , w6792 , w6793 , w6794 , w6795 , w6796 , w6797 , w6798 , w6799 , w6800 , w6801 , w6802 , w6803 , w6804 , w6805 , w6806 , w6807 , w6808 , w6809 , w6810 , w6811 , w6812 , w6813 , w6814 , w6815 , w6816 , w6817 , w6818 , w6819 , w6820 , w6821 , w6822 , w6823 , w6824 , w6825 , w6826 , w6827 , w6828 , w6829 , w6830 , w6831 , w6832 , w6833 , w6834 , w6835 , w6836 , w6837 , w6838 , w6839 , w6840 , w6841 , w6842 , w6843 , w6844 , w6845 , w6846 , w6847 , w6848 , w6849 , w6850 , w6851 , w6852 , w6853 , w6854 , w6855 , w6856 , w6857 , w6858 , w6859 , w6860 , w6861 , w6862 , w6863 , w6864 , w6865 , w6866 , w6867 , w6868 , w6869 , w6870 , w6871 , w6872 , w6873 , w6874 , w6875 , w6876 , w6877 , w6878 , w6879 , w6880 , w6881 , w6882 , w6883 , w6884 , w6885 , w6886 , w6887 , w6888 , w6889 , w6890 , w6891 , w6892 , w6893 , w6894 , w6895 , w6896 , w6897 , w6898 , w6899 , w6900 , w6901 , w6902 , w6903 , w6904 , w6905 , w6906 , w6907 , w6908 , w6909 , w6910 , w6911 , w6912 , w6913 , w6914 , w6915 , w6916 , w6917 , w6918 , w6919 , w6920 , w6921 , w6922 , w6923 , w6924 , w6925 , w6926 , w6927 , w6928 , w6929 , w6930 , w6931 , w6932 , w6933 , w6934 , w6935 , w6936 , w6937 , w6938 , w6939 , w6940 , w6941 , w6942 , w6943 , w6944 , w6945 , w6946 , w6947 , w6948 , w6949 , w6950 , w6951 , w6952 , w6953 , w6954 , w6955 , w6956 , w6957 , w6958 , w6959 , w6960 , w6961 , w6962 , w6963 , w6964 , w6965 , w6966 , w6967 , w6968 , w6969 , w6970 , w6971 , w6972 , w6973 , w6974 , w6975 , w6976 , w6977 , w6978 , w6979 , w6980 , w6981 , w6982 , w6983 , w6984 , w6985 , w6986 , w6987 , w6988 , w6989 , w6990 , w6991 , w6992 , w6993 , w6994 , w6995 , w6996 , w6997 , w6998 , w6999 , w7000 , w7001 , w7002 , w7003 , w7004 , w7005 , w7006 , w7007 , w7008 , w7009 , w7010 , w7011 , w7012 , w7013 , w7014 , w7015 , w7016 , w7017 , w7018 , w7019 , w7020 , w7021 , w7022 , w7023 , w7024 , w7025 , w7026 , w7027 , w7028 , w7029 , w7030 , w7031 , w7032 , w7033 , w7034 , w7035 , w7036 , w7037 , w7038 , w7039 , w7040 , w7041 , w7042 , w7043 , w7044 , w7045 , w7046 , w7047 , w7048 , w7049 , w7050 , w7051 , w7052 , w7053 , w7054 , w7055 , w7056 , w7057 , w7058 , w7059 , w7060 , w7061 , w7062 , w7063 , w7064 , w7065 , w7066 , w7067 , w7068 , w7069 , w7070 , w7071 , w7072 , w7073 , w7074 , w7075 , w7076 , w7077 , w7078 , w7079 , w7080 , w7081 , w7082 , w7083 , w7084 , w7085 , w7086 , w7087 , w7088 , w7089 , w7090 , w7091 , w7092 , w7093 , w7094 , w7095 , w7096 , w7097 , w7098 , w7099 , w7100 , w7101 , w7102 , w7103 , w7104 , w7105 , w7106 , w7107 , w7108 , w7109 , w7110 , w7111 , w7112 , w7113 , w7114 , w7115 , w7116 , w7117 , w7118 , w7119 , w7120 , w7121 , w7122 , w7123 , w7124 , w7125 , w7126 , w7127 , w7128 , w7129 , w7130 , w7131 , w7132 , w7133 , w7134 , w7135 , w7136 , w7137 , w7138 , w7139 , w7140 , w7141 , w7142 , w7143 , w7144 , w7145 , w7146 , w7147 , w7148 , w7149 , w7150 , w7151 , w7152 , w7153 , w7154 , w7155 , w7156 , w7157 , w7158 , w7159 , w7160 , w7161 , w7162 , w7163 , w7164 , w7165 , w7166 , w7167 , w7168 , w7169 , w7170 , w7171 , w7172 , w7173 , w7174 , w7175 , w7176 , w7177 , w7178 , w7179 , w7180 , w7181 , w7182 , w7183 , w7184 , w7185 , w7186 , w7187 , w7188 , w7189 , w7190 , w7191 , w7192 , w7193 , w7194 , w7195 , w7196 , w7197 , w7198 , w7199 , w7200 , w7201 , w7202 , w7203 , w7204 , w7205 , w7206 , w7207 , w7208 , w7209 , w7210 , w7211 , w7212 , w7213 , w7214 , w7215 , w7216 , w7217 , w7218 , w7219 , w7220 , w7221 , w7222 , w7223 , w7224 , w7225 , w7226 , w7227 , w7228 , w7229 , w7230 , w7231 , w7232 , w7233 , w7234 , w7235 , w7236 , w7237 , w7238 , w7239 , w7240 , w7241 , w7242 , w7243 , w7244 , w7245 , w7246 , w7247 , w7248 , w7249 , w7250 , w7251 , w7252 , w7253 , w7254 , w7255 , w7256 , w7257 , w7258 , w7259 , w7260 , w7261 , w7262 , w7263 , w7264 , w7265 , w7266 , w7267 , w7268 , w7269 , w7270 , w7271 , w7272 , w7273 , w7274 , w7275 , w7276 , w7277 , w7278 , w7279 , w7280 , w7281 , w7282 , w7283 , w7284 , w7285 , w7286 , w7287 , w7288 , w7289 , w7290 , w7291 , w7292 , w7293 , w7294 , w7295 , w7296 , w7297 , w7298 , w7299 , w7300 , w7301 , w7302 , w7303 , w7304 , w7305 , w7306 , w7307 , w7308 , w7309 , w7310 , w7311 , w7312 , w7313 , w7314 , w7315 , w7316 , w7317 , w7318 , w7319 , w7320 , w7321 , w7322 , w7323 , w7324 , w7325 , w7326 , w7327 , w7328 , w7329 , w7330 , w7331 , w7332 , w7333 , w7334 , w7335 , w7336 , w7337 , w7338 , w7339 , w7340 , w7341 , w7342 , w7343 , w7344 , w7345 , w7346 , w7347 , w7348 , w7349 , w7350 , w7351 , w7352 , w7353 , w7354 , w7355 , w7356 , w7357 , w7358 , w7359 , w7360 , w7361 , w7362 , w7363 , w7364 , w7365 , w7366 , w7367 , w7368 , w7369 , w7370 , w7371 , w7372 , w7373 , w7374 , w7375 , w7376 , w7377 , w7378 , w7379 , w7380 , w7381 , w7382 , w7383 , w7384 , w7385 , w7386 , w7387 , w7388 , w7389 , w7390 , w7391 , w7392 , w7393 , w7394 , w7395 , w7396 , w7397 , w7398 , w7399 , w7400 , w7401 , w7402 , w7403 , w7404 , w7405 , w7406 , w7407 , w7408 , w7409 , w7410 , w7411 , w7412 , w7413 , w7414 , w7415 , w7416 , w7417 , w7418 , w7419 , w7420 , w7421 , w7422 , w7423 , w7424 , w7425 , w7426 , w7427 , w7428 , w7429 , w7430 , w7431 , w7432 , w7433 , w7434 , w7435 , w7436 , w7437 , w7438 , w7439 , w7440 , w7441 , w7442 , w7443 , w7444 , w7445 , w7446 , w7447 , w7448 , w7449 , w7450 , w7451 , w7452 , w7453 , w7454 , w7455 , w7456 , w7457 , w7458 , w7459 , w7460 , w7461 , w7462 , w7463 , w7464 , w7465 , w7466 , w7467 , w7468 , w7469 , w7470 , w7471 , w7472 , w7473 , w7474 , w7475 , w7476 , w7477 , w7478 , w7479 , w7480 , w7481 , w7482 , w7483 , w7484 , w7485 , w7486 , w7487 , w7488 , w7489 , w7490 , w7491 , w7492 , w7493 , w7494 , w7495 , w7496 , w7497 , w7498 , w7499 , w7500 , w7501 , w7502 , w7503 , w7504 , w7505 , w7506 , w7507 , w7508 , w7509 , w7510 , w7511 , w7512 , w7513 , w7514 , w7515 , w7516 , w7517 , w7518 , w7519 , w7520 , w7521 , w7522 , w7523 , w7524 , w7525 , w7526 , w7527 , w7528 , w7529 , w7530 , w7531 , w7532 , w7533 , w7534 , w7535 , w7536 , w7537 , w7538 , w7539 , w7540 , w7541 , w7542 , w7543 , w7544 , w7545 , w7546 , w7547 , w7548 , w7549 , w7550 , w7551 , w7552 , w7553 , w7554 , w7555 , w7556 , w7557 , w7558 , w7559 , w7560 , w7561 , w7562 , w7563 , w7564 , w7565 , w7566 , w7567 , w7568 , w7569 , w7570 , w7571 , w7572 , w7573 , w7574 , w7575 , w7576 , w7577 , w7578 , w7579 , w7580 , w7581 , w7582 , w7583 , w7584 , w7585 , w7586 , w7587 , w7588 , w7589 , w7590 , w7591 , w7592 , w7593 , w7594 , w7595 , w7596 , w7597 , w7598 , w7599 , w7600 , w7601 , w7602 , w7603 , w7604 , w7605 , w7606 , w7607 , w7608 , w7609 , w7610 , w7611 , w7612 , w7613 , w7614 , w7615 , w7616 , w7617 , w7618 , w7619 , w7620 , w7621 , w7622 , w7623 , w7624 , w7625 , w7626 , w7627 , w7628 , w7629 , w7630 , w7631 , w7632 , w7633 , w7634 , w7635 , w7636 , w7637 , w7638 , w7639 , w7640 , w7641 , w7642 , w7643 , w7644 , w7645 , w7646 , w7647 , w7648 , w7649 , w7650 , w7651 , w7652 , w7653 , w7654 , w7655 , w7656 , w7657 , w7658 , w7659 , w7660 , w7661 , w7662 , w7663 , w7664 , w7665 , w7666 , w7667 , w7668 , w7669 , w7670 , w7671 , w7672 , w7673 , w7674 , w7675 , w7676 , w7677 , w7678 , w7679 , w7680 , w7681 , w7682 , w7683 , w7684 , w7685 , w7686 , w7687 , w7688 , w7689 , w7690 , w7691 , w7692 , w7693 , w7694 , w7695 , w7696 , w7697 , w7698 , w7699 , w7700 , w7701 , w7702 , w7703 , w7704 , w7705 , w7706 , w7707 , w7708 , w7709 , w7710 , w7711 , w7712 , w7713 , w7714 , w7715 , w7716 , w7717 , w7718 , w7719 , w7720 , w7721 , w7722 , w7723 , w7724 , w7725 , w7726 , w7727 , w7728 , w7729 , w7730 , w7731 , w7732 , w7733 , w7734 , w7735 , w7736 , w7737 , w7738 , w7739 , w7740 , w7741 , w7742 , w7743 , w7744 , w7745 , w7746 , w7747 , w7748 , w7749 , w7750 , w7751 , w7752 , w7753 , w7754 , w7755 , w7756 , w7757 , w7758 , w7759 , w7760 , w7761 , w7762 , w7763 , w7764 , w7765 , w7766 , w7767 , w7768 , w7769 , w7770 , w7771 , w7772 , w7773 , w7774 , w7775 , w7776 , w7777 , w7778 , w7779 , w7780 , w7781 , w7782 , w7783 , w7784 , w7785 , w7786 , w7787 , w7788 , w7789 , w7790 , w7791 , w7792 , w7793 , w7794 , w7795 , w7796 , w7797 , w7798 , w7799 , w7800 , w7801 , w7802 , w7803 , w7804 , w7805 , w7806 , w7807 , w7808 , w7809 , w7810 , w7811 , w7812 , w7813 , w7814 , w7815 , w7816 , w7817 , w7818 , w7819 , w7820 , w7821 , w7822 , w7823 , w7824 , w7825 , w7826 , w7827 , w7828 , w7829 , w7830 , w7831 , w7832 , w7833 , w7834 , w7835 , w7836 , w7837 , w7838 , w7839 , w7840 , w7841 , w7842 , w7843 , w7844 , w7845 , w7846 , w7847 , w7848 , w7849 , w7850 , w7851 , w7852 , w7853 , w7854 , w7855 , w7856 , w7857 , w7858 , w7859 , w7860 , w7861 , w7862 , w7863 , w7864 , w7865 , w7866 , w7867 , w7868 , w7869 , w7870 , w7871 , w7872 , w7873 , w7874 , w7875 , w7876 , w7877 , w7878 , w7879 , w7880 , w7881 , w7882 , w7883 , w7884 , w7885 , w7886 , w7887 , w7888 , w7889 , w7890 , w7891 , w7892 , w7893 , w7894 , w7895 , w7896 , w7897 , w7898 , w7899 , w7900 , w7901 , w7902 , w7903 , w7904 , w7905 , w7906 , w7907 , w7908 , w7909 , w7910 , w7911 , w7912 , w7913 , w7914 , w7915 , w7916 , w7917 , w7918 , w7919 , w7920 , w7921 , w7922 , w7923 , w7924 , w7925 , w7926 , w7927 , w7928 , w7929 , w7930 , w7931 , w7932 , w7933 , w7934 , w7935 , w7936 , w7937 , w7938 , w7939 , w7940 , w7941 , w7942 , w7943 , w7944 , w7945 , w7946 , w7947 , w7948 , w7949 , w7950 , w7951 , w7952 , w7953 , w7954 , w7955 , w7956 , w7957 , w7958 , w7959 , w7960 , w7961 , w7962 , w7963 , w7964 , w7965 , w7966 , w7967 , w7968 , w7969 , w7970 , w7971 , w7972 , w7973 , w7974 , w7975 , w7976 , w7977 , w7978 , w7979 , w7980 , w7981 , w7982 , w7983 , w7984 , w7985 , w7986 , w7987 , w7988 , w7989 , w7990 , w7991 , w7992 , w7993 , w7994 , w7995 , w7996 , w7997 , w7998 , w7999 , w8000 , w8001 , w8002 , w8003 , w8004 , w8005 , w8006 , w8007 , w8008 , w8009 , w8010 , w8011 , w8012 , w8013 , w8014 , w8015 , w8016 , w8017 , w8018 , w8019 , w8020 , w8021 , w8022 , w8023 , w8024 , w8025 , w8026 , w8027 , w8028 , w8029 , w8030 , w8031 , w8032 , w8033 , w8034 , w8035 , w8036 , w8037 , w8038 , w8039 , w8040 , w8041 , w8042 , w8043 , w8044 , w8045 , w8046 , w8047 , w8048 , w8049 , w8050 , w8051 , w8052 , w8053 , w8054 , w8055 , w8056 , w8057 , w8058 , w8059 , w8060 , w8061 , w8062 , w8063 , w8064 , w8065 , w8066 , w8067 , w8068 , w8069 , w8070 , w8071 , w8072 , w8073 , w8074 , w8075 , w8076 , w8077 , w8078 , w8079 , w8080 , w8081 , w8082 , w8083 , w8084 , w8085 , w8086 , w8087 , w8088 , w8089 , w8090 , w8091 , w8092 , w8093 , w8094 , w8095 , w8096 , w8097 , w8098 , w8099 , w8100 , w8101 , w8102 , w8103 , w8104 , w8105 , w8106 , w8107 , w8108 , w8109 , w8110 , w8111 , w8112 , w8113 , w8114 , w8115 , w8116 , w8117 , w8118 , w8119 , w8120 , w8121 , w8122 , w8123 , w8124 , w8125 , w8126 , w8127 , w8128 , w8129 , w8130 , w8131 , w8132 , w8133 , w8134 , w8135 , w8136 , w8137 , w8138 , w8139 , w8140 , w8141 , w8142 , w8143 , w8144 , w8145 , w8146 , w8147 , w8148 , w8149 , w8150 , w8151 , w8152 , w8153 , w8154 , w8155 , w8156 , w8157 , w8158 , w8159 , w8160 , w8161 , w8162 , w8163 , w8164 , w8165 , w8166 , w8167 , w8168 , w8169 , w8170 , w8171 , w8172 , w8173 , w8174 , w8175 , w8176 , w8177 , w8178 , w8179 , w8180 , w8181 , w8182 , w8183 , w8184 , w8185 , w8186 , w8187 , w8188 , w8189 , w8190 , w8191 , w8192 , w8193 , w8194 , w8195 , w8196 , w8197 , w8198 , w8199 , w8200 , w8201 , w8202 , w8203 , w8204 , w8205 , w8206 , w8207 , w8208 , w8209 , w8210 , w8211 , w8212 , w8213 , w8214 , w8215 , w8216 , w8217 , w8218 , w8219 , w8220 , w8221 , w8222 , w8223 , w8224 , w8225 , w8226 , w8227 , w8228 , w8229 , w8230 , w8231 , w8232 , w8233 , w8234 , w8235 , w8236 , w8237 , w8238 , w8239 , w8240 , w8241 , w8242 , w8243 , w8244 , w8245 , w8246 , w8247 , w8248 , w8249 , w8250 , w8251 , w8252 , w8253 , w8254 , w8255 , w8256 , w8257 , w8258 , w8259 , w8260 , w8261 , w8262 , w8263 , w8264 , w8265 , w8266 , w8267 , w8268 , w8269 , w8270 , w8271 , w8272 , w8273 , w8274 , w8275 , w8276 , w8277 , w8278 , w8279 , w8280 , w8281 , w8282 , w8283 , w8284 , w8285 , w8286 , w8287 , w8288 , w8289 , w8290 , w8291 , w8292 , w8293 , w8294 , w8295 , w8296 , w8297 , w8298 , w8299 , w8300 , w8301 , w8302 , w8303 , w8304 , w8305 , w8306 , w8307 , w8308 , w8309 , w8310 , w8311 , w8312 , w8313 , w8314 , w8315 , w8316 , w8317 , w8318 , w8319 , w8320 , w8321 , w8322 , w8323 , w8324 , w8325 , w8326 , w8327 , w8328 , w8329 , w8330 , w8331 , w8332 , w8333 , w8334 , w8335 , w8336 , w8337 , w8338 , w8339 , w8340 , w8341 , w8342 , w8343 , w8344 , w8345 , w8346 , w8347 , w8348 , w8349 , w8350 , w8351 , w8352 , w8353 , w8354 , w8355 , w8356 , w8357 , w8358 , w8359 , w8360 , w8361 , w8362 , w8363 , w8364 , w8365 , w8366 , w8367 , w8368 , w8369 , w8370 , w8371 , w8372 , w8373 , w8374 , w8375 , w8376 , w8377 , w8378 , w8379 , w8380 , w8381 , w8382 , w8383 , w8384 , w8385 , w8386 , w8387 , w8388 , w8389 , w8390 , w8391 , w8392 , w8393 , w8394 , w8395 , w8396 , w8397 , w8398 , w8399 , w8400 , w8401 , w8402 , w8403 , w8404 , w8405 , w8406 , w8407 , w8408 , w8409 , w8410 , w8411 , w8412 , w8413 , w8414 , w8415 , w8416 , w8417 , w8418 , w8419 , w8420 , w8421 , w8422 , w8423 , w8424 , w8425 , w8426 , w8427 , w8428 , w8429 , w8430 , w8431 , w8432 , w8433 , w8434 , w8435 , w8436 , w8437 , w8438 , w8439 , w8440 , w8441 , w8442 , w8443 , w8444 , w8445 , w8446 , w8447 , w8448 , w8449 , w8450 , w8451 , w8452 , w8453 , w8454 , w8455 , w8456 , w8457 , w8458 , w8459 , w8460 , w8461 , w8462 , w8463 , w8464 , w8465 , w8466 , w8467 , w8468 , w8469 , w8470 , w8471 , w8472 , w8473 , w8474 , w8475 , w8476 , w8477 , w8478 , w8479 , w8480 , w8481 , w8482 , w8483 , w8484 , w8485 , w8486 , w8487 , w8488 , w8489 , w8490 , w8491 , w8492 , w8493 , w8494 , w8495 , w8496 , w8497 , w8498 , w8499 , w8500 , w8501 , w8502 , w8503 , w8504 , w8505 , w8506 , w8507 , w8508 , w8509 , w8510 , w8511 , w8512 , w8513 , w8514 , w8515 , w8516 , w8517 , w8518 , w8519 , w8520 , w8521 , w8522 , w8523 , w8524 , w8525 , w8526 , w8527 , w8528 , w8529 , w8530 , w8531 , w8532 , w8533 , w8534 , w8535 , w8536 , w8537 , w8538 , w8539 , w8540 , w8541 , w8542 , w8543 , w8544 , w8545 , w8546 , w8547 , w8548 , w8549 , w8550 , w8551 , w8552 , w8553 , w8554 , w8555 , w8556 , w8557 , w8558 , w8559 , w8560 , w8561 , w8562 , w8563 , w8564 , w8565 , w8566 , w8567 , w8568 , w8569 , w8570 , w8571 , w8572 , w8573 , w8574 , w8575 , w8576 , w8577 , w8578 , w8579 , w8580 , w8581 , w8582 , w8583 , w8584 , w8585 , w8586 , w8587 , w8588 , w8589 , w8590 , w8591 , w8592 , w8593 , w8594 , w8595 , w8596 , w8597 , w8598 , w8599 , w8600 , w8601 , w8602 , w8603 , w8604 , w8605 , w8606 , w8607 , w8608 , w8609 , w8610 , w8611 , w8612 , w8613 , w8614 , w8615 , w8616 , w8617 , w8618 , w8619 , w8620 , w8621 , w8622 , w8623 , w8624 , w8625 , w8626 , w8627 , w8628 , w8629 , w8630 , w8631 , w8632 , w8633 , w8634 , w8635 , w8636 , w8637 , w8638 , w8639 , w8640 , w8641 , w8642 , w8643 , w8644 , w8645 , w8646 , w8647 , w8648 , w8649 , w8650 , w8651 , w8652 , w8653 , w8654 , w8655 , w8656 , w8657 , w8658 , w8659 , w8660 , w8661 , w8662 , w8663 , w8664 , w8665 , w8666 , w8667 , w8668 , w8669 , w8670 , w8671 , w8672 , w8673 , w8674 , w8675 , w8676 , w8677 , w8678 , w8679 , w8680 , w8681 , w8682 , w8683 , w8684 , w8685 , w8686 , w8687 , w8688 , w8689 , w8690 , w8691 , w8692 , w8693 , w8694 , w8695 , w8696 , w8697 , w8698 , w8699 , w8700 , w8701 , w8702 , w8703 , w8704 , w8705 , w8706 , w8707 , w8708 , w8709 , w8710 , w8711 , w8712 , w8713 , w8714 , w8715 , w8716 , w8717 , w8718 , w8719 , w8720 , w8721 , w8722 , w8723 , w8724 , w8725 , w8726 , w8727 , w8728 , w8729 , w8730 , w8731 , w8732 , w8733 , w8734 , w8735 , w8736 , w8737 , w8738 , w8739 , w8740 , w8741 , w8742 , w8743 , w8744 , w8745 , w8746 , w8747 , w8748 , w8749 , w8750 , w8751 , w8752 , w8753 , w8754 , w8755 , w8756 , w8757 , w8758 , w8759 , w8760 , w8761 , w8762 , w8763 , w8764 , w8765 , w8766 , w8767 , w8768 , w8769 , w8770 , w8771 , w8772 , w8773 , w8774 , w8775 , w8776 , w8777 , w8778 , w8779 , w8780 , w8781 , w8782 , w8783 , w8784 , w8785 , w8786 , w8787 , w8788 , w8789 , w8790 , w8791 , w8792 , w8793 , w8794 , w8795 , w8796 , w8797 , w8798 , w8799 , w8800 , w8801 , w8802 , w8803 , w8804 , w8805 , w8806 , w8807 , w8808 , w8809 , w8810 , w8811 , w8812 , w8813 , w8814 , w8815 , w8816 , w8817 , w8818 , w8819 , w8820 , w8821 , w8822 , w8823 , w8824 , w8825 , w8826 , w8827 , w8828 , w8829 , w8830 , w8831 , w8832 , w8833 , w8834 , w8835 , w8836 , w8837 , w8838 , w8839 , w8840 , w8841 , w8842 , w8843 , w8844 , w8845 , w8846 , w8847 , w8848 , w8849 , w8850 , w8851 , w8852 , w8853 , w8854 , w8855 , w8856 , w8857 , w8858 , w8859 , w8860 , w8861 , w8862 , w8863 , w8864 , w8865 , w8866 , w8867 , w8868 , w8869 , w8870 , w8871 , w8872 , w8873 , w8874 , w8875 , w8876 , w8877 , w8878 , w8879 , w8880 , w8881 , w8882 , w8883 , w8884 , w8885 , w8886 , w8887 , w8888 , w8889 , w8890 , w8891 , w8892 , w8893 , w8894 , w8895 , w8896 , w8897 , w8898 , w8899 , w8900 , w8901 , w8902 , w8903 , w8904 , w8905 , w8906 , w8907 , w8908 , w8909 , w8910 , w8911 , w8912 , w8913 , w8914 , w8915 , w8916 , w8917 , w8918 , w8919 , w8920 , w8921 , w8922 , w8923 , w8924 , w8925 , w8926 , w8927 , w8928 , w8929 , w8930 , w8931 , w8932 , w8933 , w8934 , w8935 , w8936 , w8937 , w8938 , w8939 , w8940 , w8941 , w8942 , w8943 , w8944 , w8945 , w8946 , w8947 , w8948 , w8949 , w8950 , w8951 , w8952 , w8953 , w8954 , w8955 , w8956 , w8957 , w8958 , w8959 , w8960 , w8961 , w8962 , w8963 , w8964 , w8965 , w8966 , w8967 , w8968 , w8969 , w8970 , w8971 , w8972 , w8973 , w8974 , w8975 , w8976 , w8977 , w8978 , w8979 , w8980 , w8981 , w8982 , w8983 , w8984 , w8985 , w8986 , w8987 , w8988 , w8989 , w8990 , w8991 , w8992 , w8993 , w8994 , w8995 , w8996 , w8997 , w8998 , w8999 , w9000 , w9001 , w9002 , w9003 , w9004 , w9005 , w9006 , w9007 , w9008 , w9009 , w9010 , w9011 , w9012 , w9013 , w9014 , w9015 , w9016 , w9017 , w9018 , w9019 , w9020 , w9021 , w9022 , w9023 , w9024 , w9025 , w9026 , w9027 , w9028 , w9029 , w9030 , w9031 , w9032 , w9033 , w9034 , w9035 , w9036 , w9037 , w9038 , w9039 , w9040 , w9041 , w9042 , w9043 , w9044 , w9045 , w9046 , w9047 , w9048 , w9049 , w9050 , w9051 , w9052 , w9053 , w9054 , w9055 , w9056 , w9057 , w9058 , w9059 , w9060 , w9061 , w9062 , w9063 , w9064 , w9065 , w9066 , w9067 , w9068 , w9069 , w9070 , w9071 , w9072 , w9073 , w9074 , w9075 , w9076 , w9077 , w9078 , w9079 , w9080 , w9081 , w9082 , w9083 , w9084 , w9085 , w9086 , w9087 , w9088 , w9089 , w9090 , w9091 , w9092 , w9093 , w9094 , w9095 , w9096 , w9097 , w9098 , w9099 , w9100 , w9101 , w9102 , w9103 , w9104 , w9105 , w9106 , w9107 , w9108 , w9109 , w9110 , w9111 , w9112 , w9113 , w9114 , w9115 , w9116 , w9117 , w9118 , w9119 , w9120 , w9121 , w9122 , w9123 , w9124 , w9125 , w9126 , w9127 , w9128 , w9129 , w9130 , w9131 , w9132 , w9133 , w9134 , w9135 , w9136 , w9137 , w9138 , w9139 , w9140 , w9141 , w9142 , w9143 , w9144 , w9145 , w9146 , w9147 , w9148 , w9149 , w9150 , w9151 , w9152 , w9153 , w9154 , w9155 , w9156 , w9157 , w9158 , w9159 , w9160 , w9161 , w9162 , w9163 , w9164 , w9165 , w9166 , w9167 , w9168 , w9169 , w9170 , w9171 , w9172 , w9173 , w9174 , w9175 , w9176 , w9177 , w9178 , w9179 , w9180 , w9181 , w9182 , w9183 , w9184 , w9185 , w9186 , w9187 , w9188 , w9189 , w9190 , w9191 , w9192 , w9193 , w9194 , w9195 , w9196 , w9197 , w9198 , w9199 , w9200 , w9201 , w9202 , w9203 , w9204 , w9205 , w9206 , w9207 , w9208 , w9209 , w9210 , w9211 , w9212 , w9213 , w9214 , w9215 , w9216 , w9217 , w9218 , w9219 , w9220 , w9221 , w9222 , w9223 , w9224 , w9225 , w9226 , w9227 , w9228 , w9229 , w9230 , w9231 , w9232 , w9233 , w9234 , w9235 , w9236 , w9237 , w9238 , w9239 , w9240 , w9241 , w9242 , w9243 , w9244 , w9245 , w9246 , w9247 , w9248 , w9249 , w9250 , w9251 , w9252 , w9253 , w9254 , w9255 , w9256 , w9257 , w9258 , w9259 , w9260 , w9261 , w9262 , w9263 , w9264 , w9265 , w9266 , w9267 , w9268 , w9269 , w9270 , w9271 , w9272 , w9273 , w9274 , w9275 , w9276 , w9277 , w9278 , w9279 , w9280 , w9281 , w9282 , w9283 , w9284 , w9285 , w9286 , w9287 , w9288 , w9289 , w9290 , w9291 , w9292 , w9293 , w9294 , w9295 , w9296 , w9297 , w9298 , w9299 , w9300 , w9301 , w9302 , w9303 , w9304 , w9305 , w9306 , w9307 , w9308 , w9309 , w9310 , w9311 , w9312 , w9313 , w9314 , w9315 , w9316 , w9317 , w9318 , w9319 , w9320 , w9321 , w9322 , w9323 , w9324 , w9325 , w9326 , w9327 , w9328 , w9329 , w9330 , w9331 , w9332 , w9333 , w9334 , w9335 , w9336 , w9337 , w9338 , w9339 , w9340 , w9341 , w9342 , w9343 , w9344 , w9345 , w9346 , w9347 , w9348 , w9349 , w9350 , w9351 , w9352 , w9353 , w9354 , w9355 , w9356 , w9357 , w9358 , w9359 , w9360 , w9361 , w9362 , w9363 , w9364 , w9365 , w9366 , w9367 , w9368 , w9369 , w9370 , w9371 , w9372 , w9373 , w9374 , w9375 , w9376 , w9377 , w9378 , w9379 , w9380 , w9381 , w9382 , w9383 , w9384 , w9385 , w9386 , w9387 , w9388 , w9389 , w9390 , w9391 , w9392 , w9393 , w9394 , w9395 , w9396 , w9397 , w9398 , w9399 , w9400 , w9401 , w9402 , w9403 , w9404 , w9405 , w9406 , w9407 , w9408 , w9409 , w9410 , w9411 , w9412 , w9413 , w9414 , w9415 , w9416 , w9417 , w9418 , w9419 , w9420 , w9421 , w9422 , w9423 , w9424 , w9425 , w9426 , w9427 , w9428 , w9429 , w9430 , w9431 , w9432 , w9433 , w9434 , w9435 , w9436 , w9437 , w9438 , w9439 , w9440 , w9441 , w9442 , w9443 , w9444 , w9445 , w9446 , w9447 , w9448 , w9449 , w9450 , w9451 , w9452 , w9453 , w9454 , w9455 , w9456 , w9457 , w9458 , w9459 , w9460 , w9461 , w9462 , w9463 , w9464 , w9465 , w9466 , w9467 , w9468 , w9469 , w9470 , w9471 , w9472 , w9473 , w9474 , w9475 , w9476 , w9477 , w9478 , w9479 , w9480 , w9481 , w9482 , w9483 , w9484 , w9485 , w9486 , w9487 , w9488 , w9489 , w9490 , w9491 , w9492 , w9493 , w9494 , w9495 , w9496 , w9497 , w9498 , w9499 , w9500 , w9501 , w9502 , w9503 , w9504 , w9505 , w9506 , w9507 , w9508 , w9509 , w9510 , w9511 , w9512 , w9513 , w9514 , w9515 , w9516 , w9517 , w9518 , w9519 , w9520 , w9521 , w9522 , w9523 , w9524 , w9525 , w9526 , w9527 , w9528 , w9529 , w9530 , w9531 , w9532 , w9533 , w9534 , w9535 , w9536 , w9537 , w9538 , w9539 , w9540 , w9541 , w9542 , w9543 , w9544 , w9545 , w9546 , w9547 , w9548 , w9549 , w9550 , w9551 , w9552 , w9553 , w9554 , w9555 , w9556 , w9557 , w9558 , w9559 , w9560 , w9561 , w9562 , w9563 , w9564 , w9565 , w9566 , w9567 , w9568 , w9569 , w9570 , w9571 , w9572 , w9573 , w9574 , w9575 , w9576 , w9577 , w9578 , w9579 , w9580 , w9581 , w9582 , w9583 , w9584 , w9585 , w9586 , w9587 , w9588 , w9589 , w9590 , w9591 , w9592 , w9593 , w9594 , w9595 , w9596 , w9597 , w9598 , w9599 , w9600 , w9601 , w9602 , w9603 , w9604 , w9605 , w9606 , w9607 , w9608 , w9609 , w9610 , w9611 , w9612 , w9613 , w9614 , w9615 , w9616 , w9617 , w9618 , w9619 , w9620 , w9621 , w9622 , w9623 , w9624 , w9625 , w9626 , w9627 , w9628 , w9629 , w9630 , w9631 , w9632 , w9633 , w9634 , w9635 , w9636 , w9637 , w9638 , w9639 , w9640 , w9641 , w9642 , w9643 , w9644 , w9645 , w9646 , w9647 , w9648 , w9649 , w9650 , w9651 , w9652 , w9653 , w9654 , w9655 , w9656 , w9657 , w9658 , w9659 , w9660 , w9661 , w9662 , w9663 , w9664 , w9665 , w9666 , w9667 , w9668 , w9669 , w9670 , w9671 , w9672 , w9673 , w9674 , w9675 , w9676 , w9677 , w9678 , w9679 , w9680 , w9681 , w9682 , w9683 , w9684 , w9685 , w9686 , w9687 , w9688 , w9689 , w9690 , w9691 , w9692 , w9693 , w9694 , w9695 , w9696 , w9697 , w9698 , w9699 , w9700 , w9701 , w9702 , w9703 , w9704 , w9705 , w9706 , w9707 , w9708 , w9709 , w9710 , w9711 , w9712 , w9713 , w9714 , w9715 , w9716 , w9717 , w9718 , w9719 , w9720 , w9721 , w9722 , w9723 , w9724 , w9725 , w9726 , w9727 , w9728 , w9729 , w9730 , w9731 , w9732 , w9733 , w9734 , w9735 , w9736 , w9737 , w9738 , w9739 , w9740 , w9741 , w9742 , w9743 , w9744 , w9745 , w9746 , w9747 , w9748 , w9749 , w9750 , w9751 , w9752 , w9753 , w9754 , w9755 , w9756 , w9757 , w9758 , w9759 , w9760 , w9761 , w9762 , w9763 , w9764 , w9765 , w9766 , w9767 , w9768 , w9769 , w9770 , w9771 , w9772 , w9773 , w9774 , w9775 , w9776 , w9777 , w9778 , w9779 , w9780 , w9781 , w9782 , w9783 , w9784 , w9785 , w9786 , w9787 , w9788 , w9789 , w9790 , w9791 , w9792 , w9793 , w9794 , w9795 , w9796 , w9797 , w9798 , w9799 , w9800 , w9801 , w9802 , w9803 , w9804 , w9805 , w9806 , w9807 , w9808 , w9809 , w9810 , w9811 , w9812 , w9813 , w9814 , w9815 , w9816 , w9817 , w9818 , w9819 , w9820 , w9821 , w9822 , w9823 , w9824 , w9825 , w9826 , w9827 , w9828 , w9829 , w9830 , w9831 , w9832 , w9833 , w9834 , w9835 , w9836 , w9837 , w9838 , w9839 , w9840 , w9841 , w9842 , w9843 , w9844 , w9845 , w9846 , w9847 , w9848 , w9849 , w9850 , w9851 , w9852 , w9853 , w9854 , w9855 , w9856 , w9857 , w9858 , w9859 , w9860 , w9861 , w9862 , w9863 , w9864 , w9865 , w9866 , w9867 , w9868 , w9869 , w9870 , w9871 , w9872 , w9873 , w9874 , w9875 , w9876 , w9877 , w9878 , w9879 , w9880 , w9881 , w9882 , w9883 , w9884 , w9885 , w9886 , w9887 , w9888 , w9889 , w9890 , w9891 , w9892 , w9893 , w9894 , w9895 , w9896 , w9897 , w9898 , w9899 , w9900 , w9901 , w9902 , w9903 , w9904 , w9905 , w9906 , w9907 , w9908 , w9909 , w9910 , w9911 , w9912 , w9913 , w9914 , w9915 , w9916 , w9917 , w9918 , w9919 , w9920 , w9921 , w9922 , w9923 , w9924 , w9925 , w9926 , w9927 , w9928 , w9929 , w9930 , w9931 , w9932 , w9933 , w9934 , w9935 , w9936 , w9937 , w9938 , w9939 , w9940 , w9941 , w9942 , w9943 , w9944 , w9945 , w9946 , w9947 , w9948 , w9949 , w9950 , w9951 , w9952 , w9953 , w9954 , w9955 , w9956 , w9957 , w9958 , w9959 , w9960 , w9961 , w9962 , w9963 , w9964 , w9965 , w9966 , w9967 , w9968 , w9969 , w9970 , w9971 , w9972 , w9973 , w9974 , w9975 , w9976 , w9977 , w9978 , w9979 , w9980 , w9981 , w9982 , w9983 , w9984 , w9985 , w9986 , w9987 , w9988 , w9989 , w9990 , w9991 , w9992 , w9993 , w9994 , w9995 , w9996 , w9997 , w9998 , w9999 , w10000 , w10001 , w10002 , w10003 , w10004 , w10005 , w10006 , w10007 , w10008 , w10009 , w10010 , w10011 , w10012 , w10013 , w10014 , w10015 , w10016 , w10017 , w10018 , w10019 , w10020 , w10021 , w10022 , w10023 , w10024 , w10025 , w10026 , w10027 , w10028 , w10029 , w10030 , w10031 , w10032 , w10033 , w10034 , w10035 , w10036 , w10037 , w10038 , w10039 , w10040 , w10041 , w10042 , w10043 , w10044 , w10045 , w10046 , w10047 , w10048 , w10049 , w10050 , w10051 , w10052 , w10053 , w10054 , w10055 , w10056 , w10057 , w10058 , w10059 , w10060 , w10061 , w10062 , w10063 , w10064 , w10065 , w10066 , w10067 , w10068 , w10069 , w10070 , w10071 , w10072 , w10073 , w10074 , w10075 , w10076 , w10077 , w10078 , w10079 , w10080 , w10081 , w10082 , w10083 , w10084 , w10085 , w10086 , w10087 , w10088 , w10089 , w10090 , w10091 , w10092 , w10093 , w10094 , w10095 , w10096 , w10097 , w10098 , w10099 , w10100 , w10101 , w10102 , w10103 , w10104 , w10105 , w10106 , w10107 , w10108 , w10109 , w10110 , w10111 , w10112 , w10113 , w10114 , w10115 , w10116 , w10117 , w10118 , w10119 , w10120 , w10121 , w10122 , w10123 , w10124 , w10125 , w10126 , w10127 , w10128 , w10129 , w10130 , w10131 , w10132 , w10133 , w10134 , w10135 , w10136 , w10137 , w10138 , w10139 , w10140 , w10141 , w10142 , w10143 , w10144 , w10145 , w10146 , w10147 , w10148 , w10149 , w10150 , w10151 , w10152 , w10153 , w10154 , w10155 , w10156 , w10157 , w10158 , w10159 , w10160 , w10161 , w10162 , w10163 , w10164 , w10165 , w10166 , w10167 , w10168 , w10169 , w10170 , w10171 , w10172 , w10173 , w10174 , w10175 , w10176 , w10177 , w10178 , w10179 , w10180 , w10181 , w10182 , w10183 , w10184 , w10185 , w10186 , w10187 , w10188 , w10189 , w10190 , w10191 , w10192 , w10193 , w10194 , w10195 , w10196 , w10197 , w10198 , w10199 , w10200 , w10201 , w10202 , w10203 , w10204 , w10205 , w10206 , w10207 , w10208 , w10209 , w10210 , w10211 , w10212 , w10213 , w10214 , w10215 , w10216 , w10217 , w10218 , w10219 , w10220 , w10221 , w10222 , w10223 , w10224 , w10225 , w10226 , w10227 , w10228 , w10229 , w10230 , w10231 , w10232 , w10233 , w10234 , w10235 , w10236 , w10237 , w10238 , w10239 , w10240 , w10241 , w10242 , w10243 , w10244 , w10245 , w10246 , w10247 , w10248 , w10249 , w10250 , w10251 , w10252 , w10253 , w10254 , w10255 , w10256 , w10257 , w10258 , w10259 , w10260 , w10261 , w10262 , w10263 , w10264 , w10265 , w10266 , w10267 , w10268 , w10269 , w10270 , w10271 , w10272 , w10273 , w10274 , w10275 , w10276 , w10277 , w10278 , w10279 , w10280 , w10281 , w10282 , w10283 , w10284 , w10285 , w10286 , w10287 , w10288 , w10289 , w10290 , w10291 , w10292 , w10293 , w10294 , w10295 , w10296 , w10297 , w10298 , w10299 , w10300 , w10301 , w10302 , w10303 , w10304 , w10305 , w10306 , w10307 , w10308 , w10309 , w10310 , w10311 , w10312 , w10313 , w10314 , w10315 , w10316 , w10317 , w10318 , w10319 , w10320 , w10321 , w10322 , w10323 , w10324 , w10325 , w10326 , w10327 , w10328 , w10329 , w10330 , w10331 , w10332 , w10333 , w10334 , w10335 , w10336 , w10337 , w10338 , w10339 , w10340 , w10341 , w10342 , w10343 , w10344 , w10345 , w10346 , w10347 , w10348 , w10349 , w10350 , w10351 , w10352 , w10353 , w10354 , w10355 , w10356 , w10357 , w10358 , w10359 , w10360 , w10361 , w10362 , w10363 , w10364 , w10365 , w10366 , w10367 , w10368 , w10369 , w10370 , w10371 , w10372 , w10373 , w10374 , w10375 , w10376 , w10377 , w10378 , w10379 , w10380 , w10381 , w10382 , w10383 , w10384 , w10385 , w10386 , w10387 , w10388 , w10389 , w10390 , w10391 , w10392 , w10393 , w10394 , w10395 , w10396 , w10397 , w10398 , w10399 , w10400 , w10401 , w10402 , w10403 , w10404 , w10405 , w10406 , w10407 , w10408 , w10409 , w10410 , w10411 , w10412 , w10413 , w10414 , w10415 , w10416 , w10417 , w10418 , w10419 , w10420 , w10421 , w10422 , w10423 , w10424 , w10425 , w10426 , w10427 , w10428 , w10429 , w10430 , w10431 , w10432 , w10433 , w10434 , w10435 , w10436 , w10437 , w10438 , w10439 , w10440 , w10441 , w10442 , w10443 , w10444 , w10445 , w10446 , w10447 , w10448 , w10449 , w10450 , w10451 , w10452 , w10453 , w10454 , w10455 , w10456 , w10457 , w10458 , w10459 , w10460 , w10461 , w10462 , w10463 , w10464 , w10465 , w10466 , w10467 , w10468 , w10469 , w10470 , w10471 , w10472 , w10473 , w10474 , w10475 , w10476 , w10477 , w10478 , w10479 , w10480 , w10481 , w10482 , w10483 , w10484 , w10485 , w10486 , w10487 , w10488 , w10489 , w10490 , w10491 , w10492 , w10493 , w10494 , w10495 , w10496 , w10497 , w10498 , w10499 , w10500 , w10501 , w10502 , w10503 , w10504 , w10505 , w10506 , w10507 , w10508 , w10509 , w10510 , w10511 , w10512 , w10513 , w10514 , w10515 , w10516 , w10517 , w10518 , w10519 , w10520 , w10521 , w10522 , w10523 , w10524 , w10525 , w10526 , w10527 , w10528 , w10529 , w10530 , w10531 , w10532 , w10533 , w10534 , w10535 , w10536 , w10537 , w10538 , w10539 , w10540 , w10541 , w10542 , w10543 , w10544 , w10545 , w10546 , w10547 , w10548 , w10549 , w10550 , w10551 , w10552 , w10553 , w10554 , w10555 , w10556 , w10557 , w10558 , w10559 , w10560 , w10561 , w10562 , w10563 , w10564 , w10565 , w10566 , w10567 , w10568 , w10569 , w10570 , w10571 , w10572 , w10573 , w10574 , w10575 , w10576 , w10577 , w10578 , w10579 , w10580 , w10581 , w10582 , w10583 , w10584 , w10585 , w10586 , w10587 , w10588 , w10589 , w10590 , w10591 , w10592 , w10593 , w10594 , w10595 , w10596 , w10597 , w10598 , w10599 , w10600 , w10601 , w10602 , w10603 , w10604 , w10605 , w10606 , w10607 , w10608 , w10609 , w10610 , w10611 , w10612 , w10613 , w10614 , w10615 , w10616 , w10617 , w10618 , w10619 , w10620 , w10621 , w10622 , w10623 , w10624 , w10625 , w10626 , w10627 , w10628 , w10629 , w10630 , w10631 , w10632 , w10633 , w10634 , w10635 , w10636 , w10637 , w10638 , w10639 , w10640 , w10641 , w10642 , w10643 , w10644 , w10645 , w10646 , w10647 , w10648 , w10649 , w10650 , w10651 , w10652 , w10653 , w10654 , w10655 , w10656 , w10657 , w10658 , w10659 , w10660 , w10661 , w10662 , w10663 , w10664 , w10665 , w10666 , w10667 , w10668 , w10669 , w10670 , w10671 , w10672 , w10673 , w10674 , w10675 , w10676 , w10677 , w10678 , w10679 , w10680 , w10681 , w10682 , w10683 , w10684 , w10685 , w10686 , w10687 , w10688 , w10689 , w10690 , w10691 , w10692 , w10693 , w10694 , w10695 , w10696 , w10697 , w10698 , w10699 , w10700 , w10701 , w10702 , w10703 , w10704 , w10705 , w10706 , w10707 , w10708 , w10709 , w10710 , w10711 , w10712 , w10713 , w10714 , w10715 , w10716 , w10717 , w10718 , w10719 , w10720 , w10721 , w10722 , w10723 , w10724 , w10725 , w10726 , w10727 , w10728 , w10729 , w10730 , w10731 , w10732 , w10733 , w10734 , w10735 , w10736 , w10737 , w10738 , w10739 , w10740 , w10741 , w10742 , w10743 , w10744 , w10745 , w10746 , w10747 , w10748 , w10749 , w10750 , w10751 , w10752 , w10753 , w10754 , w10755 , w10756 , w10757 , w10758 , w10759 , w10760 , w10761 , w10762 , w10763 , w10764 , w10765 , w10766 , w10767 , w10768 , w10769 , w10770 , w10771 , w10772 , w10773 , w10774 , w10775 , w10776 , w10777 , w10778 , w10779 , w10780 , w10781 , w10782 , w10783 , w10784 , w10785 , w10786 , w10787 , w10788 , w10789 , w10790 , w10791 , w10792 , w10793 , w10794 , w10795 , w10796 , w10797 , w10798 , w10799 , w10800 , w10801 , w10802 , w10803 , w10804 , w10805 , w10806 , w10807 , w10808 , w10809 , w10810 , w10811 , w10812 , w10813 , w10814 , w10815 , w10816 , w10817 , w10818 , w10819 , w10820 , w10821 , w10822 , w10823 , w10824 , w10825 , w10826 , w10827 , w10828 , w10829 , w10830 , w10831 , w10832 , w10833 , w10834 , w10835 , w10836 , w10837 , w10838 , w10839 , w10840 , w10841 , w10842 , w10843 , w10844 , w10845 , w10846 , w10847 , w10848 , w10849 , w10850 , w10851 , w10852 , w10853 , w10854 , w10855 , w10856 , w10857 , w10858 , w10859 , w10860 , w10861 , w10862 , w10863 , w10864 , w10865 , w10866 , w10867 , w10868 , w10869 , w10870 , w10871 , w10872 , w10873 , w10874 , w10875 , w10876 , w10877 , w10878 , w10879 , w10880 , w10881 , w10882 , w10883 , w10884 , w10885 , w10886 , w10887 , w10888 , w10889 , w10890 , w10891 , w10892 , w10893 , w10894 , w10895 , w10896 , w10897 , w10898 , w10899 , w10900 , w10901 , w10902 , w10903 , w10904 , w10905 , w10906 , w10907 , w10908 , w10909 , w10910 , w10911 , w10912 , w10913 , w10914 , w10915 , w10916 , w10917 , w10918 , w10919 , w10920 , w10921 , w10922 , w10923 , w10924 , w10925 , w10926 , w10927 , w10928 , w10929 , w10930 , w10931 , w10932 , w10933 , w10934 , w10935 , w10936 , w10937 , w10938 , w10939 , w10940 , w10941 , w10942 , w10943 , w10944 , w10945 , w10946 , w10947 , w10948 , w10949 , w10950 , w10951 , w10952 , w10953 , w10954 , w10955 , w10956 , w10957 , w10958 , w10959 , w10960 , w10961 , w10962 , w10963 , w10964 , w10965 , w10966 , w10967 , w10968 , w10969 , w10970 , w10971 , w10972 , w10973 , w10974 , w10975 , w10976 , w10977 , w10978 , w10979 , w10980 , w10981 , w10982 , w10983 , w10984 , w10985 , w10986 , w10987 , w10988 , w10989 , w10990 , w10991 , w10992 , w10993 , w10994 , w10995 , w10996 , w10997 , w10998 , w10999 , w11000 , w11001 , w11002 , w11003 , w11004 , w11005 , w11006 , w11007 , w11008 , w11009 , w11010 , w11011 , w11012 , w11013 , w11014 , w11015 , w11016 , w11017 , w11018 , w11019 , w11020 , w11021 , w11022 , w11023 , w11024 , w11025 , w11026 , w11027 , w11028 , w11029 , w11030 , w11031 , w11032 , w11033 , w11034 , w11035 , w11036 , w11037 , w11038 , w11039 , w11040 , w11041 , w11042 , w11043 , w11044 , w11045 , w11046 , w11047 , w11048 , w11049 , w11050 , w11051 , w11052 , w11053 , w11054 , w11055 , w11056 , w11057 , w11058 , w11059 , w11060 , w11061 , w11062 , w11063 , w11064 , w11065 , w11066 , w11067 , w11068 , w11069 , w11070 , w11071 , w11072 , w11073 , w11074 , w11075 , w11076 , w11077 , w11078 , w11079 , w11080 , w11081 , w11082 , w11083 , w11084 , w11085 , w11086 , w11087 , w11088 , w11089 , w11090 , w11091 , w11092 , w11093 , w11094 , w11095 , w11096 , w11097 , w11098 , w11099 , w11100 , w11101 , w11102 , w11103 , w11104 , w11105 , w11106 , w11107 , w11108 , w11109 , w11110 , w11111 , w11112 , w11113 , w11114 , w11115 , w11116 , w11117 , w11118 , w11119 , w11120 , w11121 , w11122 , w11123 , w11124 , w11125 , w11126 , w11127 , w11128 , w11129 , w11130 , w11131 , w11132 , w11133 , w11134 , w11135 , w11136 , w11137 , w11138 , w11139 , w11140 , w11141 , w11142 , w11143 , w11144 , w11145 , w11146 , w11147 , w11148 , w11149 , w11150 , w11151 , w11152 , w11153 , w11154 , w11155 , w11156 , w11157 , w11158 , w11159 , w11160 , w11161 , w11162 , w11163 , w11164 , w11165 , w11166 , w11167 , w11168 , w11169 , w11170 , w11171 , w11172 , w11173 , w11174 , w11175 , w11176 , w11177 , w11178 , w11179 , w11180 , w11181 , w11182 , w11183 , w11184 , w11185 , w11186 , w11187 , w11188 , w11189 , w11190 , w11191 , w11192 , w11193 , w11194 , w11195 , w11196 , w11197 , w11198 , w11199 , w11200 , w11201 , w11202 , w11203 , w11204 , w11205 , w11206 , w11207 , w11208 , w11209 , w11210 , w11211 , w11212 , w11213 , w11214 , w11215 , w11216 , w11217 , w11218 , w11219 , w11220 , w11221 , w11222 , w11223 , w11224 , w11225 , w11226 , w11227 , w11228 , w11229 , w11230 , w11231 , w11232 , w11233 , w11234 , w11235 , w11236 , w11237 , w11238 , w11239 , w11240 , w11241 , w11242 , w11243 , w11244 , w11245 , w11246 , w11247 , w11248 , w11249 , w11250 , w11251 , w11252 , w11253 , w11254 , w11255 , w11256 , w11257 , w11258 , w11259 , w11260 , w11261 , w11262 , w11263 , w11264 , w11265 , w11266 , w11267 , w11268 , w11269 , w11270 , w11271 , w11272 , w11273 , w11274 , w11275 , w11276 , w11277 , w11278 , w11279 , w11280 , w11281 , w11282 , w11283 , w11284 , w11285 , w11286 , w11287 , w11288 , w11289 , w11290 , w11291 , w11292 , w11293 , w11294 , w11295 , w11296 , w11297 , w11298 , w11299 , w11300 , w11301 , w11302 , w11303 , w11304 , w11305 , w11306 , w11307 , w11308 , w11309 , w11310 , w11311 , w11312 , w11313 , w11314 , w11315 , w11316 , w11317 , w11318 , w11319 , w11320 , w11321 , w11322 , w11323 , w11324 , w11325 , w11326 , w11327 , w11328 , w11329 , w11330 , w11331 , w11332 , w11333 , w11334 , w11335 , w11336 , w11337 , w11338 , w11339 , w11340 , w11341 , w11342 , w11343 , w11344 , w11345 , w11346 , w11347 , w11348 , w11349 , w11350 , w11351 , w11352 , w11353 , w11354 , w11355 , w11356 , w11357 , w11358 , w11359 , w11360 , w11361 , w11362 , w11363 , w11364 , w11365 , w11366 , w11367 , w11368 , w11369 , w11370 , w11371 , w11372 , w11373 , w11374 , w11375 , w11376 , w11377 , w11378 , w11379 , w11380 , w11381 , w11382 , w11383 , w11384 , w11385 , w11386 , w11387 , w11388 , w11389 , w11390 , w11391 , w11392 , w11393 , w11394 , w11395 , w11396 , w11397 , w11398 , w11399 , w11400 , w11401 , w11402 , w11403 , w11404 , w11405 , w11406 , w11407 , w11408 , w11409 , w11410 , w11411 , w11412 , w11413 , w11414 , w11415 , w11416 , w11417 , w11418 , w11419 , w11420 , w11421 , w11422 , w11423 , w11424 , w11425 , w11426 , w11427 , w11428 , w11429 , w11430 , w11431 , w11432 , w11433 , w11434 , w11435 , w11436 , w11437 , w11438 , w11439 , w11440 , w11441 , w11442 , w11443 , w11444 , w11445 , w11446 , w11447 , w11448 , w11449 , w11450 , w11451 , w11452 , w11453 , w11454 , w11455 , w11456 , w11457 , w11458 , w11459 , w11460 , w11461 , w11462 , w11463 , w11464 , w11465 , w11466 , w11467 , w11468 , w11469 , w11470 , w11471 , w11472 , w11473 , w11474 , w11475 , w11476 , w11477 , w11478 , w11479 , w11480 , w11481 , w11482 , w11483 , w11484 , w11485 , w11486 , w11487 , w11488 , w11489 , w11490 , w11491 , w11492 , w11493 , w11494 , w11495 , w11496 , w11497 , w11498 , w11499 , w11500 , w11501 , w11502 , w11503 , w11504 , w11505 , w11506 , w11507 , w11508 , w11509 , w11510 , w11511 , w11512 , w11513 , w11514 , w11515 , w11516 , w11517 , w11518 , w11519 , w11520 , w11521 , w11522 , w11523 , w11524 , w11525 , w11526 , w11527 , w11528 , w11529 , w11530 , w11531 , w11532 , w11533 , w11534 , w11535 , w11536 , w11537 , w11538 , w11539 , w11540 , w11541 , w11542 , w11543 , w11544 , w11545 , w11546 , w11547 , w11548 , w11549 , w11550 , w11551 , w11552 , w11553 , w11554 , w11555 , w11556 , w11557 , w11558 , w11559 , w11560 , w11561 , w11562 , w11563 , w11564 , w11565 , w11566 , w11567 , w11568 , w11569 , w11570 , w11571 , w11572 , w11573 , w11574 , w11575 , w11576 , w11577 , w11578 , w11579 , w11580 , w11581 , w11582 , w11583 , w11584 , w11585 , w11586 , w11587 , w11588 , w11589 , w11590 , w11591 , w11592 , w11593 , w11594 , w11595 , w11596 , w11597 , w11598 , w11599 , w11600 , w11601 , w11602 , w11603 , w11604 , w11605 , w11606 , w11607 , w11608 , w11609 , w11610 , w11611 , w11612 , w11613 , w11614 , w11615 , w11616 , w11617 , w11618 , w11619 , w11620 , w11621 , w11622 , w11623 , w11624 , w11625 , w11626 , w11627 , w11628 , w11629 , w11630 , w11631 , w11632 , w11633 , w11634 , w11635 , w11636 , w11637 , w11638 , w11639 , w11640 , w11641 , w11642 , w11643 , w11644 , w11645 , w11646 , w11647 , w11648 , w11649 , w11650 , w11651 , w11652 , w11653 , w11654 , w11655 , w11656 , w11657 , w11658 , w11659 , w11660 , w11661 , w11662 , w11663 , w11664 , w11665 , w11666 , w11667 , w11668 , w11669 , w11670 , w11671 , w11672 , w11673 , w11674 , w11675 , w11676 , w11677 , w11678 , w11679 , w11680 , w11681 , w11682 , w11683 , w11684 , w11685 , w11686 , w11687 , w11688 , w11689 , w11690 , w11691 , w11692 , w11693 , w11694 , w11695 , w11696 , w11697 , w11698 , w11699 , w11700 , w11701 , w11702 , w11703 , w11704 , w11705 , w11706 , w11707 , w11708 , w11709 , w11710 , w11711 , w11712 , w11713 , w11714 , w11715 , w11716 , w11717 , w11718 , w11719 , w11720 , w11721 , w11722 , w11723 , w11724 , w11725 , w11726 , w11727 , w11728 , w11729 , w11730 , w11731 , w11732 , w11733 , w11734 , w11735 , w11736 , w11737 , w11738 , w11739 , w11740 , w11741 , w11742 , w11743 , w11744 , w11745 , w11746 , w11747 , w11748 , w11749 , w11750 , w11751 , w11752 , w11753 , w11754 , w11755 , w11756 , w11757 , w11758 , w11759 , w11760 , w11761 , w11762 , w11763 , w11764 , w11765 , w11766 , w11767 , w11768 , w11769 , w11770 , w11771 , w11772 , w11773 , w11774 , w11775 , w11776 , w11777 , w11778 , w11779 , w11780 , w11781 , w11782 , w11783 , w11784 , w11785 , w11786 , w11787 , w11788 , w11789 , w11790 , w11791 , w11792 , w11793 , w11794 , w11795 , w11796 , w11797 , w11798 , w11799 , w11800 , w11801 , w11802 , w11803 , w11804 , w11805 , w11806 , w11807 , w11808 , w11809 , w11810 , w11811 , w11812 , w11813 , w11814 , w11815 , w11816 , w11817 , w11818 , w11819 , w11820 , w11821 , w11822 , w11823 , w11824 , w11825 , w11826 , w11827 , w11828 , w11829 , w11830 , w11831 , w11832 , w11833 , w11834 , w11835 , w11836 , w11837 , w11838 , w11839 , w11840 , w11841 , w11842 , w11843 , w11844 , w11845 , w11846 , w11847 , w11848 , w11849 , w11850 , w11851 , w11852 , w11853 , w11854 , w11855 , w11856 , w11857 , w11858 , w11859 , w11860 , w11861 , w11862 , w11863 , w11864 , w11865 , w11866 , w11867 , w11868 , w11869 , w11870 , w11871 , w11872 , w11873 , w11874 , w11875 , w11876 , w11877 , w11878 , w11879 , w11880 , w11881 , w11882 , w11883 , w11884 , w11885 , w11886 , w11887 , w11888 , w11889 , w11890 , w11891 , w11892 , w11893 , w11894 , w11895 , w11896 , w11897 , w11898 , w11899 , w11900 , w11901 , w11902 , w11903 , w11904 , w11905 , w11906 , w11907 , w11908 , w11909 , w11910 , w11911 , w11912 , w11913 , w11914 , w11915 , w11916 , w11917 , w11918 , w11919 , w11920 , w11921 , w11922 , w11923 , w11924 , w11925 , w11926 , w11927 , w11928 , w11929 , w11930 , w11931 , w11932 , w11933 , w11934 , w11935 , w11936 , w11937 , w11938 , w11939 , w11940 , w11941 , w11942 , w11943 , w11944 , w11945 , w11946 , w11947 , w11948 , w11949 , w11950 , w11951 , w11952 , w11953 , w11954 , w11955 , w11956 , w11957 , w11958 , w11959 , w11960 , w11961 , w11962 , w11963 , w11964 , w11965 , w11966 , w11967 , w11968 , w11969 , w11970 , w11971 , w11972 , w11973 , w11974 , w11975 , w11976 , w11977 , w11978 , w11979 , w11980 , w11981 , w11982 , w11983 , w11984 , w11985 , w11986 , w11987 , w11988 , w11989 , w11990 , w11991 , w11992 , w11993 , w11994 , w11995 , w11996 , w11997 , w11998 , w11999 , w12000 , w12001 , w12002 , w12003 , w12004 , w12005 , w12006 , w12007 , w12008 , w12009 , w12010 , w12011 , w12012 , w12013 , w12014 , w12015 , w12016 , w12017 , w12018 , w12019 , w12020 , w12021 , w12022 , w12023 , w12024 , w12025 , w12026 , w12027 , w12028 , w12029 , w12030 , w12031 , w12032 , w12033 , w12034 , w12035 , w12036 , w12037 , w12038 , w12039 , w12040 , w12041 , w12042 , w12043 , w12044 , w12045 , w12046 , w12047 , w12048 , w12049 , w12050 , w12051 , w12052 , w12053 , w12054 , w12055 , w12056 , w12057 , w12058 , w12059 , w12060 , w12061 , w12062 , w12063 , w12064 , w12065 , w12066 , w12067 , w12068 , w12069 , w12070 , w12071 , w12072 , w12073 , w12074 , w12075 , w12076 , w12077 , w12078 , w12079 , w12080 , w12081 , w12082 , w12083 , w12084 , w12085 , w12086 , w12087 , w12088 , w12089 , w12090 , w12091 , w12092 , w12093 , w12094 , w12095 , w12096 , w12097 , w12098 , w12099 , w12100 , w12101 , w12102 , w12103 , w12104 , w12105 , w12106 , w12107 , w12108 , w12109 , w12110 , w12111 , w12112 , w12113 , w12114 , w12115 , w12116 , w12117 , w12118 , w12119 , w12120 , w12121 , w12122 , w12123 , w12124 , w12125 , w12126 , w12127 , w12128 , w12129 , w12130 , w12131 , w12132 , w12133 , w12134 , w12135 , w12136 , w12137 , w12138 , w12139 , w12140 , w12141 , w12142 , w12143 , w12144 , w12145 , w12146 , w12147 , w12148 , w12149 , w12150 , w12151 , w12152 , w12153 , w12154 , w12155 , w12156 , w12157 , w12158 , w12159 , w12160 , w12161 , w12162 , w12163 , w12164 , w12165 , w12166 , w12167 , w12168 , w12169 , w12170 , w12171 , w12172 , w12173 , w12174 , w12175 , w12176 , w12177 , w12178 , w12179 , w12180 , w12181 , w12182 , w12183 , w12184 , w12185 , w12186 , w12187 , w12188 , w12189 , w12190 , w12191 , w12192 , w12193 , w12194 , w12195 , w12196 , w12197 , w12198 , w12199 , w12200 , w12201 , w12202 , w12203 , w12204 , w12205 , w12206 , w12207 , w12208 , w12209 , w12210 , w12211 , w12212 , w12213 , w12214 , w12215 , w12216 , w12217 , w12218 , w12219 , w12220 , w12221 , w12222 , w12223 , w12224 , w12225 , w12226 , w12227 , w12228 , w12229 , w12230 , w12231 , w12232 , w12233 , w12234 , w12235 , w12236 , w12237 , w12238 , w12239 , w12240 , w12241 , w12242 , w12243 , w12244 , w12245 , w12246 , w12247 , w12248 , w12249 , w12250 , w12251 , w12252 , w12253 , w12254 , w12255 , w12256 , w12257 , w12258 , w12259 , w12260 , w12261 , w12262 , w12263 , w12264 , w12265 , w12266 , w12267 , w12268 , w12269 , w12270 , w12271 , w12272 , w12273 , w12274 , w12275 , w12276 , w12277 , w12278 , w12279 , w12280 , w12281 , w12282 , w12283 , w12284 , w12285 , w12286 , w12287 , w12288 , w12289 , w12290 , w12291 , w12292 , w12293 , w12294 , w12295 , w12296 , w12297 , w12298 , w12299 , w12300 , w12301 , w12302 , w12303 , w12304 , w12305 , w12306 , w12307 , w12308 , w12309 , w12310 , w12311 , w12312 , w12313 , w12314 , w12315 , w12316 , w12317 , w12318 , w12319 , w12320 , w12321 , w12322 , w12323 , w12324 , w12325 , w12326 , w12327 , w12328 , w12329 , w12330 , w12331 , w12332 , w12333 , w12334 , w12335 , w12336 , w12337 , w12338 , w12339 , w12340 , w12341 , w12342 , w12343 , w12344 , w12345 , w12346 , w12347 , w12348 , w12349 , w12350 , w12351 , w12352 , w12353 , w12354 , w12355 , w12356 , w12357 , w12358 , w12359 , w12360 , w12361 , w12362 , w12363 , w12364 , w12365 , w12366 , w12367 , w12368 , w12369 , w12370 , w12371 , w12372 , w12373 , w12374 , w12375 , w12376 , w12377 , w12378 , w12379 , w12380 , w12381 , w12382 , w12383 , w12384 , w12385 , w12386 , w12387 , w12388 , w12389 , w12390 , w12391 , w12392 , w12393 , w12394 , w12395 , w12396 , w12397 , w12398 , w12399 , w12400 , w12401 , w12402 , w12403 , w12404 , w12405 , w12406 , w12407 , w12408 , w12409 , w12410 , w12411 , w12412 , w12413 , w12414 , w12415 , w12416 , w12417 , w12418 , w12419 , w12420 , w12421 , w12422 , w12423 , w12424 , w12425 , w12426 , w12427 , w12428 , w12429 , w12430 , w12431 , w12432 , w12433 , w12434 , w12435 , w12436 , w12437 , w12438 , w12439 , w12440 , w12441 , w12442 , w12443 , w12444 , w12445 , w12446 , w12447 , w12448 , w12449 , w12450 , w12451 , w12452 , w12453 , w12454 , w12455 , w12456 , w12457 , w12458 , w12459 , w12460 , w12461 , w12462 , w12463 , w12464 , w12465 , w12466 , w12467 , w12468 , w12469 , w12470 , w12471 , w12472 , w12473 , w12474 , w12475 , w12476 , w12477 , w12478 , w12479 , w12480 , w12481 , w12482 , w12483 , w12484 , w12485 , w12486 , w12487 , w12488 , w12489 , w12490 , w12491 , w12492 , w12493 , w12494 , w12495 , w12496 , w12497 , w12498 , w12499 , w12500 , w12501 , w12502 , w12503 , w12504 , w12505 , w12506 , w12507 , w12508 , w12509 , w12510 , w12511 , w12512 , w12513 , w12514 , w12515 , w12516 , w12517 , w12518 , w12519 , w12520 , w12521 , w12522 , w12523 , w12524 , w12525 , w12526 , w12527 , w12528 , w12529 , w12530 , w12531 , w12532 , w12533 , w12534 , w12535 , w12536 , w12537 , w12538 , w12539 , w12540 , w12541 , w12542 , w12543 , w12544 , w12545 , w12546 , w12547 , w12548 , w12549 , w12550 , w12551 , w12552 , w12553 , w12554 , w12555 , w12556 , w12557 , w12558 , w12559 , w12560 , w12561 , w12562 , w12563 , w12564 , w12565 , w12566 , w12567 , w12568 , w12569 , w12570 , w12571 , w12572 , w12573 , w12574 , w12575 , w12576 , w12577 , w12578 , w12579 , w12580 , w12581 , w12582 , w12583 , w12584 , w12585 , w12586 , w12587 , w12588 , w12589 , w12590 , w12591 , w12592 , w12593 , w12594 , w12595 , w12596 , w12597 , w12598 , w12599 , w12600 , w12601 , w12602 , w12603 , w12604 , w12605 , w12606 , w12607 , w12608 , w12609 , w12610 , w12611 , w12612 , w12613 , w12614 , w12615 , w12616 , w12617 , w12618 , w12619 , w12620 , w12621 , w12622 , w12623 , w12624 , w12625 , w12626 , w12627 , w12628 , w12629 , w12630 , w12631 , w12632 , w12633 , w12634 , w12635 , w12636 , w12637 , w12638 , w12639 , w12640 , w12641 , w12642 , w12643 , w12644 , w12645 , w12646 , w12647 , w12648 , w12649 , w12650 , w12651 , w12652 , w12653 , w12654 , w12655 , w12656 , w12657 , w12658 , w12659 , w12660 , w12661 , w12662 , w12663 , w12664 , w12665 , w12666 , w12667 , w12668 , w12669 , w12670 , w12671 , w12672 , w12673 , w12674 , w12675 , w12676 , w12677 , w12678 , w12679 , w12680 , w12681 , w12682 , w12683 , w12684 , w12685 , w12686 , w12687 , w12688 , w12689 , w12690 , w12691 , w12692 , w12693 , w12694 , w12695 , w12696 , w12697 , w12698 , w12699 , w12700 , w12701 , w12702 , w12703 , w12704 , w12705 , w12706 , w12707 , w12708 , w12709 , w12710 , w12711 , w12712 , w12713 , w12714 , w12715 , w12716 , w12717 , w12718 , w12719 , w12720 , w12721 , w12722 , w12723 , w12724 , w12725 , w12726 , w12727 , w12728 , w12729 , w12730 , w12731 , w12732 , w12733 , w12734 , w12735 , w12736 , w12737 , w12738 , w12739 , w12740 , w12741 , w12742 , w12743 , w12744 , w12745 , w12746 , w12747 , w12748 , w12749 , w12750 , w12751 , w12752 , w12753 , w12754 , w12755 , w12756 , w12757 , w12758 , w12759 , w12760 , w12761 , w12762 , w12763 , w12764 , w12765 , w12766 , w12767 , w12768 , w12769 , w12770 , w12771 , w12772 , w12773 , w12774 , w12775 , w12776 , w12777 , w12778 , w12779 , w12780 , w12781 , w12782 , w12783 , w12784 , w12785 , w12786 , w12787 , w12788 , w12789 , w12790 , w12791 , w12792 , w12793 , w12794 , w12795 , w12796 , w12797 , w12798 , w12799 , w12800 , w12801 , w12802 , w12803 , w12804 , w12805 , w12806 , w12807 , w12808 , w12809 , w12810 , w12811 , w12812 , w12813 , w12814 , w12815 , w12816 , w12817 , w12818 , w12819 , w12820 , w12821 , w12822 , w12823 , w12824 , w12825 , w12826 , w12827 , w12828 , w12829 , w12830 , w12831 , w12832 , w12833 , w12834 , w12835 , w12836 , w12837 , w12838 , w12839 , w12840 , w12841 , w12842 , w12843 , w12844 , w12845 , w12846 , w12847 , w12848 , w12849 , w12850 , w12851 , w12852 , w12853 , w12854 , w12855 , w12856 , w12857 , w12858 , w12859 , w12860 , w12861 , w12862 , w12863 , w12864 , w12865 , w12866 , w12867 , w12868 , w12869 , w12870 , w12871 , w12872 , w12873 , w12874 , w12875 , w12876 , w12877 , w12878 , w12879 , w12880 , w12881 , w12882 , w12883 , w12884 , w12885 , w12886 , w12887 , w12888 , w12889 , w12890 , w12891 , w12892 , w12893 , w12894 , w12895 , w12896 , w12897 , w12898 , w12899 , w12900 , w12901 , w12902 , w12903 , w12904 , w12905 , w12906 , w12907 , w12908 , w12909 , w12910 , w12911 , w12912 , w12913 , w12914 , w12915 , w12916 , w12917 , w12918 , w12919 , w12920 , w12921 , w12922 , w12923 , w12924 , w12925 , w12926 , w12927 , w12928 , w12929 , w12930 , w12931 , w12932 , w12933 , w12934 , w12935 , w12936 , w12937 , w12938 , w12939 , w12940 , w12941 , w12942 , w12943 , w12944 , w12945 , w12946 , w12947 , w12948 , w12949 , w12950 , w12951 , w12952 , w12953 , w12954 , w12955 , w12956 , w12957 , w12958 , w12959 , w12960 , w12961 , w12962 , w12963 , w12964 , w12965 , w12966 , w12967 , w12968 , w12969 , w12970 , w12971 , w12972 , w12973 , w12974 , w12975 , w12976 , w12977 , w12978 , w12979 , w12980 , w12981 , w12982 , w12983 , w12984 , w12985 , w12986 , w12987 , w12988 , w12989 , w12990 , w12991 , w12992 , w12993 , w12994 , w12995 , w12996 , w12997 , w12998 , w12999 , w13000 , w13001 , w13002 , w13003 , w13004 , w13005 , w13006 , w13007 , w13008 , w13009 , w13010 , w13011 , w13012 , w13013 , w13014 , w13015 , w13016 , w13017 , w13018 , w13019 , w13020 , w13021 , w13022 , w13023 , w13024 , w13025 , w13026 , w13027 , w13028 , w13029 , w13030 , w13031 , w13032 , w13033 , w13034 , w13035 , w13036 , w13037 , w13038 , w13039 , w13040 , w13041 , w13042 , w13043 , w13044 , w13045 , w13046 , w13047 , w13048 , w13049 , w13050 , w13051 , w13052 , w13053 , w13054 , w13055 , w13056 , w13057 , w13058 , w13059 , w13060 , w13061 , w13062 , w13063 , w13064 , w13065 , w13066 , w13067 , w13068 , w13069 , w13070 , w13071 , w13072 , w13073 , w13074 , w13075 , w13076 , w13077 , w13078 , w13079 , w13080 , w13081 , w13082 , w13083 , w13084 , w13085 , w13086 , w13087 , w13088 , w13089 , w13090 , w13091 , w13092 , w13093 , w13094 , w13095 , w13096 , w13097 , w13098 , w13099 , w13100 , w13101 , w13102 , w13103 , w13104 , w13105 , w13106 , w13107 , w13108 , w13109 , w13110 , w13111 , w13112 , w13113 , w13114 , w13115 , w13116 , w13117 , w13118 , w13119 , w13120 , w13121 , w13122 , w13123 , w13124 , w13125 , w13126 , w13127 , w13128 , w13129 , w13130 , w13131 , w13132 , w13133 , w13134 , w13135 , w13136 , w13137 , w13138 , w13139 , w13140 , w13141 , w13142 , w13143 , w13144 , w13145 , w13146 , w13147 , w13148 , w13149 , w13150 , w13151 , w13152 , w13153 , w13154 , w13155 , w13156 , w13157 , w13158 , w13159 , w13160 , w13161 , w13162 , w13163 , w13164 , w13165 , w13166 , w13167 , w13168 , w13169 , w13170 , w13171 , w13172 , w13173 , w13174 , w13175 , w13176 , w13177 , w13178 , w13179 , w13180 , w13181 , w13182 , w13183 , w13184 , w13185 , w13186 , w13187 , w13188 , w13189 , w13190 , w13191 , w13192 , w13193 , w13194 , w13195 , w13196 , w13197 , w13198 , w13199 , w13200 , w13201 , w13202 , w13203 , w13204 , w13205 , w13206 , w13207 , w13208 , w13209 , w13210 , w13211 , w13212 , w13213 , w13214 , w13215 , w13216 , w13217 , w13218 , w13219 , w13220 , w13221 , w13222 , w13223 , w13224 , w13225 , w13226 , w13227 , w13228 , w13229 , w13230 , w13231 , w13232 , w13233 , w13234 , w13235 , w13236 , w13237 , w13238 , w13239 , w13240 , w13241 , w13242 , w13243 , w13244 , w13245 , w13246 , w13247 , w13248 , w13249 , w13250 , w13251 , w13252 , w13253 , w13254 , w13255 , w13256 , w13257 , w13258 , w13259 , w13260 , w13261 , w13262 , w13263 , w13264 , w13265 , w13266 , w13267 , w13268 , w13269 , w13270 , w13271 , w13272 , w13273 , w13274 , w13275 , w13276 , w13277 , w13278 , w13279 , w13280 , w13281 , w13282 , w13283 , w13284 , w13285 , w13286 , w13287 , w13288 , w13289 , w13290 , w13291 , w13292 , w13293 , w13294 , w13295 , w13296 , w13297 , w13298 , w13299 , w13300 , w13301 , w13302 , w13303 , w13304 , w13305 , w13306 , w13307 , w13308 , w13309 , w13310 , w13311 , w13312 , w13313 , w13314 , w13315 , w13316 , w13317 , w13318 , w13319 , w13320 , w13321 , w13322 , w13323 , w13324 , w13325 , w13326 , w13327 , w13328 , w13329 , w13330 , w13331 , w13332 , w13333 , w13334 , w13335 , w13336 , w13337 , w13338 , w13339 , w13340 , w13341 , w13342 , w13343 , w13344 , w13345 , w13346 , w13347 , w13348 , w13349 , w13350 , w13351 , w13352 , w13353 , w13354 , w13355 , w13356 , w13357 , w13358 , w13359 , w13360 , w13361 , w13362 , w13363 , w13364 , w13365 , w13366 , w13367 , w13368 , w13369 , w13370 , w13371 , w13372 , w13373 , w13374 , w13375 , w13376 , w13377 , w13378 , w13379 , w13380 , w13381 , w13382 , w13383 , w13384 , w13385 , w13386 , w13387 , w13388 , w13389 , w13390 , w13391 , w13392 , w13393 , w13394 , w13395 , w13396 , w13397 , w13398 , w13399 , w13400 , w13401 , w13402 , w13403 , w13404 , w13405 , w13406 , w13407 , w13408 , w13409 , w13410 , w13411 , w13412 , w13413 , w13414 , w13415 , w13416 , w13417 , w13418 , w13419 , w13420 , w13421 , w13422 , w13423 , w13424 , w13425 , w13426 , w13427 , w13428 , w13429 , w13430 , w13431 , w13432 , w13433 , w13434 , w13435 , w13436 , w13437 , w13438 , w13439 , w13440 , w13441 , w13442 , w13443 , w13444 , w13445 , w13446 , w13447 , w13448 , w13449 , w13450 , w13451 , w13452 , w13453 , w13454 , w13455 , w13456 , w13457 , w13458 , w13459 , w13460 , w13461 , w13462 , w13463 , w13464 , w13465 , w13466 , w13467 , w13468 , w13469 , w13470 , w13471 , w13472 , w13473 , w13474 , w13475 , w13476 , w13477 , w13478 , w13479 , w13480 , w13481 , w13482 , w13483 , w13484 , w13485 , w13486 , w13487 , w13488 , w13489 , w13490 , w13491 , w13492 , w13493 , w13494 , w13495 , w13496 , w13497 , w13498 , w13499 , w13500 , w13501 , w13502 , w13503 , w13504 , w13505 , w13506 , w13507 , w13508 , w13509 , w13510 , w13511 , w13512 , w13513 , w13514 , w13515 , w13516 , w13517 , w13518 , w13519 , w13520 , w13521 , w13522 , w13523 , w13524 , w13525 , w13526 , w13527 , w13528 , w13529 , w13530 , w13531 , w13532 , w13533 , w13534 , w13535 , w13536 , w13537 , w13538 , w13539 , w13540 , w13541 , w13542 , w13543 , w13544 , w13545 , w13546 , w13547 , w13548 , w13549 , w13550 , w13551 , w13552 , w13553 , w13554 , w13555 , w13556 , w13557 , w13558 , w13559 , w13560 , w13561 , w13562 , w13563 , w13564 , w13565 , w13566 , w13567 , w13568 , w13569 , w13570 , w13571 , w13572 , w13573 , w13574 , w13575 , w13576 , w13577 , w13578 , w13579 , w13580 , w13581 , w13582 , w13583 , w13584 , w13585 , w13586 , w13587 , w13588 , w13589 , w13590 , w13591 , w13592 , w13593 , w13594 , w13595 , w13596 , w13597 , w13598 , w13599 , w13600 , w13601 , w13602 , w13603 , w13604 , w13605 , w13606 , w13607 , w13608 , w13609 , w13610 , w13611 , w13612 , w13613 , w13614 , w13615 , w13616 , w13617 , w13618 , w13619 , w13620 , w13621 , w13622 , w13623 , w13624 , w13625 , w13626 , w13627 , w13628 , w13629 , w13630 , w13631 , w13632 , w13633 , w13634 , w13635 , w13636 , w13637 , w13638 , w13639 , w13640 , w13641 , w13642 , w13643 , w13644 , w13645 , w13646 , w13647 , w13648 , w13649 , w13650 , w13651 , w13652 , w13653 , w13654 , w13655 , w13656 , w13657 , w13658 , w13659 , w13660 , w13661 , w13662 , w13663 , w13664 , w13665 , w13666 , w13667 , w13668 , w13669 , w13670 , w13671 , w13672 , w13673 , w13674 , w13675 , w13676 , w13677 , w13678 , w13679 , w13680 , w13681 , w13682 , w13683 , w13684 , w13685 , w13686 , w13687 , w13688 , w13689 , w13690 , w13691 , w13692 , w13693 , w13694 , w13695 , w13696 , w13697 , w13698 , w13699 , w13700 , w13701 , w13702 , w13703 , w13704 , w13705 , w13706 , w13707 , w13708 , w13709 , w13710 , w13711 , w13712 , w13713 , w13714 , w13715 , w13716 , w13717 , w13718 , w13719 , w13720 , w13721 , w13722 , w13723 , w13724 , w13725 , w13726 , w13727 , w13728 , w13729 , w13730 , w13731 , w13732 , w13733 , w13734 , w13735 , w13736 , w13737 , w13738 , w13739 , w13740 , w13741 , w13742 , w13743 , w13744 , w13745 , w13746 , w13747 , w13748 , w13749 , w13750 , w13751 , w13752 , w13753 , w13754 , w13755 , w13756 , w13757 , w13758 , w13759 , w13760 , w13761 , w13762 , w13763 , w13764 , w13765 , w13766 , w13767 , w13768 , w13769 , w13770 , w13771 , w13772 , w13773 , w13774 , w13775 , w13776 , w13777 , w13778 , w13779 , w13780 , w13781 , w13782 , w13783 , w13784 , w13785 , w13786 , w13787 , w13788 , w13789 , w13790 , w13791 , w13792 , w13793 , w13794 , w13795 , w13796 , w13797 , w13798 , w13799 , w13800 , w13801 , w13802 , w13803 , w13804 , w13805 , w13806 , w13807 , w13808 , w13809 , w13810 , w13811 , w13812 , w13813 , w13814 , w13815 , w13816 , w13817 , w13818 , w13819 , w13820 , w13821 , w13822 , w13823 , w13824 , w13825 , w13826 , w13827 , w13828 , w13829 , w13830 , w13831 , w13832 , w13833 , w13834 , w13835 , w13836 , w13837 , w13838 , w13839 , w13840 , w13841 , w13842 , w13843 , w13844 , w13845 , w13846 , w13847 , w13848 , w13849 , w13850 , w13851 , w13852 , w13853 , w13854 , w13855 , w13856 , w13857 , w13858 , w13859 , w13860 , w13861 , w13862 , w13863 , w13864 , w13865 , w13866 , w13867 , w13868 , w13869 , w13870 , w13871 , w13872 , w13873 , w13874 , w13875 , w13876 , w13877 , w13878 , w13879 , w13880 , w13881 , w13882 , w13883 , w13884 , w13885 , w13886 , w13887 , w13888 , w13889 , w13890 , w13891 , w13892 , w13893 , w13894 , w13895 , w13896 , w13897 , w13898 , w13899 , w13900 , w13901 , w13902 , w13903 , w13904 , w13905 , w13906 , w13907 , w13908 , w13909 , w13910 , w13911 , w13912 , w13913 , w13914 , w13915 , w13916 , w13917 , w13918 , w13919 , w13920 , w13921 , w13922 , w13923 , w13924 , w13925 , w13926 , w13927 , w13928 , w13929 , w13930 , w13931 , w13932 , w13933 , w13934 , w13935 , w13936 , w13937 , w13938 , w13939 , w13940 , w13941 , w13942 , w13943 , w13944 , w13945 , w13946 , w13947 , w13948 , w13949 , w13950 , w13951 , w13952 , w13953 , w13954 , w13955 , w13956 , w13957 , w13958 , w13959 , w13960 , w13961 , w13962 , w13963 , w13964 , w13965 , w13966 , w13967 , w13968 , w13969 , w13970 , w13971 , w13972 , w13973 , w13974 , w13975 , w13976 , w13977 , w13978 , w13979 , w13980 , w13981 , w13982 , w13983 , w13984 , w13985 , w13986 , w13987 , w13988 , w13989 , w13990 , w13991 , w13992 , w13993 , w13994 , w13995 , w13996 , w13997 , w13998 , w13999 , w14000 , w14001 , w14002 , w14003 , w14004 , w14005 , w14006 , w14007 , w14008 , w14009 , w14010 , w14011 , w14012 , w14013 , w14014 , w14015 , w14016 , w14017 , w14018 , w14019 , w14020 , w14021 , w14022 , w14023 , w14024 , w14025 , w14026 , w14027 , w14028 , w14029 , w14030 , w14031 , w14032 , w14033 , w14034 , w14035 , w14036 , w14037 , w14038 , w14039 , w14040 , w14041 , w14042 , w14043 , w14044 , w14045 , w14046 , w14047 , w14048 , w14049 , w14050 , w14051 , w14052 , w14053 , w14054 , w14055 , w14056 , w14057 , w14058 , w14059 , w14060 , w14061 , w14062 , w14063 , w14064 , w14065 , w14066 , w14067 , w14068 , w14069 , w14070 , w14071 , w14072 , w14073 , w14074 , w14075 , w14076 , w14077 , w14078 , w14079 , w14080 , w14081 , w14082 , w14083 , w14084 , w14085 , w14086 , w14087 , w14088 , w14089 , w14090 , w14091 , w14092 , w14093 , w14094 , w14095 , w14096 , w14097 , w14098 , w14099 , w14100 , w14101 , w14102 , w14103 , w14104 , w14105 , w14106 , w14107 , w14108 , w14109 , w14110 , w14111 , w14112 , w14113 , w14114 , w14115 , w14116 , w14117 , w14118 , w14119 , w14120 , w14121 , w14122 , w14123 , w14124 , w14125 , w14126 , w14127 , w14128 , w14129 , w14130 , w14131 , w14132 , w14133 , w14134 , w14135 , w14136 , w14137 , w14138 , w14139 , w14140 , w14141 , w14142 , w14143 , w14144 , w14145 , w14146 , w14147 , w14148 , w14149 , w14150 , w14151 , w14152 , w14153 , w14154 , w14155 , w14156 , w14157 , w14158 , w14159 , w14160 , w14161 , w14162 , w14163 , w14164 , w14165 , w14166 , w14167 , w14168 , w14169 , w14170 , w14171 , w14172 , w14173 , w14174 , w14175 , w14176 , w14177 , w14178 , w14179 , w14180 , w14181 , w14182 , w14183 , w14184 , w14185 , w14186 , w14187 , w14188 , w14189 , w14190 , w14191 , w14192 , w14193 , w14194 , w14195 , w14196 , w14197 , w14198 , w14199 , w14200 , w14201 , w14202 , w14203 , w14204 , w14205 , w14206 , w14207 , w14208 , w14209 , w14210 , w14211 , w14212 , w14213 , w14214 , w14215 , w14216 , w14217 , w14218 , w14219 , w14220 , w14221 , w14222 , w14223 , w14224 , w14225 , w14226 , w14227 , w14228 , w14229 , w14230 , w14231 , w14232 , w14233 , w14234 , w14235 , w14236 , w14237 , w14238 , w14239 , w14240 , w14241 , w14242 , w14243 , w14244 , w14245 , w14246 , w14247 , w14248 , w14249 , w14250 , w14251 , w14252 , w14253 , w14254 , w14255 , w14256 , w14257 , w14258 , w14259 , w14260 , w14261 , w14262 , w14263 , w14264 , w14265 , w14266 , w14267 , w14268 , w14269 , w14270 , w14271 , w14272 , w14273 , w14274 , w14275 , w14276 , w14277 , w14278 , w14279 , w14280 , w14281 , w14282 , w14283 , w14284 , w14285 , w14286 , w14287 , w14288 , w14289 , w14290 , w14291 , w14292 , w14293 , w14294 , w14295 , w14296 , w14297 , w14298 , w14299 , w14300 , w14301 , w14302 , w14303 , w14304 , w14305 , w14306 , w14307 , w14308 , w14309 , w14310 , w14311 , w14312 , w14313 , w14314 , w14315 , w14316 , w14317 , w14318 , w14319 , w14320 , w14321 , w14322 , w14323 , w14324 , w14325 , w14326 , w14327 , w14328 , w14329 , w14330 , w14331 , w14332 , w14333 , w14334 , w14335 , w14336 , w14337 , w14338 , w14339 , w14340 , w14341 , w14342 , w14343 , w14344 , w14345 , w14346 , w14347 , w14348 , w14349 , w14350 , w14351 , w14352 , w14353 , w14354 , w14355 , w14356 , w14357 , w14358 , w14359 , w14360 , w14361 , w14362 , w14363 , w14364 , w14365 , w14366 , w14367 , w14368 , w14369 , w14370 , w14371 , w14372 , w14373 , w14374 , w14375 , w14376 , w14377 , w14378 , w14379 , w14380 , w14381 , w14382 , w14383 , w14384 , w14385 , w14386 , w14387 , w14388 , w14389 , w14390 , w14391 , w14392 , w14393 , w14394 , w14395 , w14396 , w14397 , w14398 , w14399 , w14400 , w14401 , w14402 , w14403 , w14404 , w14405 , w14406 , w14407 , w14408 , w14409 , w14410 , w14411 , w14412 , w14413 , w14414 , w14415 , w14416 , w14417 , w14418 , w14419 , w14420 , w14421 , w14422 , w14423 , w14424 , w14425 , w14426 , w14427 , w14428 , w14429 , w14430 , w14431 , w14432 , w14433 , w14434 , w14435 , w14436 , w14437 , w14438 , w14439 , w14440 , w14441 , w14442 , w14443 , w14444 , w14445 , w14446 , w14447 , w14448 , w14449 , w14450 , w14451 , w14452 , w14453 , w14454 , w14455 , w14456 , w14457 , w14458 , w14459 , w14460 , w14461 , w14462 , w14463 , w14464 , w14465 , w14466 , w14467 , w14468 , w14469 , w14470 , w14471 , w14472 , w14473 , w14474 , w14475 , w14476 , w14477 , w14478 , w14479 , w14480 , w14481 , w14482 , w14483 , w14484 , w14485 , w14486 , w14487 , w14488 , w14489 , w14490 , w14491 , w14492 , w14493 , w14494 , w14495 , w14496 , w14497 , w14498 , w14499 , w14500 , w14501 , w14502 , w14503 , w14504 , w14505 , w14506 , w14507 , w14508 , w14509 , w14510 , w14511 , w14512 , w14513 , w14514 , w14515 , w14516 , w14517 , w14518 , w14519 , w14520 , w14521 , w14522 , w14523 , w14524 , w14525 , w14526 , w14527 , w14528 , w14529 , w14530 , w14531 , w14532 , w14533 , w14534 , w14535 , w14536 , w14537 , w14538 , w14539 , w14540 , w14541 , w14542 , w14543 , w14544 , w14545 , w14546 , w14547 , w14548 , w14549 , w14550 , w14551 , w14552 , w14553 , w14554 , w14555 , w14556 , w14557 , w14558 , w14559 , w14560 , w14561 , w14562 , w14563 , w14564 , w14565 , w14566 , w14567 , w14568 , w14569 , w14570 , w14571 , w14572 , w14573 , w14574 , w14575 , w14576 , w14577 , w14578 , w14579 , w14580 , w14581 , w14582 , w14583 , w14584 , w14585 , w14586 , w14587 , w14588 , w14589 , w14590 , w14591 , w14592 , w14593 , w14594 , w14595 , w14596 , w14597 , w14598 , w14599 , w14600 , w14601 , w14602 , w14603 , w14604 , w14605 , w14606 , w14607 , w14608 , w14609 , w14610 , w14611 , w14612 , w14613 , w14614 , w14615 , w14616 , w14617 , w14618 , w14619 , w14620 , w14621 , w14622 , w14623 , w14624 , w14625 , w14626 , w14627 , w14628 , w14629 , w14630 , w14631 , w14632 , w14633 , w14634 , w14635 , w14636 , w14637 , w14638 , w14639 , w14640 , w14641 , w14642 , w14643 , w14644 , w14645 , w14646 , w14647 , w14648 , w14649 , w14650 , w14651 , w14652 , w14653 , w14654 , w14655 , w14656 , w14657 , w14658 , w14659 , w14660 , w14661 , w14662 , w14663 , w14664 , w14665 , w14666 , w14667 , w14668 , w14669 , w14670 , w14671 , w14672 , w14673 , w14674 , w14675 , w14676 , w14677 , w14678 , w14679 , w14680 , w14681 , w14682 , w14683 , w14684 , w14685 , w14686 , w14687 , w14688 , w14689 , w14690 , w14691 , w14692 , w14693 , w14694 , w14695 , w14696 , w14697 , w14698 , w14699 , w14700 , w14701 , w14702 , w14703 , w14704 , w14705 , w14706 , w14707 , w14708 , w14709 , w14710 , w14711 , w14712 , w14713 , w14714 , w14715 , w14716 , w14717 , w14718 , w14719 , w14720 , w14721 , w14722 , w14723 , w14724 , w14725 , w14726 , w14727 , w14728 , w14729 , w14730 , w14731 , w14732 , w14733 , w14734 , w14735 , w14736 , w14737 , w14738 , w14739 , w14740 , w14741 , w14742 , w14743 , w14744 , w14745 , w14746 , w14747 , w14748 , w14749 , w14750 , w14751 , w14752 , w14753 , w14754 , w14755 , w14756 , w14757 , w14758 , w14759 , w14760 , w14761 , w14762 , w14763 , w14764 , w14765 , w14766 , w14767 , w14768 , w14769 , w14770 , w14771 , w14772 , w14773 , w14774 , w14775 , w14776 , w14777 , w14778 , w14779 , w14780 , w14781 , w14782 , w14783 , w14784 , w14785 , w14786 , w14787 , w14788 , w14789 , w14790 , w14791 , w14792 , w14793 , w14794 , w14795 , w14796 , w14797 , w14798 , w14799 , w14800 , w14801 , w14802 , w14803 , w14804 , w14805 , w14806 , w14807 , w14808 , w14809 , w14810 , w14811 , w14812 , w14813 , w14814 , w14815 , w14816 , w14817 , w14818 , w14819 , w14820 , w14821 , w14822 , w14823 , w14824 , w14825 , w14826 , w14827 , w14828 , w14829 , w14830 , w14831 , w14832 , w14833 , w14834 , w14835 , w14836 , w14837 , w14838 , w14839 , w14840 , w14841 , w14842 , w14843 , w14844 , w14845 , w14846 , w14847 , w14848 , w14849 , w14850 , w14851 , w14852 , w14853 , w14854 , w14855 , w14856 , w14857 , w14858 , w14859 , w14860 , w14861 , w14862 , w14863 , w14864 , w14865 , w14866 , w14867 , w14868 , w14869 , w14870 , w14871 , w14872 , w14873 , w14874 , w14875 , w14876 , w14877 , w14878 , w14879 , w14880 , w14881 , w14882 , w14883 , w14884 , w14885 , w14886 , w14887 , w14888 , w14889 , w14890 , w14891 , w14892 , w14893 , w14894 , w14895 , w14896 , w14897 , w14898 , w14899 , w14900 , w14901 , w14902 , w14903 , w14904 , w14905 , w14906 , w14907 , w14908 , w14909 , w14910 , w14911 , w14912 , w14913 , w14914 , w14915 , w14916 , w14917 , w14918 , w14919 , w14920 , w14921 , w14922 , w14923 , w14924 , w14925 , w14926 , w14927 , w14928 , w14929 , w14930 , w14931 , w14932 , w14933 , w14934 , w14935 , w14936 , w14937 , w14938 , w14939 , w14940 , w14941 , w14942 , w14943 , w14944 , w14945 , w14946 , w14947 , w14948 , w14949 , w14950 , w14951 , w14952 , w14953 , w14954 , w14955 , w14956 , w14957 , w14958 , w14959 , w14960 , w14961 , w14962 , w14963 , w14964 , w14965 , w14966 , w14967 , w14968 , w14969 , w14970 , w14971 , w14972 , w14973 , w14974 , w14975 , w14976 , w14977 , w14978 , w14979 , w14980 , w14981 , w14982 , w14983 , w14984 , w14985 , w14986 , w14987 , w14988 , w14989 , w14990 , w14991 , w14992 , w14993 , w14994 , w14995 , w14996 , w14997 , w14998 , w14999 , w15000 , w15001 , w15002 , w15003 , w15004 , w15005 , w15006 , w15007 , w15008 , w15009 , w15010 , w15011 , w15012 , w15013 , w15014 , w15015 , w15016 , w15017 , w15018 , w15019 , w15020 , w15021 , w15022 , w15023 , w15024 , w15025 , w15026 , w15027 , w15028 , w15029 , w15030 , w15031 , w15032 , w15033 , w15034 , w15035 , w15036 , w15037 , w15038 , w15039 , w15040 , w15041 , w15042 , w15043 , w15044 , w15045 , w15046 , w15047 , w15048 , w15049 , w15050 , w15051 , w15052 , w15053 , w15054 , w15055 , w15056 , w15057 , w15058 , w15059 , w15060 , w15061 , w15062 , w15063 , w15064 , w15065 , w15066 , w15067 , w15068 , w15069 , w15070 , w15071 , w15072 , w15073 , w15074 , w15075 , w15076 , w15077 , w15078 , w15079 , w15080 , w15081 , w15082 , w15083 , w15084 , w15085 , w15086 , w15087 , w15088 , w15089 , w15090 , w15091 , w15092 , w15093 , w15094 , w15095 , w15096 , w15097 , w15098 , w15099 , w15100 , w15101 , w15102 , w15103 , w15104 , w15105 , w15106 , w15107 , w15108 , w15109 , w15110 , w15111 , w15112 , w15113 , w15114 , w15115 , w15116 , w15117 , w15118 , w15119 , w15120 , w15121 , w15122 , w15123 , w15124 , w15125 , w15126 , w15127 , w15128 , w15129 , w15130 , w15131 , w15132 , w15133 , w15134 , w15135 , w15136 , w15137 , w15138 , w15139 , w15140 , w15141 , w15142 , w15143 , w15144 , w15145 , w15146 , w15147 , w15148 , w15149 , w15150 , w15151 , w15152 , w15153 , w15154 , w15155 , w15156 , w15157 , w15158 , w15159 , w15160 , w15161 , w15162 , w15163 , w15164 , w15165 , w15166 , w15167 , w15168 , w15169 , w15170 , w15171 , w15172 , w15173 , w15174 , w15175 , w15176 , w15177 , w15178 , w15179 , w15180 , w15181 , w15182 , w15183 , w15184 , w15185 , w15186 , w15187 , w15188 , w15189 , w15190 , w15191 , w15192 , w15193 , w15194 , w15195 , w15196 , w15197 , w15198 , w15199 , w15200 , w15201 , w15202 , w15203 , w15204 , w15205 , w15206 , w15207 , w15208 , w15209 , w15210 , w15211 , w15212 , w15213 , w15214 , w15215 , w15216 , w15217 , w15218 , w15219 , w15220 , w15221 , w15222 , w15223 , w15224 , w15225 , w15226 , w15227 , w15228 , w15229 , w15230 , w15231 , w15232 , w15233 , w15234 , w15235 , w15236 , w15237 , w15238 , w15239 , w15240 , w15241 , w15242 , w15243 , w15244 , w15245 , w15246 , w15247 , w15248 , w15249 , w15250 , w15251 , w15252 , w15253 , w15254 , w15255 , w15256 , w15257 , w15258 , w15259 , w15260 , w15261 , w15262 , w15263 , w15264 , w15265 , w15266 , w15267 , w15268 , w15269 , w15270 , w15271 , w15272 , w15273 , w15274 , w15275 , w15276 , w15277 , w15278 , w15279 , w15280 , w15281 , w15282 , w15283 , w15284 , w15285 , w15286 , w15287 , w15288 , w15289 , w15290 , w15291 , w15292 , w15293 , w15294 , w15295 , w15296 , w15297 , w15298 , w15299 , w15300 , w15301 , w15302 , w15303 , w15304 , w15305 , w15306 , w15307 , w15308 , w15309 , w15310 , w15311 , w15312 , w15313 , w15314 , w15315 , w15316 , w15317 , w15318 , w15319 , w15320 , w15321 , w15322 , w15323 , w15324 , w15325 , w15326 , w15327 , w15328 , w15329 , w15330 , w15331 , w15332 , w15333 , w15334 , w15335 , w15336 , w15337 , w15338 , w15339 , w15340 , w15341 , w15342 , w15343 , w15344 , w15345 , w15346 , w15347 , w15348 , w15349 , w15350 , w15351 , w15352 , w15353 , w15354 , w15355 , w15356 , w15357 , w15358 , w15359 , w15360 , w15361 , w15362 , w15363 , w15364 , w15365 , w15366 , w15367 , w15368 , w15369 , w15370 , w15371 , w15372 , w15373 , w15374 , w15375 , w15376 , w15377 , w15378 , w15379 , w15380 , w15381 , w15382 , w15383 , w15384 , w15385 , w15386 , w15387 , w15388 , w15389 , w15390 , w15391 , w15392 , w15393 , w15394 , w15395 , w15396 , w15397 , w15398 , w15399 , w15400 , w15401 , w15402 , w15403 , w15404 , w15405 , w15406 , w15407 , w15408 , w15409 , w15410 , w15411 , w15412 , w15413 , w15414 , w15415 , w15416 , w15417 , w15418 , w15419 , w15420 , w15421 , w15422 , w15423 , w15424 , w15425 , w15426 , w15427 , w15428 , w15429 , w15430 , w15431 , w15432 , w15433 , w15434 , w15435 , w15436 , w15437 , w15438 , w15439 , w15440 , w15441 , w15442 , w15443 , w15444 , w15445 , w15446 , w15447 , w15448 , w15449 , w15450 , w15451 , w15452 , w15453 , w15454 , w15455 , w15456 , w15457 , w15458 , w15459 , w15460 , w15461 , w15462 , w15463 , w15464 , w15465 , w15466 , w15467 , w15468 , w15469 , w15470 , w15471 , w15472 , w15473 , w15474 , w15475 , w15476 , w15477 , w15478 , w15479 , w15480 , w15481 , w15482 , w15483 , w15484 , w15485 , w15486 , w15487 , w15488 , w15489 , w15490 , w15491 , w15492 , w15493 , w15494 , w15495 , w15496 , w15497 , w15498 , w15499 , w15500 , w15501 , w15502 , w15503 , w15504 , w15505 , w15506 , w15507 , w15508 , w15509 , w15510 , w15511 , w15512 , w15513 , w15514 , w15515 , w15516 , w15517 , w15518 , w15519 , w15520 , w15521 , w15522 , w15523 , w15524 , w15525 , w15526 , w15527 , w15528 , w15529 , w15530 , w15531 , w15532 , w15533 , w15534 , w15535 , w15536 , w15537 , w15538 , w15539 , w15540 , w15541 , w15542 , w15543 , w15544 , w15545 , w15546 , w15547 , w15548 , w15549 , w15550 , w15551 , w15552 , w15553 , w15554 , w15555 , w15556 , w15557 , w15558 , w15559 , w15560 , w15561 , w15562 , w15563 , w15564 , w15565 , w15566 , w15567 , w15568 , w15569 , w15570 , w15571 , w15572 , w15573 , w15574 , w15575 , w15576 , w15577 , w15578 , w15579 , w15580 , w15581 , w15582 , w15583 , w15584 , w15585 , w15586 , w15587 , w15588 , w15589 , w15590 , w15591 , w15592 , w15593 , w15594 , w15595 , w15596 , w15597 , w15598 , w15599 , w15600 , w15601 , w15602 , w15603 , w15604 , w15605 , w15606 , w15607 , w15608 , w15609 , w15610 , w15611 , w15612 , w15613 , w15614 , w15615 , w15616 , w15617 , w15618 , w15619 , w15620 , w15621 , w15622 , w15623 , w15624 , w15625 , w15626 , w15627 , w15628 , w15629 , w15630 , w15631 , w15632 , w15633 , w15634 , w15635 , w15636 , w15637 , w15638 , w15639 , w15640 , w15641 , w15642 , w15643 , w15644 , w15645 , w15646 , w15647 , w15648 , w15649 , w15650 , w15651 , w15652 , w15653 , w15654 , w15655 , w15656 , w15657 , w15658 , w15659 , w15660 , w15661 , w15662 , w15663 , w15664 , w15665 , w15666 , w15667 , w15668 , w15669 , w15670 , w15671 , w15672 , w15673 , w15674 , w15675 , w15676 , w15677 , w15678 , w15679 , w15680 , w15681 , w15682 , w15683 , w15684 , w15685 , w15686 , w15687 , w15688 , w15689 , w15690 , w15691 , w15692 , w15693 , w15694 , w15695 , w15696 , w15697 , w15698 , w15699 , w15700 , w15701 , w15702 , w15703 , w15704 , w15705 , w15706 , w15707 , w15708 , w15709 , w15710 , w15711 , w15712 , w15713 , w15714 , w15715 , w15716 , w15717 , w15718 , w15719 , w15720 , w15721 , w15722 , w15723 , w15724 , w15725 , w15726 , w15727 , w15728 , w15729 , w15730 , w15731 , w15732 , w15733 , w15734 , w15735 , w15736 , w15737 , w15738 , w15739 , w15740 , w15741 , w15742 , w15743 , w15744 , w15745 , w15746 , w15747 , w15748 , w15749 , w15750 , w15751 , w15752 , w15753 , w15754 , w15755 , w15756 , w15757 , w15758 , w15759 , w15760 , w15761 , w15762 , w15763 , w15764 , w15765 , w15766 , w15767 , w15768 , w15769 , w15770 , w15771 , w15772 , w15773 , w15774 , w15775 , w15776 , w15777 , w15778 , w15779 , w15780 , w15781 , w15782 , w15783 , w15784 , w15785 , w15786 , w15787 , w15788 , w15789 , w15790 , w15791 , w15792 , w15793 , w15794 , w15795 , w15796 , w15797 , w15798 , w15799 , w15800 , w15801 , w15802 , w15803 , w15804 , w15805 , w15806 , w15807 , w15808 , w15809 , w15810 , w15811 , w15812 , w15813 , w15814 , w15815 , w15816 , w15817 , w15818 , w15819 , w15820 , w15821 , w15822 , w15823 , w15824 , w15825 , w15826 , w15827 , w15828 , w15829 , w15830 , w15831 , w15832 , w15833 , w15834 , w15835 , w15836 , w15837 , w15838 , w15839 , w15840 , w15841 , w15842 , w15843 , w15844 , w15845 , w15846 , w15847 , w15848 , w15849 , w15850 , w15851 , w15852 , w15853 , w15854 , w15855 , w15856 , w15857 , w15858 , w15859 , w15860 , w15861 , w15862 , w15863 , w15864 , w15865 , w15866 , w15867 , w15868 , w15869 , w15870 , w15871 , w15872 , w15873 , w15874 , w15875 , w15876 , w15877 , w15878 , w15879 , w15880 , w15881 , w15882 , w15883 , w15884 , w15885 , w15886 , w15887 , w15888 , w15889 , w15890 , w15891 , w15892 , w15893 , w15894 , w15895 , w15896 , w15897 , w15898 , w15899 , w15900 , w15901 , w15902 , w15903 , w15904 , w15905 , w15906 , w15907 , w15908 , w15909 , w15910 , w15911 , w15912 , w15913 , w15914 , w15915 , w15916 , w15917 , w15918 , w15919 , w15920 , w15921 , w15922 , w15923 , w15924 , w15925 , w15926 , w15927 , w15928 , w15929 , w15930 , w15931 , w15932 , w15933 , w15934 , w15935 , w15936 , w15937 , w15938 , w15939 , w15940 , w15941 , w15942 , w15943 , w15944 , w15945 , w15946 , w15947 , w15948 , w15949 , w15950 , w15951 , w15952 , w15953 , w15954 , w15955 , w15956 , w15957 , w15958 , w15959 , w15960 , w15961 , w15962 , w15963 , w15964 , w15965 , w15966 , w15967 , w15968 , w15969 , w15970 , w15971 , w15972 , w15973 , w15974 , w15975 , w15976 , w15977 , w15978 , w15979 , w15980 , w15981 , w15982 , w15983 , w15984 , w15985 , w15986 , w15987 , w15988 , w15989 , w15990 , w15991 , w15992 , w15993 , w15994 , w15995 , w15996 , w15997 , w15998 , w15999 , w16000 , w16001 , w16002 , w16003 , w16004 , w16005 , w16006 , w16007 , w16008 , w16009 , w16010 , w16011 , w16012 , w16013 , w16014 , w16015 , w16016 , w16017 , w16018 , w16019 , w16020 , w16021 , w16022 , w16023 , w16024 , w16025 , w16026 , w16027 , w16028 , w16029 , w16030 , w16031 , w16032 , w16033 , w16034 , w16035 , w16036 , w16037 , w16038 , w16039 , w16040 , w16041 , w16042 , w16043 , w16044 , w16045 , w16046 , w16047 , w16048 , w16049 , w16050 , w16051 , w16052 , w16053 , w16054 , w16055 , w16056 , w16057 , w16058 , w16059 , w16060 , w16061 , w16062 , w16063 , w16064 , w16065 , w16066 , w16067 , w16068 , w16069 , w16070 , w16071 , w16072 , w16073 , w16074 , w16075 , w16076 , w16077 , w16078 , w16079 , w16080 , w16081 , w16082 , w16083 , w16084 , w16085 , w16086 , w16087 , w16088 , w16089 , w16090 , w16091 , w16092 , w16093 , w16094 , w16095 , w16096 , w16097 , w16098 , w16099 , w16100 , w16101 , w16102 , w16103 , w16104 , w16105 , w16106 , w16107 , w16108 , w16109 , w16110 , w16111 , w16112 , w16113 , w16114 , w16115 , w16116 , w16117 , w16118 , w16119 , w16120 , w16121 , w16122 , w16123 , w16124 , w16125 , w16126 , w16127 , w16128 , w16129 , w16130 , w16131 , w16132 , w16133 , w16134 , w16135 , w16136 , w16137 , w16138 , w16139 , w16140 , w16141 , w16142 , w16143 , w16144 , w16145 , w16146 , w16147 , w16148 , w16149 , w16150 , w16151 , w16152 , w16153 , w16154 , w16155 , w16156 , w16157 , w16158 , w16159 , w16160 , w16161 , w16162 , w16163 , w16164 , w16165 , w16166 , w16167 , w16168 , w16169 , w16170 , w16171 , w16172 , w16173 , w16174 , w16175 , w16176 , w16177 , w16178 , w16179 , w16180 , w16181 , w16182 , w16183 , w16184 , w16185 , w16186 , w16187 , w16188 , w16189 , w16190 , w16191 , w16192 , w16193 , w16194 , w16195 , w16196 , w16197 , w16198 , w16199 , w16200 , w16201 , w16202 , w16203 , w16204 , w16205 , w16206 , w16207 , w16208 , w16209 , w16210 , w16211 , w16212 , w16213 , w16214 , w16215 , w16216 , w16217 , w16218 , w16219 , w16220 , w16221 , w16222 , w16223 , w16224 , w16225 , w16226 , w16227 , w16228 , w16229 , w16230 , w16231 , w16232 , w16233 , w16234 , w16235 , w16236 , w16237 , w16238 , w16239 , w16240 , w16241 , w16242 , w16243 , w16244 , w16245 , w16246 , w16247 , w16248 , w16249 , w16250 , w16251 , w16252 , w16253 , w16254 , w16255 , w16256 , w16257 , w16258 , w16259 , w16260 , w16261 , w16262 , w16263 , w16264 , w16265 , w16266 , w16267 , w16268 , w16269 , w16270 , w16271 , w16272 , w16273 , w16274 , w16275 , w16276 , w16277 , w16278 , w16279 , w16280 , w16281 , w16282 , w16283 , w16284 , w16285 , w16286 , w16287 , w16288 , w16289 , w16290 , w16291 , w16292 , w16293 , w16294 , w16295 , w16296 , w16297 , w16298 , w16299 , w16300 , w16301 , w16302 , w16303 , w16304 , w16305 , w16306 , w16307 , w16308 , w16309 , w16310 , w16311 , w16312 , w16313 , w16314 , w16315 , w16316 , w16317 , w16318 , w16319 , w16320 , w16321 , w16322 , w16323 , w16324 , w16325 , w16326 , w16327 , w16328 , w16329 , w16330 , w16331 , w16332 , w16333 , w16334 , w16335 , w16336 , w16337 , w16338 , w16339 , w16340 , w16341 , w16342 , w16343 , w16344 , w16345 , w16346 , w16347 , w16348 , w16349 , w16350 , w16351 , w16352 , w16353 , w16354 , w16355 , w16356 , w16357 , w16358 , w16359 , w16360 , w16361 , w16362 , w16363 , w16364 , w16365 , w16366 , w16367 , w16368 , w16369 , w16370 , w16371 , w16372 , w16373 , w16374 , w16375 , w16376 , w16377 , w16378 , w16379 , w16380 , w16381 , w16382 , w16383 , w16384 , w16385 , w16386 , w16387 , w16388 , w16389 , w16390 , w16391 , w16392 , w16393 , w16394 , w16395 , w16396 , w16397 , w16398 , w16399 , w16400 , w16401 , w16402 , w16403 , w16404 , w16405 , w16406 , w16407 , w16408 , w16409 , w16410 , w16411 , w16412 , w16413 , w16414 , w16415 , w16416 , w16417 , w16418 , w16419 , w16420 , w16421 , w16422 , w16423 , w16424 , w16425 , w16426 , w16427 , w16428 , w16429 , w16430 , w16431 , w16432 , w16433 , w16434 , w16435 , w16436 , w16437 , w16438 , w16439 , w16440 , w16441 , w16442 , w16443 , w16444 , w16445 , w16446 , w16447 , w16448 , w16449 , w16450 , w16451 , w16452 , w16453 , w16454 , w16455 , w16456 , w16457 , w16458 , w16459 , w16460 , w16461 , w16462 , w16463 , w16464 , w16465 , w16466 , w16467 , w16468 , w16469 , w16470 , w16471 , w16472 , w16473 , w16474 , w16475 , w16476 , w16477 , w16478 , w16479 , w16480 , w16481 , w16482 , w16483 , w16484 , w16485 , w16486 , w16487 , w16488 , w16489 , w16490 , w16491 , w16492 , w16493 , w16494 , w16495 , w16496 , w16497 , w16498 , w16499 , w16500 , w16501 , w16502 , w16503 , w16504 , w16505 , w16506 , w16507 , w16508 , w16509 , w16510 , w16511 , w16512 , w16513 , w16514 , w16515 , w16516 , w16517 , w16518 , w16519 , w16520 , w16521 , w16522 , w16523 , w16524 , w16525 , w16526 , w16527 , w16528 , w16529 , w16530 , w16531 , w16532 , w16533 , w16534 , w16535 , w16536 , w16537 , w16538 , w16539 , w16540 , w16541 , w16542 , w16543 , w16544 , w16545 , w16546 , w16547 , w16548 , w16549 , w16550 , w16551 , w16552 , w16553 , w16554 , w16555 , w16556 , w16557 , w16558 , w16559 , w16560 , w16561 , w16562 , w16563 , w16564 , w16565 , w16566 , w16567 , w16568 , w16569 , w16570 , w16571 , w16572 , w16573 , w16574 , w16575 , w16576 , w16577 , w16578 , w16579 , w16580 , w16581 , w16582 , w16583 , w16584 , w16585 , w16586 , w16587 , w16588 , w16589 , w16590 , w16591 , w16592 , w16593 , w16594 , w16595 , w16596 , w16597 , w16598 , w16599 , w16600 , w16601 , w16602 , w16603 , w16604 , w16605 , w16606 , w16607 , w16608 , w16609 , w16610 , w16611 , w16612 , w16613 , w16614 , w16615 , w16616 , w16617 , w16618 , w16619 , w16620 , w16621 , w16622 , w16623 , w16624 , w16625 , w16626 , w16627 , w16628 , w16629 , w16630 , w16631 , w16632 , w16633 , w16634 , w16635 , w16636 , w16637 , w16638 , w16639 , w16640 , w16641 , w16642 , w16643 , w16644 , w16645 , w16646 , w16647 , w16648 , w16649 , w16650 , w16651 , w16652 , w16653 , w16654 , w16655 , w16656 , w16657 , w16658 , w16659 , w16660 , w16661 , w16662 , w16663 , w16664 , w16665 , w16666 , w16667 , w16668 , w16669 , w16670 , w16671 , w16672 , w16673 , w16674 , w16675 , w16676 , w16677 , w16678 , w16679 , w16680 , w16681 , w16682 , w16683 , w16684 , w16685 , w16686 , w16687 , w16688 , w16689 , w16690 , w16691 , w16692 , w16693 , w16694 , w16695 , w16696 , w16697 , w16698 , w16699 , w16700 , w16701 , w16702 , w16703 ;
  assign zero = 0;
  assign w129 = \pi000 & \pi064 ;
  assign w130 = \pi000 & \pi065 ;
  assign w131 = \pi001 & \pi064 ;
  assign w132 = w130 ^ w131 ;
  assign w133 = ~\pi064 & \pi065 ;
  assign w134 = \pi066 ^ w133 ;
  assign w135 = \pi001 ^ \pi065 ;
  assign w136 = ( \pi001 & \pi066 ) | ( \pi001 & ~w135 ) | ( \pi066 & ~w135 ) ;
  assign w137 = ( \pi000 & \pi065 ) | ( \pi000 & w136 ) | ( \pi065 & w136 ) ;
  assign w138 = ( \pi002 & \pi064 ) | ( \pi002 & ~w137 ) | ( \pi064 & ~w137 ) ;
  assign w139 = ~\pi064 & w138 ;
  assign w140 = \pi001 & \pi065 ;
  assign w141 = \pi064 & w140 ;
  assign w142 = \pi066 ^ w141 ;
  assign w143 = \pi000 & w142 ;
  assign w144 = \pi002 & w141 ;
  assign w145 = \pi066 & w144 ;
  assign w146 = ( \pi002 & \pi064 ) | ( \pi002 & w145 ) | ( \pi064 & w145 ) ;
  assign w147 = w140 ^ w146 ;
  assign w148 = w143 ^ w147 ;
  assign w149 = ( ~\pi002 & \pi066 ) | ( ~\pi002 & \pi067 ) | ( \pi066 & \pi067 ) ;
  assign w150 = \pi000 ^ w149 ;
  assign w151 = ( \pi002 & \pi067 ) | ( \pi002 & ~w150 ) | ( \pi067 & ~w150 ) ;
  assign w152 = ( \pi002 & \pi066 ) | ( \pi002 & w150 ) | ( \pi066 & w150 ) ;
  assign w153 = \pi001 & w152 ;
  assign w154 = ( ~\pi000 & \pi065 ) | ( ~\pi000 & w153 ) | ( \pi065 & w153 ) ;
  assign w155 = ( \pi001 & \pi002 ) | ( \pi001 & ~w154 ) | ( \pi002 & ~w154 ) ;
  assign w156 = ( w151 & w153 ) | ( w151 & ~w155 ) | ( w153 & ~w155 ) ;
  assign w157 = \pi066 ^ \pi067 ;
  assign w158 = \pi065 & \pi066 ;
  assign w159 = ( \pi064 & \pi065 ) | ( \pi064 & w158 ) | ( \pi065 & w158 ) ;
  assign w160 = w157 ^ w159 ;
  assign w161 = \pi002 ^ w156 ;
  assign w162 = ~w156 & w160 ;
  assign w163 = \pi000 & w162 ;
  assign w164 = \pi001 ^ w163 ;
  assign w165 = ( \pi001 & w161 ) | ( \pi001 & ~w164 ) | ( w161 & ~w164 ) ;
  assign w166 = w139 ^ w165 ;
  assign w167 = \pi002 ^ \pi003 ;
  assign w168 = \pi064 & w167 ;
  assign w169 = w166 ^ w168 ;
  assign w170 = ( ~\pi002 & \pi067 ) | ( ~\pi002 & \pi068 ) | ( \pi067 & \pi068 ) ;
  assign w171 = \pi000 ^ w170 ;
  assign w172 = ( \pi002 & \pi068 ) | ( \pi002 & ~w171 ) | ( \pi068 & ~w171 ) ;
  assign w173 = ( \pi002 & \pi067 ) | ( \pi002 & w171 ) | ( \pi067 & w171 ) ;
  assign w174 = \pi001 & w173 ;
  assign w175 = ( ~\pi000 & \pi066 ) | ( ~\pi000 & w174 ) | ( \pi066 & w174 ) ;
  assign w176 = ( \pi001 & \pi002 ) | ( \pi001 & ~w175 ) | ( \pi002 & ~w175 ) ;
  assign w177 = ( w172 & w174 ) | ( w172 & ~w176 ) | ( w174 & ~w176 ) ;
  assign w178 = ( ~\pi065 & \pi066 ) | ( ~\pi065 & \pi067 ) | ( \pi066 & \pi067 ) ;
  assign w179 = ~\pi064 & \pi067 ;
  assign w180 = w178 | w179 ;
  assign w181 = \pi066 ^ \pi068 ;
  assign w182 = w180 ^ w181 ;
  assign w183 = \pi002 ^ w177 ;
  assign w184 = ~w177 & w182 ;
  assign w185 = \pi000 & w184 ;
  assign w186 = \pi001 ^ w185 ;
  assign w187 = ( \pi001 & w183 ) | ( \pi001 & ~w186 ) | ( w183 & ~w186 ) ;
  assign w188 = ( \pi002 & \pi003 ) | ( \pi002 & \pi004 ) | ( \pi003 & \pi004 ) ;
  assign w189 = \pi004 ^ w188 ;
  assign w190 = \pi004 ^ \pi005 ;
  assign w191 = w167 & ~w190 ;
  assign w192 = w167 & w190 ;
  assign w193 = ( \pi002 & \pi003 ) | ( \pi002 & ~\pi005 ) | ( \pi003 & ~\pi005 ) ;
  assign w194 = \pi005 & ~\pi064 ;
  assign w195 = ~\pi065 & w194 ;
  assign w196 = ( \pi002 & \pi003 ) | ( \pi002 & ~w195 ) | ( \pi003 & ~w195 ) ;
  assign w197 = ( \pi004 & \pi005 ) | ( \pi004 & ~w196 ) | ( \pi005 & ~w196 ) ;
  assign w198 = ( \pi004 & ~w194 ) | ( \pi004 & w196 ) | ( ~w194 & w196 ) ;
  assign w199 = ( w193 & w197 ) | ( w193 & ~w198 ) | ( w197 & ~w198 ) ;
  assign w200 = ( \pi002 & \pi003 ) | ( \pi002 & \pi065 ) | ( \pi003 & \pi065 ) ;
  assign w201 = \pi002 & \pi003 ;
  assign w202 = \pi064 ^ w201 ;
  assign w203 = ( \pi004 & w201 ) | ( \pi004 & w202 ) | ( w201 & w202 ) ;
  assign w204 = w200 ^ w203 ;
  assign w205 = ( w139 & w165 ) | ( w139 & w168 ) | ( w165 & w168 ) ;
  assign w206 = w187 ^ w205 ;
  assign w207 = w204 ^ w206 ;
  assign w208 = ( ~\pi002 & \pi068 ) | ( ~\pi002 & \pi069 ) | ( \pi068 & \pi069 ) ;
  assign w209 = \pi000 ^ w208 ;
  assign w210 = ( \pi002 & \pi069 ) | ( \pi002 & ~w209 ) | ( \pi069 & ~w209 ) ;
  assign w211 = ( \pi002 & \pi068 ) | ( \pi002 & w209 ) | ( \pi068 & w209 ) ;
  assign w212 = \pi001 & w211 ;
  assign w213 = ( ~\pi000 & \pi067 ) | ( ~\pi000 & w212 ) | ( \pi067 & w212 ) ;
  assign w214 = ( \pi001 & \pi002 ) | ( \pi001 & ~w213 ) | ( \pi002 & ~w213 ) ;
  assign w215 = ( w210 & w212 ) | ( w210 & ~w214 ) | ( w212 & ~w214 ) ;
  assign w216 = \pi067 ^ \pi069 ;
  assign w217 = ( ~\pi066 & \pi067 ) | ( ~\pi066 & \pi068 ) | ( \pi067 & \pi068 ) ;
  assign w218 = ( ~\pi065 & \pi068 ) | ( ~\pi065 & w217 ) | ( \pi068 & w217 ) ;
  assign w219 = w217 | w218 ;
  assign w220 = ( ~\pi064 & w218 ) | ( ~\pi064 & w219 ) | ( w218 & w219 ) ;
  assign w221 = w216 ^ w220 ;
  assign w222 = \pi002 ^ w215 ;
  assign w223 = ~w215 & w221 ;
  assign w224 = \pi000 & w223 ;
  assign w225 = \pi001 ^ w224 ;
  assign w226 = ( \pi001 & w222 ) | ( \pi001 & ~w225 ) | ( w222 & ~w225 ) ;
  assign w227 = ( \pi003 & ~\pi004 ) | ( \pi003 & \pi005 ) | ( ~\pi004 & \pi005 ) ;
  assign w228 = ( \pi002 & \pi003 ) | ( \pi002 & w227 ) | ( \pi003 & w227 ) ;
  assign w229 = w227 ^ w228 ;
  assign w230 = \pi064 & w229 ;
  assign w231 = ( \pi066 & w191 ) | ( \pi066 & w230 ) | ( w191 & w230 ) ;
  assign w232 = \pi065 | w231 ;
  assign w233 = ( w189 & w231 ) | ( w189 & w232 ) | ( w231 & w232 ) ;
  assign w234 = w230 | w233 ;
  assign w235 = ~w134 & w192 ;
  assign w236 = ( w192 & w234 ) | ( w192 & ~w235 ) | ( w234 & ~w235 ) ;
  assign w237 = \pi005 ^ w236 ;
  assign w238 = w199 & w237 ;
  assign w239 = ( w187 & w204 ) | ( w187 & w205 ) | ( w204 & w205 ) ;
  assign w240 = w199 ^ w226 ;
  assign w241 = w239 ^ w240 ;
  assign w242 = w237 ^ w241 ;
  assign w243 = w199 ^ w237 ;
  assign w244 = ( w226 & w239 ) | ( w226 & w243 ) | ( w239 & w243 ) ;
  assign w245 = ~\pi066 & w189 ;
  assign w246 = \pi065 & w229 ;
  assign w247 = ( w189 & ~w245 ) | ( w189 & w246 ) | ( ~w245 & w246 ) ;
  assign w248 = ~\pi067 & w191 ;
  assign w249 = w160 | w247 ;
  assign w250 = ( w192 & w247 ) | ( w192 & w249 ) | ( w247 & w249 ) ;
  assign w251 = ( w191 & ~w248 ) | ( w191 & w250 ) | ( ~w248 & w250 ) ;
  assign w252 = \pi005 ^ w251 ;
  assign w253 = w238 ^ w252 ;
  assign w254 = \pi005 ^ \pi006 ;
  assign w255 = \pi064 & w254 ;
  assign w256 = w253 ^ w255 ;
  assign w257 = ( ~\pi002 & \pi069 ) | ( ~\pi002 & \pi070 ) | ( \pi069 & \pi070 ) ;
  assign w258 = \pi000 ^ w257 ;
  assign w259 = ( \pi002 & \pi070 ) | ( \pi002 & ~w258 ) | ( \pi070 & ~w258 ) ;
  assign w260 = ( \pi002 & \pi069 ) | ( \pi002 & w258 ) | ( \pi069 & w258 ) ;
  assign w261 = \pi001 & w260 ;
  assign w262 = ( ~\pi000 & \pi068 ) | ( ~\pi000 & w261 ) | ( \pi068 & w261 ) ;
  assign w263 = ( \pi001 & \pi002 ) | ( \pi001 & ~w262 ) | ( \pi002 & ~w262 ) ;
  assign w264 = ( w259 & w261 ) | ( w259 & ~w263 ) | ( w261 & ~w263 ) ;
  assign w265 = ( \pi067 & \pi068 ) | ( \pi067 & \pi069 ) | ( \pi068 & \pi069 ) ;
  assign w266 = \pi065 & \pi068 ;
  assign w267 = ( \pi064 & \pi065 ) | ( \pi064 & w266 ) | ( \pi065 & w266 ) ;
  assign w268 = ( \pi066 & ~\pi068 ) | ( \pi066 & w267 ) | ( ~\pi068 & w267 ) ;
  assign w269 = ( \pi068 & w265 ) | ( \pi068 & w268 ) | ( w265 & w268 ) ;
  assign w270 = \pi069 ^ w269 ;
  assign w271 = \pi070 ^ w270 ;
  assign w272 = \pi002 ^ w264 ;
  assign w273 = \pi000 & ~w264 ;
  assign w274 = w271 & w273 ;
  assign w275 = \pi001 ^ w274 ;
  assign w276 = ( \pi001 & w272 ) | ( \pi001 & ~w275 ) | ( w272 & ~w275 ) ;
  assign w277 = w244 ^ w256 ;
  assign w278 = w276 ^ w277 ;
  assign w279 = ( w244 & w256 ) | ( w244 & w276 ) | ( w256 & w276 ) ;
  assign w280 = ( ~\pi002 & \pi070 ) | ( ~\pi002 & \pi071 ) | ( \pi070 & \pi071 ) ;
  assign w281 = \pi000 ^ w280 ;
  assign w282 = ( \pi002 & \pi071 ) | ( \pi002 & ~w281 ) | ( \pi071 & ~w281 ) ;
  assign w283 = ( \pi002 & \pi070 ) | ( \pi002 & w281 ) | ( \pi070 & w281 ) ;
  assign w284 = \pi001 & w283 ;
  assign w285 = ( ~\pi000 & \pi069 ) | ( ~\pi000 & w284 ) | ( \pi069 & w284 ) ;
  assign w286 = ( \pi001 & \pi002 ) | ( \pi001 & ~w285 ) | ( \pi002 & ~w285 ) ;
  assign w287 = ( w282 & w284 ) | ( w282 & ~w286 ) | ( w284 & ~w286 ) ;
  assign w288 = ( \pi069 & \pi070 ) | ( \pi069 & w269 ) | ( \pi070 & w269 ) ;
  assign w289 = \pi070 ^ w288 ;
  assign w290 = \pi071 ^ w289 ;
  assign w291 = \pi002 ^ w287 ;
  assign w292 = \pi000 & ~w287 ;
  assign w293 = w290 & w292 ;
  assign w294 = \pi001 ^ w293 ;
  assign w295 = ( \pi001 & w291 ) | ( \pi001 & ~w294 ) | ( w291 & ~w294 ) ;
  assign w296 = ~\pi067 & w189 ;
  assign w297 = \pi066 & w229 ;
  assign w298 = ( w189 & ~w296 ) | ( w189 & w297 ) | ( ~w296 & w297 ) ;
  assign w299 = ~\pi068 & w191 ;
  assign w300 = w182 | w298 ;
  assign w301 = ( w192 & w298 ) | ( w192 & w300 ) | ( w298 & w300 ) ;
  assign w302 = ( w191 & ~w299 ) | ( w191 & w301 ) | ( ~w299 & w301 ) ;
  assign w303 = \pi005 ^ w302 ;
  assign w304 = ( \pi005 & \pi006 ) | ( \pi005 & \pi007 ) | ( \pi006 & \pi007 ) ;
  assign w305 = \pi007 ^ w304 ;
  assign w306 = \pi007 ^ \pi008 ;
  assign w307 = w254 & ~w306 ;
  assign w308 = w254 & w306 ;
  assign w309 = ( \pi005 & \pi006 ) | ( \pi005 & ~\pi008 ) | ( \pi006 & ~\pi008 ) ;
  assign w310 = \pi008 & ~\pi064 ;
  assign w311 = ~\pi065 & w310 ;
  assign w312 = ( \pi005 & \pi006 ) | ( \pi005 & ~w311 ) | ( \pi006 & ~w311 ) ;
  assign w313 = ( \pi007 & \pi008 ) | ( \pi007 & ~w312 ) | ( \pi008 & ~w312 ) ;
  assign w314 = ( \pi007 & ~w310 ) | ( \pi007 & w312 ) | ( ~w310 & w312 ) ;
  assign w315 = ( w309 & w313 ) | ( w309 & ~w314 ) | ( w313 & ~w314 ) ;
  assign w316 = ( \pi005 & \pi006 ) | ( \pi005 & \pi065 ) | ( \pi006 & \pi065 ) ;
  assign w317 = \pi005 & \pi006 ;
  assign w318 = \pi064 ^ w317 ;
  assign w319 = ( \pi007 & w317 ) | ( \pi007 & w318 ) | ( w317 & w318 ) ;
  assign w320 = w316 ^ w319 ;
  assign w321 = ( w238 & w252 ) | ( w238 & w255 ) | ( w252 & w255 ) ;
  assign w322 = w303 ^ w321 ;
  assign w323 = w320 ^ w322 ;
  assign w324 = w279 ^ w323 ;
  assign w325 = w295 ^ w324 ;
  assign w326 = ( \pi006 & ~\pi007 ) | ( \pi006 & \pi008 ) | ( ~\pi007 & \pi008 ) ;
  assign w327 = ( \pi005 & \pi006 ) | ( \pi005 & w326 ) | ( \pi006 & w326 ) ;
  assign w328 = w326 ^ w327 ;
  assign w329 = \pi064 & w328 ;
  assign w330 = ( \pi066 & w307 ) | ( \pi066 & w329 ) | ( w307 & w329 ) ;
  assign w331 = \pi065 | w330 ;
  assign w332 = ( w305 & w330 ) | ( w305 & w331 ) | ( w330 & w331 ) ;
  assign w333 = w329 | w332 ;
  assign w334 = ~w134 & w308 ;
  assign w335 = ( w308 & w333 ) | ( w308 & ~w334 ) | ( w333 & ~w334 ) ;
  assign w336 = \pi008 ^ w335 ;
  assign w337 = w315 & w336 ;
  assign w338 = w315 ^ w336 ;
  assign w339 = ~\pi068 & w189 ;
  assign w340 = \pi067 & w229 ;
  assign w341 = ( w189 & ~w339 ) | ( w189 & w340 ) | ( ~w339 & w340 ) ;
  assign w342 = ~\pi069 & w191 ;
  assign w343 = w192 | w341 ;
  assign w344 = ( w221 & w341 ) | ( w221 & w343 ) | ( w341 & w343 ) ;
  assign w345 = ( w191 & ~w342 ) | ( w191 & w344 ) | ( ~w342 & w344 ) ;
  assign w346 = \pi005 ^ w345 ;
  assign w347 = ( w303 & w320 ) | ( w303 & w321 ) | ( w320 & w321 ) ;
  assign w348 = w338 ^ w347 ;
  assign w349 = w346 ^ w348 ;
  assign w350 = ( ~\pi002 & \pi071 ) | ( ~\pi002 & \pi072 ) | ( \pi071 & \pi072 ) ;
  assign w351 = \pi000 ^ w350 ;
  assign w352 = ( \pi002 & \pi072 ) | ( \pi002 & ~w351 ) | ( \pi072 & ~w351 ) ;
  assign w353 = ( \pi002 & \pi071 ) | ( \pi002 & w351 ) | ( \pi071 & w351 ) ;
  assign w354 = \pi001 & w353 ;
  assign w355 = ( ~\pi000 & \pi070 ) | ( ~\pi000 & w354 ) | ( \pi070 & w354 ) ;
  assign w356 = ( \pi001 & \pi002 ) | ( \pi001 & ~w355 ) | ( \pi002 & ~w355 ) ;
  assign w357 = ( w352 & w354 ) | ( w352 & ~w356 ) | ( w354 & ~w356 ) ;
  assign w358 = ( \pi069 & ~\pi071 ) | ( \pi069 & w269 ) | ( ~\pi071 & w269 ) ;
  assign w359 = ( ~\pi070 & \pi071 ) | ( ~\pi070 & w358 ) | ( \pi071 & w358 ) ;
  assign w360 = \pi072 ^ w358 ;
  assign w361 = w359 ^ w360 ;
  assign w362 = \pi002 ^ w357 ;
  assign w363 = \pi000 & ~w357 ;
  assign w364 = w361 & w363 ;
  assign w365 = \pi001 ^ w364 ;
  assign w366 = ( \pi001 & w362 ) | ( \pi001 & ~w365 ) | ( w362 & ~w365 ) ;
  assign w367 = ( w279 & w295 ) | ( w279 & w323 ) | ( w295 & w323 ) ;
  assign w368 = w349 ^ w367 ;
  assign w369 = w366 ^ w368 ;
  assign w370 = ~\pi069 & w189 ;
  assign w371 = \pi068 & w229 ;
  assign w372 = ( w189 & ~w370 ) | ( w189 & w371 ) | ( ~w370 & w371 ) ;
  assign w373 = ~\pi070 & w191 ;
  assign w374 = w271 | w372 ;
  assign w375 = ( w192 & w372 ) | ( w192 & w374 ) | ( w372 & w374 ) ;
  assign w376 = ( w191 & ~w373 ) | ( w191 & w375 ) | ( ~w373 & w375 ) ;
  assign w377 = \pi005 ^ w376 ;
  assign w378 = ~\pi066 & w305 ;
  assign w379 = \pi065 & w328 ;
  assign w380 = ( w305 & ~w378 ) | ( w305 & w379 ) | ( ~w378 & w379 ) ;
  assign w381 = ~\pi067 & w307 ;
  assign w382 = w160 | w380 ;
  assign w383 = ( w308 & w380 ) | ( w308 & w382 ) | ( w380 & w382 ) ;
  assign w384 = ( w307 & ~w381 ) | ( w307 & w383 ) | ( ~w381 & w383 ) ;
  assign w385 = \pi008 ^ w384 ;
  assign w386 = w337 ^ w385 ;
  assign w387 = \pi008 ^ \pi009 ;
  assign w388 = \pi064 & w387 ;
  assign w389 = w386 ^ w388 ;
  assign w390 = ( w338 & w346 ) | ( w338 & w347 ) | ( w346 & w347 ) ;
  assign w391 = w389 ^ w390 ;
  assign w392 = w377 ^ w391 ;
  assign w393 = ( ~\pi002 & \pi072 ) | ( ~\pi002 & \pi073 ) | ( \pi072 & \pi073 ) ;
  assign w394 = \pi000 ^ w393 ;
  assign w395 = ( \pi002 & \pi073 ) | ( \pi002 & ~w394 ) | ( \pi073 & ~w394 ) ;
  assign w396 = ( \pi002 & \pi072 ) | ( \pi002 & w394 ) | ( \pi072 & w394 ) ;
  assign w397 = \pi001 & w396 ;
  assign w398 = ( ~\pi000 & \pi071 ) | ( ~\pi000 & w397 ) | ( \pi071 & w397 ) ;
  assign w399 = ( \pi001 & \pi002 ) | ( \pi001 & ~w398 ) | ( \pi002 & ~w398 ) ;
  assign w400 = ( w395 & w397 ) | ( w395 & ~w399 ) | ( w397 & ~w399 ) ;
  assign w401 = ( \pi070 & \pi071 ) | ( \pi070 & \pi072 ) | ( \pi071 & \pi072 ) ;
  assign w402 = ( \pi071 & w288 ) | ( \pi071 & w401 ) | ( w288 & w401 ) ;
  assign w403 = \pi072 ^ \pi073 ;
  assign w404 = w402 ^ w403 ;
  assign w405 = \pi002 ^ w400 ;
  assign w406 = \pi000 & ~w400 ;
  assign w407 = w404 & w406 ;
  assign w408 = \pi001 ^ w407 ;
  assign w409 = ( \pi001 & w405 ) | ( \pi001 & ~w408 ) | ( w405 & ~w408 ) ;
  assign w410 = ( w349 & w366 ) | ( w349 & w367 ) | ( w366 & w367 ) ;
  assign w411 = w392 ^ w410 ;
  assign w412 = w409 ^ w411 ;
  assign w413 = ( w392 & w409 ) | ( w392 & w410 ) | ( w409 & w410 ) ;
  assign w414 = ~\pi070 & w189 ;
  assign w415 = \pi069 & w229 ;
  assign w416 = ( w189 & ~w414 ) | ( w189 & w415 ) | ( ~w414 & w415 ) ;
  assign w417 = ~\pi071 & w191 ;
  assign w418 = w290 | w416 ;
  assign w419 = ( w192 & w416 ) | ( w192 & w418 ) | ( w416 & w418 ) ;
  assign w420 = ( w191 & ~w417 ) | ( w191 & w419 ) | ( ~w417 & w419 ) ;
  assign w421 = \pi005 ^ w420 ;
  assign w422 = ( w337 & w385 ) | ( w337 & w388 ) | ( w385 & w388 ) ;
  assign w423 = ~\pi067 & w305 ;
  assign w424 = \pi066 & w328 ;
  assign w425 = ( w305 & ~w423 ) | ( w305 & w424 ) | ( ~w423 & w424 ) ;
  assign w426 = ~\pi068 & w307 ;
  assign w427 = w182 | w425 ;
  assign w428 = ( w308 & w425 ) | ( w308 & w427 ) | ( w425 & w427 ) ;
  assign w429 = ( w307 & ~w426 ) | ( w307 & w428 ) | ( ~w426 & w428 ) ;
  assign w430 = \pi008 ^ w429 ;
  assign w431 = ( \pi008 & \pi009 ) | ( \pi008 & \pi010 ) | ( \pi009 & \pi010 ) ;
  assign w432 = \pi010 ^ w431 ;
  assign w433 = \pi010 ^ \pi011 ;
  assign w434 = w387 & ~w433 ;
  assign w435 = w387 & w433 ;
  assign w436 = ( \pi008 & \pi009 ) | ( \pi008 & ~\pi011 ) | ( \pi009 & ~\pi011 ) ;
  assign w437 = \pi011 & ~\pi064 ;
  assign w438 = ~\pi065 & w437 ;
  assign w439 = ( \pi008 & \pi009 ) | ( \pi008 & ~w438 ) | ( \pi009 & ~w438 ) ;
  assign w440 = ( \pi010 & \pi011 ) | ( \pi010 & ~w439 ) | ( \pi011 & ~w439 ) ;
  assign w441 = ( \pi010 & ~w437 ) | ( \pi010 & w439 ) | ( ~w437 & w439 ) ;
  assign w442 = ( w436 & w440 ) | ( w436 & ~w441 ) | ( w440 & ~w441 ) ;
  assign w443 = ( \pi008 & \pi009 ) | ( \pi008 & \pi065 ) | ( \pi009 & \pi065 ) ;
  assign w444 = \pi008 & \pi009 ;
  assign w445 = \pi064 ^ w444 ;
  assign w446 = ( \pi010 & w444 ) | ( \pi010 & w445 ) | ( w444 & w445 ) ;
  assign w447 = w443 ^ w446 ;
  assign w448 = w422 ^ w430 ;
  assign w449 = w447 ^ w448 ;
  assign w450 = ( w377 & w389 ) | ( w377 & w390 ) | ( w389 & w390 ) ;
  assign w451 = w449 ^ w450 ;
  assign w452 = w421 ^ w451 ;
  assign w453 = ( ~\pi002 & \pi073 ) | ( ~\pi002 & \pi074 ) | ( \pi073 & \pi074 ) ;
  assign w454 = \pi000 ^ w453 ;
  assign w455 = ( \pi002 & \pi074 ) | ( \pi002 & ~w454 ) | ( \pi074 & ~w454 ) ;
  assign w456 = ( \pi002 & \pi073 ) | ( \pi002 & w454 ) | ( \pi073 & w454 ) ;
  assign w457 = \pi001 & w456 ;
  assign w458 = ( ~\pi000 & \pi072 ) | ( ~\pi000 & w457 ) | ( \pi072 & w457 ) ;
  assign w459 = ( \pi001 & \pi002 ) | ( \pi001 & ~w458 ) | ( \pi002 & ~w458 ) ;
  assign w460 = ( w455 & w457 ) | ( w455 & ~w459 ) | ( w457 & ~w459 ) ;
  assign w461 = ( \pi070 & \pi071 ) | ( \pi070 & ~\pi073 ) | ( \pi071 & ~\pi073 ) ;
  assign w462 = ( \pi071 & w288 ) | ( \pi071 & w461 ) | ( w288 & w461 ) ;
  assign w463 = ( \pi072 & \pi073 ) | ( \pi072 & w462 ) | ( \pi073 & w462 ) ;
  assign w464 = \pi073 ^ w463 ;
  assign w465 = \pi074 ^ w464 ;
  assign w466 = \pi002 ^ w460 ;
  assign w467 = \pi000 & ~w460 ;
  assign w468 = w465 & w467 ;
  assign w469 = \pi001 ^ w468 ;
  assign w470 = ( \pi001 & w466 ) | ( \pi001 & ~w469 ) | ( w466 & ~w469 ) ;
  assign w471 = w413 ^ w452 ;
  assign w472 = w470 ^ w471 ;
  assign w473 = ( w413 & w452 ) | ( w413 & w470 ) | ( w452 & w470 ) ;
  assign w474 = ( w421 & w449 ) | ( w421 & w450 ) | ( w449 & w450 ) ;
  assign w475 = ~\pi071 & w189 ;
  assign w476 = \pi070 & w229 ;
  assign w477 = ( w189 & ~w475 ) | ( w189 & w476 ) | ( ~w475 & w476 ) ;
  assign w478 = ~\pi072 & w191 ;
  assign w479 = w361 | w477 ;
  assign w480 = ( w192 & w477 ) | ( w192 & w479 ) | ( w477 & w479 ) ;
  assign w481 = ( w191 & ~w478 ) | ( w191 & w480 ) | ( ~w478 & w480 ) ;
  assign w482 = \pi005 ^ w481 ;
  assign w483 = ( w422 & w430 ) | ( w422 & w447 ) | ( w430 & w447 ) ;
  assign w484 = ( \pi009 & ~\pi010 ) | ( \pi009 & \pi011 ) | ( ~\pi010 & \pi011 ) ;
  assign w485 = ( \pi008 & \pi009 ) | ( \pi008 & w484 ) | ( \pi009 & w484 ) ;
  assign w486 = w484 ^ w485 ;
  assign w487 = \pi064 & w486 ;
  assign w488 = ( \pi066 & w434 ) | ( \pi066 & w487 ) | ( w434 & w487 ) ;
  assign w489 = \pi065 | w488 ;
  assign w490 = ( w432 & w488 ) | ( w432 & w489 ) | ( w488 & w489 ) ;
  assign w491 = w487 | w490 ;
  assign w492 = ~w134 & w435 ;
  assign w493 = ( w435 & w491 ) | ( w435 & ~w492 ) | ( w491 & ~w492 ) ;
  assign w494 = \pi011 ^ w493 ;
  assign w495 = w442 & w494 ;
  assign w496 = w442 ^ w494 ;
  assign w497 = ~\pi068 & w305 ;
  assign w498 = \pi067 & w328 ;
  assign w499 = ( w305 & ~w497 ) | ( w305 & w498 ) | ( ~w497 & w498 ) ;
  assign w500 = ~\pi069 & w307 ;
  assign w501 = w221 | w499 ;
  assign w502 = ( w308 & w499 ) | ( w308 & w501 ) | ( w499 & w501 ) ;
  assign w503 = ( w307 & ~w500 ) | ( w307 & w502 ) | ( ~w500 & w502 ) ;
  assign w504 = \pi008 ^ w503 ;
  assign w505 = w483 ^ w496 ;
  assign w506 = w504 ^ w505 ;
  assign w507 = w474 ^ w506 ;
  assign w508 = w482 ^ w507 ;
  assign w509 = ( ~\pi002 & \pi074 ) | ( ~\pi002 & \pi075 ) | ( \pi074 & \pi075 ) ;
  assign w510 = \pi000 ^ w509 ;
  assign w511 = ( \pi002 & \pi075 ) | ( \pi002 & ~w510 ) | ( \pi075 & ~w510 ) ;
  assign w512 = ( \pi002 & \pi074 ) | ( \pi002 & w510 ) | ( \pi074 & w510 ) ;
  assign w513 = \pi001 & w512 ;
  assign w514 = ( ~\pi000 & \pi073 ) | ( ~\pi000 & w513 ) | ( \pi073 & w513 ) ;
  assign w515 = ( \pi001 & \pi002 ) | ( \pi001 & ~w514 ) | ( \pi002 & ~w514 ) ;
  assign w516 = ( w511 & w513 ) | ( w511 & ~w515 ) | ( w513 & ~w515 ) ;
  assign w517 = ( \pi073 & \pi074 ) | ( \pi073 & w463 ) | ( \pi074 & w463 ) ;
  assign w518 = \pi074 ^ w517 ;
  assign w519 = \pi075 ^ w518 ;
  assign w520 = \pi002 ^ w516 ;
  assign w521 = \pi000 & ~w516 ;
  assign w522 = w519 & w521 ;
  assign w523 = \pi001 ^ w522 ;
  assign w524 = ( \pi001 & w520 ) | ( \pi001 & ~w523 ) | ( w520 & ~w523 ) ;
  assign w525 = w473 ^ w508 ;
  assign w526 = w524 ^ w525 ;
  assign w527 = ( ~\pi002 & \pi075 ) | ( ~\pi002 & \pi076 ) | ( \pi075 & \pi076 ) ;
  assign w528 = \pi000 ^ w527 ;
  assign w529 = ( \pi002 & \pi076 ) | ( \pi002 & ~w528 ) | ( \pi076 & ~w528 ) ;
  assign w530 = ( \pi002 & \pi075 ) | ( \pi002 & w528 ) | ( \pi075 & w528 ) ;
  assign w531 = \pi001 & w530 ;
  assign w532 = ( ~\pi000 & \pi074 ) | ( ~\pi000 & w531 ) | ( \pi074 & w531 ) ;
  assign w533 = ( \pi001 & \pi002 ) | ( \pi001 & ~w532 ) | ( \pi002 & ~w532 ) ;
  assign w534 = ( w529 & w531 ) | ( w529 & ~w533 ) | ( w531 & ~w533 ) ;
  assign w535 = ( \pi073 & ~\pi075 ) | ( \pi073 & w463 ) | ( ~\pi075 & w463 ) ;
  assign w536 = ( ~\pi074 & \pi075 ) | ( ~\pi074 & w535 ) | ( \pi075 & w535 ) ;
  assign w537 = \pi076 ^ w535 ;
  assign w538 = w536 ^ w537 ;
  assign w539 = \pi002 ^ w534 ;
  assign w540 = \pi000 & ~w534 ;
  assign w541 = w538 & w540 ;
  assign w542 = \pi001 ^ w541 ;
  assign w543 = ( \pi001 & w539 ) | ( \pi001 & ~w542 ) | ( w539 & ~w542 ) ;
  assign w544 = ~\pi069 & w305 ;
  assign w545 = \pi068 & w328 ;
  assign w546 = ( w305 & ~w544 ) | ( w305 & w545 ) | ( ~w544 & w545 ) ;
  assign w547 = ~\pi070 & w307 ;
  assign w548 = w271 | w546 ;
  assign w549 = ( w308 & w546 ) | ( w308 & w548 ) | ( w546 & w548 ) ;
  assign w550 = ( w307 & ~w547 ) | ( w307 & w549 ) | ( ~w547 & w549 ) ;
  assign w551 = \pi008 ^ w550 ;
  assign w552 = ~\pi066 & w432 ;
  assign w553 = \pi065 & w486 ;
  assign w554 = ( w432 & ~w552 ) | ( w432 & w553 ) | ( ~w552 & w553 ) ;
  assign w555 = ~\pi067 & w434 ;
  assign w556 = w160 | w554 ;
  assign w557 = ( w435 & w554 ) | ( w435 & w556 ) | ( w554 & w556 ) ;
  assign w558 = ( w434 & ~w555 ) | ( w434 & w557 ) | ( ~w555 & w557 ) ;
  assign w559 = \pi011 ^ w558 ;
  assign w560 = w495 ^ w559 ;
  assign w561 = \pi011 ^ \pi012 ;
  assign w562 = \pi064 & w561 ;
  assign w563 = w560 ^ w562 ;
  assign w564 = ( w483 & w496 ) | ( w483 & w504 ) | ( w496 & w504 ) ;
  assign w565 = w563 ^ w564 ;
  assign w566 = w551 ^ w565 ;
  assign w567 = ~\pi072 & w189 ;
  assign w568 = \pi071 & w229 ;
  assign w569 = ( w189 & ~w567 ) | ( w189 & w568 ) | ( ~w567 & w568 ) ;
  assign w570 = ~\pi073 & w191 ;
  assign w571 = w404 | w569 ;
  assign w572 = ( w192 & w569 ) | ( w192 & w571 ) | ( w569 & w571 ) ;
  assign w573 = ( w191 & ~w570 ) | ( w191 & w572 ) | ( ~w570 & w572 ) ;
  assign w574 = \pi005 ^ w573 ;
  assign w575 = ( w474 & w482 ) | ( w474 & w506 ) | ( w482 & w506 ) ;
  assign w576 = w566 ^ w575 ;
  assign w577 = w574 ^ w576 ;
  assign w578 = ( w473 & w508 ) | ( w473 & w524 ) | ( w508 & w524 ) ;
  assign w579 = w577 ^ w578 ;
  assign w580 = w543 ^ w579 ;
  assign w581 = ( w543 & w577 ) | ( w543 & w578 ) | ( w577 & w578 ) ;
  assign w582 = ( w566 & w574 ) | ( w566 & w575 ) | ( w574 & w575 ) ;
  assign w583 = ~\pi070 & w305 ;
  assign w584 = \pi069 & w328 ;
  assign w585 = ( w305 & ~w583 ) | ( w305 & w584 ) | ( ~w583 & w584 ) ;
  assign w586 = ~\pi071 & w307 ;
  assign w587 = w290 | w585 ;
  assign w588 = ( w308 & w585 ) | ( w308 & w587 ) | ( w585 & w587 ) ;
  assign w589 = ( w307 & ~w586 ) | ( w307 & w588 ) | ( ~w586 & w588 ) ;
  assign w590 = \pi008 ^ w589 ;
  assign w591 = ( w495 & w559 ) | ( w495 & w562 ) | ( w559 & w562 ) ;
  assign w592 = ~\pi067 & w432 ;
  assign w593 = \pi066 & w486 ;
  assign w594 = ( w432 & ~w592 ) | ( w432 & w593 ) | ( ~w592 & w593 ) ;
  assign w595 = ~\pi068 & w434 ;
  assign w596 = w182 | w594 ;
  assign w597 = ( w435 & w594 ) | ( w435 & w596 ) | ( w594 & w596 ) ;
  assign w598 = ( w434 & ~w595 ) | ( w434 & w597 ) | ( ~w595 & w597 ) ;
  assign w599 = \pi011 ^ w598 ;
  assign w600 = ( \pi011 & \pi012 ) | ( \pi011 & \pi013 ) | ( \pi012 & \pi013 ) ;
  assign w601 = \pi013 ^ w600 ;
  assign w602 = \pi013 ^ \pi014 ;
  assign w603 = w561 & ~w602 ;
  assign w604 = w561 & w602 ;
  assign w605 = ( \pi011 & \pi012 ) | ( \pi011 & ~\pi014 ) | ( \pi012 & ~\pi014 ) ;
  assign w606 = \pi014 & ~\pi064 ;
  assign w607 = ~\pi065 & w606 ;
  assign w608 = ( \pi011 & \pi012 ) | ( \pi011 & ~w607 ) | ( \pi012 & ~w607 ) ;
  assign w609 = ( \pi013 & \pi014 ) | ( \pi013 & ~w608 ) | ( \pi014 & ~w608 ) ;
  assign w610 = ( \pi013 & ~w606 ) | ( \pi013 & w608 ) | ( ~w606 & w608 ) ;
  assign w611 = ( w605 & w609 ) | ( w605 & ~w610 ) | ( w609 & ~w610 ) ;
  assign w612 = ( \pi011 & \pi012 ) | ( \pi011 & \pi065 ) | ( \pi012 & \pi065 ) ;
  assign w613 = \pi011 & \pi012 ;
  assign w614 = \pi064 ^ w613 ;
  assign w615 = ( \pi013 & w613 ) | ( \pi013 & w614 ) | ( w613 & w614 ) ;
  assign w616 = w612 ^ w615 ;
  assign w617 = w591 ^ w599 ;
  assign w618 = w616 ^ w617 ;
  assign w619 = ( w551 & w563 ) | ( w551 & w564 ) | ( w563 & w564 ) ;
  assign w620 = w618 ^ w619 ;
  assign w621 = w590 ^ w620 ;
  assign w622 = ~\pi073 & w189 ;
  assign w623 = \pi072 & w229 ;
  assign w624 = ( w189 & ~w622 ) | ( w189 & w623 ) | ( ~w622 & w623 ) ;
  assign w625 = ~\pi074 & w191 ;
  assign w626 = w465 | w624 ;
  assign w627 = ( w192 & w624 ) | ( w192 & w626 ) | ( w624 & w626 ) ;
  assign w628 = ( w191 & ~w625 ) | ( w191 & w627 ) | ( ~w625 & w627 ) ;
  assign w629 = \pi005 ^ w628 ;
  assign w630 = ( w582 & w621 ) | ( w582 & w629 ) | ( w621 & w629 ) ;
  assign w631 = w582 ^ w621 ;
  assign w632 = w629 ^ w631 ;
  assign w633 = ( ~\pi002 & \pi076 ) | ( ~\pi002 & \pi077 ) | ( \pi076 & \pi077 ) ;
  assign w634 = \pi000 ^ w633 ;
  assign w635 = ( \pi002 & \pi077 ) | ( \pi002 & ~w634 ) | ( \pi077 & ~w634 ) ;
  assign w636 = ( \pi002 & \pi076 ) | ( \pi002 & w634 ) | ( \pi076 & w634 ) ;
  assign w637 = \pi001 & w636 ;
  assign w638 = ( ~\pi000 & \pi075 ) | ( ~\pi000 & w637 ) | ( \pi075 & w637 ) ;
  assign w639 = ( \pi001 & \pi002 ) | ( \pi001 & ~w638 ) | ( \pi002 & ~w638 ) ;
  assign w640 = ( w635 & w637 ) | ( w635 & ~w639 ) | ( w637 & ~w639 ) ;
  assign w641 = ( \pi074 & \pi075 ) | ( \pi074 & \pi076 ) | ( \pi075 & \pi076 ) ;
  assign w642 = ( \pi075 & w517 ) | ( \pi075 & w641 ) | ( w517 & w641 ) ;
  assign w643 = \pi076 ^ \pi077 ;
  assign w644 = w642 ^ w643 ;
  assign w645 = \pi002 ^ w640 ;
  assign w646 = \pi000 & ~w640 ;
  assign w647 = w644 & w646 ;
  assign w648 = \pi001 ^ w647 ;
  assign w649 = ( \pi001 & w645 ) | ( \pi001 & ~w648 ) | ( w645 & ~w648 ) ;
  assign w650 = w581 ^ w632 ;
  assign w651 = w649 ^ w650 ;
  assign w652 = ( w581 & w632 ) | ( w581 & w649 ) | ( w632 & w649 ) ;
  assign w653 = ( ~\pi002 & \pi077 ) | ( ~\pi002 & \pi078 ) | ( \pi077 & \pi078 ) ;
  assign w654 = \pi000 ^ w653 ;
  assign w655 = ( \pi002 & \pi078 ) | ( \pi002 & ~w654 ) | ( \pi078 & ~w654 ) ;
  assign w656 = ( \pi002 & \pi077 ) | ( \pi002 & w654 ) | ( \pi077 & w654 ) ;
  assign w657 = \pi001 & w656 ;
  assign w658 = ( ~\pi000 & \pi076 ) | ( ~\pi000 & w657 ) | ( \pi076 & w657 ) ;
  assign w659 = ( \pi001 & \pi002 ) | ( \pi001 & ~w658 ) | ( \pi002 & ~w658 ) ;
  assign w660 = ( w655 & w657 ) | ( w655 & ~w659 ) | ( w657 & ~w659 ) ;
  assign w661 = ( \pi074 & \pi075 ) | ( \pi074 & ~\pi077 ) | ( \pi075 & ~\pi077 ) ;
  assign w662 = ( \pi075 & w517 ) | ( \pi075 & w661 ) | ( w517 & w661 ) ;
  assign w663 = ( \pi076 & \pi077 ) | ( \pi076 & w662 ) | ( \pi077 & w662 ) ;
  assign w664 = \pi077 ^ w663 ;
  assign w665 = \pi078 ^ w664 ;
  assign w666 = \pi002 ^ w660 ;
  assign w667 = \pi000 & ~w660 ;
  assign w668 = w665 & w667 ;
  assign w669 = \pi001 ^ w668 ;
  assign w670 = ( \pi001 & w666 ) | ( \pi001 & ~w669 ) | ( w666 & ~w669 ) ;
  assign w671 = ~\pi074 & w189 ;
  assign w672 = \pi073 & w229 ;
  assign w673 = ( w189 & ~w671 ) | ( w189 & w672 ) | ( ~w671 & w672 ) ;
  assign w674 = ~\pi075 & w191 ;
  assign w675 = w519 | w673 ;
  assign w676 = ( w192 & w673 ) | ( w192 & w675 ) | ( w673 & w675 ) ;
  assign w677 = ( w191 & ~w674 ) | ( w191 & w676 ) | ( ~w674 & w676 ) ;
  assign w678 = \pi005 ^ w677 ;
  assign w679 = ( w590 & w618 ) | ( w590 & w619 ) | ( w618 & w619 ) ;
  assign w680 = ( w591 & w599 ) | ( w591 & w616 ) | ( w599 & w616 ) ;
  assign w681 = ( \pi012 & ~\pi013 ) | ( \pi012 & \pi014 ) | ( ~\pi013 & \pi014 ) ;
  assign w682 = ( \pi011 & \pi012 ) | ( \pi011 & w681 ) | ( \pi012 & w681 ) ;
  assign w683 = w681 ^ w682 ;
  assign w684 = \pi064 & w683 ;
  assign w685 = ( \pi066 & w603 ) | ( \pi066 & w684 ) | ( w603 & w684 ) ;
  assign w686 = \pi065 | w685 ;
  assign w687 = ( w601 & w685 ) | ( w601 & w686 ) | ( w685 & w686 ) ;
  assign w688 = w684 | w687 ;
  assign w689 = ~w134 & w604 ;
  assign w690 = ( w604 & w688 ) | ( w604 & ~w689 ) | ( w688 & ~w689 ) ;
  assign w691 = \pi014 ^ w690 ;
  assign w692 = w611 & w691 ;
  assign w693 = w611 ^ w691 ;
  assign w694 = ~\pi068 & w432 ;
  assign w695 = \pi067 & w486 ;
  assign w696 = ( w432 & ~w694 ) | ( w432 & w695 ) | ( ~w694 & w695 ) ;
  assign w697 = ~\pi069 & w434 ;
  assign w698 = w221 | w696 ;
  assign w699 = ( w435 & w696 ) | ( w435 & w698 ) | ( w696 & w698 ) ;
  assign w700 = ( w434 & ~w697 ) | ( w434 & w699 ) | ( ~w697 & w699 ) ;
  assign w701 = \pi011 ^ w700 ;
  assign w702 = ( w680 & w693 ) | ( w680 & w701 ) | ( w693 & w701 ) ;
  assign w703 = w680 ^ w693 ;
  assign w704 = w701 ^ w703 ;
  assign w705 = ~\pi071 & w305 ;
  assign w706 = \pi070 & w328 ;
  assign w707 = ( w305 & ~w705 ) | ( w305 & w706 ) | ( ~w705 & w706 ) ;
  assign w708 = ~\pi072 & w307 ;
  assign w709 = w361 | w707 ;
  assign w710 = ( w308 & w707 ) | ( w308 & w709 ) | ( w707 & w709 ) ;
  assign w711 = ( w307 & ~w708 ) | ( w307 & w710 ) | ( ~w708 & w710 ) ;
  assign w712 = \pi008 ^ w711 ;
  assign w713 = w679 ^ w704 ;
  assign w714 = w712 ^ w713 ;
  assign w715 = w630 ^ w714 ;
  assign w716 = w678 ^ w715 ;
  assign w717 = w652 ^ w716 ;
  assign w718 = w670 ^ w717 ;
  assign w719 = ( w652 & w670 ) | ( w652 & w716 ) | ( w670 & w716 ) ;
  assign w720 = ( ~\pi002 & \pi078 ) | ( ~\pi002 & \pi079 ) | ( \pi078 & \pi079 ) ;
  assign w721 = \pi000 ^ w720 ;
  assign w722 = ( \pi002 & \pi079 ) | ( \pi002 & ~w721 ) | ( \pi079 & ~w721 ) ;
  assign w723 = ( \pi002 & \pi078 ) | ( \pi002 & w721 ) | ( \pi078 & w721 ) ;
  assign w724 = \pi001 & w723 ;
  assign w725 = ( ~\pi000 & \pi077 ) | ( ~\pi000 & w724 ) | ( \pi077 & w724 ) ;
  assign w726 = ( \pi001 & \pi002 ) | ( \pi001 & ~w725 ) | ( \pi002 & ~w725 ) ;
  assign w727 = ( w722 & w724 ) | ( w722 & ~w726 ) | ( w724 & ~w726 ) ;
  assign w728 = ( \pi077 & \pi078 ) | ( \pi077 & w663 ) | ( \pi078 & w663 ) ;
  assign w729 = \pi078 ^ w728 ;
  assign w730 = \pi079 ^ w729 ;
  assign w731 = \pi002 ^ w727 ;
  assign w732 = \pi000 & ~w727 ;
  assign w733 = w730 & w732 ;
  assign w734 = \pi001 ^ w733 ;
  assign w735 = ( \pi001 & w731 ) | ( \pi001 & ~w734 ) | ( w731 & ~w734 ) ;
  assign w736 = ( w630 & w678 ) | ( w630 & w714 ) | ( w678 & w714 ) ;
  assign w737 = ~\pi075 & w189 ;
  assign w738 = \pi074 & w229 ;
  assign w739 = ( w189 & ~w737 ) | ( w189 & w738 ) | ( ~w737 & w738 ) ;
  assign w740 = ~\pi076 & w191 ;
  assign w741 = w538 | w739 ;
  assign w742 = ( w192 & w739 ) | ( w192 & w741 ) | ( w739 & w741 ) ;
  assign w743 = ( w191 & ~w740 ) | ( w191 & w742 ) | ( ~w740 & w742 ) ;
  assign w744 = \pi005 ^ w743 ;
  assign w745 = ( w679 & w704 ) | ( w679 & w712 ) | ( w704 & w712 ) ;
  assign w746 = ~\pi072 & w305 ;
  assign w747 = \pi071 & w328 ;
  assign w748 = ( w305 & ~w746 ) | ( w305 & w747 ) | ( ~w746 & w747 ) ;
  assign w749 = ~\pi073 & w307 ;
  assign w750 = w404 | w748 ;
  assign w751 = ( w308 & w748 ) | ( w308 & w750 ) | ( w748 & w750 ) ;
  assign w752 = ( w307 & ~w749 ) | ( w307 & w751 ) | ( ~w749 & w751 ) ;
  assign w753 = \pi008 ^ w752 ;
  assign w754 = ~\pi069 & w432 ;
  assign w755 = \pi068 & w486 ;
  assign w756 = ( w432 & ~w754 ) | ( w432 & w755 ) | ( ~w754 & w755 ) ;
  assign w757 = ~\pi070 & w434 ;
  assign w758 = w271 | w756 ;
  assign w759 = ( w435 & w756 ) | ( w435 & w758 ) | ( w756 & w758 ) ;
  assign w760 = ( w434 & ~w757 ) | ( w434 & w759 ) | ( ~w757 & w759 ) ;
  assign w761 = \pi011 ^ w760 ;
  assign w762 = ~\pi066 & w601 ;
  assign w763 = \pi065 & w683 ;
  assign w764 = ( w601 & ~w762 ) | ( w601 & w763 ) | ( ~w762 & w763 ) ;
  assign w765 = ~\pi067 & w603 ;
  assign w766 = w160 | w764 ;
  assign w767 = ( w604 & w764 ) | ( w604 & w766 ) | ( w764 & w766 ) ;
  assign w768 = ( w603 & ~w765 ) | ( w603 & w767 ) | ( ~w765 & w767 ) ;
  assign w769 = \pi014 ^ w768 ;
  assign w770 = w692 ^ w769 ;
  assign w771 = \pi014 ^ \pi015 ;
  assign w772 = \pi064 & w771 ;
  assign w773 = w770 ^ w772 ;
  assign w774 = w702 ^ w773 ;
  assign w775 = w761 ^ w774 ;
  assign w776 = w745 ^ w775 ;
  assign w777 = w753 ^ w776 ;
  assign w778 = w736 ^ w777 ;
  assign w779 = w744 ^ w778 ;
  assign w780 = w719 ^ w779 ;
  assign w781 = w735 ^ w780 ;
  assign w782 = ( w719 & w735 ) | ( w719 & w779 ) | ( w735 & w779 ) ;
  assign w783 = ( ~\pi002 & \pi079 ) | ( ~\pi002 & \pi080 ) | ( \pi079 & \pi080 ) ;
  assign w784 = \pi000 ^ w783 ;
  assign w785 = ( \pi002 & \pi080 ) | ( \pi002 & ~w784 ) | ( \pi080 & ~w784 ) ;
  assign w786 = ( \pi002 & \pi079 ) | ( \pi002 & w784 ) | ( \pi079 & w784 ) ;
  assign w787 = \pi001 & w786 ;
  assign w788 = ( ~\pi000 & \pi078 ) | ( ~\pi000 & w787 ) | ( \pi078 & w787 ) ;
  assign w789 = ( \pi001 & \pi002 ) | ( \pi001 & ~w788 ) | ( \pi002 & ~w788 ) ;
  assign w790 = ( w785 & w787 ) | ( w785 & ~w789 ) | ( w787 & ~w789 ) ;
  assign w791 = ( \pi077 & ~\pi079 ) | ( \pi077 & w663 ) | ( ~\pi079 & w663 ) ;
  assign w792 = ( ~\pi078 & \pi079 ) | ( ~\pi078 & w791 ) | ( \pi079 & w791 ) ;
  assign w793 = \pi080 ^ w791 ;
  assign w794 = w792 ^ w793 ;
  assign w795 = \pi002 ^ w790 ;
  assign w796 = \pi000 & ~w790 ;
  assign w797 = w794 & w796 ;
  assign w798 = \pi001 ^ w797 ;
  assign w799 = ( \pi001 & w795 ) | ( \pi001 & ~w798 ) | ( w795 & ~w798 ) ;
  assign w800 = ( w736 & w744 ) | ( w736 & w777 ) | ( w744 & w777 ) ;
  assign w801 = ~\pi076 & w189 ;
  assign w802 = \pi075 & w229 ;
  assign w803 = ( w189 & ~w801 ) | ( w189 & w802 ) | ( ~w801 & w802 ) ;
  assign w804 = ~\pi077 & w191 ;
  assign w805 = w644 | w803 ;
  assign w806 = ( w192 & w803 ) | ( w192 & w805 ) | ( w803 & w805 ) ;
  assign w807 = ( w191 & ~w804 ) | ( w191 & w806 ) | ( ~w804 & w806 ) ;
  assign w808 = \pi005 ^ w807 ;
  assign w809 = ( w745 & w753 ) | ( w745 & w775 ) | ( w753 & w775 ) ;
  assign w810 = ~\pi073 & w305 ;
  assign w811 = \pi072 & w328 ;
  assign w812 = ( w305 & ~w810 ) | ( w305 & w811 ) | ( ~w810 & w811 ) ;
  assign w813 = ~\pi074 & w307 ;
  assign w814 = w465 | w812 ;
  assign w815 = ( w308 & w812 ) | ( w308 & w814 ) | ( w812 & w814 ) ;
  assign w816 = ( w307 & ~w813 ) | ( w307 & w815 ) | ( ~w813 & w815 ) ;
  assign w817 = \pi008 ^ w816 ;
  assign w818 = ( w702 & w761 ) | ( w702 & w773 ) | ( w761 & w773 ) ;
  assign w819 = ~\pi070 & w432 ;
  assign w820 = \pi069 & w486 ;
  assign w821 = ( w432 & ~w819 ) | ( w432 & w820 ) | ( ~w819 & w820 ) ;
  assign w822 = ~\pi071 & w434 ;
  assign w823 = w290 | w821 ;
  assign w824 = ( w435 & w821 ) | ( w435 & w823 ) | ( w821 & w823 ) ;
  assign w825 = ( w434 & ~w822 ) | ( w434 & w824 ) | ( ~w822 & w824 ) ;
  assign w826 = \pi011 ^ w825 ;
  assign w827 = ( w692 & w769 ) | ( w692 & w772 ) | ( w769 & w772 ) ;
  assign w828 = ~\pi067 & w601 ;
  assign w829 = \pi066 & w683 ;
  assign w830 = ( w601 & ~w828 ) | ( w601 & w829 ) | ( ~w828 & w829 ) ;
  assign w831 = ~\pi068 & w603 ;
  assign w832 = w182 | w830 ;
  assign w833 = ( w604 & w830 ) | ( w604 & w832 ) | ( w830 & w832 ) ;
  assign w834 = ( w603 & ~w831 ) | ( w603 & w833 ) | ( ~w831 & w833 ) ;
  assign w835 = \pi014 ^ w834 ;
  assign w836 = ( \pi014 & \pi015 ) | ( \pi014 & \pi016 ) | ( \pi015 & \pi016 ) ;
  assign w837 = \pi016 ^ w836 ;
  assign w838 = \pi016 ^ \pi017 ;
  assign w839 = w771 & ~w838 ;
  assign w840 = w771 & w838 ;
  assign w841 = ( \pi014 & \pi015 ) | ( \pi014 & ~\pi017 ) | ( \pi015 & ~\pi017 ) ;
  assign w842 = \pi017 & ~\pi064 ;
  assign w843 = ~\pi065 & w842 ;
  assign w844 = ( \pi014 & \pi015 ) | ( \pi014 & ~w843 ) | ( \pi015 & ~w843 ) ;
  assign w845 = ( \pi016 & \pi017 ) | ( \pi016 & ~w844 ) | ( \pi017 & ~w844 ) ;
  assign w846 = ( \pi016 & ~w842 ) | ( \pi016 & w844 ) | ( ~w842 & w844 ) ;
  assign w847 = ( w841 & w845 ) | ( w841 & ~w846 ) | ( w845 & ~w846 ) ;
  assign w848 = ( \pi014 & \pi015 ) | ( \pi014 & \pi065 ) | ( \pi015 & \pi065 ) ;
  assign w849 = \pi014 & \pi015 ;
  assign w850 = \pi064 ^ w849 ;
  assign w851 = ( \pi016 & w849 ) | ( \pi016 & w850 ) | ( w849 & w850 ) ;
  assign w852 = w848 ^ w851 ;
  assign w853 = w827 ^ w835 ;
  assign w854 = w852 ^ w853 ;
  assign w855 = w818 ^ w854 ;
  assign w856 = w826 ^ w855 ;
  assign w857 = w809 ^ w856 ;
  assign w858 = w817 ^ w857 ;
  assign w859 = w800 ^ w858 ;
  assign w860 = w808 ^ w859 ;
  assign w861 = w782 ^ w860 ;
  assign w862 = w799 ^ w861 ;
  assign w863 = ( ~\pi002 & \pi080 ) | ( ~\pi002 & \pi081 ) | ( \pi080 & \pi081 ) ;
  assign w864 = \pi000 ^ w863 ;
  assign w865 = ( \pi002 & \pi081 ) | ( \pi002 & ~w864 ) | ( \pi081 & ~w864 ) ;
  assign w866 = ( \pi002 & \pi080 ) | ( \pi002 & w864 ) | ( \pi080 & w864 ) ;
  assign w867 = \pi001 & w866 ;
  assign w868 = ( ~\pi000 & \pi079 ) | ( ~\pi000 & w867 ) | ( \pi079 & w867 ) ;
  assign w869 = ( \pi001 & \pi002 ) | ( \pi001 & ~w868 ) | ( \pi002 & ~w868 ) ;
  assign w870 = ( w865 & w867 ) | ( w865 & ~w869 ) | ( w867 & ~w869 ) ;
  assign w871 = ( \pi078 & \pi079 ) | ( \pi078 & \pi080 ) | ( \pi079 & \pi080 ) ;
  assign w872 = ( \pi079 & w728 ) | ( \pi079 & w871 ) | ( w728 & w871 ) ;
  assign w873 = \pi080 ^ \pi081 ;
  assign w874 = w872 ^ w873 ;
  assign w875 = \pi002 ^ w870 ;
  assign w876 = \pi000 & ~w870 ;
  assign w877 = w874 & w876 ;
  assign w878 = \pi001 ^ w877 ;
  assign w879 = ( \pi001 & w875 ) | ( \pi001 & ~w878 ) | ( w875 & ~w878 ) ;
  assign w880 = ( w800 & w808 ) | ( w800 & w858 ) | ( w808 & w858 ) ;
  assign w881 = ~\pi077 & w189 ;
  assign w882 = \pi076 & w229 ;
  assign w883 = ( w189 & ~w881 ) | ( w189 & w882 ) | ( ~w881 & w882 ) ;
  assign w884 = ~\pi078 & w191 ;
  assign w885 = w665 | w883 ;
  assign w886 = ( w192 & w883 ) | ( w192 & w885 ) | ( w883 & w885 ) ;
  assign w887 = ( w191 & ~w884 ) | ( w191 & w886 ) | ( ~w884 & w886 ) ;
  assign w888 = \pi005 ^ w887 ;
  assign w889 = ( w809 & w817 ) | ( w809 & w856 ) | ( w817 & w856 ) ;
  assign w890 = ~\pi074 & w305 ;
  assign w891 = \pi073 & w328 ;
  assign w892 = ( w305 & ~w890 ) | ( w305 & w891 ) | ( ~w890 & w891 ) ;
  assign w893 = ~\pi075 & w307 ;
  assign w894 = w519 | w892 ;
  assign w895 = ( w308 & w892 ) | ( w308 & w894 ) | ( w892 & w894 ) ;
  assign w896 = ( w307 & ~w893 ) | ( w307 & w895 ) | ( ~w893 & w895 ) ;
  assign w897 = \pi008 ^ w896 ;
  assign w898 = ( w818 & w826 ) | ( w818 & w854 ) | ( w826 & w854 ) ;
  assign w899 = ( w827 & w835 ) | ( w827 & w852 ) | ( w835 & w852 ) ;
  assign w900 = ( \pi015 & ~\pi016 ) | ( \pi015 & \pi017 ) | ( ~\pi016 & \pi017 ) ;
  assign w901 = ( \pi014 & \pi015 ) | ( \pi014 & w900 ) | ( \pi015 & w900 ) ;
  assign w902 = w900 ^ w901 ;
  assign w903 = \pi064 & w902 ;
  assign w904 = ( \pi066 & w839 ) | ( \pi066 & w903 ) | ( w839 & w903 ) ;
  assign w905 = \pi065 | w904 ;
  assign w906 = ( w837 & w904 ) | ( w837 & w905 ) | ( w904 & w905 ) ;
  assign w907 = w903 | w906 ;
  assign w908 = ~w134 & w840 ;
  assign w909 = ( w840 & w907 ) | ( w840 & ~w908 ) | ( w907 & ~w908 ) ;
  assign w910 = \pi017 ^ w909 ;
  assign w911 = w847 & w910 ;
  assign w912 = w847 ^ w910 ;
  assign w913 = ~\pi068 & w601 ;
  assign w914 = \pi067 & w683 ;
  assign w915 = ( w601 & ~w913 ) | ( w601 & w914 ) | ( ~w913 & w914 ) ;
  assign w916 = ~\pi069 & w603 ;
  assign w917 = w221 | w915 ;
  assign w918 = ( w604 & w915 ) | ( w604 & w917 ) | ( w915 & w917 ) ;
  assign w919 = ( w603 & ~w916 ) | ( w603 & w918 ) | ( ~w916 & w918 ) ;
  assign w920 = \pi014 ^ w919 ;
  assign w921 = ( w899 & w912 ) | ( w899 & w920 ) | ( w912 & w920 ) ;
  assign w922 = w899 ^ w912 ;
  assign w923 = w920 ^ w922 ;
  assign w924 = ~\pi071 & w432 ;
  assign w925 = \pi070 & w486 ;
  assign w926 = ( w432 & ~w924 ) | ( w432 & w925 ) | ( ~w924 & w925 ) ;
  assign w927 = ~\pi072 & w434 ;
  assign w928 = w361 | w926 ;
  assign w929 = ( w435 & w926 ) | ( w435 & w928 ) | ( w926 & w928 ) ;
  assign w930 = ( w434 & ~w927 ) | ( w434 & w929 ) | ( ~w927 & w929 ) ;
  assign w931 = \pi011 ^ w930 ;
  assign w932 = w898 ^ w923 ;
  assign w933 = w931 ^ w932 ;
  assign w934 = w889 ^ w933 ;
  assign w935 = w897 ^ w934 ;
  assign w936 = w880 ^ w935 ;
  assign w937 = w888 ^ w936 ;
  assign w938 = ( w782 & w799 ) | ( w782 & w860 ) | ( w799 & w860 ) ;
  assign w939 = w937 ^ w938 ;
  assign w940 = w879 ^ w939 ;
  assign w941 = ( w880 & w888 ) | ( w880 & w935 ) | ( w888 & w935 ) ;
  assign w942 = ~\pi078 & w189 ;
  assign w943 = \pi077 & w229 ;
  assign w944 = ( w189 & ~w942 ) | ( w189 & w943 ) | ( ~w942 & w943 ) ;
  assign w945 = ~\pi079 & w191 ;
  assign w946 = w730 | w944 ;
  assign w947 = ( w192 & w944 ) | ( w192 & w946 ) | ( w944 & w946 ) ;
  assign w948 = ( w191 & ~w945 ) | ( w191 & w947 ) | ( ~w945 & w947 ) ;
  assign w949 = \pi005 ^ w948 ;
  assign w950 = ( w889 & w897 ) | ( w889 & w933 ) | ( w897 & w933 ) ;
  assign w951 = ~\pi075 & w305 ;
  assign w952 = \pi074 & w328 ;
  assign w953 = ( w305 & ~w951 ) | ( w305 & w952 ) | ( ~w951 & w952 ) ;
  assign w954 = ~\pi076 & w307 ;
  assign w955 = w538 | w953 ;
  assign w956 = ( w308 & w953 ) | ( w308 & w955 ) | ( w953 & w955 ) ;
  assign w957 = ( w307 & ~w954 ) | ( w307 & w956 ) | ( ~w954 & w956 ) ;
  assign w958 = \pi008 ^ w957 ;
  assign w959 = ( w898 & w923 ) | ( w898 & w931 ) | ( w923 & w931 ) ;
  assign w960 = ~\pi069 & w601 ;
  assign w961 = \pi068 & w683 ;
  assign w962 = ( w601 & ~w960 ) | ( w601 & w961 ) | ( ~w960 & w961 ) ;
  assign w963 = ~\pi070 & w603 ;
  assign w964 = w271 | w962 ;
  assign w965 = ( w604 & w962 ) | ( w604 & w964 ) | ( w962 & w964 ) ;
  assign w966 = ( w603 & ~w963 ) | ( w603 & w965 ) | ( ~w963 & w965 ) ;
  assign w967 = \pi014 ^ w966 ;
  assign w968 = ~\pi066 & w837 ;
  assign w969 = \pi065 & w902 ;
  assign w970 = ( w837 & ~w968 ) | ( w837 & w969 ) | ( ~w968 & w969 ) ;
  assign w971 = ~\pi067 & w839 ;
  assign w972 = w160 | w970 ;
  assign w973 = ( w840 & w970 ) | ( w840 & w972 ) | ( w970 & w972 ) ;
  assign w974 = ( w839 & ~w971 ) | ( w839 & w973 ) | ( ~w971 & w973 ) ;
  assign w975 = \pi017 ^ w974 ;
  assign w976 = w911 ^ w975 ;
  assign w977 = \pi017 ^ \pi018 ;
  assign w978 = \pi064 & w977 ;
  assign w979 = w976 ^ w978 ;
  assign w980 = w921 ^ w979 ;
  assign w981 = w967 ^ w980 ;
  assign w982 = ~\pi072 & w432 ;
  assign w983 = \pi071 & w486 ;
  assign w984 = ( w432 & ~w982 ) | ( w432 & w983 ) | ( ~w982 & w983 ) ;
  assign w985 = ~\pi073 & w434 ;
  assign w986 = w404 | w984 ;
  assign w987 = ( w435 & w984 ) | ( w435 & w986 ) | ( w984 & w986 ) ;
  assign w988 = ( w434 & ~w985 ) | ( w434 & w987 ) | ( ~w985 & w987 ) ;
  assign w989 = \pi011 ^ w988 ;
  assign w990 = w959 ^ w981 ;
  assign w991 = w989 ^ w990 ;
  assign w992 = w950 ^ w991 ;
  assign w993 = w958 ^ w992 ;
  assign w994 = w941 ^ w993 ;
  assign w995 = w949 ^ w994 ;
  assign w996 = ( ~\pi002 & \pi081 ) | ( ~\pi002 & \pi082 ) | ( \pi081 & \pi082 ) ;
  assign w997 = \pi000 ^ w996 ;
  assign w998 = ( \pi002 & \pi082 ) | ( \pi002 & ~w997 ) | ( \pi082 & ~w997 ) ;
  assign w999 = ( \pi002 & \pi081 ) | ( \pi002 & w997 ) | ( \pi081 & w997 ) ;
  assign w1000 = \pi001 & w999 ;
  assign w1001 = ( ~\pi000 & \pi080 ) | ( ~\pi000 & w1000 ) | ( \pi080 & w1000 ) ;
  assign w1002 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1001 ) | ( \pi002 & ~w1001 ) ;
  assign w1003 = ( w998 & w1000 ) | ( w998 & ~w1002 ) | ( w1000 & ~w1002 ) ;
  assign w1004 = ( \pi078 & \pi079 ) | ( \pi078 & ~\pi081 ) | ( \pi079 & ~\pi081 ) ;
  assign w1005 = ( \pi079 & w728 ) | ( \pi079 & w1004 ) | ( w728 & w1004 ) ;
  assign w1006 = ( \pi080 & \pi081 ) | ( \pi080 & w1005 ) | ( \pi081 & w1005 ) ;
  assign w1007 = \pi081 ^ w1006 ;
  assign w1008 = \pi082 ^ w1007 ;
  assign w1009 = \pi002 ^ w1003 ;
  assign w1010 = \pi000 & ~w1003 ;
  assign w1011 = w1008 & w1010 ;
  assign w1012 = \pi001 ^ w1011 ;
  assign w1013 = ( \pi001 & w1009 ) | ( \pi001 & ~w1012 ) | ( w1009 & ~w1012 ) ;
  assign w1014 = ( w879 & w937 ) | ( w879 & w938 ) | ( w937 & w938 ) ;
  assign w1015 = w995 ^ w1014 ;
  assign w1016 = w1013 ^ w1015 ;
  assign w1017 = ~\pi079 & w189 ;
  assign w1018 = \pi078 & w229 ;
  assign w1019 = ( w189 & ~w1017 ) | ( w189 & w1018 ) | ( ~w1017 & w1018 ) ;
  assign w1020 = ~\pi080 & w191 ;
  assign w1021 = w794 | w1019 ;
  assign w1022 = ( w192 & w1019 ) | ( w192 & w1021 ) | ( w1019 & w1021 ) ;
  assign w1023 = ( w191 & ~w1020 ) | ( w191 & w1022 ) | ( ~w1020 & w1022 ) ;
  assign w1024 = \pi005 ^ w1023 ;
  assign w1025 = ( w921 & w967 ) | ( w921 & w979 ) | ( w967 & w979 ) ;
  assign w1026 = ~\pi070 & w601 ;
  assign w1027 = \pi069 & w683 ;
  assign w1028 = ( w601 & ~w1026 ) | ( w601 & w1027 ) | ( ~w1026 & w1027 ) ;
  assign w1029 = ~\pi071 & w603 ;
  assign w1030 = w290 | w1028 ;
  assign w1031 = ( w604 & w1028 ) | ( w604 & w1030 ) | ( w1028 & w1030 ) ;
  assign w1032 = ( w603 & ~w1029 ) | ( w603 & w1031 ) | ( ~w1029 & w1031 ) ;
  assign w1033 = \pi014 ^ w1032 ;
  assign w1034 = ( w911 & w975 ) | ( w911 & w978 ) | ( w975 & w978 ) ;
  assign w1035 = ~\pi067 & w837 ;
  assign w1036 = \pi066 & w902 ;
  assign w1037 = ( w837 & ~w1035 ) | ( w837 & w1036 ) | ( ~w1035 & w1036 ) ;
  assign w1038 = ~\pi068 & w839 ;
  assign w1039 = w182 | w1037 ;
  assign w1040 = ( w840 & w1037 ) | ( w840 & w1039 ) | ( w1037 & w1039 ) ;
  assign w1041 = ( w839 & ~w1038 ) | ( w839 & w1040 ) | ( ~w1038 & w1040 ) ;
  assign w1042 = \pi017 ^ w1041 ;
  assign w1043 = ( \pi017 & \pi018 ) | ( \pi017 & \pi019 ) | ( \pi018 & \pi019 ) ;
  assign w1044 = \pi019 ^ w1043 ;
  assign w1045 = \pi019 ^ \pi020 ;
  assign w1046 = w977 & ~w1045 ;
  assign w1047 = w977 & w1045 ;
  assign w1048 = ( \pi017 & \pi018 ) | ( \pi017 & ~\pi020 ) | ( \pi018 & ~\pi020 ) ;
  assign w1049 = \pi020 & ~\pi064 ;
  assign w1050 = ~\pi065 & w1049 ;
  assign w1051 = ( \pi017 & \pi018 ) | ( \pi017 & ~w1050 ) | ( \pi018 & ~w1050 ) ;
  assign w1052 = ( \pi019 & \pi020 ) | ( \pi019 & ~w1051 ) | ( \pi020 & ~w1051 ) ;
  assign w1053 = ( \pi019 & ~w1049 ) | ( \pi019 & w1051 ) | ( ~w1049 & w1051 ) ;
  assign w1054 = ( w1048 & w1052 ) | ( w1048 & ~w1053 ) | ( w1052 & ~w1053 ) ;
  assign w1055 = ( \pi017 & \pi018 ) | ( \pi017 & \pi065 ) | ( \pi018 & \pi065 ) ;
  assign w1056 = \pi017 & \pi018 ;
  assign w1057 = \pi064 ^ w1056 ;
  assign w1058 = ( \pi019 & w1056 ) | ( \pi019 & w1057 ) | ( w1056 & w1057 ) ;
  assign w1059 = w1055 ^ w1058 ;
  assign w1060 = w1034 ^ w1042 ;
  assign w1061 = w1059 ^ w1060 ;
  assign w1062 = w1025 ^ w1061 ;
  assign w1063 = w1033 ^ w1062 ;
  assign w1064 = ~\pi073 & w432 ;
  assign w1065 = \pi072 & w486 ;
  assign w1066 = ( w432 & ~w1064 ) | ( w432 & w1065 ) | ( ~w1064 & w1065 ) ;
  assign w1067 = ~\pi074 & w434 ;
  assign w1068 = w465 | w1066 ;
  assign w1069 = ( w435 & w1066 ) | ( w435 & w1068 ) | ( w1066 & w1068 ) ;
  assign w1070 = ( w434 & ~w1067 ) | ( w434 & w1069 ) | ( ~w1067 & w1069 ) ;
  assign w1071 = \pi011 ^ w1070 ;
  assign w1072 = ( w959 & w981 ) | ( w959 & w989 ) | ( w981 & w989 ) ;
  assign w1073 = w1063 ^ w1072 ;
  assign w1074 = w1071 ^ w1073 ;
  assign w1075 = ~\pi076 & w305 ;
  assign w1076 = \pi075 & w328 ;
  assign w1077 = ( w305 & ~w1075 ) | ( w305 & w1076 ) | ( ~w1075 & w1076 ) ;
  assign w1078 = ~\pi077 & w307 ;
  assign w1079 = w644 | w1077 ;
  assign w1080 = ( w308 & w1077 ) | ( w308 & w1079 ) | ( w1077 & w1079 ) ;
  assign w1081 = ( w307 & ~w1078 ) | ( w307 & w1080 ) | ( ~w1078 & w1080 ) ;
  assign w1082 = \pi008 ^ w1081 ;
  assign w1083 = ( w950 & w958 ) | ( w950 & w991 ) | ( w958 & w991 ) ;
  assign w1084 = w1074 ^ w1083 ;
  assign w1085 = w1082 ^ w1084 ;
  assign w1086 = ( w941 & w949 ) | ( w941 & w993 ) | ( w949 & w993 ) ;
  assign w1087 = w1085 ^ w1086 ;
  assign w1088 = w1024 ^ w1087 ;
  assign w1089 = ( ~\pi002 & \pi082 ) | ( ~\pi002 & \pi083 ) | ( \pi082 & \pi083 ) ;
  assign w1090 = \pi000 ^ w1089 ;
  assign w1091 = ( \pi002 & \pi083 ) | ( \pi002 & ~w1090 ) | ( \pi083 & ~w1090 ) ;
  assign w1092 = ( \pi002 & \pi082 ) | ( \pi002 & w1090 ) | ( \pi082 & w1090 ) ;
  assign w1093 = \pi001 & w1092 ;
  assign w1094 = ( ~\pi000 & \pi081 ) | ( ~\pi000 & w1093 ) | ( \pi081 & w1093 ) ;
  assign w1095 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1094 ) | ( \pi002 & ~w1094 ) ;
  assign w1096 = ( w1091 & w1093 ) | ( w1091 & ~w1095 ) | ( w1093 & ~w1095 ) ;
  assign w1097 = ( \pi081 & \pi082 ) | ( \pi081 & w1006 ) | ( \pi082 & w1006 ) ;
  assign w1098 = \pi082 ^ w1097 ;
  assign w1099 = \pi083 ^ w1098 ;
  assign w1100 = \pi002 ^ w1096 ;
  assign w1101 = \pi000 & ~w1096 ;
  assign w1102 = w1099 & w1101 ;
  assign w1103 = \pi001 ^ w1102 ;
  assign w1104 = ( \pi001 & w1100 ) | ( \pi001 & ~w1103 ) | ( w1100 & ~w1103 ) ;
  assign w1105 = ( w995 & w1013 ) | ( w995 & w1014 ) | ( w1013 & w1014 ) ;
  assign w1106 = w1088 ^ w1105 ;
  assign w1107 = w1104 ^ w1106 ;
  assign w1108 = ( w1024 & w1085 ) | ( w1024 & w1086 ) | ( w1085 & w1086 ) ;
  assign w1109 = ~\pi080 & w189 ;
  assign w1110 = \pi079 & w229 ;
  assign w1111 = ( w189 & ~w1109 ) | ( w189 & w1110 ) | ( ~w1109 & w1110 ) ;
  assign w1112 = ~\pi081 & w191 ;
  assign w1113 = w874 | w1111 ;
  assign w1114 = ( w192 & w1111 ) | ( w192 & w1113 ) | ( w1111 & w1113 ) ;
  assign w1115 = ( w191 & ~w1112 ) | ( w191 & w1114 ) | ( ~w1112 & w1114 ) ;
  assign w1116 = \pi005 ^ w1115 ;
  assign w1117 = ~\pi077 & w305 ;
  assign w1118 = \pi076 & w328 ;
  assign w1119 = ( w305 & ~w1117 ) | ( w305 & w1118 ) | ( ~w1117 & w1118 ) ;
  assign w1120 = ~\pi078 & w307 ;
  assign w1121 = w665 | w1119 ;
  assign w1122 = ( w308 & w1119 ) | ( w308 & w1121 ) | ( w1119 & w1121 ) ;
  assign w1123 = ( w307 & ~w1120 ) | ( w307 & w1122 ) | ( ~w1120 & w1122 ) ;
  assign w1124 = \pi008 ^ w1123 ;
  assign w1125 = ( w1063 & w1071 ) | ( w1063 & w1072 ) | ( w1071 & w1072 ) ;
  assign w1126 = ~\pi074 & w432 ;
  assign w1127 = \pi073 & w486 ;
  assign w1128 = ( w432 & ~w1126 ) | ( w432 & w1127 ) | ( ~w1126 & w1127 ) ;
  assign w1129 = ~\pi075 & w434 ;
  assign w1130 = w519 | w1128 ;
  assign w1131 = ( w435 & w1128 ) | ( w435 & w1130 ) | ( w1128 & w1130 ) ;
  assign w1132 = ( w434 & ~w1129 ) | ( w434 & w1131 ) | ( ~w1129 & w1131 ) ;
  assign w1133 = \pi011 ^ w1132 ;
  assign w1134 = ( w1025 & w1033 ) | ( w1025 & w1061 ) | ( w1033 & w1061 ) ;
  assign w1135 = ( w1034 & w1042 ) | ( w1034 & w1059 ) | ( w1042 & w1059 ) ;
  assign w1136 = ( \pi018 & ~\pi019 ) | ( \pi018 & \pi020 ) | ( ~\pi019 & \pi020 ) ;
  assign w1137 = ( \pi017 & \pi018 ) | ( \pi017 & w1136 ) | ( \pi018 & w1136 ) ;
  assign w1138 = w1136 ^ w1137 ;
  assign w1139 = \pi064 & w1138 ;
  assign w1140 = ( \pi066 & w1046 ) | ( \pi066 & w1139 ) | ( w1046 & w1139 ) ;
  assign w1141 = \pi065 | w1140 ;
  assign w1142 = ( w1044 & w1140 ) | ( w1044 & w1141 ) | ( w1140 & w1141 ) ;
  assign w1143 = w1139 | w1142 ;
  assign w1144 = ~w134 & w1047 ;
  assign w1145 = ( w1047 & w1143 ) | ( w1047 & ~w1144 ) | ( w1143 & ~w1144 ) ;
  assign w1146 = \pi020 ^ w1145 ;
  assign w1147 = w1054 & w1146 ;
  assign w1148 = w1054 ^ w1146 ;
  assign w1149 = ~\pi068 & w837 ;
  assign w1150 = \pi067 & w902 ;
  assign w1151 = ( w837 & ~w1149 ) | ( w837 & w1150 ) | ( ~w1149 & w1150 ) ;
  assign w1152 = ~\pi069 & w839 ;
  assign w1153 = w221 | w1151 ;
  assign w1154 = ( w840 & w1151 ) | ( w840 & w1153 ) | ( w1151 & w1153 ) ;
  assign w1155 = ( w839 & ~w1152 ) | ( w839 & w1154 ) | ( ~w1152 & w1154 ) ;
  assign w1156 = \pi017 ^ w1155 ;
  assign w1157 = ( w1135 & w1148 ) | ( w1135 & w1156 ) | ( w1148 & w1156 ) ;
  assign w1158 = w1135 ^ w1148 ;
  assign w1159 = w1156 ^ w1158 ;
  assign w1160 = ~\pi071 & w601 ;
  assign w1161 = \pi070 & w683 ;
  assign w1162 = ( w601 & ~w1160 ) | ( w601 & w1161 ) | ( ~w1160 & w1161 ) ;
  assign w1163 = ~\pi072 & w603 ;
  assign w1164 = w361 | w1162 ;
  assign w1165 = ( w604 & w1162 ) | ( w604 & w1164 ) | ( w1162 & w1164 ) ;
  assign w1166 = ( w603 & ~w1163 ) | ( w603 & w1165 ) | ( ~w1163 & w1165 ) ;
  assign w1167 = \pi014 ^ w1166 ;
  assign w1168 = w1134 ^ w1159 ;
  assign w1169 = w1167 ^ w1168 ;
  assign w1170 = w1125 ^ w1169 ;
  assign w1171 = w1133 ^ w1170 ;
  assign w1172 = ( w1074 & w1082 ) | ( w1074 & w1083 ) | ( w1082 & w1083 ) ;
  assign w1173 = w1171 ^ w1172 ;
  assign w1174 = w1124 ^ w1173 ;
  assign w1175 = w1108 ^ w1174 ;
  assign w1176 = w1116 ^ w1175 ;
  assign w1177 = ( ~\pi002 & \pi083 ) | ( ~\pi002 & \pi084 ) | ( \pi083 & \pi084 ) ;
  assign w1178 = \pi000 ^ w1177 ;
  assign w1179 = ( \pi002 & \pi084 ) | ( \pi002 & ~w1178 ) | ( \pi084 & ~w1178 ) ;
  assign w1180 = ( \pi002 & \pi083 ) | ( \pi002 & w1178 ) | ( \pi083 & w1178 ) ;
  assign w1181 = \pi001 & w1180 ;
  assign w1182 = ( ~\pi000 & \pi082 ) | ( ~\pi000 & w1181 ) | ( \pi082 & w1181 ) ;
  assign w1183 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1182 ) | ( \pi002 & ~w1182 ) ;
  assign w1184 = ( w1179 & w1181 ) | ( w1179 & ~w1183 ) | ( w1181 & ~w1183 ) ;
  assign w1185 = ( \pi081 & ~\pi083 ) | ( \pi081 & w1006 ) | ( ~\pi083 & w1006 ) ;
  assign w1186 = ( ~\pi082 & \pi083 ) | ( ~\pi082 & w1185 ) | ( \pi083 & w1185 ) ;
  assign w1187 = \pi084 ^ w1185 ;
  assign w1188 = w1186 ^ w1187 ;
  assign w1189 = \pi002 ^ w1184 ;
  assign w1190 = \pi000 & ~w1184 ;
  assign w1191 = w1188 & w1190 ;
  assign w1192 = \pi001 ^ w1191 ;
  assign w1193 = ( \pi001 & w1189 ) | ( \pi001 & ~w1192 ) | ( w1189 & ~w1192 ) ;
  assign w1194 = ( w1088 & w1104 ) | ( w1088 & w1105 ) | ( w1104 & w1105 ) ;
  assign w1195 = w1176 ^ w1194 ;
  assign w1196 = w1193 ^ w1195 ;
  assign w1197 = ( w1124 & w1171 ) | ( w1124 & w1172 ) | ( w1171 & w1172 ) ;
  assign w1198 = ~\pi078 & w305 ;
  assign w1199 = \pi077 & w328 ;
  assign w1200 = ( w305 & ~w1198 ) | ( w305 & w1199 ) | ( ~w1198 & w1199 ) ;
  assign w1201 = ~\pi079 & w307 ;
  assign w1202 = w730 | w1200 ;
  assign w1203 = ( w308 & w1200 ) | ( w308 & w1202 ) | ( w1200 & w1202 ) ;
  assign w1204 = ( w307 & ~w1201 ) | ( w307 & w1203 ) | ( ~w1201 & w1203 ) ;
  assign w1205 = \pi008 ^ w1204 ;
  assign w1206 = ( w1125 & w1133 ) | ( w1125 & w1169 ) | ( w1133 & w1169 ) ;
  assign w1207 = ~\pi075 & w432 ;
  assign w1208 = \pi074 & w486 ;
  assign w1209 = ( w432 & ~w1207 ) | ( w432 & w1208 ) | ( ~w1207 & w1208 ) ;
  assign w1210 = ~\pi076 & w434 ;
  assign w1211 = w538 | w1209 ;
  assign w1212 = ( w435 & w1209 ) | ( w435 & w1211 ) | ( w1209 & w1211 ) ;
  assign w1213 = ( w434 & ~w1210 ) | ( w434 & w1212 ) | ( ~w1210 & w1212 ) ;
  assign w1214 = \pi011 ^ w1213 ;
  assign w1215 = ( w1134 & w1159 ) | ( w1134 & w1167 ) | ( w1159 & w1167 ) ;
  assign w1216 = ~\pi069 & w837 ;
  assign w1217 = \pi068 & w902 ;
  assign w1218 = ( w837 & ~w1216 ) | ( w837 & w1217 ) | ( ~w1216 & w1217 ) ;
  assign w1219 = ~\pi070 & w839 ;
  assign w1220 = w271 | w1218 ;
  assign w1221 = ( w840 & w1218 ) | ( w840 & w1220 ) | ( w1218 & w1220 ) ;
  assign w1222 = ( w839 & ~w1219 ) | ( w839 & w1221 ) | ( ~w1219 & w1221 ) ;
  assign w1223 = \pi017 ^ w1222 ;
  assign w1224 = ~\pi066 & w1044 ;
  assign w1225 = \pi065 & w1138 ;
  assign w1226 = ( w1044 & ~w1224 ) | ( w1044 & w1225 ) | ( ~w1224 & w1225 ) ;
  assign w1227 = ~\pi067 & w1046 ;
  assign w1228 = w160 | w1226 ;
  assign w1229 = ( w1047 & w1226 ) | ( w1047 & w1228 ) | ( w1226 & w1228 ) ;
  assign w1230 = ( w1046 & ~w1227 ) | ( w1046 & w1229 ) | ( ~w1227 & w1229 ) ;
  assign w1231 = \pi020 ^ w1230 ;
  assign w1232 = w1147 ^ w1231 ;
  assign w1233 = \pi020 ^ \pi021 ;
  assign w1234 = \pi064 & w1233 ;
  assign w1235 = w1232 ^ w1234 ;
  assign w1236 = w1157 ^ w1235 ;
  assign w1237 = w1223 ^ w1236 ;
  assign w1238 = ~\pi072 & w601 ;
  assign w1239 = \pi071 & w683 ;
  assign w1240 = ( w601 & ~w1238 ) | ( w601 & w1239 ) | ( ~w1238 & w1239 ) ;
  assign w1241 = ~\pi073 & w603 ;
  assign w1242 = w404 | w1240 ;
  assign w1243 = ( w604 & w1240 ) | ( w604 & w1242 ) | ( w1240 & w1242 ) ;
  assign w1244 = ( w603 & ~w1241 ) | ( w603 & w1243 ) | ( ~w1241 & w1243 ) ;
  assign w1245 = \pi014 ^ w1244 ;
  assign w1246 = w1215 ^ w1237 ;
  assign w1247 = w1245 ^ w1246 ;
  assign w1248 = w1206 ^ w1247 ;
  assign w1249 = w1214 ^ w1248 ;
  assign w1250 = w1197 ^ w1249 ;
  assign w1251 = w1205 ^ w1250 ;
  assign w1252 = ~\pi081 & w189 ;
  assign w1253 = \pi080 & w229 ;
  assign w1254 = ( w189 & ~w1252 ) | ( w189 & w1253 ) | ( ~w1252 & w1253 ) ;
  assign w1255 = ~\pi082 & w191 ;
  assign w1256 = w1008 | w1254 ;
  assign w1257 = ( w192 & w1254 ) | ( w192 & w1256 ) | ( w1254 & w1256 ) ;
  assign w1258 = ( w191 & ~w1255 ) | ( w191 & w1257 ) | ( ~w1255 & w1257 ) ;
  assign w1259 = \pi005 ^ w1258 ;
  assign w1260 = ( w1108 & w1116 ) | ( w1108 & w1174 ) | ( w1116 & w1174 ) ;
  assign w1261 = w1251 ^ w1260 ;
  assign w1262 = w1259 ^ w1261 ;
  assign w1263 = ( ~\pi002 & \pi084 ) | ( ~\pi002 & \pi085 ) | ( \pi084 & \pi085 ) ;
  assign w1264 = \pi000 ^ w1263 ;
  assign w1265 = ( \pi002 & \pi085 ) | ( \pi002 & ~w1264 ) | ( \pi085 & ~w1264 ) ;
  assign w1266 = ( \pi002 & \pi084 ) | ( \pi002 & w1264 ) | ( \pi084 & w1264 ) ;
  assign w1267 = \pi001 & w1266 ;
  assign w1268 = ( ~\pi000 & \pi083 ) | ( ~\pi000 & w1267 ) | ( \pi083 & w1267 ) ;
  assign w1269 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1268 ) | ( \pi002 & ~w1268 ) ;
  assign w1270 = ( w1265 & w1267 ) | ( w1265 & ~w1269 ) | ( w1267 & ~w1269 ) ;
  assign w1271 = ( \pi082 & \pi083 ) | ( \pi082 & \pi084 ) | ( \pi083 & \pi084 ) ;
  assign w1272 = ( \pi083 & w1097 ) | ( \pi083 & w1271 ) | ( w1097 & w1271 ) ;
  assign w1273 = \pi084 ^ \pi085 ;
  assign w1274 = w1272 ^ w1273 ;
  assign w1275 = \pi002 ^ w1270 ;
  assign w1276 = \pi000 & ~w1270 ;
  assign w1277 = w1274 & w1276 ;
  assign w1278 = \pi001 ^ w1277 ;
  assign w1279 = ( \pi001 & w1275 ) | ( \pi001 & ~w1278 ) | ( w1275 & ~w1278 ) ;
  assign w1280 = ( w1176 & w1193 ) | ( w1176 & w1194 ) | ( w1193 & w1194 ) ;
  assign w1281 = w1262 ^ w1280 ;
  assign w1282 = w1279 ^ w1281 ;
  assign w1283 = ( w1262 & w1279 ) | ( w1262 & w1280 ) | ( w1279 & w1280 ) ;
  assign w1284 = ( w1197 & w1205 ) | ( w1197 & w1249 ) | ( w1205 & w1249 ) ;
  assign w1285 = ~\pi079 & w305 ;
  assign w1286 = \pi078 & w328 ;
  assign w1287 = ( w305 & ~w1285 ) | ( w305 & w1286 ) | ( ~w1285 & w1286 ) ;
  assign w1288 = ~\pi080 & w307 ;
  assign w1289 = w794 | w1287 ;
  assign w1290 = ( w308 & w1287 ) | ( w308 & w1289 ) | ( w1287 & w1289 ) ;
  assign w1291 = ( w307 & ~w1288 ) | ( w307 & w1290 ) | ( ~w1288 & w1290 ) ;
  assign w1292 = \pi008 ^ w1291 ;
  assign w1293 = ( w1206 & w1214 ) | ( w1206 & w1247 ) | ( w1214 & w1247 ) ;
  assign w1294 = ( w1157 & w1223 ) | ( w1157 & w1235 ) | ( w1223 & w1235 ) ;
  assign w1295 = ~\pi070 & w837 ;
  assign w1296 = \pi069 & w902 ;
  assign w1297 = ( w837 & ~w1295 ) | ( w837 & w1296 ) | ( ~w1295 & w1296 ) ;
  assign w1298 = ~\pi071 & w839 ;
  assign w1299 = w290 | w1297 ;
  assign w1300 = ( w840 & w1297 ) | ( w840 & w1299 ) | ( w1297 & w1299 ) ;
  assign w1301 = ( w839 & ~w1298 ) | ( w839 & w1300 ) | ( ~w1298 & w1300 ) ;
  assign w1302 = \pi017 ^ w1301 ;
  assign w1303 = ( w1147 & w1231 ) | ( w1147 & w1234 ) | ( w1231 & w1234 ) ;
  assign w1304 = ~\pi067 & w1044 ;
  assign w1305 = \pi066 & w1138 ;
  assign w1306 = ( w1044 & ~w1304 ) | ( w1044 & w1305 ) | ( ~w1304 & w1305 ) ;
  assign w1307 = ~\pi068 & w1046 ;
  assign w1308 = w182 | w1306 ;
  assign w1309 = ( w1047 & w1306 ) | ( w1047 & w1308 ) | ( w1306 & w1308 ) ;
  assign w1310 = ( w1046 & ~w1307 ) | ( w1046 & w1309 ) | ( ~w1307 & w1309 ) ;
  assign w1311 = \pi020 ^ w1310 ;
  assign w1312 = ( \pi020 & \pi021 ) | ( \pi020 & \pi022 ) | ( \pi021 & \pi022 ) ;
  assign w1313 = \pi022 ^ w1312 ;
  assign w1314 = \pi022 ^ \pi023 ;
  assign w1315 = w1233 & ~w1314 ;
  assign w1316 = w1233 & w1314 ;
  assign w1317 = ( \pi020 & \pi021 ) | ( \pi020 & ~\pi023 ) | ( \pi021 & ~\pi023 ) ;
  assign w1318 = \pi023 & ~\pi064 ;
  assign w1319 = ~\pi065 & w1318 ;
  assign w1320 = ( \pi020 & \pi021 ) | ( \pi020 & ~w1319 ) | ( \pi021 & ~w1319 ) ;
  assign w1321 = ( \pi022 & \pi023 ) | ( \pi022 & ~w1320 ) | ( \pi023 & ~w1320 ) ;
  assign w1322 = ( \pi022 & ~w1318 ) | ( \pi022 & w1320 ) | ( ~w1318 & w1320 ) ;
  assign w1323 = ( w1317 & w1321 ) | ( w1317 & ~w1322 ) | ( w1321 & ~w1322 ) ;
  assign w1324 = ( \pi020 & \pi021 ) | ( \pi020 & \pi065 ) | ( \pi021 & \pi065 ) ;
  assign w1325 = \pi020 & \pi021 ;
  assign w1326 = \pi064 ^ w1325 ;
  assign w1327 = ( \pi022 & w1325 ) | ( \pi022 & w1326 ) | ( w1325 & w1326 ) ;
  assign w1328 = w1324 ^ w1327 ;
  assign w1329 = w1303 ^ w1311 ;
  assign w1330 = w1328 ^ w1329 ;
  assign w1331 = w1294 ^ w1330 ;
  assign w1332 = w1302 ^ w1331 ;
  assign w1333 = ~\pi073 & w601 ;
  assign w1334 = \pi072 & w683 ;
  assign w1335 = ( w601 & ~w1333 ) | ( w601 & w1334 ) | ( ~w1333 & w1334 ) ;
  assign w1336 = ~\pi074 & w603 ;
  assign w1337 = w465 | w1335 ;
  assign w1338 = ( w604 & w1335 ) | ( w604 & w1337 ) | ( w1335 & w1337 ) ;
  assign w1339 = ( w603 & ~w1336 ) | ( w603 & w1338 ) | ( ~w1336 & w1338 ) ;
  assign w1340 = \pi014 ^ w1339 ;
  assign w1341 = ( w1215 & w1237 ) | ( w1215 & w1245 ) | ( w1237 & w1245 ) ;
  assign w1342 = w1332 ^ w1341 ;
  assign w1343 = w1340 ^ w1342 ;
  assign w1344 = ~\pi076 & w432 ;
  assign w1345 = \pi075 & w486 ;
  assign w1346 = ( w432 & ~w1344 ) | ( w432 & w1345 ) | ( ~w1344 & w1345 ) ;
  assign w1347 = ~\pi077 & w434 ;
  assign w1348 = w644 | w1346 ;
  assign w1349 = ( w435 & w1346 ) | ( w435 & w1348 ) | ( w1346 & w1348 ) ;
  assign w1350 = ( w434 & ~w1347 ) | ( w434 & w1349 ) | ( ~w1347 & w1349 ) ;
  assign w1351 = \pi011 ^ w1350 ;
  assign w1352 = w1293 ^ w1343 ;
  assign w1353 = w1351 ^ w1352 ;
  assign w1354 = w1284 ^ w1353 ;
  assign w1355 = w1292 ^ w1354 ;
  assign w1356 = ~\pi082 & w189 ;
  assign w1357 = \pi081 & w229 ;
  assign w1358 = ( w189 & ~w1356 ) | ( w189 & w1357 ) | ( ~w1356 & w1357 ) ;
  assign w1359 = ~\pi083 & w191 ;
  assign w1360 = w1099 | w1358 ;
  assign w1361 = ( w192 & w1358 ) | ( w192 & w1360 ) | ( w1358 & w1360 ) ;
  assign w1362 = ( w191 & ~w1359 ) | ( w191 & w1361 ) | ( ~w1359 & w1361 ) ;
  assign w1363 = \pi005 ^ w1362 ;
  assign w1364 = ( w1251 & w1259 ) | ( w1251 & w1260 ) | ( w1259 & w1260 ) ;
  assign w1365 = w1355 ^ w1364 ;
  assign w1366 = w1363 ^ w1365 ;
  assign w1367 = ( ~\pi002 & \pi085 ) | ( ~\pi002 & \pi086 ) | ( \pi085 & \pi086 ) ;
  assign w1368 = \pi000 ^ w1367 ;
  assign w1369 = ( \pi002 & \pi086 ) | ( \pi002 & ~w1368 ) | ( \pi086 & ~w1368 ) ;
  assign w1370 = ( \pi002 & \pi085 ) | ( \pi002 & w1368 ) | ( \pi085 & w1368 ) ;
  assign w1371 = \pi001 & w1370 ;
  assign w1372 = ( ~\pi000 & \pi084 ) | ( ~\pi000 & w1371 ) | ( \pi084 & w1371 ) ;
  assign w1373 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1372 ) | ( \pi002 & ~w1372 ) ;
  assign w1374 = ( w1369 & w1371 ) | ( w1369 & ~w1373 ) | ( w1371 & ~w1373 ) ;
  assign w1375 = ( \pi082 & \pi083 ) | ( \pi082 & ~\pi085 ) | ( \pi083 & ~\pi085 ) ;
  assign w1376 = ( \pi083 & w1097 ) | ( \pi083 & w1375 ) | ( w1097 & w1375 ) ;
  assign w1377 = ( \pi084 & \pi085 ) | ( \pi084 & w1376 ) | ( \pi085 & w1376 ) ;
  assign w1378 = \pi085 ^ w1377 ;
  assign w1379 = \pi086 ^ w1378 ;
  assign w1380 = \pi002 ^ w1374 ;
  assign w1381 = \pi000 & ~w1374 ;
  assign w1382 = w1379 & w1381 ;
  assign w1383 = \pi001 ^ w1382 ;
  assign w1384 = ( \pi001 & w1380 ) | ( \pi001 & ~w1383 ) | ( w1380 & ~w1383 ) ;
  assign w1385 = w1283 ^ w1366 ;
  assign w1386 = w1384 ^ w1385 ;
  assign w1387 = ( w1284 & w1292 ) | ( w1284 & w1353 ) | ( w1292 & w1353 ) ;
  assign w1388 = ~\pi080 & w305 ;
  assign w1389 = \pi079 & w328 ;
  assign w1390 = ( w305 & ~w1388 ) | ( w305 & w1389 ) | ( ~w1388 & w1389 ) ;
  assign w1391 = ~\pi081 & w307 ;
  assign w1392 = w874 | w1390 ;
  assign w1393 = ( w308 & w1390 ) | ( w308 & w1392 ) | ( w1390 & w1392 ) ;
  assign w1394 = ( w307 & ~w1391 ) | ( w307 & w1393 ) | ( ~w1391 & w1393 ) ;
  assign w1395 = \pi008 ^ w1394 ;
  assign w1396 = ~\pi077 & w432 ;
  assign w1397 = \pi076 & w486 ;
  assign w1398 = ( w432 & ~w1396 ) | ( w432 & w1397 ) | ( ~w1396 & w1397 ) ;
  assign w1399 = ~\pi078 & w434 ;
  assign w1400 = w665 | w1398 ;
  assign w1401 = ( w435 & w1398 ) | ( w435 & w1400 ) | ( w1398 & w1400 ) ;
  assign w1402 = ( w434 & ~w1399 ) | ( w434 & w1401 ) | ( ~w1399 & w1401 ) ;
  assign w1403 = \pi011 ^ w1402 ;
  assign w1404 = ( w1332 & w1340 ) | ( w1332 & w1341 ) | ( w1340 & w1341 ) ;
  assign w1405 = ~\pi074 & w601 ;
  assign w1406 = \pi073 & w683 ;
  assign w1407 = ( w601 & ~w1405 ) | ( w601 & w1406 ) | ( ~w1405 & w1406 ) ;
  assign w1408 = ~\pi075 & w603 ;
  assign w1409 = w519 | w1407 ;
  assign w1410 = ( w604 & w1407 ) | ( w604 & w1409 ) | ( w1407 & w1409 ) ;
  assign w1411 = ( w603 & ~w1408 ) | ( w603 & w1410 ) | ( ~w1408 & w1410 ) ;
  assign w1412 = \pi014 ^ w1411 ;
  assign w1413 = ( w1294 & w1302 ) | ( w1294 & w1330 ) | ( w1302 & w1330 ) ;
  assign w1414 = ( w1303 & w1311 ) | ( w1303 & w1328 ) | ( w1311 & w1328 ) ;
  assign w1415 = ( \pi021 & ~\pi022 ) | ( \pi021 & \pi023 ) | ( ~\pi022 & \pi023 ) ;
  assign w1416 = ( \pi020 & \pi021 ) | ( \pi020 & w1415 ) | ( \pi021 & w1415 ) ;
  assign w1417 = w1415 ^ w1416 ;
  assign w1418 = \pi064 & w1417 ;
  assign w1419 = ( \pi066 & w1315 ) | ( \pi066 & w1418 ) | ( w1315 & w1418 ) ;
  assign w1420 = \pi065 | w1419 ;
  assign w1421 = ( w1313 & w1419 ) | ( w1313 & w1420 ) | ( w1419 & w1420 ) ;
  assign w1422 = w1418 | w1421 ;
  assign w1423 = ~w134 & w1316 ;
  assign w1424 = ( w1316 & w1422 ) | ( w1316 & ~w1423 ) | ( w1422 & ~w1423 ) ;
  assign w1425 = \pi023 ^ w1424 ;
  assign w1426 = w1323 & w1425 ;
  assign w1427 = w1323 ^ w1425 ;
  assign w1428 = ~\pi068 & w1044 ;
  assign w1429 = \pi067 & w1138 ;
  assign w1430 = ( w1044 & ~w1428 ) | ( w1044 & w1429 ) | ( ~w1428 & w1429 ) ;
  assign w1431 = ~\pi069 & w1046 ;
  assign w1432 = w221 | w1430 ;
  assign w1433 = ( w1047 & w1430 ) | ( w1047 & w1432 ) | ( w1430 & w1432 ) ;
  assign w1434 = ( w1046 & ~w1431 ) | ( w1046 & w1433 ) | ( ~w1431 & w1433 ) ;
  assign w1435 = \pi020 ^ w1434 ;
  assign w1436 = ( w1414 & w1427 ) | ( w1414 & w1435 ) | ( w1427 & w1435 ) ;
  assign w1437 = w1414 ^ w1427 ;
  assign w1438 = w1435 ^ w1437 ;
  assign w1439 = ~\pi071 & w837 ;
  assign w1440 = \pi070 & w902 ;
  assign w1441 = ( w837 & ~w1439 ) | ( w837 & w1440 ) | ( ~w1439 & w1440 ) ;
  assign w1442 = ~\pi072 & w839 ;
  assign w1443 = w361 | w1441 ;
  assign w1444 = ( w840 & w1441 ) | ( w840 & w1443 ) | ( w1441 & w1443 ) ;
  assign w1445 = ( w839 & ~w1442 ) | ( w839 & w1444 ) | ( ~w1442 & w1444 ) ;
  assign w1446 = \pi017 ^ w1445 ;
  assign w1447 = w1413 ^ w1438 ;
  assign w1448 = w1446 ^ w1447 ;
  assign w1449 = w1404 ^ w1448 ;
  assign w1450 = w1412 ^ w1449 ;
  assign w1451 = ( w1293 & w1343 ) | ( w1293 & w1351 ) | ( w1343 & w1351 ) ;
  assign w1452 = w1450 ^ w1451 ;
  assign w1453 = w1403 ^ w1452 ;
  assign w1454 = w1387 ^ w1453 ;
  assign w1455 = w1395 ^ w1454 ;
  assign w1456 = ~\pi083 & w189 ;
  assign w1457 = \pi082 & w229 ;
  assign w1458 = ( w189 & ~w1456 ) | ( w189 & w1457 ) | ( ~w1456 & w1457 ) ;
  assign w1459 = ~\pi084 & w191 ;
  assign w1460 = w1188 | w1458 ;
  assign w1461 = ( w192 & w1458 ) | ( w192 & w1460 ) | ( w1458 & w1460 ) ;
  assign w1462 = ( w191 & ~w1459 ) | ( w191 & w1461 ) | ( ~w1459 & w1461 ) ;
  assign w1463 = \pi005 ^ w1462 ;
  assign w1464 = ( w1355 & w1363 ) | ( w1355 & w1364 ) | ( w1363 & w1364 ) ;
  assign w1465 = w1455 ^ w1464 ;
  assign w1466 = w1463 ^ w1465 ;
  assign w1467 = ( ~\pi002 & \pi086 ) | ( ~\pi002 & \pi087 ) | ( \pi086 & \pi087 ) ;
  assign w1468 = \pi000 ^ w1467 ;
  assign w1469 = ( \pi002 & \pi087 ) | ( \pi002 & ~w1468 ) | ( \pi087 & ~w1468 ) ;
  assign w1470 = ( \pi002 & \pi086 ) | ( \pi002 & w1468 ) | ( \pi086 & w1468 ) ;
  assign w1471 = \pi001 & w1470 ;
  assign w1472 = ( ~\pi000 & \pi085 ) | ( ~\pi000 & w1471 ) | ( \pi085 & w1471 ) ;
  assign w1473 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1472 ) | ( \pi002 & ~w1472 ) ;
  assign w1474 = ( w1469 & w1471 ) | ( w1469 & ~w1473 ) | ( w1471 & ~w1473 ) ;
  assign w1475 = ( \pi085 & \pi086 ) | ( \pi085 & w1377 ) | ( \pi086 & w1377 ) ;
  assign w1476 = \pi086 ^ w1475 ;
  assign w1477 = \pi087 ^ w1476 ;
  assign w1478 = \pi002 ^ w1474 ;
  assign w1479 = \pi000 & ~w1474 ;
  assign w1480 = w1477 & w1479 ;
  assign w1481 = \pi001 ^ w1480 ;
  assign w1482 = ( \pi001 & w1478 ) | ( \pi001 & ~w1481 ) | ( w1478 & ~w1481 ) ;
  assign w1483 = ( w1283 & w1366 ) | ( w1283 & w1384 ) | ( w1366 & w1384 ) ;
  assign w1484 = w1466 ^ w1483 ;
  assign w1485 = w1482 ^ w1484 ;
  assign w1486 = ( w1455 & w1463 ) | ( w1455 & w1464 ) | ( w1463 & w1464 ) ;
  assign w1487 = ~\pi084 & w189 ;
  assign w1488 = \pi083 & w229 ;
  assign w1489 = ( w189 & ~w1487 ) | ( w189 & w1488 ) | ( ~w1487 & w1488 ) ;
  assign w1490 = ~\pi085 & w191 ;
  assign w1491 = w1274 | w1489 ;
  assign w1492 = ( w192 & w1489 ) | ( w192 & w1491 ) | ( w1489 & w1491 ) ;
  assign w1493 = ( w191 & ~w1490 ) | ( w191 & w1492 ) | ( ~w1490 & w1492 ) ;
  assign w1494 = \pi005 ^ w1493 ;
  assign w1495 = ( w1387 & w1395 ) | ( w1387 & w1453 ) | ( w1395 & w1453 ) ;
  assign w1496 = ~\pi078 & w432 ;
  assign w1497 = \pi077 & w486 ;
  assign w1498 = ( w432 & ~w1496 ) | ( w432 & w1497 ) | ( ~w1496 & w1497 ) ;
  assign w1499 = ~\pi079 & w434 ;
  assign w1500 = w730 | w1498 ;
  assign w1501 = ( w435 & w1498 ) | ( w435 & w1500 ) | ( w1498 & w1500 ) ;
  assign w1502 = ( w434 & ~w1499 ) | ( w434 & w1501 ) | ( ~w1499 & w1501 ) ;
  assign w1503 = \pi011 ^ w1502 ;
  assign w1504 = ( w1404 & w1412 ) | ( w1404 & w1448 ) | ( w1412 & w1448 ) ;
  assign w1505 = ~\pi075 & w601 ;
  assign w1506 = \pi074 & w683 ;
  assign w1507 = ( w601 & ~w1505 ) | ( w601 & w1506 ) | ( ~w1505 & w1506 ) ;
  assign w1508 = ~\pi076 & w603 ;
  assign w1509 = w538 | w1507 ;
  assign w1510 = ( w604 & w1507 ) | ( w604 & w1509 ) | ( w1507 & w1509 ) ;
  assign w1511 = ( w603 & ~w1508 ) | ( w603 & w1510 ) | ( ~w1508 & w1510 ) ;
  assign w1512 = \pi014 ^ w1511 ;
  assign w1513 = ( w1413 & w1438 ) | ( w1413 & w1446 ) | ( w1438 & w1446 ) ;
  assign w1514 = ~\pi069 & w1044 ;
  assign w1515 = \pi068 & w1138 ;
  assign w1516 = ( w1044 & ~w1514 ) | ( w1044 & w1515 ) | ( ~w1514 & w1515 ) ;
  assign w1517 = ~\pi070 & w1046 ;
  assign w1518 = w271 | w1516 ;
  assign w1519 = ( w1047 & w1516 ) | ( w1047 & w1518 ) | ( w1516 & w1518 ) ;
  assign w1520 = ( w1046 & ~w1517 ) | ( w1046 & w1519 ) | ( ~w1517 & w1519 ) ;
  assign w1521 = \pi020 ^ w1520 ;
  assign w1522 = ~\pi066 & w1313 ;
  assign w1523 = \pi065 & w1417 ;
  assign w1524 = ( w1313 & ~w1522 ) | ( w1313 & w1523 ) | ( ~w1522 & w1523 ) ;
  assign w1525 = ~\pi067 & w1315 ;
  assign w1526 = w160 | w1524 ;
  assign w1527 = ( w1316 & w1524 ) | ( w1316 & w1526 ) | ( w1524 & w1526 ) ;
  assign w1528 = ( w1315 & ~w1525 ) | ( w1315 & w1527 ) | ( ~w1525 & w1527 ) ;
  assign w1529 = \pi023 ^ w1528 ;
  assign w1530 = w1426 ^ w1529 ;
  assign w1531 = \pi023 ^ \pi024 ;
  assign w1532 = \pi064 & w1531 ;
  assign w1533 = w1530 ^ w1532 ;
  assign w1534 = w1436 ^ w1533 ;
  assign w1535 = w1521 ^ w1534 ;
  assign w1536 = ~\pi072 & w837 ;
  assign w1537 = \pi071 & w902 ;
  assign w1538 = ( w837 & ~w1536 ) | ( w837 & w1537 ) | ( ~w1536 & w1537 ) ;
  assign w1539 = ~\pi073 & w839 ;
  assign w1540 = w404 | w1538 ;
  assign w1541 = ( w840 & w1538 ) | ( w840 & w1540 ) | ( w1538 & w1540 ) ;
  assign w1542 = ( w839 & ~w1539 ) | ( w839 & w1541 ) | ( ~w1539 & w1541 ) ;
  assign w1543 = \pi017 ^ w1542 ;
  assign w1544 = w1513 ^ w1535 ;
  assign w1545 = w1543 ^ w1544 ;
  assign w1546 = w1504 ^ w1545 ;
  assign w1547 = w1512 ^ w1546 ;
  assign w1548 = ( w1403 & w1450 ) | ( w1403 & w1451 ) | ( w1450 & w1451 ) ;
  assign w1549 = w1547 ^ w1548 ;
  assign w1550 = w1503 ^ w1549 ;
  assign w1551 = ~\pi081 & w305 ;
  assign w1552 = \pi080 & w328 ;
  assign w1553 = ( w305 & ~w1551 ) | ( w305 & w1552 ) | ( ~w1551 & w1552 ) ;
  assign w1554 = ~\pi082 & w307 ;
  assign w1555 = w1008 | w1553 ;
  assign w1556 = ( w308 & w1553 ) | ( w308 & w1555 ) | ( w1553 & w1555 ) ;
  assign w1557 = ( w307 & ~w1554 ) | ( w307 & w1556 ) | ( ~w1554 & w1556 ) ;
  assign w1558 = \pi008 ^ w1557 ;
  assign w1559 = w1495 ^ w1550 ;
  assign w1560 = w1558 ^ w1559 ;
  assign w1561 = w1486 ^ w1560 ;
  assign w1562 = w1494 ^ w1561 ;
  assign w1563 = ( ~\pi002 & \pi087 ) | ( ~\pi002 & \pi088 ) | ( \pi087 & \pi088 ) ;
  assign w1564 = \pi000 ^ w1563 ;
  assign w1565 = ( \pi002 & \pi088 ) | ( \pi002 & ~w1564 ) | ( \pi088 & ~w1564 ) ;
  assign w1566 = ( \pi002 & \pi087 ) | ( \pi002 & w1564 ) | ( \pi087 & w1564 ) ;
  assign w1567 = \pi001 & w1566 ;
  assign w1568 = ( ~\pi000 & \pi086 ) | ( ~\pi000 & w1567 ) | ( \pi086 & w1567 ) ;
  assign w1569 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1568 ) | ( \pi002 & ~w1568 ) ;
  assign w1570 = ( w1565 & w1567 ) | ( w1565 & ~w1569 ) | ( w1567 & ~w1569 ) ;
  assign w1571 = ( \pi085 & ~\pi087 ) | ( \pi085 & w1377 ) | ( ~\pi087 & w1377 ) ;
  assign w1572 = ( ~\pi086 & \pi087 ) | ( ~\pi086 & w1571 ) | ( \pi087 & w1571 ) ;
  assign w1573 = \pi088 ^ w1571 ;
  assign w1574 = w1572 ^ w1573 ;
  assign w1575 = \pi002 ^ w1570 ;
  assign w1576 = \pi000 & ~w1570 ;
  assign w1577 = w1574 & w1576 ;
  assign w1578 = \pi001 ^ w1577 ;
  assign w1579 = ( \pi001 & w1575 ) | ( \pi001 & ~w1578 ) | ( w1575 & ~w1578 ) ;
  assign w1580 = ( w1466 & w1482 ) | ( w1466 & w1483 ) | ( w1482 & w1483 ) ;
  assign w1581 = w1562 ^ w1580 ;
  assign w1582 = w1579 ^ w1581 ;
  assign w1583 = ( w1562 & w1579 ) | ( w1562 & w1580 ) | ( w1579 & w1580 ) ;
  assign w1584 = ( ~\pi002 & \pi088 ) | ( ~\pi002 & \pi089 ) | ( \pi088 & \pi089 ) ;
  assign w1585 = \pi000 ^ w1584 ;
  assign w1586 = ( \pi002 & \pi089 ) | ( \pi002 & ~w1585 ) | ( \pi089 & ~w1585 ) ;
  assign w1587 = ( \pi002 & \pi088 ) | ( \pi002 & w1585 ) | ( \pi088 & w1585 ) ;
  assign w1588 = \pi001 & w1587 ;
  assign w1589 = ( ~\pi000 & \pi087 ) | ( ~\pi000 & w1588 ) | ( \pi087 & w1588 ) ;
  assign w1590 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1589 ) | ( \pi002 & ~w1589 ) ;
  assign w1591 = ( w1586 & w1588 ) | ( w1586 & ~w1590 ) | ( w1588 & ~w1590 ) ;
  assign w1592 = ( \pi086 & \pi087 ) | ( \pi086 & \pi088 ) | ( \pi087 & \pi088 ) ;
  assign w1593 = ( \pi087 & w1475 ) | ( \pi087 & w1592 ) | ( w1475 & w1592 ) ;
  assign w1594 = \pi088 ^ \pi089 ;
  assign w1595 = w1593 ^ w1594 ;
  assign w1596 = \pi002 ^ w1591 ;
  assign w1597 = \pi000 & ~w1591 ;
  assign w1598 = w1595 & w1597 ;
  assign w1599 = \pi001 ^ w1598 ;
  assign w1600 = ( \pi001 & w1596 ) | ( \pi001 & ~w1599 ) | ( w1596 & ~w1599 ) ;
  assign w1601 = ( w1486 & w1494 ) | ( w1486 & w1560 ) | ( w1494 & w1560 ) ;
  assign w1602 = ~\pi079 & w432 ;
  assign w1603 = \pi078 & w486 ;
  assign w1604 = ( w432 & ~w1602 ) | ( w432 & w1603 ) | ( ~w1602 & w1603 ) ;
  assign w1605 = ~\pi080 & w434 ;
  assign w1606 = w794 | w1604 ;
  assign w1607 = ( w435 & w1604 ) | ( w435 & w1606 ) | ( w1604 & w1606 ) ;
  assign w1608 = ( w434 & ~w1605 ) | ( w434 & w1607 ) | ( ~w1605 & w1607 ) ;
  assign w1609 = \pi011 ^ w1608 ;
  assign w1610 = ( w1436 & w1521 ) | ( w1436 & w1533 ) | ( w1521 & w1533 ) ;
  assign w1611 = ~\pi070 & w1044 ;
  assign w1612 = \pi069 & w1138 ;
  assign w1613 = ( w1044 & ~w1611 ) | ( w1044 & w1612 ) | ( ~w1611 & w1612 ) ;
  assign w1614 = ~\pi071 & w1046 ;
  assign w1615 = w290 | w1613 ;
  assign w1616 = ( w1047 & w1613 ) | ( w1047 & w1615 ) | ( w1613 & w1615 ) ;
  assign w1617 = ( w1046 & ~w1614 ) | ( w1046 & w1616 ) | ( ~w1614 & w1616 ) ;
  assign w1618 = \pi020 ^ w1617 ;
  assign w1619 = ( w1426 & w1529 ) | ( w1426 & w1532 ) | ( w1529 & w1532 ) ;
  assign w1620 = ~\pi067 & w1313 ;
  assign w1621 = \pi066 & w1417 ;
  assign w1622 = ( w1313 & ~w1620 ) | ( w1313 & w1621 ) | ( ~w1620 & w1621 ) ;
  assign w1623 = ~\pi068 & w1315 ;
  assign w1624 = w182 | w1622 ;
  assign w1625 = ( w1316 & w1622 ) | ( w1316 & w1624 ) | ( w1622 & w1624 ) ;
  assign w1626 = ( w1315 & ~w1623 ) | ( w1315 & w1625 ) | ( ~w1623 & w1625 ) ;
  assign w1627 = \pi023 ^ w1626 ;
  assign w1628 = ( \pi023 & \pi024 ) | ( \pi023 & \pi025 ) | ( \pi024 & \pi025 ) ;
  assign w1629 = \pi025 ^ w1628 ;
  assign w1630 = \pi025 ^ \pi026 ;
  assign w1631 = w1531 & ~w1630 ;
  assign w1632 = w1531 & w1630 ;
  assign w1633 = ( \pi023 & \pi024 ) | ( \pi023 & ~\pi026 ) | ( \pi024 & ~\pi026 ) ;
  assign w1634 = \pi026 & ~\pi064 ;
  assign w1635 = ~\pi065 & w1634 ;
  assign w1636 = ( \pi023 & \pi024 ) | ( \pi023 & ~w1635 ) | ( \pi024 & ~w1635 ) ;
  assign w1637 = ( \pi025 & \pi026 ) | ( \pi025 & ~w1636 ) | ( \pi026 & ~w1636 ) ;
  assign w1638 = ( \pi025 & ~w1634 ) | ( \pi025 & w1636 ) | ( ~w1634 & w1636 ) ;
  assign w1639 = ( w1633 & w1637 ) | ( w1633 & ~w1638 ) | ( w1637 & ~w1638 ) ;
  assign w1640 = ( \pi023 & \pi024 ) | ( \pi023 & \pi065 ) | ( \pi024 & \pi065 ) ;
  assign w1641 = \pi023 & \pi024 ;
  assign w1642 = \pi064 ^ w1641 ;
  assign w1643 = ( \pi025 & w1641 ) | ( \pi025 & w1642 ) | ( w1641 & w1642 ) ;
  assign w1644 = w1640 ^ w1643 ;
  assign w1645 = w1619 ^ w1627 ;
  assign w1646 = w1644 ^ w1645 ;
  assign w1647 = w1610 ^ w1646 ;
  assign w1648 = w1618 ^ w1647 ;
  assign w1649 = ~\pi073 & w837 ;
  assign w1650 = \pi072 & w902 ;
  assign w1651 = ( w837 & ~w1649 ) | ( w837 & w1650 ) | ( ~w1649 & w1650 ) ;
  assign w1652 = ~\pi074 & w839 ;
  assign w1653 = w465 | w1651 ;
  assign w1654 = ( w840 & w1651 ) | ( w840 & w1653 ) | ( w1651 & w1653 ) ;
  assign w1655 = ( w839 & ~w1652 ) | ( w839 & w1654 ) | ( ~w1652 & w1654 ) ;
  assign w1656 = \pi017 ^ w1655 ;
  assign w1657 = ( w1513 & w1535 ) | ( w1513 & w1543 ) | ( w1535 & w1543 ) ;
  assign w1658 = w1648 ^ w1657 ;
  assign w1659 = w1656 ^ w1658 ;
  assign w1660 = ~\pi076 & w601 ;
  assign w1661 = \pi075 & w683 ;
  assign w1662 = ( w601 & ~w1660 ) | ( w601 & w1661 ) | ( ~w1660 & w1661 ) ;
  assign w1663 = ~\pi077 & w603 ;
  assign w1664 = w644 | w1662 ;
  assign w1665 = ( w604 & w1662 ) | ( w604 & w1664 ) | ( w1662 & w1664 ) ;
  assign w1666 = ( w603 & ~w1663 ) | ( w603 & w1665 ) | ( ~w1663 & w1665 ) ;
  assign w1667 = \pi014 ^ w1666 ;
  assign w1668 = ( w1504 & w1512 ) | ( w1504 & w1545 ) | ( w1512 & w1545 ) ;
  assign w1669 = w1659 ^ w1668 ;
  assign w1670 = w1667 ^ w1669 ;
  assign w1671 = ( w1503 & w1547 ) | ( w1503 & w1548 ) | ( w1547 & w1548 ) ;
  assign w1672 = w1670 ^ w1671 ;
  assign w1673 = w1609 ^ w1672 ;
  assign w1674 = ~\pi082 & w305 ;
  assign w1675 = \pi081 & w328 ;
  assign w1676 = ( w305 & ~w1674 ) | ( w305 & w1675 ) | ( ~w1674 & w1675 ) ;
  assign w1677 = ~\pi083 & w307 ;
  assign w1678 = w1099 | w1676 ;
  assign w1679 = ( w308 & w1676 ) | ( w308 & w1678 ) | ( w1676 & w1678 ) ;
  assign w1680 = ( w307 & ~w1677 ) | ( w307 & w1679 ) | ( ~w1677 & w1679 ) ;
  assign w1681 = \pi008 ^ w1680 ;
  assign w1682 = ( w1495 & w1550 ) | ( w1495 & w1558 ) | ( w1550 & w1558 ) ;
  assign w1683 = w1673 ^ w1682 ;
  assign w1684 = w1681 ^ w1683 ;
  assign w1685 = ~\pi085 & w189 ;
  assign w1686 = \pi084 & w229 ;
  assign w1687 = ( w189 & ~w1685 ) | ( w189 & w1686 ) | ( ~w1685 & w1686 ) ;
  assign w1688 = ~\pi086 & w191 ;
  assign w1689 = w1379 | w1687 ;
  assign w1690 = ( w192 & w1687 ) | ( w192 & w1689 ) | ( w1687 & w1689 ) ;
  assign w1691 = ( w191 & ~w1688 ) | ( w191 & w1690 ) | ( ~w1688 & w1690 ) ;
  assign w1692 = \pi005 ^ w1691 ;
  assign w1693 = w1601 ^ w1684 ;
  assign w1694 = w1692 ^ w1693 ;
  assign w1695 = w1583 ^ w1694 ;
  assign w1696 = w1600 ^ w1695 ;
  assign w1697 = ( w1583 & w1600 ) | ( w1583 & w1694 ) | ( w1600 & w1694 ) ;
  assign w1698 = ( w1601 & w1684 ) | ( w1601 & w1692 ) | ( w1684 & w1692 ) ;
  assign w1699 = ( w1609 & w1670 ) | ( w1609 & w1671 ) | ( w1670 & w1671 ) ;
  assign w1700 = ( w1659 & w1667 ) | ( w1659 & w1668 ) | ( w1667 & w1668 ) ;
  assign w1701 = ~\pi077 & w601 ;
  assign w1702 = \pi076 & w683 ;
  assign w1703 = ( w601 & ~w1701 ) | ( w601 & w1702 ) | ( ~w1701 & w1702 ) ;
  assign w1704 = ~\pi078 & w603 ;
  assign w1705 = w665 | w1703 ;
  assign w1706 = ( w604 & w1703 ) | ( w604 & w1705 ) | ( w1703 & w1705 ) ;
  assign w1707 = ( w603 & ~w1704 ) | ( w603 & w1706 ) | ( ~w1704 & w1706 ) ;
  assign w1708 = \pi014 ^ w1707 ;
  assign w1709 = ( w1648 & w1656 ) | ( w1648 & w1657 ) | ( w1656 & w1657 ) ;
  assign w1710 = ~\pi074 & w837 ;
  assign w1711 = \pi073 & w902 ;
  assign w1712 = ( w837 & ~w1710 ) | ( w837 & w1711 ) | ( ~w1710 & w1711 ) ;
  assign w1713 = ~\pi075 & w839 ;
  assign w1714 = w519 | w1712 ;
  assign w1715 = ( w840 & w1712 ) | ( w840 & w1714 ) | ( w1712 & w1714 ) ;
  assign w1716 = ( w839 & ~w1713 ) | ( w839 & w1715 ) | ( ~w1713 & w1715 ) ;
  assign w1717 = \pi017 ^ w1716 ;
  assign w1718 = ( w1610 & w1618 ) | ( w1610 & w1646 ) | ( w1618 & w1646 ) ;
  assign w1719 = ( w1619 & w1627 ) | ( w1619 & w1644 ) | ( w1627 & w1644 ) ;
  assign w1720 = ( \pi024 & ~\pi025 ) | ( \pi024 & \pi026 ) | ( ~\pi025 & \pi026 ) ;
  assign w1721 = ( \pi023 & \pi024 ) | ( \pi023 & w1720 ) | ( \pi024 & w1720 ) ;
  assign w1722 = w1720 ^ w1721 ;
  assign w1723 = \pi064 & w1722 ;
  assign w1724 = ( \pi066 & w1631 ) | ( \pi066 & w1723 ) | ( w1631 & w1723 ) ;
  assign w1725 = \pi065 | w1724 ;
  assign w1726 = ( w1629 & w1724 ) | ( w1629 & w1725 ) | ( w1724 & w1725 ) ;
  assign w1727 = w1723 | w1726 ;
  assign w1728 = ~w134 & w1632 ;
  assign w1729 = ( w1632 & w1727 ) | ( w1632 & ~w1728 ) | ( w1727 & ~w1728 ) ;
  assign w1730 = \pi026 ^ w1729 ;
  assign w1731 = w1639 & w1730 ;
  assign w1732 = w1639 ^ w1730 ;
  assign w1733 = ~\pi068 & w1313 ;
  assign w1734 = \pi067 & w1417 ;
  assign w1735 = ( w1313 & ~w1733 ) | ( w1313 & w1734 ) | ( ~w1733 & w1734 ) ;
  assign w1736 = ~\pi069 & w1315 ;
  assign w1737 = w221 | w1735 ;
  assign w1738 = ( w1316 & w1735 ) | ( w1316 & w1737 ) | ( w1735 & w1737 ) ;
  assign w1739 = ( w1315 & ~w1736 ) | ( w1315 & w1738 ) | ( ~w1736 & w1738 ) ;
  assign w1740 = \pi023 ^ w1739 ;
  assign w1741 = ( w1719 & w1732 ) | ( w1719 & w1740 ) | ( w1732 & w1740 ) ;
  assign w1742 = w1719 ^ w1732 ;
  assign w1743 = w1740 ^ w1742 ;
  assign w1744 = ~\pi071 & w1044 ;
  assign w1745 = \pi070 & w1138 ;
  assign w1746 = ( w1044 & ~w1744 ) | ( w1044 & w1745 ) | ( ~w1744 & w1745 ) ;
  assign w1747 = ~\pi072 & w1046 ;
  assign w1748 = w361 | w1746 ;
  assign w1749 = ( w1047 & w1746 ) | ( w1047 & w1748 ) | ( w1746 & w1748 ) ;
  assign w1750 = ( w1046 & ~w1747 ) | ( w1046 & w1749 ) | ( ~w1747 & w1749 ) ;
  assign w1751 = \pi020 ^ w1750 ;
  assign w1752 = w1718 ^ w1743 ;
  assign w1753 = w1751 ^ w1752 ;
  assign w1754 = w1709 ^ w1753 ;
  assign w1755 = w1717 ^ w1754 ;
  assign w1756 = w1700 ^ w1755 ;
  assign w1757 = w1708 ^ w1756 ;
  assign w1758 = ~\pi080 & w432 ;
  assign w1759 = \pi079 & w486 ;
  assign w1760 = ( w432 & ~w1758 ) | ( w432 & w1759 ) | ( ~w1758 & w1759 ) ;
  assign w1761 = ~\pi081 & w434 ;
  assign w1762 = w874 | w1760 ;
  assign w1763 = ( w435 & w1760 ) | ( w435 & w1762 ) | ( w1760 & w1762 ) ;
  assign w1764 = ( w434 & ~w1761 ) | ( w434 & w1763 ) | ( ~w1761 & w1763 ) ;
  assign w1765 = \pi011 ^ w1764 ;
  assign w1766 = w1699 ^ w1757 ;
  assign w1767 = w1765 ^ w1766 ;
  assign w1768 = ~\pi083 & w305 ;
  assign w1769 = \pi082 & w328 ;
  assign w1770 = ( w305 & ~w1768 ) | ( w305 & w1769 ) | ( ~w1768 & w1769 ) ;
  assign w1771 = ~\pi084 & w307 ;
  assign w1772 = w1188 | w1770 ;
  assign w1773 = ( w308 & w1770 ) | ( w308 & w1772 ) | ( w1770 & w1772 ) ;
  assign w1774 = ( w307 & ~w1771 ) | ( w307 & w1773 ) | ( ~w1771 & w1773 ) ;
  assign w1775 = \pi008 ^ w1774 ;
  assign w1776 = ( w1673 & w1681 ) | ( w1673 & w1682 ) | ( w1681 & w1682 ) ;
  assign w1777 = w1767 ^ w1776 ;
  assign w1778 = w1775 ^ w1777 ;
  assign w1779 = ~\pi086 & w189 ;
  assign w1780 = \pi085 & w229 ;
  assign w1781 = ( w189 & ~w1779 ) | ( w189 & w1780 ) | ( ~w1779 & w1780 ) ;
  assign w1782 = ~\pi087 & w191 ;
  assign w1783 = w1477 | w1781 ;
  assign w1784 = ( w192 & w1781 ) | ( w192 & w1783 ) | ( w1781 & w1783 ) ;
  assign w1785 = ( w191 & ~w1782 ) | ( w191 & w1784 ) | ( ~w1782 & w1784 ) ;
  assign w1786 = \pi005 ^ w1785 ;
  assign w1787 = w1698 ^ w1778 ;
  assign w1788 = w1786 ^ w1787 ;
  assign w1789 = ( ~\pi002 & \pi089 ) | ( ~\pi002 & \pi090 ) | ( \pi089 & \pi090 ) ;
  assign w1790 = \pi000 ^ w1789 ;
  assign w1791 = ( \pi002 & \pi090 ) | ( \pi002 & ~w1790 ) | ( \pi090 & ~w1790 ) ;
  assign w1792 = ( \pi002 & \pi089 ) | ( \pi002 & w1790 ) | ( \pi089 & w1790 ) ;
  assign w1793 = \pi001 & w1792 ;
  assign w1794 = ( ~\pi000 & \pi088 ) | ( ~\pi000 & w1793 ) | ( \pi088 & w1793 ) ;
  assign w1795 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1794 ) | ( \pi002 & ~w1794 ) ;
  assign w1796 = ( w1791 & w1793 ) | ( w1791 & ~w1795 ) | ( w1793 & ~w1795 ) ;
  assign w1797 = ( \pi086 & \pi087 ) | ( \pi086 & ~\pi089 ) | ( \pi087 & ~\pi089 ) ;
  assign w1798 = ( \pi087 & w1475 ) | ( \pi087 & w1797 ) | ( w1475 & w1797 ) ;
  assign w1799 = ( \pi088 & \pi089 ) | ( \pi088 & w1798 ) | ( \pi089 & w1798 ) ;
  assign w1800 = \pi089 ^ w1799 ;
  assign w1801 = \pi090 ^ w1800 ;
  assign w1802 = \pi002 ^ w1796 ;
  assign w1803 = \pi000 & ~w1796 ;
  assign w1804 = w1801 & w1803 ;
  assign w1805 = \pi001 ^ w1804 ;
  assign w1806 = ( \pi001 & w1802 ) | ( \pi001 & ~w1805 ) | ( w1802 & ~w1805 ) ;
  assign w1807 = w1697 ^ w1788 ;
  assign w1808 = w1806 ^ w1807 ;
  assign w1809 = ( w1697 & w1788 ) | ( w1697 & w1806 ) | ( w1788 & w1806 ) ;
  assign w1810 = ~\pi087 & w189 ;
  assign w1811 = \pi086 & w229 ;
  assign w1812 = ( w189 & ~w1810 ) | ( w189 & w1811 ) | ( ~w1810 & w1811 ) ;
  assign w1813 = ~\pi088 & w191 ;
  assign w1814 = w1574 | w1812 ;
  assign w1815 = ( w192 & w1812 ) | ( w192 & w1814 ) | ( w1812 & w1814 ) ;
  assign w1816 = ( w191 & ~w1813 ) | ( w191 & w1815 ) | ( ~w1813 & w1815 ) ;
  assign w1817 = \pi005 ^ w1816 ;
  assign w1818 = ~\pi078 & w601 ;
  assign w1819 = \pi077 & w683 ;
  assign w1820 = ( w601 & ~w1818 ) | ( w601 & w1819 ) | ( ~w1818 & w1819 ) ;
  assign w1821 = ~\pi079 & w603 ;
  assign w1822 = w730 | w1820 ;
  assign w1823 = ( w604 & w1820 ) | ( w604 & w1822 ) | ( w1820 & w1822 ) ;
  assign w1824 = ( w603 & ~w1821 ) | ( w603 & w1823 ) | ( ~w1821 & w1823 ) ;
  assign w1825 = \pi014 ^ w1824 ;
  assign w1826 = ( w1709 & w1717 ) | ( w1709 & w1753 ) | ( w1717 & w1753 ) ;
  assign w1827 = ~\pi075 & w837 ;
  assign w1828 = \pi074 & w902 ;
  assign w1829 = ( w837 & ~w1827 ) | ( w837 & w1828 ) | ( ~w1827 & w1828 ) ;
  assign w1830 = ~\pi076 & w839 ;
  assign w1831 = w538 | w1829 ;
  assign w1832 = ( w840 & w1829 ) | ( w840 & w1831 ) | ( w1829 & w1831 ) ;
  assign w1833 = ( w839 & ~w1830 ) | ( w839 & w1832 ) | ( ~w1830 & w1832 ) ;
  assign w1834 = \pi017 ^ w1833 ;
  assign w1835 = ( w1718 & w1743 ) | ( w1718 & w1751 ) | ( w1743 & w1751 ) ;
  assign w1836 = ~\pi069 & w1313 ;
  assign w1837 = \pi068 & w1417 ;
  assign w1838 = ( w1313 & ~w1836 ) | ( w1313 & w1837 ) | ( ~w1836 & w1837 ) ;
  assign w1839 = ~\pi070 & w1315 ;
  assign w1840 = w271 | w1838 ;
  assign w1841 = ( w1316 & w1838 ) | ( w1316 & w1840 ) | ( w1838 & w1840 ) ;
  assign w1842 = ( w1315 & ~w1839 ) | ( w1315 & w1841 ) | ( ~w1839 & w1841 ) ;
  assign w1843 = \pi023 ^ w1842 ;
  assign w1844 = ~\pi066 & w1629 ;
  assign w1845 = \pi065 & w1722 ;
  assign w1846 = ( w1629 & ~w1844 ) | ( w1629 & w1845 ) | ( ~w1844 & w1845 ) ;
  assign w1847 = ~\pi067 & w1631 ;
  assign w1848 = w160 | w1846 ;
  assign w1849 = ( w1632 & w1846 ) | ( w1632 & w1848 ) | ( w1846 & w1848 ) ;
  assign w1850 = ( w1631 & ~w1847 ) | ( w1631 & w1849 ) | ( ~w1847 & w1849 ) ;
  assign w1851 = \pi026 ^ w1850 ;
  assign w1852 = w1731 ^ w1851 ;
  assign w1853 = \pi026 ^ \pi027 ;
  assign w1854 = \pi064 & w1853 ;
  assign w1855 = w1852 ^ w1854 ;
  assign w1856 = w1741 ^ w1855 ;
  assign w1857 = w1843 ^ w1856 ;
  assign w1858 = ~\pi072 & w1044 ;
  assign w1859 = \pi071 & w1138 ;
  assign w1860 = ( w1044 & ~w1858 ) | ( w1044 & w1859 ) | ( ~w1858 & w1859 ) ;
  assign w1861 = ~\pi073 & w1046 ;
  assign w1862 = w404 | w1860 ;
  assign w1863 = ( w1047 & w1860 ) | ( w1047 & w1862 ) | ( w1860 & w1862 ) ;
  assign w1864 = ( w1046 & ~w1861 ) | ( w1046 & w1863 ) | ( ~w1861 & w1863 ) ;
  assign w1865 = \pi020 ^ w1864 ;
  assign w1866 = w1835 ^ w1857 ;
  assign w1867 = w1865 ^ w1866 ;
  assign w1868 = w1826 ^ w1867 ;
  assign w1869 = w1834 ^ w1868 ;
  assign w1870 = ( w1700 & w1708 ) | ( w1700 & w1755 ) | ( w1708 & w1755 ) ;
  assign w1871 = w1869 ^ w1870 ;
  assign w1872 = w1825 ^ w1871 ;
  assign w1873 = ~\pi081 & w432 ;
  assign w1874 = \pi080 & w486 ;
  assign w1875 = ( w432 & ~w1873 ) | ( w432 & w1874 ) | ( ~w1873 & w1874 ) ;
  assign w1876 = ~\pi082 & w434 ;
  assign w1877 = w1008 | w1875 ;
  assign w1878 = ( w435 & w1875 ) | ( w435 & w1877 ) | ( w1875 & w1877 ) ;
  assign w1879 = ( w434 & ~w1876 ) | ( w434 & w1878 ) | ( ~w1876 & w1878 ) ;
  assign w1880 = \pi011 ^ w1879 ;
  assign w1881 = ( w1699 & w1757 ) | ( w1699 & w1765 ) | ( w1757 & w1765 ) ;
  assign w1882 = w1872 ^ w1881 ;
  assign w1883 = w1880 ^ w1882 ;
  assign w1884 = ~\pi084 & w305 ;
  assign w1885 = \pi083 & w328 ;
  assign w1886 = ( w305 & ~w1884 ) | ( w305 & w1885 ) | ( ~w1884 & w1885 ) ;
  assign w1887 = ~\pi085 & w307 ;
  assign w1888 = w1274 | w1886 ;
  assign w1889 = ( w308 & w1886 ) | ( w308 & w1888 ) | ( w1886 & w1888 ) ;
  assign w1890 = ( w307 & ~w1887 ) | ( w307 & w1889 ) | ( ~w1887 & w1889 ) ;
  assign w1891 = \pi008 ^ w1890 ;
  assign w1892 = ( w1767 & w1775 ) | ( w1767 & w1776 ) | ( w1775 & w1776 ) ;
  assign w1893 = w1883 ^ w1892 ;
  assign w1894 = w1891 ^ w1893 ;
  assign w1895 = ( w1698 & w1778 ) | ( w1698 & w1786 ) | ( w1778 & w1786 ) ;
  assign w1896 = w1894 ^ w1895 ;
  assign w1897 = w1817 ^ w1896 ;
  assign w1898 = ( ~\pi002 & \pi090 ) | ( ~\pi002 & \pi091 ) | ( \pi090 & \pi091 ) ;
  assign w1899 = \pi000 ^ w1898 ;
  assign w1900 = ( \pi002 & \pi091 ) | ( \pi002 & ~w1899 ) | ( \pi091 & ~w1899 ) ;
  assign w1901 = ( \pi002 & \pi090 ) | ( \pi002 & w1899 ) | ( \pi090 & w1899 ) ;
  assign w1902 = \pi001 & w1901 ;
  assign w1903 = ( ~\pi000 & \pi089 ) | ( ~\pi000 & w1902 ) | ( \pi089 & w1902 ) ;
  assign w1904 = ( \pi001 & \pi002 ) | ( \pi001 & ~w1903 ) | ( \pi002 & ~w1903 ) ;
  assign w1905 = ( w1900 & w1902 ) | ( w1900 & ~w1904 ) | ( w1902 & ~w1904 ) ;
  assign w1906 = ( \pi089 & \pi090 ) | ( \pi089 & w1799 ) | ( \pi090 & w1799 ) ;
  assign w1907 = \pi090 ^ w1906 ;
  assign w1908 = \pi091 ^ w1907 ;
  assign w1909 = \pi002 ^ w1905 ;
  assign w1910 = \pi000 & ~w1905 ;
  assign w1911 = w1908 & w1910 ;
  assign w1912 = \pi001 ^ w1911 ;
  assign w1913 = ( \pi001 & w1909 ) | ( \pi001 & ~w1912 ) | ( w1909 & ~w1912 ) ;
  assign w1914 = w1809 ^ w1897 ;
  assign w1915 = w1913 ^ w1914 ;
  assign w1916 = ( w1809 & w1897 ) | ( w1809 & w1913 ) | ( w1897 & w1913 ) ;
  assign w1917 = ~\pi088 & w189 ;
  assign w1918 = \pi087 & w229 ;
  assign w1919 = ( w189 & ~w1917 ) | ( w189 & w1918 ) | ( ~w1917 & w1918 ) ;
  assign w1920 = ~\pi089 & w191 ;
  assign w1921 = w1595 | w1919 ;
  assign w1922 = ( w192 & w1919 ) | ( w192 & w1921 ) | ( w1919 & w1921 ) ;
  assign w1923 = ( w191 & ~w1920 ) | ( w191 & w1922 ) | ( ~w1920 & w1922 ) ;
  assign w1924 = \pi005 ^ w1923 ;
  assign w1925 = ( w1741 & w1843 ) | ( w1741 & w1855 ) | ( w1843 & w1855 ) ;
  assign w1926 = ~\pi070 & w1313 ;
  assign w1927 = \pi069 & w1417 ;
  assign w1928 = ( w1313 & ~w1926 ) | ( w1313 & w1927 ) | ( ~w1926 & w1927 ) ;
  assign w1929 = ~\pi071 & w1315 ;
  assign w1930 = w290 | w1928 ;
  assign w1931 = ( w1316 & w1928 ) | ( w1316 & w1930 ) | ( w1928 & w1930 ) ;
  assign w1932 = ( w1315 & ~w1929 ) | ( w1315 & w1931 ) | ( ~w1929 & w1931 ) ;
  assign w1933 = \pi023 ^ w1932 ;
  assign w1934 = ( w1731 & w1851 ) | ( w1731 & w1854 ) | ( w1851 & w1854 ) ;
  assign w1935 = ~\pi067 & w1629 ;
  assign w1936 = \pi066 & w1722 ;
  assign w1937 = ( w1629 & ~w1935 ) | ( w1629 & w1936 ) | ( ~w1935 & w1936 ) ;
  assign w1938 = ~\pi068 & w1631 ;
  assign w1939 = w182 | w1937 ;
  assign w1940 = ( w1632 & w1937 ) | ( w1632 & w1939 ) | ( w1937 & w1939 ) ;
  assign w1941 = ( w1631 & ~w1938 ) | ( w1631 & w1940 ) | ( ~w1938 & w1940 ) ;
  assign w1942 = \pi026 ^ w1941 ;
  assign w1943 = ( \pi026 & \pi027 ) | ( \pi026 & \pi028 ) | ( \pi027 & \pi028 ) ;
  assign w1944 = \pi028 ^ w1943 ;
  assign w1945 = \pi028 ^ \pi029 ;
  assign w1946 = w1853 & ~w1945 ;
  assign w1947 = w1853 & w1945 ;
  assign w1948 = ( \pi026 & \pi027 ) | ( \pi026 & ~\pi029 ) | ( \pi027 & ~\pi029 ) ;
  assign w1949 = \pi029 & ~\pi064 ;
  assign w1950 = ~\pi065 & w1949 ;
  assign w1951 = ( \pi026 & \pi027 ) | ( \pi026 & ~w1950 ) | ( \pi027 & ~w1950 ) ;
  assign w1952 = ( \pi028 & \pi029 ) | ( \pi028 & ~w1951 ) | ( \pi029 & ~w1951 ) ;
  assign w1953 = ( \pi028 & ~w1949 ) | ( \pi028 & w1951 ) | ( ~w1949 & w1951 ) ;
  assign w1954 = ( w1948 & w1952 ) | ( w1948 & ~w1953 ) | ( w1952 & ~w1953 ) ;
  assign w1955 = ( \pi026 & \pi027 ) | ( \pi026 & \pi065 ) | ( \pi027 & \pi065 ) ;
  assign w1956 = \pi026 & \pi027 ;
  assign w1957 = \pi064 ^ w1956 ;
  assign w1958 = ( \pi028 & w1956 ) | ( \pi028 & w1957 ) | ( w1956 & w1957 ) ;
  assign w1959 = w1955 ^ w1958 ;
  assign w1960 = w1934 ^ w1942 ;
  assign w1961 = w1959 ^ w1960 ;
  assign w1962 = w1925 ^ w1961 ;
  assign w1963 = w1933 ^ w1962 ;
  assign w1964 = ~\pi073 & w1044 ;
  assign w1965 = \pi072 & w1138 ;
  assign w1966 = ( w1044 & ~w1964 ) | ( w1044 & w1965 ) | ( ~w1964 & w1965 ) ;
  assign w1967 = ~\pi074 & w1046 ;
  assign w1968 = w465 | w1966 ;
  assign w1969 = ( w1047 & w1966 ) | ( w1047 & w1968 ) | ( w1966 & w1968 ) ;
  assign w1970 = ( w1046 & ~w1967 ) | ( w1046 & w1969 ) | ( ~w1967 & w1969 ) ;
  assign w1971 = \pi020 ^ w1970 ;
  assign w1972 = ( w1835 & w1857 ) | ( w1835 & w1865 ) | ( w1857 & w1865 ) ;
  assign w1973 = w1963 ^ w1972 ;
  assign w1974 = w1971 ^ w1973 ;
  assign w1975 = ~\pi076 & w837 ;
  assign w1976 = \pi075 & w902 ;
  assign w1977 = ( w837 & ~w1975 ) | ( w837 & w1976 ) | ( ~w1975 & w1976 ) ;
  assign w1978 = ~\pi077 & w839 ;
  assign w1979 = w644 | w1977 ;
  assign w1980 = ( w840 & w1977 ) | ( w840 & w1979 ) | ( w1977 & w1979 ) ;
  assign w1981 = ( w839 & ~w1978 ) | ( w839 & w1980 ) | ( ~w1978 & w1980 ) ;
  assign w1982 = \pi017 ^ w1981 ;
  assign w1983 = ( w1826 & w1834 ) | ( w1826 & w1867 ) | ( w1834 & w1867 ) ;
  assign w1984 = w1974 ^ w1983 ;
  assign w1985 = w1982 ^ w1984 ;
  assign w1986 = ~\pi079 & w601 ;
  assign w1987 = \pi078 & w683 ;
  assign w1988 = ( w601 & ~w1986 ) | ( w601 & w1987 ) | ( ~w1986 & w1987 ) ;
  assign w1989 = ~\pi080 & w603 ;
  assign w1990 = w794 | w1988 ;
  assign w1991 = ( w604 & w1988 ) | ( w604 & w1990 ) | ( w1988 & w1990 ) ;
  assign w1992 = ( w603 & ~w1989 ) | ( w603 & w1991 ) | ( ~w1989 & w1991 ) ;
  assign w1993 = \pi014 ^ w1992 ;
  assign w1994 = ( w1825 & w1869 ) | ( w1825 & w1870 ) | ( w1869 & w1870 ) ;
  assign w1995 = w1985 ^ w1994 ;
  assign w1996 = w1993 ^ w1995 ;
  assign w1997 = ~\pi082 & w432 ;
  assign w1998 = \pi081 & w486 ;
  assign w1999 = ( w432 & ~w1997 ) | ( w432 & w1998 ) | ( ~w1997 & w1998 ) ;
  assign w2000 = ~\pi083 & w434 ;
  assign w2001 = w1099 | w1999 ;
  assign w2002 = ( w435 & w1999 ) | ( w435 & w2001 ) | ( w1999 & w2001 ) ;
  assign w2003 = ( w434 & ~w2000 ) | ( w434 & w2002 ) | ( ~w2000 & w2002 ) ;
  assign w2004 = \pi011 ^ w2003 ;
  assign w2005 = ( w1872 & w1880 ) | ( w1872 & w1881 ) | ( w1880 & w1881 ) ;
  assign w2006 = w1996 ^ w2005 ;
  assign w2007 = w2004 ^ w2006 ;
  assign w2008 = ~\pi085 & w305 ;
  assign w2009 = \pi084 & w328 ;
  assign w2010 = ( w305 & ~w2008 ) | ( w305 & w2009 ) | ( ~w2008 & w2009 ) ;
  assign w2011 = ~\pi086 & w307 ;
  assign w2012 = w1379 | w2010 ;
  assign w2013 = ( w308 & w2010 ) | ( w308 & w2012 ) | ( w2010 & w2012 ) ;
  assign w2014 = ( w307 & ~w2011 ) | ( w307 & w2013 ) | ( ~w2011 & w2013 ) ;
  assign w2015 = \pi008 ^ w2014 ;
  assign w2016 = ( w1883 & w1891 ) | ( w1883 & w1892 ) | ( w1891 & w1892 ) ;
  assign w2017 = w2007 ^ w2016 ;
  assign w2018 = w2015 ^ w2017 ;
  assign w2019 = ( w1817 & w1894 ) | ( w1817 & w1895 ) | ( w1894 & w1895 ) ;
  assign w2020 = w2018 ^ w2019 ;
  assign w2021 = w1924 ^ w2020 ;
  assign w2022 = ( ~\pi002 & \pi091 ) | ( ~\pi002 & \pi092 ) | ( \pi091 & \pi092 ) ;
  assign w2023 = \pi000 ^ w2022 ;
  assign w2024 = ( \pi002 & \pi092 ) | ( \pi002 & ~w2023 ) | ( \pi092 & ~w2023 ) ;
  assign w2025 = ( \pi002 & \pi091 ) | ( \pi002 & w2023 ) | ( \pi091 & w2023 ) ;
  assign w2026 = \pi001 & w2025 ;
  assign w2027 = ( ~\pi000 & \pi090 ) | ( ~\pi000 & w2026 ) | ( \pi090 & w2026 ) ;
  assign w2028 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2027 ) | ( \pi002 & ~w2027 ) ;
  assign w2029 = ( w2024 & w2026 ) | ( w2024 & ~w2028 ) | ( w2026 & ~w2028 ) ;
  assign w2030 = ( \pi089 & ~\pi091 ) | ( \pi089 & w1799 ) | ( ~\pi091 & w1799 ) ;
  assign w2031 = ( ~\pi090 & \pi091 ) | ( ~\pi090 & w2030 ) | ( \pi091 & w2030 ) ;
  assign w2032 = \pi092 ^ w2030 ;
  assign w2033 = w2031 ^ w2032 ;
  assign w2034 = \pi002 ^ w2029 ;
  assign w2035 = \pi000 & ~w2029 ;
  assign w2036 = w2033 & w2035 ;
  assign w2037 = \pi001 ^ w2036 ;
  assign w2038 = ( \pi001 & w2034 ) | ( \pi001 & ~w2037 ) | ( w2034 & ~w2037 ) ;
  assign w2039 = w1916 ^ w2021 ;
  assign w2040 = w2038 ^ w2039 ;
  assign w2041 = ( w1924 & w2018 ) | ( w1924 & w2019 ) | ( w2018 & w2019 ) ;
  assign w2042 = ~\pi089 & w189 ;
  assign w2043 = \pi088 & w229 ;
  assign w2044 = ( w189 & ~w2042 ) | ( w189 & w2043 ) | ( ~w2042 & w2043 ) ;
  assign w2045 = ~\pi090 & w191 ;
  assign w2046 = w1801 | w2044 ;
  assign w2047 = ( w192 & w2044 ) | ( w192 & w2046 ) | ( w2044 & w2046 ) ;
  assign w2048 = ( w191 & ~w2045 ) | ( w191 & w2047 ) | ( ~w2045 & w2047 ) ;
  assign w2049 = \pi005 ^ w2048 ;
  assign w2050 = ( w1996 & w2004 ) | ( w1996 & w2005 ) | ( w2004 & w2005 ) ;
  assign w2051 = ~\pi077 & w837 ;
  assign w2052 = \pi076 & w902 ;
  assign w2053 = ( w837 & ~w2051 ) | ( w837 & w2052 ) | ( ~w2051 & w2052 ) ;
  assign w2054 = ~\pi078 & w839 ;
  assign w2055 = w665 | w2053 ;
  assign w2056 = ( w840 & w2053 ) | ( w840 & w2055 ) | ( w2053 & w2055 ) ;
  assign w2057 = ( w839 & ~w2054 ) | ( w839 & w2056 ) | ( ~w2054 & w2056 ) ;
  assign w2058 = \pi017 ^ w2057 ;
  assign w2059 = ( w1963 & w1971 ) | ( w1963 & w1972 ) | ( w1971 & w1972 ) ;
  assign w2060 = ~\pi074 & w1044 ;
  assign w2061 = \pi073 & w1138 ;
  assign w2062 = ( w1044 & ~w2060 ) | ( w1044 & w2061 ) | ( ~w2060 & w2061 ) ;
  assign w2063 = ~\pi075 & w1046 ;
  assign w2064 = w519 | w2062 ;
  assign w2065 = ( w1047 & w2062 ) | ( w1047 & w2064 ) | ( w2062 & w2064 ) ;
  assign w2066 = ( w1046 & ~w2063 ) | ( w1046 & w2065 ) | ( ~w2063 & w2065 ) ;
  assign w2067 = \pi020 ^ w2066 ;
  assign w2068 = ( w1925 & w1933 ) | ( w1925 & w1961 ) | ( w1933 & w1961 ) ;
  assign w2069 = ( w1934 & w1942 ) | ( w1934 & w1959 ) | ( w1942 & w1959 ) ;
  assign w2070 = ( \pi027 & ~\pi028 ) | ( \pi027 & \pi029 ) | ( ~\pi028 & \pi029 ) ;
  assign w2071 = ( \pi026 & \pi027 ) | ( \pi026 & w2070 ) | ( \pi027 & w2070 ) ;
  assign w2072 = w2070 ^ w2071 ;
  assign w2073 = \pi064 & w2072 ;
  assign w2074 = ( \pi066 & w1946 ) | ( \pi066 & w2073 ) | ( w1946 & w2073 ) ;
  assign w2075 = \pi065 | w2074 ;
  assign w2076 = ( w1944 & w2074 ) | ( w1944 & w2075 ) | ( w2074 & w2075 ) ;
  assign w2077 = w2073 | w2076 ;
  assign w2078 = ~w134 & w1947 ;
  assign w2079 = ( w1947 & w2077 ) | ( w1947 & ~w2078 ) | ( w2077 & ~w2078 ) ;
  assign w2080 = \pi029 ^ w2079 ;
  assign w2081 = w1954 & w2080 ;
  assign w2082 = w1954 ^ w2080 ;
  assign w2083 = ~\pi068 & w1629 ;
  assign w2084 = \pi067 & w1722 ;
  assign w2085 = ( w1629 & ~w2083 ) | ( w1629 & w2084 ) | ( ~w2083 & w2084 ) ;
  assign w2086 = ~\pi069 & w1631 ;
  assign w2087 = w221 | w2085 ;
  assign w2088 = ( w1632 & w2085 ) | ( w1632 & w2087 ) | ( w2085 & w2087 ) ;
  assign w2089 = ( w1631 & ~w2086 ) | ( w1631 & w2088 ) | ( ~w2086 & w2088 ) ;
  assign w2090 = \pi026 ^ w2089 ;
  assign w2091 = ( w2069 & w2082 ) | ( w2069 & w2090 ) | ( w2082 & w2090 ) ;
  assign w2092 = w2069 ^ w2082 ;
  assign w2093 = w2090 ^ w2092 ;
  assign w2094 = ~\pi071 & w1313 ;
  assign w2095 = \pi070 & w1417 ;
  assign w2096 = ( w1313 & ~w2094 ) | ( w1313 & w2095 ) | ( ~w2094 & w2095 ) ;
  assign w2097 = ~\pi072 & w1315 ;
  assign w2098 = w361 | w2096 ;
  assign w2099 = ( w1316 & w2096 ) | ( w1316 & w2098 ) | ( w2096 & w2098 ) ;
  assign w2100 = ( w1315 & ~w2097 ) | ( w1315 & w2099 ) | ( ~w2097 & w2099 ) ;
  assign w2101 = \pi023 ^ w2100 ;
  assign w2102 = w2068 ^ w2093 ;
  assign w2103 = w2101 ^ w2102 ;
  assign w2104 = w2059 ^ w2103 ;
  assign w2105 = w2067 ^ w2104 ;
  assign w2106 = ( w1974 & w1982 ) | ( w1974 & w1983 ) | ( w1982 & w1983 ) ;
  assign w2107 = w2105 ^ w2106 ;
  assign w2108 = w2058 ^ w2107 ;
  assign w2109 = ~\pi080 & w601 ;
  assign w2110 = \pi079 & w683 ;
  assign w2111 = ( w601 & ~w2109 ) | ( w601 & w2110 ) | ( ~w2109 & w2110 ) ;
  assign w2112 = ~\pi081 & w603 ;
  assign w2113 = w874 | w2111 ;
  assign w2114 = ( w604 & w2111 ) | ( w604 & w2113 ) | ( w2111 & w2113 ) ;
  assign w2115 = ( w603 & ~w2112 ) | ( w603 & w2114 ) | ( ~w2112 & w2114 ) ;
  assign w2116 = \pi014 ^ w2115 ;
  assign w2117 = ( w1985 & w1993 ) | ( w1985 & w1994 ) | ( w1993 & w1994 ) ;
  assign w2118 = w2108 ^ w2117 ;
  assign w2119 = w2116 ^ w2118 ;
  assign w2120 = ~\pi083 & w432 ;
  assign w2121 = \pi082 & w486 ;
  assign w2122 = ( w432 & ~w2120 ) | ( w432 & w2121 ) | ( ~w2120 & w2121 ) ;
  assign w2123 = ~\pi084 & w434 ;
  assign w2124 = w1188 | w2122 ;
  assign w2125 = ( w435 & w2122 ) | ( w435 & w2124 ) | ( w2122 & w2124 ) ;
  assign w2126 = ( w434 & ~w2123 ) | ( w434 & w2125 ) | ( ~w2123 & w2125 ) ;
  assign w2127 = \pi011 ^ w2126 ;
  assign w2128 = ( w2050 & w2119 ) | ( w2050 & w2127 ) | ( w2119 & w2127 ) ;
  assign w2129 = w2050 ^ w2119 ;
  assign w2130 = w2127 ^ w2129 ;
  assign w2131 = ~\pi086 & w305 ;
  assign w2132 = \pi085 & w328 ;
  assign w2133 = ( w305 & ~w2131 ) | ( w305 & w2132 ) | ( ~w2131 & w2132 ) ;
  assign w2134 = ~\pi087 & w307 ;
  assign w2135 = w1477 | w2133 ;
  assign w2136 = ( w308 & w2133 ) | ( w308 & w2135 ) | ( w2133 & w2135 ) ;
  assign w2137 = ( w307 & ~w2134 ) | ( w307 & w2136 ) | ( ~w2134 & w2136 ) ;
  assign w2138 = \pi008 ^ w2137 ;
  assign w2139 = ( w2007 & w2015 ) | ( w2007 & w2016 ) | ( w2015 & w2016 ) ;
  assign w2140 = w2130 ^ w2139 ;
  assign w2141 = w2138 ^ w2140 ;
  assign w2142 = w2041 ^ w2141 ;
  assign w2143 = w2049 ^ w2142 ;
  assign w2144 = ( ~\pi002 & \pi092 ) | ( ~\pi002 & \pi093 ) | ( \pi092 & \pi093 ) ;
  assign w2145 = \pi000 ^ w2144 ;
  assign w2146 = ( \pi002 & \pi093 ) | ( \pi002 & ~w2145 ) | ( \pi093 & ~w2145 ) ;
  assign w2147 = ( \pi002 & \pi092 ) | ( \pi002 & w2145 ) | ( \pi092 & w2145 ) ;
  assign w2148 = \pi001 & w2147 ;
  assign w2149 = ( ~\pi000 & \pi091 ) | ( ~\pi000 & w2148 ) | ( \pi091 & w2148 ) ;
  assign w2150 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2149 ) | ( \pi002 & ~w2149 ) ;
  assign w2151 = ( w2146 & w2148 ) | ( w2146 & ~w2150 ) | ( w2148 & ~w2150 ) ;
  assign w2152 = ( \pi090 & \pi091 ) | ( \pi090 & \pi092 ) | ( \pi091 & \pi092 ) ;
  assign w2153 = ( \pi091 & w1906 ) | ( \pi091 & w2152 ) | ( w1906 & w2152 ) ;
  assign w2154 = \pi092 ^ \pi093 ;
  assign w2155 = w2153 ^ w2154 ;
  assign w2156 = \pi002 ^ w2151 ;
  assign w2157 = \pi000 & ~w2151 ;
  assign w2158 = w2155 & w2157 ;
  assign w2159 = \pi001 ^ w2158 ;
  assign w2160 = ( \pi001 & w2156 ) | ( \pi001 & ~w2159 ) | ( w2156 & ~w2159 ) ;
  assign w2161 = ( w1916 & w2021 ) | ( w1916 & w2038 ) | ( w2021 & w2038 ) ;
  assign w2162 = w2143 ^ w2161 ;
  assign w2163 = w2160 ^ w2162 ;
  assign w2164 = ( w2130 & w2138 ) | ( w2130 & w2139 ) | ( w2138 & w2139 ) ;
  assign w2165 = ~\pi078 & w837 ;
  assign w2166 = \pi077 & w902 ;
  assign w2167 = ( w837 & ~w2165 ) | ( w837 & w2166 ) | ( ~w2165 & w2166 ) ;
  assign w2168 = ~\pi079 & w839 ;
  assign w2169 = w730 | w2167 ;
  assign w2170 = ( w840 & w2167 ) | ( w840 & w2169 ) | ( w2167 & w2169 ) ;
  assign w2171 = ( w839 & ~w2168 ) | ( w839 & w2170 ) | ( ~w2168 & w2170 ) ;
  assign w2172 = \pi017 ^ w2171 ;
  assign w2173 = ( w2059 & w2067 ) | ( w2059 & w2103 ) | ( w2067 & w2103 ) ;
  assign w2174 = ~\pi075 & w1044 ;
  assign w2175 = \pi074 & w1138 ;
  assign w2176 = ( w1044 & ~w2174 ) | ( w1044 & w2175 ) | ( ~w2174 & w2175 ) ;
  assign w2177 = ~\pi076 & w1046 ;
  assign w2178 = w538 | w2176 ;
  assign w2179 = ( w1047 & w2176 ) | ( w1047 & w2178 ) | ( w2176 & w2178 ) ;
  assign w2180 = ( w1046 & ~w2177 ) | ( w1046 & w2179 ) | ( ~w2177 & w2179 ) ;
  assign w2181 = \pi020 ^ w2180 ;
  assign w2182 = ( w2068 & w2093 ) | ( w2068 & w2101 ) | ( w2093 & w2101 ) ;
  assign w2183 = ~\pi069 & w1629 ;
  assign w2184 = \pi068 & w1722 ;
  assign w2185 = ( w1629 & ~w2183 ) | ( w1629 & w2184 ) | ( ~w2183 & w2184 ) ;
  assign w2186 = ~\pi070 & w1631 ;
  assign w2187 = w271 | w2185 ;
  assign w2188 = ( w1632 & w2185 ) | ( w1632 & w2187 ) | ( w2185 & w2187 ) ;
  assign w2189 = ( w1631 & ~w2186 ) | ( w1631 & w2188 ) | ( ~w2186 & w2188 ) ;
  assign w2190 = \pi026 ^ w2189 ;
  assign w2191 = ~\pi066 & w1944 ;
  assign w2192 = \pi065 & w2072 ;
  assign w2193 = ( w1944 & ~w2191 ) | ( w1944 & w2192 ) | ( ~w2191 & w2192 ) ;
  assign w2194 = ~\pi067 & w1946 ;
  assign w2195 = w160 | w2193 ;
  assign w2196 = ( w1947 & w2193 ) | ( w1947 & w2195 ) | ( w2193 & w2195 ) ;
  assign w2197 = ( w1946 & ~w2194 ) | ( w1946 & w2196 ) | ( ~w2194 & w2196 ) ;
  assign w2198 = \pi029 ^ w2197 ;
  assign w2199 = w2081 ^ w2198 ;
  assign w2200 = \pi029 ^ \pi030 ;
  assign w2201 = \pi064 & w2200 ;
  assign w2202 = w2199 ^ w2201 ;
  assign w2203 = w2091 ^ w2202 ;
  assign w2204 = w2190 ^ w2203 ;
  assign w2205 = ~\pi072 & w1313 ;
  assign w2206 = \pi071 & w1417 ;
  assign w2207 = ( w1313 & ~w2205 ) | ( w1313 & w2206 ) | ( ~w2205 & w2206 ) ;
  assign w2208 = ~\pi073 & w1315 ;
  assign w2209 = w404 | w2207 ;
  assign w2210 = ( w1316 & w2207 ) | ( w1316 & w2209 ) | ( w2207 & w2209 ) ;
  assign w2211 = ( w1315 & ~w2208 ) | ( w1315 & w2210 ) | ( ~w2208 & w2210 ) ;
  assign w2212 = \pi023 ^ w2211 ;
  assign w2213 = w2182 ^ w2204 ;
  assign w2214 = w2212 ^ w2213 ;
  assign w2215 = w2173 ^ w2214 ;
  assign w2216 = w2181 ^ w2215 ;
  assign w2217 = ( w2058 & w2105 ) | ( w2058 & w2106 ) | ( w2105 & w2106 ) ;
  assign w2218 = w2216 ^ w2217 ;
  assign w2219 = w2172 ^ w2218 ;
  assign w2220 = ~\pi081 & w601 ;
  assign w2221 = \pi080 & w683 ;
  assign w2222 = ( w601 & ~w2220 ) | ( w601 & w2221 ) | ( ~w2220 & w2221 ) ;
  assign w2223 = ~\pi082 & w603 ;
  assign w2224 = w1008 | w2222 ;
  assign w2225 = ( w604 & w2222 ) | ( w604 & w2224 ) | ( w2222 & w2224 ) ;
  assign w2226 = ( w603 & ~w2223 ) | ( w603 & w2225 ) | ( ~w2223 & w2225 ) ;
  assign w2227 = \pi014 ^ w2226 ;
  assign w2228 = ( w2108 & w2116 ) | ( w2108 & w2117 ) | ( w2116 & w2117 ) ;
  assign w2229 = w2219 ^ w2228 ;
  assign w2230 = w2227 ^ w2229 ;
  assign w2231 = ~\pi084 & w432 ;
  assign w2232 = \pi083 & w486 ;
  assign w2233 = ( w432 & ~w2231 ) | ( w432 & w2232 ) | ( ~w2231 & w2232 ) ;
  assign w2234 = ~\pi085 & w434 ;
  assign w2235 = w1274 | w2233 ;
  assign w2236 = ( w435 & w2233 ) | ( w435 & w2235 ) | ( w2233 & w2235 ) ;
  assign w2237 = ( w434 & ~w2234 ) | ( w434 & w2236 ) | ( ~w2234 & w2236 ) ;
  assign w2238 = \pi011 ^ w2237 ;
  assign w2239 = w2128 ^ w2230 ;
  assign w2240 = w2238 ^ w2239 ;
  assign w2241 = ~\pi087 & w305 ;
  assign w2242 = \pi086 & w328 ;
  assign w2243 = ( w305 & ~w2241 ) | ( w305 & w2242 ) | ( ~w2241 & w2242 ) ;
  assign w2244 = ~\pi088 & w307 ;
  assign w2245 = w1574 | w2243 ;
  assign w2246 = ( w308 & w2243 ) | ( w308 & w2245 ) | ( w2243 & w2245 ) ;
  assign w2247 = ( w307 & ~w2244 ) | ( w307 & w2246 ) | ( ~w2244 & w2246 ) ;
  assign w2248 = \pi008 ^ w2247 ;
  assign w2249 = w2164 ^ w2240 ;
  assign w2250 = w2248 ^ w2249 ;
  assign w2251 = ~\pi090 & w189 ;
  assign w2252 = \pi089 & w229 ;
  assign w2253 = ( w189 & ~w2251 ) | ( w189 & w2252 ) | ( ~w2251 & w2252 ) ;
  assign w2254 = ~\pi091 & w191 ;
  assign w2255 = w1908 | w2253 ;
  assign w2256 = ( w192 & w2253 ) | ( w192 & w2255 ) | ( w2253 & w2255 ) ;
  assign w2257 = ( w191 & ~w2254 ) | ( w191 & w2256 ) | ( ~w2254 & w2256 ) ;
  assign w2258 = \pi005 ^ w2257 ;
  assign w2259 = ( w2041 & w2049 ) | ( w2041 & w2141 ) | ( w2049 & w2141 ) ;
  assign w2260 = w2250 ^ w2259 ;
  assign w2261 = w2258 ^ w2260 ;
  assign w2262 = ( ~\pi002 & \pi093 ) | ( ~\pi002 & \pi094 ) | ( \pi093 & \pi094 ) ;
  assign w2263 = \pi000 ^ w2262 ;
  assign w2264 = ( \pi002 & \pi094 ) | ( \pi002 & ~w2263 ) | ( \pi094 & ~w2263 ) ;
  assign w2265 = ( \pi002 & \pi093 ) | ( \pi002 & w2263 ) | ( \pi093 & w2263 ) ;
  assign w2266 = \pi001 & w2265 ;
  assign w2267 = ( ~\pi000 & \pi092 ) | ( ~\pi000 & w2266 ) | ( \pi092 & w2266 ) ;
  assign w2268 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2267 ) | ( \pi002 & ~w2267 ) ;
  assign w2269 = ( w2264 & w2266 ) | ( w2264 & ~w2268 ) | ( w2266 & ~w2268 ) ;
  assign w2270 = ( \pi090 & \pi091 ) | ( \pi090 & ~\pi093 ) | ( \pi091 & ~\pi093 ) ;
  assign w2271 = ( \pi091 & w1906 ) | ( \pi091 & w2270 ) | ( w1906 & w2270 ) ;
  assign w2272 = ( \pi092 & \pi093 ) | ( \pi092 & w2271 ) | ( \pi093 & w2271 ) ;
  assign w2273 = \pi093 ^ w2272 ;
  assign w2274 = \pi094 ^ w2273 ;
  assign w2275 = \pi002 ^ w2269 ;
  assign w2276 = \pi000 & ~w2269 ;
  assign w2277 = w2274 & w2276 ;
  assign w2278 = \pi001 ^ w2277 ;
  assign w2279 = ( \pi001 & w2275 ) | ( \pi001 & ~w2278 ) | ( w2275 & ~w2278 ) ;
  assign w2280 = ( w2143 & w2160 ) | ( w2143 & w2161 ) | ( w2160 & w2161 ) ;
  assign w2281 = w2261 ^ w2280 ;
  assign w2282 = w2279 ^ w2281 ;
  assign w2283 = ~\pi079 & w837 ;
  assign w2284 = \pi078 & w902 ;
  assign w2285 = ( w837 & ~w2283 ) | ( w837 & w2284 ) | ( ~w2283 & w2284 ) ;
  assign w2286 = ~\pi080 & w839 ;
  assign w2287 = w794 | w2285 ;
  assign w2288 = ( w840 & w2285 ) | ( w840 & w2287 ) | ( w2285 & w2287 ) ;
  assign w2289 = ( w839 & ~w2286 ) | ( w839 & w2288 ) | ( ~w2286 & w2288 ) ;
  assign w2290 = \pi017 ^ w2289 ;
  assign w2291 = ( w2091 & w2190 ) | ( w2091 & w2202 ) | ( w2190 & w2202 ) ;
  assign w2292 = ~\pi070 & w1629 ;
  assign w2293 = \pi069 & w1722 ;
  assign w2294 = ( w1629 & ~w2292 ) | ( w1629 & w2293 ) | ( ~w2292 & w2293 ) ;
  assign w2295 = ~\pi071 & w1631 ;
  assign w2296 = w290 | w2294 ;
  assign w2297 = ( w1632 & w2294 ) | ( w1632 & w2296 ) | ( w2294 & w2296 ) ;
  assign w2298 = ( w1631 & ~w2295 ) | ( w1631 & w2297 ) | ( ~w2295 & w2297 ) ;
  assign w2299 = \pi026 ^ w2298 ;
  assign w2300 = ( w2081 & w2198 ) | ( w2081 & w2201 ) | ( w2198 & w2201 ) ;
  assign w2301 = ~\pi067 & w1944 ;
  assign w2302 = \pi066 & w2072 ;
  assign w2303 = ( w1944 & ~w2301 ) | ( w1944 & w2302 ) | ( ~w2301 & w2302 ) ;
  assign w2304 = ~\pi068 & w1946 ;
  assign w2305 = w182 | w2303 ;
  assign w2306 = ( w1947 & w2303 ) | ( w1947 & w2305 ) | ( w2303 & w2305 ) ;
  assign w2307 = ( w1946 & ~w2304 ) | ( w1946 & w2306 ) | ( ~w2304 & w2306 ) ;
  assign w2308 = \pi029 ^ w2307 ;
  assign w2309 = ( \pi029 & \pi030 ) | ( \pi029 & \pi031 ) | ( \pi030 & \pi031 ) ;
  assign w2310 = \pi031 ^ w2309 ;
  assign w2311 = \pi031 ^ \pi032 ;
  assign w2312 = w2200 & ~w2311 ;
  assign w2313 = w2200 & w2311 ;
  assign w2314 = ( \pi029 & \pi030 ) | ( \pi029 & ~\pi032 ) | ( \pi030 & ~\pi032 ) ;
  assign w2315 = \pi032 & ~\pi064 ;
  assign w2316 = ~\pi065 & w2315 ;
  assign w2317 = ( \pi029 & \pi030 ) | ( \pi029 & ~w2316 ) | ( \pi030 & ~w2316 ) ;
  assign w2318 = ( \pi031 & \pi032 ) | ( \pi031 & ~w2317 ) | ( \pi032 & ~w2317 ) ;
  assign w2319 = ( \pi031 & ~w2315 ) | ( \pi031 & w2317 ) | ( ~w2315 & w2317 ) ;
  assign w2320 = ( w2314 & w2318 ) | ( w2314 & ~w2319 ) | ( w2318 & ~w2319 ) ;
  assign w2321 = ( \pi029 & \pi030 ) | ( \pi029 & \pi065 ) | ( \pi030 & \pi065 ) ;
  assign w2322 = \pi029 & \pi030 ;
  assign w2323 = \pi064 ^ w2322 ;
  assign w2324 = ( \pi031 & w2322 ) | ( \pi031 & w2323 ) | ( w2322 & w2323 ) ;
  assign w2325 = w2321 ^ w2324 ;
  assign w2326 = w2300 ^ w2308 ;
  assign w2327 = w2325 ^ w2326 ;
  assign w2328 = w2291 ^ w2327 ;
  assign w2329 = w2299 ^ w2328 ;
  assign w2330 = ~\pi073 & w1313 ;
  assign w2331 = \pi072 & w1417 ;
  assign w2332 = ( w1313 & ~w2330 ) | ( w1313 & w2331 ) | ( ~w2330 & w2331 ) ;
  assign w2333 = ~\pi074 & w1315 ;
  assign w2334 = w465 | w2332 ;
  assign w2335 = ( w1316 & w2332 ) | ( w1316 & w2334 ) | ( w2332 & w2334 ) ;
  assign w2336 = ( w1315 & ~w2333 ) | ( w1315 & w2335 ) | ( ~w2333 & w2335 ) ;
  assign w2337 = \pi023 ^ w2336 ;
  assign w2338 = ( w2182 & w2204 ) | ( w2182 & w2212 ) | ( w2204 & w2212 ) ;
  assign w2339 = w2329 ^ w2338 ;
  assign w2340 = w2337 ^ w2339 ;
  assign w2341 = ~\pi076 & w1044 ;
  assign w2342 = \pi075 & w1138 ;
  assign w2343 = ( w1044 & ~w2341 ) | ( w1044 & w2342 ) | ( ~w2341 & w2342 ) ;
  assign w2344 = ~\pi077 & w1046 ;
  assign w2345 = w644 | w2343 ;
  assign w2346 = ( w1047 & w2343 ) | ( w1047 & w2345 ) | ( w2343 & w2345 ) ;
  assign w2347 = ( w1046 & ~w2344 ) | ( w1046 & w2346 ) | ( ~w2344 & w2346 ) ;
  assign w2348 = \pi020 ^ w2347 ;
  assign w2349 = ( w2173 & w2181 ) | ( w2173 & w2214 ) | ( w2181 & w2214 ) ;
  assign w2350 = w2340 ^ w2349 ;
  assign w2351 = w2348 ^ w2350 ;
  assign w2352 = ( w2172 & w2216 ) | ( w2172 & w2217 ) | ( w2216 & w2217 ) ;
  assign w2353 = w2351 ^ w2352 ;
  assign w2354 = w2290 ^ w2353 ;
  assign w2355 = ~\pi082 & w601 ;
  assign w2356 = \pi081 & w683 ;
  assign w2357 = ( w601 & ~w2355 ) | ( w601 & w2356 ) | ( ~w2355 & w2356 ) ;
  assign w2358 = ~\pi083 & w603 ;
  assign w2359 = w1099 | w2357 ;
  assign w2360 = ( w604 & w2357 ) | ( w604 & w2359 ) | ( w2357 & w2359 ) ;
  assign w2361 = ( w603 & ~w2358 ) | ( w603 & w2360 ) | ( ~w2358 & w2360 ) ;
  assign w2362 = \pi014 ^ w2361 ;
  assign w2363 = ( w2219 & w2227 ) | ( w2219 & w2228 ) | ( w2227 & w2228 ) ;
  assign w2364 = w2354 ^ w2363 ;
  assign w2365 = w2362 ^ w2364 ;
  assign w2366 = ~\pi085 & w432 ;
  assign w2367 = \pi084 & w486 ;
  assign w2368 = ( w432 & ~w2366 ) | ( w432 & w2367 ) | ( ~w2366 & w2367 ) ;
  assign w2369 = ~\pi086 & w434 ;
  assign w2370 = w1379 | w2368 ;
  assign w2371 = ( w435 & w2368 ) | ( w435 & w2370 ) | ( w2368 & w2370 ) ;
  assign w2372 = ( w434 & ~w2369 ) | ( w434 & w2371 ) | ( ~w2369 & w2371 ) ;
  assign w2373 = \pi011 ^ w2372 ;
  assign w2374 = ( w2128 & w2230 ) | ( w2128 & w2238 ) | ( w2230 & w2238 ) ;
  assign w2375 = w2365 ^ w2374 ;
  assign w2376 = w2373 ^ w2375 ;
  assign w2377 = ~\pi088 & w305 ;
  assign w2378 = \pi087 & w328 ;
  assign w2379 = ( w305 & ~w2377 ) | ( w305 & w2378 ) | ( ~w2377 & w2378 ) ;
  assign w2380 = ~\pi089 & w307 ;
  assign w2381 = w1595 | w2379 ;
  assign w2382 = ( w308 & w2379 ) | ( w308 & w2381 ) | ( w2379 & w2381 ) ;
  assign w2383 = ( w307 & ~w2380 ) | ( w307 & w2382 ) | ( ~w2380 & w2382 ) ;
  assign w2384 = \pi008 ^ w2383 ;
  assign w2385 = ( w2164 & w2240 ) | ( w2164 & w2248 ) | ( w2240 & w2248 ) ;
  assign w2386 = w2376 ^ w2385 ;
  assign w2387 = w2384 ^ w2386 ;
  assign w2388 = ~\pi091 & w189 ;
  assign w2389 = \pi090 & w229 ;
  assign w2390 = ( w189 & ~w2388 ) | ( w189 & w2389 ) | ( ~w2388 & w2389 ) ;
  assign w2391 = ~\pi092 & w191 ;
  assign w2392 = w2033 | w2390 ;
  assign w2393 = ( w192 & w2390 ) | ( w192 & w2392 ) | ( w2390 & w2392 ) ;
  assign w2394 = ( w191 & ~w2391 ) | ( w191 & w2393 ) | ( ~w2391 & w2393 ) ;
  assign w2395 = \pi005 ^ w2394 ;
  assign w2396 = ( w2250 & w2258 ) | ( w2250 & w2259 ) | ( w2258 & w2259 ) ;
  assign w2397 = w2387 ^ w2396 ;
  assign w2398 = w2395 ^ w2397 ;
  assign w2399 = ( ~\pi002 & \pi094 ) | ( ~\pi002 & \pi095 ) | ( \pi094 & \pi095 ) ;
  assign w2400 = \pi000 ^ w2399 ;
  assign w2401 = ( \pi002 & \pi095 ) | ( \pi002 & ~w2400 ) | ( \pi095 & ~w2400 ) ;
  assign w2402 = ( \pi002 & \pi094 ) | ( \pi002 & w2400 ) | ( \pi094 & w2400 ) ;
  assign w2403 = \pi001 & w2402 ;
  assign w2404 = ( ~\pi000 & \pi093 ) | ( ~\pi000 & w2403 ) | ( \pi093 & w2403 ) ;
  assign w2405 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2404 ) | ( \pi002 & ~w2404 ) ;
  assign w2406 = ( w2401 & w2403 ) | ( w2401 & ~w2405 ) | ( w2403 & ~w2405 ) ;
  assign w2407 = ( \pi093 & \pi094 ) | ( \pi093 & w2272 ) | ( \pi094 & w2272 ) ;
  assign w2408 = \pi094 ^ w2407 ;
  assign w2409 = \pi095 ^ w2408 ;
  assign w2410 = \pi002 ^ w2406 ;
  assign w2411 = \pi000 & ~w2406 ;
  assign w2412 = w2409 & w2411 ;
  assign w2413 = \pi001 ^ w2412 ;
  assign w2414 = ( \pi001 & w2410 ) | ( \pi001 & ~w2413 ) | ( w2410 & ~w2413 ) ;
  assign w2415 = ( w2261 & w2279 ) | ( w2261 & w2280 ) | ( w2279 & w2280 ) ;
  assign w2416 = w2398 ^ w2415 ;
  assign w2417 = w2414 ^ w2416 ;
  assign w2418 = ( w2398 & w2414 ) | ( w2398 & w2415 ) | ( w2414 & w2415 ) ;
  assign w2419 = ( w2387 & w2395 ) | ( w2387 & w2396 ) | ( w2395 & w2396 ) ;
  assign w2420 = ~\pi089 & w305 ;
  assign w2421 = \pi088 & w328 ;
  assign w2422 = ( w305 & ~w2420 ) | ( w305 & w2421 ) | ( ~w2420 & w2421 ) ;
  assign w2423 = ~\pi090 & w307 ;
  assign w2424 = w1801 | w2422 ;
  assign w2425 = ( w308 & w2422 ) | ( w308 & w2424 ) | ( w2422 & w2424 ) ;
  assign w2426 = ( w307 & ~w2423 ) | ( w307 & w2425 ) | ( ~w2423 & w2425 ) ;
  assign w2427 = \pi008 ^ w2426 ;
  assign w2428 = ( w2365 & w2373 ) | ( w2365 & w2374 ) | ( w2373 & w2374 ) ;
  assign w2429 = ( w2354 & w2362 ) | ( w2354 & w2363 ) | ( w2362 & w2363 ) ;
  assign w2430 = ~\pi080 & w837 ;
  assign w2431 = \pi079 & w902 ;
  assign w2432 = ( w837 & ~w2430 ) | ( w837 & w2431 ) | ( ~w2430 & w2431 ) ;
  assign w2433 = ~\pi081 & w839 ;
  assign w2434 = w874 | w2432 ;
  assign w2435 = ( w840 & w2432 ) | ( w840 & w2434 ) | ( w2432 & w2434 ) ;
  assign w2436 = ( w839 & ~w2433 ) | ( w839 & w2435 ) | ( ~w2433 & w2435 ) ;
  assign w2437 = \pi017 ^ w2436 ;
  assign w2438 = ( w2340 & w2348 ) | ( w2340 & w2349 ) | ( w2348 & w2349 ) ;
  assign w2439 = ( w2329 & w2337 ) | ( w2329 & w2338 ) | ( w2337 & w2338 ) ;
  assign w2440 = ( w2300 & w2308 ) | ( w2300 & w2325 ) | ( w2308 & w2325 ) ;
  assign w2441 = ( \pi030 & ~\pi031 ) | ( \pi030 & \pi032 ) | ( ~\pi031 & \pi032 ) ;
  assign w2442 = ( \pi029 & \pi030 ) | ( \pi029 & w2441 ) | ( \pi030 & w2441 ) ;
  assign w2443 = w2441 ^ w2442 ;
  assign w2444 = \pi064 & w2443 ;
  assign w2445 = ( \pi066 & w2312 ) | ( \pi066 & w2444 ) | ( w2312 & w2444 ) ;
  assign w2446 = \pi065 | w2445 ;
  assign w2447 = ( w2310 & w2445 ) | ( w2310 & w2446 ) | ( w2445 & w2446 ) ;
  assign w2448 = w2444 | w2447 ;
  assign w2449 = ~w134 & w2313 ;
  assign w2450 = ( w2313 & w2448 ) | ( w2313 & ~w2449 ) | ( w2448 & ~w2449 ) ;
  assign w2451 = \pi032 ^ w2450 ;
  assign w2452 = w2320 & w2451 ;
  assign w2453 = w2320 ^ w2451 ;
  assign w2454 = ~\pi068 & w1944 ;
  assign w2455 = \pi067 & w2072 ;
  assign w2456 = ( w1944 & ~w2454 ) | ( w1944 & w2455 ) | ( ~w2454 & w2455 ) ;
  assign w2457 = ~\pi069 & w1946 ;
  assign w2458 = w221 | w2456 ;
  assign w2459 = ( w1947 & w2456 ) | ( w1947 & w2458 ) | ( w2456 & w2458 ) ;
  assign w2460 = ( w1946 & ~w2457 ) | ( w1946 & w2459 ) | ( ~w2457 & w2459 ) ;
  assign w2461 = \pi029 ^ w2460 ;
  assign w2462 = ( w2440 & w2453 ) | ( w2440 & w2461 ) | ( w2453 & w2461 ) ;
  assign w2463 = w2440 ^ w2453 ;
  assign w2464 = w2461 ^ w2463 ;
  assign w2465 = ~\pi071 & w1629 ;
  assign w2466 = \pi070 & w1722 ;
  assign w2467 = ( w1629 & ~w2465 ) | ( w1629 & w2466 ) | ( ~w2465 & w2466 ) ;
  assign w2468 = ~\pi072 & w1631 ;
  assign w2469 = w361 | w2467 ;
  assign w2470 = ( w1632 & w2467 ) | ( w1632 & w2469 ) | ( w2467 & w2469 ) ;
  assign w2471 = ( w1631 & ~w2468 ) | ( w1631 & w2470 ) | ( ~w2468 & w2470 ) ;
  assign w2472 = \pi026 ^ w2471 ;
  assign w2473 = ( w2291 & w2299 ) | ( w2291 & w2327 ) | ( w2299 & w2327 ) ;
  assign w2474 = w2464 ^ w2473 ;
  assign w2475 = w2472 ^ w2474 ;
  assign w2476 = ~\pi074 & w1313 ;
  assign w2477 = \pi073 & w1417 ;
  assign w2478 = ( w1313 & ~w2476 ) | ( w1313 & w2477 ) | ( ~w2476 & w2477 ) ;
  assign w2479 = ~\pi075 & w1315 ;
  assign w2480 = w519 | w2478 ;
  assign w2481 = ( w1316 & w2478 ) | ( w1316 & w2480 ) | ( w2478 & w2480 ) ;
  assign w2482 = ( w1315 & ~w2479 ) | ( w1315 & w2481 ) | ( ~w2479 & w2481 ) ;
  assign w2483 = \pi023 ^ w2482 ;
  assign w2484 = ( w2439 & w2475 ) | ( w2439 & w2483 ) | ( w2475 & w2483 ) ;
  assign w2485 = w2439 ^ w2475 ;
  assign w2486 = w2483 ^ w2485 ;
  assign w2487 = ~\pi077 & w1044 ;
  assign w2488 = \pi076 & w1138 ;
  assign w2489 = ( w1044 & ~w2487 ) | ( w1044 & w2488 ) | ( ~w2487 & w2488 ) ;
  assign w2490 = ~\pi078 & w1046 ;
  assign w2491 = w665 | w2489 ;
  assign w2492 = ( w1047 & w2489 ) | ( w1047 & w2491 ) | ( w2489 & w2491 ) ;
  assign w2493 = ( w1046 & ~w2490 ) | ( w1046 & w2492 ) | ( ~w2490 & w2492 ) ;
  assign w2494 = \pi020 ^ w2493 ;
  assign w2495 = w2438 ^ w2486 ;
  assign w2496 = w2494 ^ w2495 ;
  assign w2497 = ( w2290 & w2351 ) | ( w2290 & w2352 ) | ( w2351 & w2352 ) ;
  assign w2498 = w2496 ^ w2497 ;
  assign w2499 = w2437 ^ w2498 ;
  assign w2500 = ~\pi083 & w601 ;
  assign w2501 = \pi082 & w683 ;
  assign w2502 = ( w601 & ~w2500 ) | ( w601 & w2501 ) | ( ~w2500 & w2501 ) ;
  assign w2503 = ~\pi084 & w603 ;
  assign w2504 = w1188 | w2502 ;
  assign w2505 = ( w604 & w2502 ) | ( w604 & w2504 ) | ( w2502 & w2504 ) ;
  assign w2506 = ( w603 & ~w2503 ) | ( w603 & w2505 ) | ( ~w2503 & w2505 ) ;
  assign w2507 = \pi014 ^ w2506 ;
  assign w2508 = ( w2429 & w2499 ) | ( w2429 & w2507 ) | ( w2499 & w2507 ) ;
  assign w2509 = w2429 ^ w2499 ;
  assign w2510 = w2507 ^ w2509 ;
  assign w2511 = ~\pi086 & w432 ;
  assign w2512 = \pi085 & w486 ;
  assign w2513 = ( w432 & ~w2511 ) | ( w432 & w2512 ) | ( ~w2511 & w2512 ) ;
  assign w2514 = ~\pi087 & w434 ;
  assign w2515 = w1477 | w2513 ;
  assign w2516 = ( w435 & w2513 ) | ( w435 & w2515 ) | ( w2513 & w2515 ) ;
  assign w2517 = ( w434 & ~w2514 ) | ( w434 & w2516 ) | ( ~w2514 & w2516 ) ;
  assign w2518 = \pi011 ^ w2517 ;
  assign w2519 = w2428 ^ w2510 ;
  assign w2520 = w2518 ^ w2519 ;
  assign w2521 = ( w2376 & w2384 ) | ( w2376 & w2385 ) | ( w2384 & w2385 ) ;
  assign w2522 = w2520 ^ w2521 ;
  assign w2523 = w2427 ^ w2522 ;
  assign w2524 = ~\pi092 & w189 ;
  assign w2525 = \pi091 & w229 ;
  assign w2526 = ( w189 & ~w2524 ) | ( w189 & w2525 ) | ( ~w2524 & w2525 ) ;
  assign w2527 = ~\pi093 & w191 ;
  assign w2528 = w2155 | w2526 ;
  assign w2529 = ( w192 & w2526 ) | ( w192 & w2528 ) | ( w2526 & w2528 ) ;
  assign w2530 = ( w191 & ~w2527 ) | ( w191 & w2529 ) | ( ~w2527 & w2529 ) ;
  assign w2531 = \pi005 ^ w2530 ;
  assign w2532 = ( w2419 & w2523 ) | ( w2419 & w2531 ) | ( w2523 & w2531 ) ;
  assign w2533 = w2419 ^ w2523 ;
  assign w2534 = w2531 ^ w2533 ;
  assign w2535 = ( ~\pi002 & \pi095 ) | ( ~\pi002 & \pi096 ) | ( \pi095 & \pi096 ) ;
  assign w2536 = \pi000 ^ w2535 ;
  assign w2537 = ( \pi002 & \pi096 ) | ( \pi002 & ~w2536 ) | ( \pi096 & ~w2536 ) ;
  assign w2538 = ( \pi002 & \pi095 ) | ( \pi002 & w2536 ) | ( \pi095 & w2536 ) ;
  assign w2539 = \pi001 & w2538 ;
  assign w2540 = ( ~\pi000 & \pi094 ) | ( ~\pi000 & w2539 ) | ( \pi094 & w2539 ) ;
  assign w2541 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2540 ) | ( \pi002 & ~w2540 ) ;
  assign w2542 = ( w2537 & w2539 ) | ( w2537 & ~w2541 ) | ( w2539 & ~w2541 ) ;
  assign w2543 = ( \pi093 & ~\pi095 ) | ( \pi093 & w2272 ) | ( ~\pi095 & w2272 ) ;
  assign w2544 = ( ~\pi094 & \pi095 ) | ( ~\pi094 & w2543 ) | ( \pi095 & w2543 ) ;
  assign w2545 = \pi096 ^ w2543 ;
  assign w2546 = w2544 ^ w2545 ;
  assign w2547 = \pi002 ^ w2542 ;
  assign w2548 = \pi000 & ~w2542 ;
  assign w2549 = w2546 & w2548 ;
  assign w2550 = \pi001 ^ w2549 ;
  assign w2551 = ( \pi001 & w2547 ) | ( \pi001 & ~w2550 ) | ( w2547 & ~w2550 ) ;
  assign w2552 = w2418 ^ w2534 ;
  assign w2553 = w2551 ^ w2552 ;
  assign w2554 = ( w2418 & w2534 ) | ( w2418 & w2551 ) | ( w2534 & w2551 ) ;
  assign w2555 = ~\pi090 & w305 ;
  assign w2556 = \pi089 & w328 ;
  assign w2557 = ( w305 & ~w2555 ) | ( w305 & w2556 ) | ( ~w2555 & w2556 ) ;
  assign w2558 = ~\pi091 & w307 ;
  assign w2559 = w1908 | w2557 ;
  assign w2560 = ( w308 & w2557 ) | ( w308 & w2559 ) | ( w2557 & w2559 ) ;
  assign w2561 = ( w307 & ~w2558 ) | ( w307 & w2560 ) | ( ~w2558 & w2560 ) ;
  assign w2562 = \pi008 ^ w2561 ;
  assign w2563 = ( w2428 & w2510 ) | ( w2428 & w2518 ) | ( w2510 & w2518 ) ;
  assign w2564 = ( w2437 & w2496 ) | ( w2437 & w2497 ) | ( w2496 & w2497 ) ;
  assign w2565 = ( w2438 & w2486 ) | ( w2438 & w2494 ) | ( w2486 & w2494 ) ;
  assign w2566 = ~\pi078 & w1044 ;
  assign w2567 = \pi077 & w1138 ;
  assign w2568 = ( w1044 & ~w2566 ) | ( w1044 & w2567 ) | ( ~w2566 & w2567 ) ;
  assign w2569 = ~\pi079 & w1046 ;
  assign w2570 = w730 | w2568 ;
  assign w2571 = ( w1047 & w2568 ) | ( w1047 & w2570 ) | ( w2568 & w2570 ) ;
  assign w2572 = ( w1046 & ~w2569 ) | ( w1046 & w2571 ) | ( ~w2569 & w2571 ) ;
  assign w2573 = \pi020 ^ w2572 ;
  assign w2574 = ( w2464 & w2472 ) | ( w2464 & w2473 ) | ( w2472 & w2473 ) ;
  assign w2575 = ~\pi069 & w1944 ;
  assign w2576 = \pi068 & w2072 ;
  assign w2577 = ( w1944 & ~w2575 ) | ( w1944 & w2576 ) | ( ~w2575 & w2576 ) ;
  assign w2578 = ~\pi070 & w1946 ;
  assign w2579 = w271 | w2577 ;
  assign w2580 = ( w1947 & w2577 ) | ( w1947 & w2579 ) | ( w2577 & w2579 ) ;
  assign w2581 = ( w1946 & ~w2578 ) | ( w1946 & w2580 ) | ( ~w2578 & w2580 ) ;
  assign w2582 = \pi029 ^ w2581 ;
  assign w2583 = ~\pi066 & w2310 ;
  assign w2584 = \pi065 & w2443 ;
  assign w2585 = ( w2310 & ~w2583 ) | ( w2310 & w2584 ) | ( ~w2583 & w2584 ) ;
  assign w2586 = ~\pi067 & w2312 ;
  assign w2587 = w160 | w2585 ;
  assign w2588 = ( w2313 & w2585 ) | ( w2313 & w2587 ) | ( w2585 & w2587 ) ;
  assign w2589 = ( w2312 & ~w2586 ) | ( w2312 & w2588 ) | ( ~w2586 & w2588 ) ;
  assign w2590 = \pi032 ^ w2589 ;
  assign w2591 = w2452 ^ w2590 ;
  assign w2592 = \pi032 ^ \pi033 ;
  assign w2593 = \pi064 & w2592 ;
  assign w2594 = w2591 ^ w2593 ;
  assign w2595 = w2462 ^ w2594 ;
  assign w2596 = w2582 ^ w2595 ;
  assign w2597 = ~\pi072 & w1629 ;
  assign w2598 = \pi071 & w1722 ;
  assign w2599 = ( w1629 & ~w2597 ) | ( w1629 & w2598 ) | ( ~w2597 & w2598 ) ;
  assign w2600 = ~\pi073 & w1631 ;
  assign w2601 = w404 | w2599 ;
  assign w2602 = ( w1632 & w2599 ) | ( w1632 & w2601 ) | ( w2599 & w2601 ) ;
  assign w2603 = ( w1631 & ~w2600 ) | ( w1631 & w2602 ) | ( ~w2600 & w2602 ) ;
  assign w2604 = \pi026 ^ w2603 ;
  assign w2605 = w2574 ^ w2596 ;
  assign w2606 = w2604 ^ w2605 ;
  assign w2607 = ~\pi075 & w1313 ;
  assign w2608 = \pi074 & w1417 ;
  assign w2609 = ( w1313 & ~w2607 ) | ( w1313 & w2608 ) | ( ~w2607 & w2608 ) ;
  assign w2610 = ~\pi076 & w1315 ;
  assign w2611 = w538 | w2609 ;
  assign w2612 = ( w1316 & w2609 ) | ( w1316 & w2611 ) | ( w2609 & w2611 ) ;
  assign w2613 = ( w1315 & ~w2610 ) | ( w1315 & w2612 ) | ( ~w2610 & w2612 ) ;
  assign w2614 = \pi023 ^ w2613 ;
  assign w2615 = w2484 ^ w2606 ;
  assign w2616 = w2614 ^ w2615 ;
  assign w2617 = w2565 ^ w2616 ;
  assign w2618 = w2573 ^ w2617 ;
  assign w2619 = ~\pi081 & w837 ;
  assign w2620 = \pi080 & w902 ;
  assign w2621 = ( w837 & ~w2619 ) | ( w837 & w2620 ) | ( ~w2619 & w2620 ) ;
  assign w2622 = ~\pi082 & w839 ;
  assign w2623 = w1008 | w2621 ;
  assign w2624 = ( w840 & w2621 ) | ( w840 & w2623 ) | ( w2621 & w2623 ) ;
  assign w2625 = ( w839 & ~w2622 ) | ( w839 & w2624 ) | ( ~w2622 & w2624 ) ;
  assign w2626 = \pi017 ^ w2625 ;
  assign w2627 = w2564 ^ w2618 ;
  assign w2628 = w2626 ^ w2627 ;
  assign w2629 = ~\pi084 & w601 ;
  assign w2630 = \pi083 & w683 ;
  assign w2631 = ( w601 & ~w2629 ) | ( w601 & w2630 ) | ( ~w2629 & w2630 ) ;
  assign w2632 = ~\pi085 & w603 ;
  assign w2633 = w1274 | w2631 ;
  assign w2634 = ( w604 & w2631 ) | ( w604 & w2633 ) | ( w2631 & w2633 ) ;
  assign w2635 = ( w603 & ~w2632 ) | ( w603 & w2634 ) | ( ~w2632 & w2634 ) ;
  assign w2636 = \pi014 ^ w2635 ;
  assign w2637 = w2508 ^ w2628 ;
  assign w2638 = w2636 ^ w2637 ;
  assign w2639 = ~\pi087 & w432 ;
  assign w2640 = \pi086 & w486 ;
  assign w2641 = ( w432 & ~w2639 ) | ( w432 & w2640 ) | ( ~w2639 & w2640 ) ;
  assign w2642 = ~\pi088 & w434 ;
  assign w2643 = w1574 | w2641 ;
  assign w2644 = ( w435 & w2641 ) | ( w435 & w2643 ) | ( w2641 & w2643 ) ;
  assign w2645 = ( w434 & ~w2642 ) | ( w434 & w2644 ) | ( ~w2642 & w2644 ) ;
  assign w2646 = \pi011 ^ w2645 ;
  assign w2647 = w2563 ^ w2638 ;
  assign w2648 = w2646 ^ w2647 ;
  assign w2649 = ( w2427 & w2520 ) | ( w2427 & w2521 ) | ( w2520 & w2521 ) ;
  assign w2650 = w2648 ^ w2649 ;
  assign w2651 = w2562 ^ w2650 ;
  assign w2652 = ~\pi093 & w189 ;
  assign w2653 = \pi092 & w229 ;
  assign w2654 = ( w189 & ~w2652 ) | ( w189 & w2653 ) | ( ~w2652 & w2653 ) ;
  assign w2655 = ~\pi094 & w191 ;
  assign w2656 = w2274 | w2654 ;
  assign w2657 = ( w192 & w2654 ) | ( w192 & w2656 ) | ( w2654 & w2656 ) ;
  assign w2658 = ( w191 & ~w2655 ) | ( w191 & w2657 ) | ( ~w2655 & w2657 ) ;
  assign w2659 = \pi005 ^ w2658 ;
  assign w2660 = w2532 ^ w2651 ;
  assign w2661 = w2659 ^ w2660 ;
  assign w2662 = ( ~\pi002 & \pi096 ) | ( ~\pi002 & \pi097 ) | ( \pi096 & \pi097 ) ;
  assign w2663 = \pi000 ^ w2662 ;
  assign w2664 = ( \pi002 & \pi097 ) | ( \pi002 & ~w2663 ) | ( \pi097 & ~w2663 ) ;
  assign w2665 = ( \pi002 & \pi096 ) | ( \pi002 & w2663 ) | ( \pi096 & w2663 ) ;
  assign w2666 = \pi001 & w2665 ;
  assign w2667 = ( ~\pi000 & \pi095 ) | ( ~\pi000 & w2666 ) | ( \pi095 & w2666 ) ;
  assign w2668 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2667 ) | ( \pi002 & ~w2667 ) ;
  assign w2669 = ( w2664 & w2666 ) | ( w2664 & ~w2668 ) | ( w2666 & ~w2668 ) ;
  assign w2670 = ( \pi094 & \pi095 ) | ( \pi094 & \pi096 ) | ( \pi095 & \pi096 ) ;
  assign w2671 = ( \pi095 & w2407 ) | ( \pi095 & w2670 ) | ( w2407 & w2670 ) ;
  assign w2672 = \pi096 ^ \pi097 ;
  assign w2673 = w2671 ^ w2672 ;
  assign w2674 = \pi002 ^ w2669 ;
  assign w2675 = \pi000 & ~w2669 ;
  assign w2676 = w2673 & w2675 ;
  assign w2677 = \pi001 ^ w2676 ;
  assign w2678 = ( \pi001 & w2674 ) | ( \pi001 & ~w2677 ) | ( w2674 & ~w2677 ) ;
  assign w2679 = w2554 ^ w2661 ;
  assign w2680 = w2678 ^ w2679 ;
  assign w2681 = ( w2554 & w2661 ) | ( w2554 & w2678 ) | ( w2661 & w2678 ) ;
  assign w2682 = ( w2532 & w2651 ) | ( w2532 & w2659 ) | ( w2651 & w2659 ) ;
  assign w2683 = ( w2563 & w2638 ) | ( w2563 & w2646 ) | ( w2638 & w2646 ) ;
  assign w2684 = ( w2484 & w2606 ) | ( w2484 & w2614 ) | ( w2606 & w2614 ) ;
  assign w2685 = ~\pi073 & w1629 ;
  assign w2686 = \pi072 & w1722 ;
  assign w2687 = ( w1629 & ~w2685 ) | ( w1629 & w2686 ) | ( ~w2685 & w2686 ) ;
  assign w2688 = ~\pi074 & w1631 ;
  assign w2689 = w465 | w2687 ;
  assign w2690 = ( w1632 & w2687 ) | ( w1632 & w2689 ) | ( w2687 & w2689 ) ;
  assign w2691 = ( w1631 & ~w2688 ) | ( w1631 & w2690 ) | ( ~w2688 & w2690 ) ;
  assign w2692 = \pi026 ^ w2691 ;
  assign w2693 = ( w2462 & w2582 ) | ( w2462 & w2594 ) | ( w2582 & w2594 ) ;
  assign w2694 = ~\pi070 & w1944 ;
  assign w2695 = \pi069 & w2072 ;
  assign w2696 = ( w1944 & ~w2694 ) | ( w1944 & w2695 ) | ( ~w2694 & w2695 ) ;
  assign w2697 = ~\pi071 & w1946 ;
  assign w2698 = w290 | w2696 ;
  assign w2699 = ( w1947 & w2696 ) | ( w1947 & w2698 ) | ( w2696 & w2698 ) ;
  assign w2700 = ( w1946 & ~w2697 ) | ( w1946 & w2699 ) | ( ~w2697 & w2699 ) ;
  assign w2701 = \pi029 ^ w2700 ;
  assign w2702 = ( w2452 & w2590 ) | ( w2452 & w2593 ) | ( w2590 & w2593 ) ;
  assign w2703 = ~\pi067 & w2310 ;
  assign w2704 = \pi066 & w2443 ;
  assign w2705 = ( w2310 & ~w2703 ) | ( w2310 & w2704 ) | ( ~w2703 & w2704 ) ;
  assign w2706 = ~\pi068 & w2312 ;
  assign w2707 = w182 | w2705 ;
  assign w2708 = ( w2313 & w2705 ) | ( w2313 & w2707 ) | ( w2705 & w2707 ) ;
  assign w2709 = ( w2312 & ~w2706 ) | ( w2312 & w2708 ) | ( ~w2706 & w2708 ) ;
  assign w2710 = \pi032 ^ w2709 ;
  assign w2711 = ( \pi032 & \pi033 ) | ( \pi032 & \pi034 ) | ( \pi033 & \pi034 ) ;
  assign w2712 = \pi034 ^ w2711 ;
  assign w2713 = \pi034 ^ \pi035 ;
  assign w2714 = w2592 & ~w2713 ;
  assign w2715 = w2592 & w2713 ;
  assign w2716 = ( \pi032 & \pi033 ) | ( \pi032 & ~\pi035 ) | ( \pi033 & ~\pi035 ) ;
  assign w2717 = \pi035 & ~\pi064 ;
  assign w2718 = ~\pi065 & w2717 ;
  assign w2719 = ( \pi032 & \pi033 ) | ( \pi032 & ~w2718 ) | ( \pi033 & ~w2718 ) ;
  assign w2720 = ( \pi034 & \pi035 ) | ( \pi034 & ~w2719 ) | ( \pi035 & ~w2719 ) ;
  assign w2721 = ( \pi034 & ~w2717 ) | ( \pi034 & w2719 ) | ( ~w2717 & w2719 ) ;
  assign w2722 = ( w2716 & w2720 ) | ( w2716 & ~w2721 ) | ( w2720 & ~w2721 ) ;
  assign w2723 = ( \pi032 & \pi033 ) | ( \pi032 & \pi065 ) | ( \pi033 & \pi065 ) ;
  assign w2724 = \pi032 & \pi033 ;
  assign w2725 = \pi064 ^ w2724 ;
  assign w2726 = ( \pi034 & w2724 ) | ( \pi034 & w2725 ) | ( w2724 & w2725 ) ;
  assign w2727 = w2723 ^ w2726 ;
  assign w2728 = w2702 ^ w2710 ;
  assign w2729 = w2727 ^ w2728 ;
  assign w2730 = w2693 ^ w2729 ;
  assign w2731 = w2701 ^ w2730 ;
  assign w2732 = ( w2574 & w2596 ) | ( w2574 & w2604 ) | ( w2596 & w2604 ) ;
  assign w2733 = w2731 ^ w2732 ;
  assign w2734 = w2692 ^ w2733 ;
  assign w2735 = ~\pi076 & w1313 ;
  assign w2736 = \pi075 & w1417 ;
  assign w2737 = ( w1313 & ~w2735 ) | ( w1313 & w2736 ) | ( ~w2735 & w2736 ) ;
  assign w2738 = ~\pi077 & w1315 ;
  assign w2739 = w644 | w2737 ;
  assign w2740 = ( w1316 & w2737 ) | ( w1316 & w2739 ) | ( w2737 & w2739 ) ;
  assign w2741 = ( w1315 & ~w2738 ) | ( w1315 & w2740 ) | ( ~w2738 & w2740 ) ;
  assign w2742 = \pi023 ^ w2741 ;
  assign w2743 = ( w2684 & w2734 ) | ( w2684 & w2742 ) | ( w2734 & w2742 ) ;
  assign w2744 = w2684 ^ w2734 ;
  assign w2745 = w2742 ^ w2744 ;
  assign w2746 = ~\pi079 & w1044 ;
  assign w2747 = \pi078 & w1138 ;
  assign w2748 = ( w1044 & ~w2746 ) | ( w1044 & w2747 ) | ( ~w2746 & w2747 ) ;
  assign w2749 = ~\pi080 & w1046 ;
  assign w2750 = w794 | w2748 ;
  assign w2751 = ( w1047 & w2748 ) | ( w1047 & w2750 ) | ( w2748 & w2750 ) ;
  assign w2752 = ( w1046 & ~w2749 ) | ( w1046 & w2751 ) | ( ~w2749 & w2751 ) ;
  assign w2753 = \pi020 ^ w2752 ;
  assign w2754 = ( w2565 & w2573 ) | ( w2565 & w2616 ) | ( w2573 & w2616 ) ;
  assign w2755 = w2745 ^ w2754 ;
  assign w2756 = w2753 ^ w2755 ;
  assign w2757 = ~\pi082 & w837 ;
  assign w2758 = \pi081 & w902 ;
  assign w2759 = ( w837 & ~w2757 ) | ( w837 & w2758 ) | ( ~w2757 & w2758 ) ;
  assign w2760 = ~\pi083 & w839 ;
  assign w2761 = w1099 | w2759 ;
  assign w2762 = ( w840 & w2759 ) | ( w840 & w2761 ) | ( w2759 & w2761 ) ;
  assign w2763 = ( w839 & ~w2760 ) | ( w839 & w2762 ) | ( ~w2760 & w2762 ) ;
  assign w2764 = \pi017 ^ w2763 ;
  assign w2765 = ( w2564 & w2618 ) | ( w2564 & w2626 ) | ( w2618 & w2626 ) ;
  assign w2766 = w2756 ^ w2765 ;
  assign w2767 = w2764 ^ w2766 ;
  assign w2768 = ~\pi085 & w601 ;
  assign w2769 = \pi084 & w683 ;
  assign w2770 = ( w601 & ~w2768 ) | ( w601 & w2769 ) | ( ~w2768 & w2769 ) ;
  assign w2771 = ~\pi086 & w603 ;
  assign w2772 = w1379 | w2770 ;
  assign w2773 = ( w604 & w2770 ) | ( w604 & w2772 ) | ( w2770 & w2772 ) ;
  assign w2774 = ( w603 & ~w2771 ) | ( w603 & w2773 ) | ( ~w2771 & w2773 ) ;
  assign w2775 = \pi014 ^ w2774 ;
  assign w2776 = ( w2508 & w2628 ) | ( w2508 & w2636 ) | ( w2628 & w2636 ) ;
  assign w2777 = w2767 ^ w2776 ;
  assign w2778 = w2775 ^ w2777 ;
  assign w2779 = ~\pi088 & w432 ;
  assign w2780 = \pi087 & w486 ;
  assign w2781 = ( w432 & ~w2779 ) | ( w432 & w2780 ) | ( ~w2779 & w2780 ) ;
  assign w2782 = ~\pi089 & w434 ;
  assign w2783 = w1595 | w2781 ;
  assign w2784 = ( w435 & w2781 ) | ( w435 & w2783 ) | ( w2781 & w2783 ) ;
  assign w2785 = ( w434 & ~w2782 ) | ( w434 & w2784 ) | ( ~w2782 & w2784 ) ;
  assign w2786 = \pi011 ^ w2785 ;
  assign w2787 = ( w2683 & w2778 ) | ( w2683 & w2786 ) | ( w2778 & w2786 ) ;
  assign w2788 = w2683 ^ w2778 ;
  assign w2789 = w2786 ^ w2788 ;
  assign w2790 = ~\pi091 & w305 ;
  assign w2791 = \pi090 & w328 ;
  assign w2792 = ( w305 & ~w2790 ) | ( w305 & w2791 ) | ( ~w2790 & w2791 ) ;
  assign w2793 = ~\pi092 & w307 ;
  assign w2794 = w2033 | w2792 ;
  assign w2795 = ( w308 & w2792 ) | ( w308 & w2794 ) | ( w2792 & w2794 ) ;
  assign w2796 = ( w307 & ~w2793 ) | ( w307 & w2795 ) | ( ~w2793 & w2795 ) ;
  assign w2797 = \pi008 ^ w2796 ;
  assign w2798 = ( w2562 & w2648 ) | ( w2562 & w2649 ) | ( w2648 & w2649 ) ;
  assign w2799 = w2789 ^ w2798 ;
  assign w2800 = w2797 ^ w2799 ;
  assign w2801 = ~\pi094 & w189 ;
  assign w2802 = \pi093 & w229 ;
  assign w2803 = ( w189 & ~w2801 ) | ( w189 & w2802 ) | ( ~w2801 & w2802 ) ;
  assign w2804 = ~\pi095 & w191 ;
  assign w2805 = w2409 | w2803 ;
  assign w2806 = ( w192 & w2803 ) | ( w192 & w2805 ) | ( w2803 & w2805 ) ;
  assign w2807 = ( w191 & ~w2804 ) | ( w191 & w2806 ) | ( ~w2804 & w2806 ) ;
  assign w2808 = \pi005 ^ w2807 ;
  assign w2809 = ( w2682 & w2800 ) | ( w2682 & w2808 ) | ( w2800 & w2808 ) ;
  assign w2810 = w2682 ^ w2800 ;
  assign w2811 = w2808 ^ w2810 ;
  assign w2812 = ( ~\pi002 & \pi097 ) | ( ~\pi002 & \pi098 ) | ( \pi097 & \pi098 ) ;
  assign w2813 = \pi000 ^ w2812 ;
  assign w2814 = ( \pi002 & \pi098 ) | ( \pi002 & ~w2813 ) | ( \pi098 & ~w2813 ) ;
  assign w2815 = ( \pi002 & \pi097 ) | ( \pi002 & w2813 ) | ( \pi097 & w2813 ) ;
  assign w2816 = \pi001 & w2815 ;
  assign w2817 = ( ~\pi000 & \pi096 ) | ( ~\pi000 & w2816 ) | ( \pi096 & w2816 ) ;
  assign w2818 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2817 ) | ( \pi002 & ~w2817 ) ;
  assign w2819 = ( w2814 & w2816 ) | ( w2814 & ~w2818 ) | ( w2816 & ~w2818 ) ;
  assign w2820 = ( \pi094 & \pi095 ) | ( \pi094 & ~\pi097 ) | ( \pi095 & ~\pi097 ) ;
  assign w2821 = ( \pi095 & w2407 ) | ( \pi095 & w2820 ) | ( w2407 & w2820 ) ;
  assign w2822 = ( \pi096 & \pi097 ) | ( \pi096 & w2821 ) | ( \pi097 & w2821 ) ;
  assign w2823 = \pi097 ^ w2822 ;
  assign w2824 = \pi098 ^ w2823 ;
  assign w2825 = \pi002 ^ w2819 ;
  assign w2826 = \pi000 & ~w2819 ;
  assign w2827 = w2824 & w2826 ;
  assign w2828 = \pi001 ^ w2827 ;
  assign w2829 = ( \pi001 & w2825 ) | ( \pi001 & ~w2828 ) | ( w2825 & ~w2828 ) ;
  assign w2830 = w2681 ^ w2811 ;
  assign w2831 = w2829 ^ w2830 ;
  assign w2832 = ( w2681 & w2811 ) | ( w2681 & w2829 ) | ( w2811 & w2829 ) ;
  assign w2833 = ~\pi092 & w305 ;
  assign w2834 = \pi091 & w328 ;
  assign w2835 = ( w305 & ~w2833 ) | ( w305 & w2834 ) | ( ~w2833 & w2834 ) ;
  assign w2836 = ~\pi093 & w307 ;
  assign w2837 = w2155 | w2835 ;
  assign w2838 = ( w308 & w2835 ) | ( w308 & w2837 ) | ( w2835 & w2837 ) ;
  assign w2839 = ( w307 & ~w2836 ) | ( w307 & w2838 ) | ( ~w2836 & w2838 ) ;
  assign w2840 = \pi008 ^ w2839 ;
  assign w2841 = ~\pi089 & w432 ;
  assign w2842 = \pi088 & w486 ;
  assign w2843 = ( w432 & ~w2841 ) | ( w432 & w2842 ) | ( ~w2841 & w2842 ) ;
  assign w2844 = ~\pi090 & w434 ;
  assign w2845 = w1801 | w2843 ;
  assign w2846 = ( w435 & w2843 ) | ( w435 & w2845 ) | ( w2843 & w2845 ) ;
  assign w2847 = ( w434 & ~w2844 ) | ( w434 & w2846 ) | ( ~w2844 & w2846 ) ;
  assign w2848 = \pi011 ^ w2847 ;
  assign w2849 = ( w2767 & w2775 ) | ( w2767 & w2776 ) | ( w2775 & w2776 ) ;
  assign w2850 = ( w2756 & w2764 ) | ( w2756 & w2765 ) | ( w2764 & w2765 ) ;
  assign w2851 = ~\pi080 & w1044 ;
  assign w2852 = \pi079 & w1138 ;
  assign w2853 = ( w1044 & ~w2851 ) | ( w1044 & w2852 ) | ( ~w2851 & w2852 ) ;
  assign w2854 = ~\pi081 & w1046 ;
  assign w2855 = w874 | w2853 ;
  assign w2856 = ( w1047 & w2853 ) | ( w1047 & w2855 ) | ( w2853 & w2855 ) ;
  assign w2857 = ( w1046 & ~w2854 ) | ( w1046 & w2856 ) | ( ~w2854 & w2856 ) ;
  assign w2858 = \pi020 ^ w2857 ;
  assign w2859 = ( w2692 & w2731 ) | ( w2692 & w2732 ) | ( w2731 & w2732 ) ;
  assign w2860 = ~\pi074 & w1629 ;
  assign w2861 = \pi073 & w1722 ;
  assign w2862 = ( w1629 & ~w2860 ) | ( w1629 & w2861 ) | ( ~w2860 & w2861 ) ;
  assign w2863 = ~\pi075 & w1631 ;
  assign w2864 = w519 | w2862 ;
  assign w2865 = ( w1632 & w2862 ) | ( w1632 & w2864 ) | ( w2862 & w2864 ) ;
  assign w2866 = ( w1631 & ~w2863 ) | ( w1631 & w2865 ) | ( ~w2863 & w2865 ) ;
  assign w2867 = \pi026 ^ w2866 ;
  assign w2868 = ( w2693 & w2701 ) | ( w2693 & w2729 ) | ( w2701 & w2729 ) ;
  assign w2869 = ( w2702 & w2710 ) | ( w2702 & w2727 ) | ( w2710 & w2727 ) ;
  assign w2870 = ( \pi033 & ~\pi034 ) | ( \pi033 & \pi035 ) | ( ~\pi034 & \pi035 ) ;
  assign w2871 = ( \pi032 & \pi033 ) | ( \pi032 & w2870 ) | ( \pi033 & w2870 ) ;
  assign w2872 = w2870 ^ w2871 ;
  assign w2873 = \pi064 & w2872 ;
  assign w2874 = ( \pi066 & w2714 ) | ( \pi066 & w2873 ) | ( w2714 & w2873 ) ;
  assign w2875 = \pi065 | w2874 ;
  assign w2876 = ( w2712 & w2874 ) | ( w2712 & w2875 ) | ( w2874 & w2875 ) ;
  assign w2877 = w2873 | w2876 ;
  assign w2878 = ~w134 & w2715 ;
  assign w2879 = ( w2715 & w2877 ) | ( w2715 & ~w2878 ) | ( w2877 & ~w2878 ) ;
  assign w2880 = \pi035 ^ w2879 ;
  assign w2881 = w2722 & w2880 ;
  assign w2882 = w2722 ^ w2880 ;
  assign w2883 = ~\pi068 & w2310 ;
  assign w2884 = \pi067 & w2443 ;
  assign w2885 = ( w2310 & ~w2883 ) | ( w2310 & w2884 ) | ( ~w2883 & w2884 ) ;
  assign w2886 = ~\pi069 & w2312 ;
  assign w2887 = w221 | w2885 ;
  assign w2888 = ( w2313 & w2885 ) | ( w2313 & w2887 ) | ( w2885 & w2887 ) ;
  assign w2889 = ( w2312 & ~w2886 ) | ( w2312 & w2888 ) | ( ~w2886 & w2888 ) ;
  assign w2890 = \pi032 ^ w2889 ;
  assign w2891 = ( w2869 & w2882 ) | ( w2869 & w2890 ) | ( w2882 & w2890 ) ;
  assign w2892 = w2869 ^ w2882 ;
  assign w2893 = w2890 ^ w2892 ;
  assign w2894 = ~\pi071 & w1944 ;
  assign w2895 = \pi070 & w2072 ;
  assign w2896 = ( w1944 & ~w2894 ) | ( w1944 & w2895 ) | ( ~w2894 & w2895 ) ;
  assign w2897 = ~\pi072 & w1946 ;
  assign w2898 = w361 | w2896 ;
  assign w2899 = ( w1947 & w2896 ) | ( w1947 & w2898 ) | ( w2896 & w2898 ) ;
  assign w2900 = ( w1946 & ~w2897 ) | ( w1946 & w2899 ) | ( ~w2897 & w2899 ) ;
  assign w2901 = \pi029 ^ w2900 ;
  assign w2902 = w2868 ^ w2893 ;
  assign w2903 = w2901 ^ w2902 ;
  assign w2904 = w2859 ^ w2903 ;
  assign w2905 = w2867 ^ w2904 ;
  assign w2906 = ~\pi077 & w1313 ;
  assign w2907 = \pi076 & w1417 ;
  assign w2908 = ( w1313 & ~w2906 ) | ( w1313 & w2907 ) | ( ~w2906 & w2907 ) ;
  assign w2909 = ~\pi078 & w1315 ;
  assign w2910 = w665 | w2908 ;
  assign w2911 = ( w1316 & w2908 ) | ( w1316 & w2910 ) | ( w2908 & w2910 ) ;
  assign w2912 = ( w1315 & ~w2909 ) | ( w1315 & w2911 ) | ( ~w2909 & w2911 ) ;
  assign w2913 = \pi023 ^ w2912 ;
  assign w2914 = w2743 ^ w2905 ;
  assign w2915 = w2913 ^ w2914 ;
  assign w2916 = ( w2745 & w2753 ) | ( w2745 & w2754 ) | ( w2753 & w2754 ) ;
  assign w2917 = w2915 ^ w2916 ;
  assign w2918 = w2858 ^ w2917 ;
  assign w2919 = ~\pi083 & w837 ;
  assign w2920 = \pi082 & w902 ;
  assign w2921 = ( w837 & ~w2919 ) | ( w837 & w2920 ) | ( ~w2919 & w2920 ) ;
  assign w2922 = ~\pi084 & w839 ;
  assign w2923 = w1188 | w2921 ;
  assign w2924 = ( w840 & w2921 ) | ( w840 & w2923 ) | ( w2921 & w2923 ) ;
  assign w2925 = ( w839 & ~w2922 ) | ( w839 & w2924 ) | ( ~w2922 & w2924 ) ;
  assign w2926 = \pi017 ^ w2925 ;
  assign w2927 = ( w2850 & w2918 ) | ( w2850 & w2926 ) | ( w2918 & w2926 ) ;
  assign w2928 = w2850 ^ w2918 ;
  assign w2929 = w2926 ^ w2928 ;
  assign w2930 = ~\pi086 & w601 ;
  assign w2931 = \pi085 & w683 ;
  assign w2932 = ( w601 & ~w2930 ) | ( w601 & w2931 ) | ( ~w2930 & w2931 ) ;
  assign w2933 = ~\pi087 & w603 ;
  assign w2934 = w1477 | w2932 ;
  assign w2935 = ( w604 & w2932 ) | ( w604 & w2934 ) | ( w2932 & w2934 ) ;
  assign w2936 = ( w603 & ~w2933 ) | ( w603 & w2935 ) | ( ~w2933 & w2935 ) ;
  assign w2937 = \pi014 ^ w2936 ;
  assign w2938 = w2849 ^ w2929 ;
  assign w2939 = w2937 ^ w2938 ;
  assign w2940 = w2787 ^ w2939 ;
  assign w2941 = w2848 ^ w2940 ;
  assign w2942 = ( w2789 & w2797 ) | ( w2789 & w2798 ) | ( w2797 & w2798 ) ;
  assign w2943 = w2941 ^ w2942 ;
  assign w2944 = w2840 ^ w2943 ;
  assign w2945 = ~\pi095 & w189 ;
  assign w2946 = \pi094 & w229 ;
  assign w2947 = ( w189 & ~w2945 ) | ( w189 & w2946 ) | ( ~w2945 & w2946 ) ;
  assign w2948 = ~\pi096 & w191 ;
  assign w2949 = w2546 | w2947 ;
  assign w2950 = ( w192 & w2947 ) | ( w192 & w2949 ) | ( w2947 & w2949 ) ;
  assign w2951 = ( w191 & ~w2948 ) | ( w191 & w2950 ) | ( ~w2948 & w2950 ) ;
  assign w2952 = \pi005 ^ w2951 ;
  assign w2953 = ( w2809 & w2944 ) | ( w2809 & w2952 ) | ( w2944 & w2952 ) ;
  assign w2954 = w2809 ^ w2944 ;
  assign w2955 = w2952 ^ w2954 ;
  assign w2956 = ( ~\pi002 & \pi098 ) | ( ~\pi002 & \pi099 ) | ( \pi098 & \pi099 ) ;
  assign w2957 = \pi000 ^ w2956 ;
  assign w2958 = ( \pi002 & \pi099 ) | ( \pi002 & ~w2957 ) | ( \pi099 & ~w2957 ) ;
  assign w2959 = ( \pi002 & \pi098 ) | ( \pi002 & w2957 ) | ( \pi098 & w2957 ) ;
  assign w2960 = \pi001 & w2959 ;
  assign w2961 = ( ~\pi000 & \pi097 ) | ( ~\pi000 & w2960 ) | ( \pi097 & w2960 ) ;
  assign w2962 = ( \pi001 & \pi002 ) | ( \pi001 & ~w2961 ) | ( \pi002 & ~w2961 ) ;
  assign w2963 = ( w2958 & w2960 ) | ( w2958 & ~w2962 ) | ( w2960 & ~w2962 ) ;
  assign w2964 = ( \pi097 & \pi098 ) | ( \pi097 & w2822 ) | ( \pi098 & w2822 ) ;
  assign w2965 = \pi098 ^ w2964 ;
  assign w2966 = \pi099 ^ w2965 ;
  assign w2967 = \pi002 ^ w2963 ;
  assign w2968 = \pi000 & ~w2963 ;
  assign w2969 = w2966 & w2968 ;
  assign w2970 = \pi001 ^ w2969 ;
  assign w2971 = ( \pi001 & w2967 ) | ( \pi001 & ~w2970 ) | ( w2967 & ~w2970 ) ;
  assign w2972 = w2832 ^ w2955 ;
  assign w2973 = w2971 ^ w2972 ;
  assign w2974 = ~\pi096 & w189 ;
  assign w2975 = \pi095 & w229 ;
  assign w2976 = ( w189 & ~w2974 ) | ( w189 & w2975 ) | ( ~w2974 & w2975 ) ;
  assign w2977 = ~\pi097 & w191 ;
  assign w2978 = w2673 | w2976 ;
  assign w2979 = ( w192 & w2976 ) | ( w192 & w2978 ) | ( w2976 & w2978 ) ;
  assign w2980 = ( w191 & ~w2977 ) | ( w191 & w2979 ) | ( ~w2977 & w2979 ) ;
  assign w2981 = \pi005 ^ w2980 ;
  assign w2982 = ( w2840 & w2941 ) | ( w2840 & w2942 ) | ( w2941 & w2942 ) ;
  assign w2983 = ( w2787 & w2848 ) | ( w2787 & w2939 ) | ( w2848 & w2939 ) ;
  assign w2984 = ~\pi090 & w432 ;
  assign w2985 = \pi089 & w486 ;
  assign w2986 = ( w432 & ~w2984 ) | ( w432 & w2985 ) | ( ~w2984 & w2985 ) ;
  assign w2987 = ~\pi091 & w434 ;
  assign w2988 = w1908 | w2986 ;
  assign w2989 = ( w435 & w2986 ) | ( w435 & w2988 ) | ( w2986 & w2988 ) ;
  assign w2990 = ( w434 & ~w2987 ) | ( w434 & w2989 ) | ( ~w2987 & w2989 ) ;
  assign w2991 = \pi011 ^ w2990 ;
  assign w2992 = ( w2849 & w2929 ) | ( w2849 & w2937 ) | ( w2929 & w2937 ) ;
  assign w2993 = ( w2858 & w2915 ) | ( w2858 & w2916 ) | ( w2915 & w2916 ) ;
  assign w2994 = ( w2743 & w2905 ) | ( w2743 & w2913 ) | ( w2905 & w2913 ) ;
  assign w2995 = ~\pi078 & w1313 ;
  assign w2996 = \pi077 & w1417 ;
  assign w2997 = ( w1313 & ~w2995 ) | ( w1313 & w2996 ) | ( ~w2995 & w2996 ) ;
  assign w2998 = ~\pi079 & w1315 ;
  assign w2999 = w730 | w2997 ;
  assign w3000 = ( w1316 & w2997 ) | ( w1316 & w2999 ) | ( w2997 & w2999 ) ;
  assign w3001 = ( w1315 & ~w2998 ) | ( w1315 & w3000 ) | ( ~w2998 & w3000 ) ;
  assign w3002 = \pi023 ^ w3001 ;
  assign w3003 = ( w2868 & w2893 ) | ( w2868 & w2901 ) | ( w2893 & w2901 ) ;
  assign w3004 = ~\pi069 & w2310 ;
  assign w3005 = \pi068 & w2443 ;
  assign w3006 = ( w2310 & ~w3004 ) | ( w2310 & w3005 ) | ( ~w3004 & w3005 ) ;
  assign w3007 = ~\pi070 & w2312 ;
  assign w3008 = w271 | w3006 ;
  assign w3009 = ( w2313 & w3006 ) | ( w2313 & w3008 ) | ( w3006 & w3008 ) ;
  assign w3010 = ( w2312 & ~w3007 ) | ( w2312 & w3009 ) | ( ~w3007 & w3009 ) ;
  assign w3011 = \pi032 ^ w3010 ;
  assign w3012 = ~\pi066 & w2712 ;
  assign w3013 = \pi065 & w2872 ;
  assign w3014 = ( w2712 & ~w3012 ) | ( w2712 & w3013 ) | ( ~w3012 & w3013 ) ;
  assign w3015 = ~\pi067 & w2714 ;
  assign w3016 = w160 | w3014 ;
  assign w3017 = ( w2715 & w3014 ) | ( w2715 & w3016 ) | ( w3014 & w3016 ) ;
  assign w3018 = ( w2714 & ~w3015 ) | ( w2714 & w3017 ) | ( ~w3015 & w3017 ) ;
  assign w3019 = \pi035 ^ w3018 ;
  assign w3020 = w2881 ^ w3019 ;
  assign w3021 = \pi035 ^ \pi036 ;
  assign w3022 = \pi064 & w3021 ;
  assign w3023 = w3020 ^ w3022 ;
  assign w3024 = w2891 ^ w3023 ;
  assign w3025 = w3011 ^ w3024 ;
  assign w3026 = ~\pi072 & w1944 ;
  assign w3027 = \pi071 & w2072 ;
  assign w3028 = ( w1944 & ~w3026 ) | ( w1944 & w3027 ) | ( ~w3026 & w3027 ) ;
  assign w3029 = ~\pi073 & w1946 ;
  assign w3030 = w404 | w3028 ;
  assign w3031 = ( w1947 & w3028 ) | ( w1947 & w3030 ) | ( w3028 & w3030 ) ;
  assign w3032 = ( w1946 & ~w3029 ) | ( w1946 & w3031 ) | ( ~w3029 & w3031 ) ;
  assign w3033 = \pi029 ^ w3032 ;
  assign w3034 = w3003 ^ w3025 ;
  assign w3035 = w3033 ^ w3034 ;
  assign w3036 = ~\pi075 & w1629 ;
  assign w3037 = \pi074 & w1722 ;
  assign w3038 = ( w1629 & ~w3036 ) | ( w1629 & w3037 ) | ( ~w3036 & w3037 ) ;
  assign w3039 = ~\pi076 & w1631 ;
  assign w3040 = w538 | w3038 ;
  assign w3041 = ( w1632 & w3038 ) | ( w1632 & w3040 ) | ( w3038 & w3040 ) ;
  assign w3042 = ( w1631 & ~w3039 ) | ( w1631 & w3041 ) | ( ~w3039 & w3041 ) ;
  assign w3043 = \pi026 ^ w3042 ;
  assign w3044 = ( w2859 & w2867 ) | ( w2859 & w2903 ) | ( w2867 & w2903 ) ;
  assign w3045 = w3035 ^ w3044 ;
  assign w3046 = w3043 ^ w3045 ;
  assign w3047 = w2994 ^ w3046 ;
  assign w3048 = w3002 ^ w3047 ;
  assign w3049 = ~\pi081 & w1044 ;
  assign w3050 = \pi080 & w1138 ;
  assign w3051 = ( w1044 & ~w3049 ) | ( w1044 & w3050 ) | ( ~w3049 & w3050 ) ;
  assign w3052 = ~\pi082 & w1046 ;
  assign w3053 = w1008 | w3051 ;
  assign w3054 = ( w1047 & w3051 ) | ( w1047 & w3053 ) | ( w3051 & w3053 ) ;
  assign w3055 = ( w1046 & ~w3052 ) | ( w1046 & w3054 ) | ( ~w3052 & w3054 ) ;
  assign w3056 = \pi020 ^ w3055 ;
  assign w3057 = w2993 ^ w3048 ;
  assign w3058 = w3056 ^ w3057 ;
  assign w3059 = ~\pi084 & w837 ;
  assign w3060 = \pi083 & w902 ;
  assign w3061 = ( w837 & ~w3059 ) | ( w837 & w3060 ) | ( ~w3059 & w3060 ) ;
  assign w3062 = ~\pi085 & w839 ;
  assign w3063 = w1274 | w3061 ;
  assign w3064 = ( w840 & w3061 ) | ( w840 & w3063 ) | ( w3061 & w3063 ) ;
  assign w3065 = ( w839 & ~w3062 ) | ( w839 & w3064 ) | ( ~w3062 & w3064 ) ;
  assign w3066 = \pi017 ^ w3065 ;
  assign w3067 = w2927 ^ w3058 ;
  assign w3068 = w3066 ^ w3067 ;
  assign w3069 = ~\pi087 & w601 ;
  assign w3070 = \pi086 & w683 ;
  assign w3071 = ( w601 & ~w3069 ) | ( w601 & w3070 ) | ( ~w3069 & w3070 ) ;
  assign w3072 = ~\pi088 & w603 ;
  assign w3073 = w1574 | w3071 ;
  assign w3074 = ( w604 & w3071 ) | ( w604 & w3073 ) | ( w3071 & w3073 ) ;
  assign w3075 = ( w603 & ~w3072 ) | ( w603 & w3074 ) | ( ~w3072 & w3074 ) ;
  assign w3076 = \pi014 ^ w3075 ;
  assign w3077 = w2992 ^ w3068 ;
  assign w3078 = w3076 ^ w3077 ;
  assign w3079 = w2983 ^ w3078 ;
  assign w3080 = w2991 ^ w3079 ;
  assign w3081 = ~\pi093 & w305 ;
  assign w3082 = \pi092 & w328 ;
  assign w3083 = ( w305 & ~w3081 ) | ( w305 & w3082 ) | ( ~w3081 & w3082 ) ;
  assign w3084 = ~\pi094 & w307 ;
  assign w3085 = w2274 | w3083 ;
  assign w3086 = ( w308 & w3083 ) | ( w308 & w3085 ) | ( w3083 & w3085 ) ;
  assign w3087 = ( w307 & ~w3084 ) | ( w307 & w3086 ) | ( ~w3084 & w3086 ) ;
  assign w3088 = \pi008 ^ w3087 ;
  assign w3089 = w2982 ^ w3080 ;
  assign w3090 = w3088 ^ w3089 ;
  assign w3091 = w2953 ^ w3090 ;
  assign w3092 = w2981 ^ w3091 ;
  assign w3093 = ( ~\pi002 & \pi099 ) | ( ~\pi002 & \pi100 ) | ( \pi099 & \pi100 ) ;
  assign w3094 = \pi000 ^ w3093 ;
  assign w3095 = ( \pi002 & \pi100 ) | ( \pi002 & ~w3094 ) | ( \pi100 & ~w3094 ) ;
  assign w3096 = ( \pi002 & \pi099 ) | ( \pi002 & w3094 ) | ( \pi099 & w3094 ) ;
  assign w3097 = \pi001 & w3096 ;
  assign w3098 = ( ~\pi000 & \pi098 ) | ( ~\pi000 & w3097 ) | ( \pi098 & w3097 ) ;
  assign w3099 = ( \pi001 & \pi002 ) | ( \pi001 & ~w3098 ) | ( \pi002 & ~w3098 ) ;
  assign w3100 = ( w3095 & w3097 ) | ( w3095 & ~w3099 ) | ( w3097 & ~w3099 ) ;
  assign w3101 = ( \pi097 & ~\pi099 ) | ( \pi097 & w2822 ) | ( ~\pi099 & w2822 ) ;
  assign w3102 = ( ~\pi098 & \pi099 ) | ( ~\pi098 & w3101 ) | ( \pi099 & w3101 ) ;
  assign w3103 = \pi100 ^ w3101 ;
  assign w3104 = w3102 ^ w3103 ;
  assign w3105 = \pi002 ^ w3100 ;
  assign w3106 = \pi000 & ~w3100 ;
  assign w3107 = w3104 & w3106 ;
  assign w3108 = \pi001 ^ w3107 ;
  assign w3109 = ( \pi001 & w3105 ) | ( \pi001 & ~w3108 ) | ( w3105 & ~w3108 ) ;
  assign w3110 = ( w2832 & w2955 ) | ( w2832 & w2971 ) | ( w2955 & w2971 ) ;
  assign w3111 = w3092 ^ w3110 ;
  assign w3112 = w3109 ^ w3111 ;
  assign w3113 = ( w3092 & w3109 ) | ( w3092 & w3110 ) | ( w3109 & w3110 ) ;
  assign w3114 = ~\pi097 & w189 ;
  assign w3115 = \pi096 & w229 ;
  assign w3116 = ( w189 & ~w3114 ) | ( w189 & w3115 ) | ( ~w3114 & w3115 ) ;
  assign w3117 = ~\pi098 & w191 ;
  assign w3118 = w2824 | w3116 ;
  assign w3119 = ( w192 & w3116 ) | ( w192 & w3118 ) | ( w3116 & w3118 ) ;
  assign w3120 = ( w191 & ~w3117 ) | ( w191 & w3119 ) | ( ~w3117 & w3119 ) ;
  assign w3121 = \pi005 ^ w3120 ;
  assign w3122 = ( w2982 & w3080 ) | ( w2982 & w3088 ) | ( w3080 & w3088 ) ;
  assign w3123 = ~\pi094 & w305 ;
  assign w3124 = \pi093 & w328 ;
  assign w3125 = ( w305 & ~w3123 ) | ( w305 & w3124 ) | ( ~w3123 & w3124 ) ;
  assign w3126 = ~\pi095 & w307 ;
  assign w3127 = w2409 | w3125 ;
  assign w3128 = ( w308 & w3125 ) | ( w308 & w3127 ) | ( w3125 & w3127 ) ;
  assign w3129 = ( w307 & ~w3126 ) | ( w307 & w3128 ) | ( ~w3126 & w3128 ) ;
  assign w3130 = \pi008 ^ w3129 ;
  assign w3131 = ( w2983 & w2991 ) | ( w2983 & w3078 ) | ( w2991 & w3078 ) ;
  assign w3132 = ( w2992 & w3068 ) | ( w2992 & w3076 ) | ( w3068 & w3076 ) ;
  assign w3133 = ~\pi079 & w1313 ;
  assign w3134 = \pi078 & w1417 ;
  assign w3135 = ( w1313 & ~w3133 ) | ( w1313 & w3134 ) | ( ~w3133 & w3134 ) ;
  assign w3136 = ~\pi080 & w1315 ;
  assign w3137 = w794 | w3135 ;
  assign w3138 = ( w1316 & w3135 ) | ( w1316 & w3137 ) | ( w3135 & w3137 ) ;
  assign w3139 = ( w1315 & ~w3136 ) | ( w1315 & w3138 ) | ( ~w3136 & w3138 ) ;
  assign w3140 = \pi023 ^ w3139 ;
  assign w3141 = ( w3035 & w3043 ) | ( w3035 & w3044 ) | ( w3043 & w3044 ) ;
  assign w3142 = ~\pi076 & w1629 ;
  assign w3143 = \pi075 & w1722 ;
  assign w3144 = ( w1629 & ~w3142 ) | ( w1629 & w3143 ) | ( ~w3142 & w3143 ) ;
  assign w3145 = ~\pi077 & w1631 ;
  assign w3146 = w644 | w3144 ;
  assign w3147 = ( w1632 & w3144 ) | ( w1632 & w3146 ) | ( w3144 & w3146 ) ;
  assign w3148 = ( w1631 & ~w3145 ) | ( w1631 & w3147 ) | ( ~w3145 & w3147 ) ;
  assign w3149 = \pi026 ^ w3148 ;
  assign w3150 = ( w3003 & w3025 ) | ( w3003 & w3033 ) | ( w3025 & w3033 ) ;
  assign w3151 = ~\pi073 & w1944 ;
  assign w3152 = \pi072 & w2072 ;
  assign w3153 = ( w1944 & ~w3151 ) | ( w1944 & w3152 ) | ( ~w3151 & w3152 ) ;
  assign w3154 = ~\pi074 & w1946 ;
  assign w3155 = w465 | w3153 ;
  assign w3156 = ( w1947 & w3153 ) | ( w1947 & w3155 ) | ( w3153 & w3155 ) ;
  assign w3157 = ( w1946 & ~w3154 ) | ( w1946 & w3156 ) | ( ~w3154 & w3156 ) ;
  assign w3158 = \pi029 ^ w3157 ;
  assign w3159 = ( w2891 & w3011 ) | ( w2891 & w3023 ) | ( w3011 & w3023 ) ;
  assign w3160 = ~\pi070 & w2310 ;
  assign w3161 = \pi069 & w2443 ;
  assign w3162 = ( w2310 & ~w3160 ) | ( w2310 & w3161 ) | ( ~w3160 & w3161 ) ;
  assign w3163 = ~\pi071 & w2312 ;
  assign w3164 = w290 | w3162 ;
  assign w3165 = ( w2313 & w3162 ) | ( w2313 & w3164 ) | ( w3162 & w3164 ) ;
  assign w3166 = ( w2312 & ~w3163 ) | ( w2312 & w3165 ) | ( ~w3163 & w3165 ) ;
  assign w3167 = \pi032 ^ w3166 ;
  assign w3168 = ( w2881 & w3019 ) | ( w2881 & w3022 ) | ( w3019 & w3022 ) ;
  assign w3169 = ~\pi067 & w2712 ;
  assign w3170 = \pi066 & w2872 ;
  assign w3171 = ( w2712 & ~w3169 ) | ( w2712 & w3170 ) | ( ~w3169 & w3170 ) ;
  assign w3172 = ~\pi068 & w2714 ;
  assign w3173 = w182 | w3171 ;
  assign w3174 = ( w2715 & w3171 ) | ( w2715 & w3173 ) | ( w3171 & w3173 ) ;
  assign w3175 = ( w2714 & ~w3172 ) | ( w2714 & w3174 ) | ( ~w3172 & w3174 ) ;
  assign w3176 = \pi035 ^ w3175 ;
  assign w3177 = ( \pi035 & \pi036 ) | ( \pi035 & \pi037 ) | ( \pi036 & \pi037 ) ;
  assign w3178 = \pi037 ^ w3177 ;
  assign w3179 = \pi037 ^ \pi038 ;
  assign w3180 = w3021 & ~w3179 ;
  assign w3181 = w3021 & w3179 ;
  assign w3182 = ( \pi035 & \pi036 ) | ( \pi035 & ~\pi038 ) | ( \pi036 & ~\pi038 ) ;
  assign w3183 = \pi038 & ~\pi064 ;
  assign w3184 = ~\pi065 & w3183 ;
  assign w3185 = ( \pi035 & \pi036 ) | ( \pi035 & ~w3184 ) | ( \pi036 & ~w3184 ) ;
  assign w3186 = ( \pi037 & \pi038 ) | ( \pi037 & ~w3185 ) | ( \pi038 & ~w3185 ) ;
  assign w3187 = ( \pi037 & ~w3183 ) | ( \pi037 & w3185 ) | ( ~w3183 & w3185 ) ;
  assign w3188 = ( w3182 & w3186 ) | ( w3182 & ~w3187 ) | ( w3186 & ~w3187 ) ;
  assign w3189 = ( \pi035 & \pi036 ) | ( \pi035 & \pi065 ) | ( \pi036 & \pi065 ) ;
  assign w3190 = \pi035 & \pi036 ;
  assign w3191 = \pi064 ^ w3190 ;
  assign w3192 = ( \pi037 & w3190 ) | ( \pi037 & w3191 ) | ( w3190 & w3191 ) ;
  assign w3193 = w3189 ^ w3192 ;
  assign w3194 = w3168 ^ w3176 ;
  assign w3195 = w3193 ^ w3194 ;
  assign w3196 = w3159 ^ w3195 ;
  assign w3197 = w3167 ^ w3196 ;
  assign w3198 = w3150 ^ w3197 ;
  assign w3199 = w3158 ^ w3198 ;
  assign w3200 = w3141 ^ w3199 ;
  assign w3201 = w3149 ^ w3200 ;
  assign w3202 = ( w2994 & w3002 ) | ( w2994 & w3046 ) | ( w3002 & w3046 ) ;
  assign w3203 = w3201 ^ w3202 ;
  assign w3204 = w3140 ^ w3203 ;
  assign w3205 = ~\pi082 & w1044 ;
  assign w3206 = \pi081 & w1138 ;
  assign w3207 = ( w1044 & ~w3205 ) | ( w1044 & w3206 ) | ( ~w3205 & w3206 ) ;
  assign w3208 = ~\pi083 & w1046 ;
  assign w3209 = w1099 | w3207 ;
  assign w3210 = ( w1047 & w3207 ) | ( w1047 & w3209 ) | ( w3207 & w3209 ) ;
  assign w3211 = ( w1046 & ~w3208 ) | ( w1046 & w3210 ) | ( ~w3208 & w3210 ) ;
  assign w3212 = \pi020 ^ w3211 ;
  assign w3213 = ( w2993 & w3048 ) | ( w2993 & w3056 ) | ( w3048 & w3056 ) ;
  assign w3214 = w3204 ^ w3213 ;
  assign w3215 = w3212 ^ w3214 ;
  assign w3216 = ~\pi085 & w837 ;
  assign w3217 = \pi084 & w902 ;
  assign w3218 = ( w837 & ~w3216 ) | ( w837 & w3217 ) | ( ~w3216 & w3217 ) ;
  assign w3219 = ~\pi086 & w839 ;
  assign w3220 = w1379 | w3218 ;
  assign w3221 = ( w840 & w3218 ) | ( w840 & w3220 ) | ( w3218 & w3220 ) ;
  assign w3222 = ( w839 & ~w3219 ) | ( w839 & w3221 ) | ( ~w3219 & w3221 ) ;
  assign w3223 = \pi017 ^ w3222 ;
  assign w3224 = ( w2927 & w3058 ) | ( w2927 & w3066 ) | ( w3058 & w3066 ) ;
  assign w3225 = w3215 ^ w3224 ;
  assign w3226 = w3223 ^ w3225 ;
  assign w3227 = ~\pi088 & w601 ;
  assign w3228 = \pi087 & w683 ;
  assign w3229 = ( w601 & ~w3227 ) | ( w601 & w3228 ) | ( ~w3227 & w3228 ) ;
  assign w3230 = ~\pi089 & w603 ;
  assign w3231 = w1595 | w3229 ;
  assign w3232 = ( w604 & w3229 ) | ( w604 & w3231 ) | ( w3229 & w3231 ) ;
  assign w3233 = ( w603 & ~w3230 ) | ( w603 & w3232 ) | ( ~w3230 & w3232 ) ;
  assign w3234 = \pi014 ^ w3233 ;
  assign w3235 = ( w3132 & w3226 ) | ( w3132 & w3234 ) | ( w3226 & w3234 ) ;
  assign w3236 = w3132 ^ w3226 ;
  assign w3237 = w3234 ^ w3236 ;
  assign w3238 = ~\pi091 & w432 ;
  assign w3239 = \pi090 & w486 ;
  assign w3240 = ( w432 & ~w3238 ) | ( w432 & w3239 ) | ( ~w3238 & w3239 ) ;
  assign w3241 = ~\pi092 & w434 ;
  assign w3242 = w2033 | w3240 ;
  assign w3243 = ( w435 & w3240 ) | ( w435 & w3242 ) | ( w3240 & w3242 ) ;
  assign w3244 = ( w434 & ~w3241 ) | ( w434 & w3243 ) | ( ~w3241 & w3243 ) ;
  assign w3245 = \pi011 ^ w3244 ;
  assign w3246 = w3131 ^ w3237 ;
  assign w3247 = w3245 ^ w3246 ;
  assign w3248 = w3122 ^ w3247 ;
  assign w3249 = w3130 ^ w3248 ;
  assign w3250 = ( w2953 & w2981 ) | ( w2953 & w3090 ) | ( w2981 & w3090 ) ;
  assign w3251 = w3249 ^ w3250 ;
  assign w3252 = w3121 ^ w3251 ;
  assign w3253 = ( ~\pi002 & \pi100 ) | ( ~\pi002 & \pi101 ) | ( \pi100 & \pi101 ) ;
  assign w3254 = \pi000 ^ w3253 ;
  assign w3255 = ( \pi002 & \pi101 ) | ( \pi002 & ~w3254 ) | ( \pi101 & ~w3254 ) ;
  assign w3256 = ( \pi002 & \pi100 ) | ( \pi002 & w3254 ) | ( \pi100 & w3254 ) ;
  assign w3257 = \pi001 & w3256 ;
  assign w3258 = ( ~\pi000 & \pi099 ) | ( ~\pi000 & w3257 ) | ( \pi099 & w3257 ) ;
  assign w3259 = ( \pi001 & \pi002 ) | ( \pi001 & ~w3258 ) | ( \pi002 & ~w3258 ) ;
  assign w3260 = ( w3255 & w3257 ) | ( w3255 & ~w3259 ) | ( w3257 & ~w3259 ) ;
  assign w3261 = ( \pi098 & \pi099 ) | ( \pi098 & \pi100 ) | ( \pi099 & \pi100 ) ;
  assign w3262 = ( \pi099 & w2964 ) | ( \pi099 & w3261 ) | ( w2964 & w3261 ) ;
  assign w3263 = \pi100 ^ \pi101 ;
  assign w3264 = w3262 ^ w3263 ;
  assign w3265 = \pi002 ^ w3260 ;
  assign w3266 = \pi000 & ~w3260 ;
  assign w3267 = w3264 & w3266 ;
  assign w3268 = \pi001 ^ w3267 ;
  assign w3269 = ( \pi001 & w3265 ) | ( \pi001 & ~w3268 ) | ( w3265 & ~w3268 ) ;
  assign w3270 = w3113 ^ w3252 ;
  assign w3271 = w3269 ^ w3270 ;
  assign w3272 = ( ~\pi002 & \pi101 ) | ( ~\pi002 & \pi102 ) | ( \pi101 & \pi102 ) ;
  assign w3273 = \pi000 ^ w3272 ;
  assign w3274 = ( \pi002 & \pi102 ) | ( \pi002 & ~w3273 ) | ( \pi102 & ~w3273 ) ;
  assign w3275 = ( \pi002 & \pi101 ) | ( \pi002 & w3273 ) | ( \pi101 & w3273 ) ;
  assign w3276 = \pi001 & w3275 ;
  assign w3277 = ( ~\pi000 & \pi100 ) | ( ~\pi000 & w3276 ) | ( \pi100 & w3276 ) ;
  assign w3278 = ( \pi001 & \pi002 ) | ( \pi001 & ~w3277 ) | ( \pi002 & ~w3277 ) ;
  assign w3279 = ( w3274 & w3276 ) | ( w3274 & ~w3278 ) | ( w3276 & ~w3278 ) ;
  assign w3280 = ( \pi098 & \pi099 ) | ( \pi098 & ~\pi101 ) | ( \pi099 & ~\pi101 ) ;
  assign w3281 = ( \pi099 & w2964 ) | ( \pi099 & w3280 ) | ( w2964 & w3280 ) ;
  assign w3282 = ( \pi100 & \pi101 ) | ( \pi100 & w3281 ) | ( \pi101 & w3281 ) ;
  assign w3283 = \pi101 ^ w3282 ;
  assign w3284 = \pi102 ^ w3283 ;
  assign w3285 = \pi002 ^ w3279 ;
  assign w3286 = \pi000 & ~w3279 ;
  assign w3287 = w3284 & w3286 ;
  assign w3288 = \pi001 ^ w3287 ;
  assign w3289 = ( \pi001 & w3285 ) | ( \pi001 & ~w3288 ) | ( w3285 & ~w3288 ) ;
  assign w3290 = ( w3121 & w3249 ) | ( w3121 & w3250 ) | ( w3249 & w3250 ) ;
  assign w3291 = ~\pi098 & w189 ;
  assign w3292 = \pi097 & w229 ;
  assign w3293 = ( w189 & ~w3291 ) | ( w189 & w3292 ) | ( ~w3291 & w3292 ) ;
  assign w3294 = ~\pi099 & w191 ;
  assign w3295 = w2966 | w3293 ;
  assign w3296 = ( w192 & w3293 ) | ( w192 & w3295 ) | ( w3293 & w3295 ) ;
  assign w3297 = ( w191 & ~w3294 ) | ( w191 & w3296 ) | ( ~w3294 & w3296 ) ;
  assign w3298 = \pi005 ^ w3297 ;
  assign w3299 = ( w3122 & w3130 ) | ( w3122 & w3247 ) | ( w3130 & w3247 ) ;
  assign w3300 = ~\pi095 & w305 ;
  assign w3301 = \pi094 & w328 ;
  assign w3302 = ( w305 & ~w3300 ) | ( w305 & w3301 ) | ( ~w3300 & w3301 ) ;
  assign w3303 = ~\pi096 & w307 ;
  assign w3304 = w2546 | w3302 ;
  assign w3305 = ( w308 & w3302 ) | ( w308 & w3304 ) | ( w3302 & w3304 ) ;
  assign w3306 = ( w307 & ~w3303 ) | ( w307 & w3305 ) | ( ~w3303 & w3305 ) ;
  assign w3307 = \pi008 ^ w3306 ;
  assign w3308 = ( w3131 & w3237 ) | ( w3131 & w3245 ) | ( w3237 & w3245 ) ;
  assign w3309 = ~\pi092 & w432 ;
  assign w3310 = \pi091 & w486 ;
  assign w3311 = ( w432 & ~w3309 ) | ( w432 & w3310 ) | ( ~w3309 & w3310 ) ;
  assign w3312 = ~\pi093 & w434 ;
  assign w3313 = w2155 | w3311 ;
  assign w3314 = ( w435 & w3311 ) | ( w435 & w3313 ) | ( w3311 & w3313 ) ;
  assign w3315 = ( w434 & ~w3312 ) | ( w434 & w3314 ) | ( ~w3312 & w3314 ) ;
  assign w3316 = \pi011 ^ w3315 ;
  assign w3317 = ( w3215 & w3223 ) | ( w3215 & w3224 ) | ( w3223 & w3224 ) ;
  assign w3318 = ~\pi080 & w1313 ;
  assign w3319 = \pi079 & w1417 ;
  assign w3320 = ( w1313 & ~w3318 ) | ( w1313 & w3319 ) | ( ~w3318 & w3319 ) ;
  assign w3321 = ~\pi081 & w1315 ;
  assign w3322 = w874 | w3320 ;
  assign w3323 = ( w1316 & w3320 ) | ( w1316 & w3322 ) | ( w3320 & w3322 ) ;
  assign w3324 = ( w1315 & ~w3321 ) | ( w1315 & w3323 ) | ( ~w3321 & w3323 ) ;
  assign w3325 = \pi023 ^ w3324 ;
  assign w3326 = ( w3141 & w3149 ) | ( w3141 & w3199 ) | ( w3149 & w3199 ) ;
  assign w3327 = ( w3150 & w3158 ) | ( w3150 & w3197 ) | ( w3158 & w3197 ) ;
  assign w3328 = ~\pi074 & w1944 ;
  assign w3329 = \pi073 & w2072 ;
  assign w3330 = ( w1944 & ~w3328 ) | ( w1944 & w3329 ) | ( ~w3328 & w3329 ) ;
  assign w3331 = ~\pi075 & w1946 ;
  assign w3332 = w519 | w3330 ;
  assign w3333 = ( w1947 & w3330 ) | ( w1947 & w3332 ) | ( w3330 & w3332 ) ;
  assign w3334 = ( w1946 & ~w3331 ) | ( w1946 & w3333 ) | ( ~w3331 & w3333 ) ;
  assign w3335 = \pi029 ^ w3334 ;
  assign w3336 = ( w3159 & w3167 ) | ( w3159 & w3195 ) | ( w3167 & w3195 ) ;
  assign w3337 = ( w3168 & w3176 ) | ( w3168 & w3193 ) | ( w3176 & w3193 ) ;
  assign w3338 = ( \pi036 & ~\pi037 ) | ( \pi036 & \pi038 ) | ( ~\pi037 & \pi038 ) ;
  assign w3339 = ( \pi035 & \pi036 ) | ( \pi035 & w3338 ) | ( \pi036 & w3338 ) ;
  assign w3340 = w3338 ^ w3339 ;
  assign w3341 = \pi064 & w3340 ;
  assign w3342 = ( \pi066 & w3180 ) | ( \pi066 & w3341 ) | ( w3180 & w3341 ) ;
  assign w3343 = \pi065 | w3342 ;
  assign w3344 = ( w3178 & w3342 ) | ( w3178 & w3343 ) | ( w3342 & w3343 ) ;
  assign w3345 = w3341 | w3344 ;
  assign w3346 = ~w134 & w3181 ;
  assign w3347 = ( w3181 & w3345 ) | ( w3181 & ~w3346 ) | ( w3345 & ~w3346 ) ;
  assign w3348 = \pi038 ^ w3347 ;
  assign w3349 = w3188 & w3348 ;
  assign w3350 = w3188 ^ w3348 ;
  assign w3351 = ~\pi068 & w2712 ;
  assign w3352 = \pi067 & w2872 ;
  assign w3353 = ( w2712 & ~w3351 ) | ( w2712 & w3352 ) | ( ~w3351 & w3352 ) ;
  assign w3354 = ~\pi069 & w2714 ;
  assign w3355 = w221 | w3353 ;
  assign w3356 = ( w2715 & w3353 ) | ( w2715 & w3355 ) | ( w3353 & w3355 ) ;
  assign w3357 = ( w2714 & ~w3354 ) | ( w2714 & w3356 ) | ( ~w3354 & w3356 ) ;
  assign w3358 = \pi035 ^ w3357 ;
  assign w3359 = w3337 ^ w3350 ;
  assign w3360 = w3358 ^ w3359 ;
  assign w3361 = ~\pi071 & w2310 ;
  assign w3362 = \pi070 & w2443 ;
  assign w3363 = ( w2310 & ~w3361 ) | ( w2310 & w3362 ) | ( ~w3361 & w3362 ) ;
  assign w3364 = ~\pi072 & w2312 ;
  assign w3365 = w361 | w3363 ;
  assign w3366 = ( w2313 & w3363 ) | ( w2313 & w3365 ) | ( w3363 & w3365 ) ;
  assign w3367 = ( w2312 & ~w3364 ) | ( w2312 & w3366 ) | ( ~w3364 & w3366 ) ;
  assign w3368 = \pi032 ^ w3367 ;
  assign w3369 = w3336 ^ w3360 ;
  assign w3370 = w3368 ^ w3369 ;
  assign w3371 = w3327 ^ w3370 ;
  assign w3372 = w3335 ^ w3371 ;
  assign w3373 = ~\pi077 & w1629 ;
  assign w3374 = \pi076 & w1722 ;
  assign w3375 = ( w1629 & ~w3373 ) | ( w1629 & w3374 ) | ( ~w3373 & w3374 ) ;
  assign w3376 = ~\pi078 & w1631 ;
  assign w3377 = w665 | w3375 ;
  assign w3378 = ( w1632 & w3375 ) | ( w1632 & w3377 ) | ( w3375 & w3377 ) ;
  assign w3379 = ( w1631 & ~w3376 ) | ( w1631 & w3378 ) | ( ~w3376 & w3378 ) ;
  assign w3380 = \pi026 ^ w3379 ;
  assign w3381 = w3326 ^ w3372 ;
  assign w3382 = w3380 ^ w3381 ;
  assign w3383 = ( w3140 & w3201 ) | ( w3140 & w3202 ) | ( w3201 & w3202 ) ;
  assign w3384 = w3382 ^ w3383 ;
  assign w3385 = w3325 ^ w3384 ;
  assign w3386 = ~\pi083 & w1044 ;
  assign w3387 = \pi082 & w1138 ;
  assign w3388 = ( w1044 & ~w3386 ) | ( w1044 & w3387 ) | ( ~w3386 & w3387 ) ;
  assign w3389 = ~\pi084 & w1046 ;
  assign w3390 = w1188 | w3388 ;
  assign w3391 = ( w1047 & w3388 ) | ( w1047 & w3390 ) | ( w3388 & w3390 ) ;
  assign w3392 = ( w1046 & ~w3389 ) | ( w1046 & w3391 ) | ( ~w3389 & w3391 ) ;
  assign w3393 = \pi020 ^ w3392 ;
  assign w3394 = ( w3204 & w3212 ) | ( w3204 & w3213 ) | ( w3212 & w3213 ) ;
  assign w3395 = w3385 ^ w3394 ;
  assign w3396 = w3393 ^ w3395 ;
  assign w3397 = ~\pi086 & w837 ;
  assign w3398 = \pi085 & w902 ;
  assign w3399 = ( w837 & ~w3397 ) | ( w837 & w3398 ) | ( ~w3397 & w3398 ) ;
  assign w3400 = ~\pi087 & w839 ;
  assign w3401 = w1477 | w3399 ;
  assign w3402 = ( w840 & w3399 ) | ( w840 & w3401 ) | ( w3399 & w3401 ) ;
  assign w3403 = ( w839 & ~w3400 ) | ( w839 & w3402 ) | ( ~w3400 & w3402 ) ;
  assign w3404 = \pi017 ^ w3403 ;
  assign w3405 = ( w3317 & w3396 ) | ( w3317 & w3404 ) | ( w3396 & w3404 ) ;
  assign w3406 = w3317 ^ w3396 ;
  assign w3407 = w3404 ^ w3406 ;
  assign w3408 = ~\pi089 & w601 ;
  assign w3409 = \pi088 & w683 ;
  assign w3410 = ( w601 & ~w3408 ) | ( w601 & w3409 ) | ( ~w3408 & w3409 ) ;
  assign w3411 = ~\pi090 & w603 ;
  assign w3412 = w1801 | w3410 ;
  assign w3413 = ( w604 & w3410 ) | ( w604 & w3412 ) | ( w3410 & w3412 ) ;
  assign w3414 = ( w603 & ~w3411 ) | ( w603 & w3413 ) | ( ~w3411 & w3413 ) ;
  assign w3415 = \pi014 ^ w3414 ;
  assign w3416 = w3235 ^ w3407 ;
  assign w3417 = w3415 ^ w3416 ;
  assign w3418 = w3308 ^ w3417 ;
  assign w3419 = w3316 ^ w3418 ;
  assign w3420 = w3299 ^ w3419 ;
  assign w3421 = w3307 ^ w3420 ;
  assign w3422 = w3290 ^ w3421 ;
  assign w3423 = w3298 ^ w3422 ;
  assign w3424 = ( w3113 & w3252 ) | ( w3113 & w3269 ) | ( w3252 & w3269 ) ;
  assign w3425 = w3423 ^ w3424 ;
  assign w3426 = w3289 ^ w3425 ;
  assign w3427 = ( ~\pi002 & \pi102 ) | ( ~\pi002 & \pi103 ) | ( \pi102 & \pi103 ) ;
  assign w3428 = \pi000 ^ w3427 ;
  assign w3429 = ( \pi002 & \pi103 ) | ( \pi002 & ~w3428 ) | ( \pi103 & ~w3428 ) ;
  assign w3430 = ( \pi002 & \pi102 ) | ( \pi002 & w3428 ) | ( \pi102 & w3428 ) ;
  assign w3431 = \pi001 & w3430 ;
  assign w3432 = ( ~\pi000 & \pi101 ) | ( ~\pi000 & w3431 ) | ( \pi101 & w3431 ) ;
  assign w3433 = ( \pi001 & \pi002 ) | ( \pi001 & ~w3432 ) | ( \pi002 & ~w3432 ) ;
  assign w3434 = ( w3429 & w3431 ) | ( w3429 & ~w3433 ) | ( w3431 & ~w3433 ) ;
  assign w3435 = ( \pi101 & \pi102 ) | ( \pi101 & w3282 ) | ( \pi102 & w3282 ) ;
  assign w3436 = \pi102 ^ w3435 ;
  assign w3437 = \pi103 ^ w3436 ;
  assign w3438 = \pi002 ^ w3434 ;
  assign w3439 = \pi000 & ~w3434 ;
  assign w3440 = w3437 & w3439 ;
  assign w3441 = \pi001 ^ w3440 ;
  assign w3442 = ( \pi001 & w3438 ) | ( \pi001 & ~w3441 ) | ( w3438 & ~w3441 ) ;
  assign w3443 = ( w3290 & w3298 ) | ( w3290 & w3421 ) | ( w3298 & w3421 ) ;
  assign w3444 = ( w3299 & w3307 ) | ( w3299 & w3419 ) | ( w3307 & w3419 ) ;
  assign w3445 = ~\pi096 & w305 ;
  assign w3446 = \pi095 & w328 ;
  assign w3447 = ( w305 & ~w3445 ) | ( w305 & w3446 ) | ( ~w3445 & w3446 ) ;
  assign w3448 = ~\pi097 & w307 ;
  assign w3449 = w2673 | w3447 ;
  assign w3450 = ( w308 & w3447 ) | ( w308 & w3449 ) | ( w3447 & w3449 ) ;
  assign w3451 = ( w307 & ~w3448 ) | ( w307 & w3450 ) | ( ~w3448 & w3450 ) ;
  assign w3452 = \pi008 ^ w3451 ;
  assign w3453 = ( w3308 & w3316 ) | ( w3308 & w3417 ) | ( w3316 & w3417 ) ;
  assign w3454 = ( w3235 & w3407 ) | ( w3235 & w3415 ) | ( w3407 & w3415 ) ;
  assign w3455 = ~\pi090 & w601 ;
  assign w3456 = \pi089 & w683 ;
  assign w3457 = ( w601 & ~w3455 ) | ( w601 & w3456 ) | ( ~w3455 & w3456 ) ;
  assign w3458 = ~\pi091 & w603 ;
  assign w3459 = w1908 | w3457 ;
  assign w3460 = ( w604 & w3457 ) | ( w604 & w3459 ) | ( w3457 & w3459 ) ;
  assign w3461 = ( w603 & ~w3458 ) | ( w603 & w3460 ) | ( ~w3458 & w3460 ) ;
  assign w3462 = \pi014 ^ w3461 ;
  assign w3463 = ( w3325 & w3382 ) | ( w3325 & w3383 ) | ( w3382 & w3383 ) ;
  assign w3464 = ( w3326 & w3372 ) | ( w3326 & w3380 ) | ( w3372 & w3380 ) ;
  assign w3465 = ~\pi078 & w1629 ;
  assign w3466 = \pi077 & w1722 ;
  assign w3467 = ( w1629 & ~w3465 ) | ( w1629 & w3466 ) | ( ~w3465 & w3466 ) ;
  assign w3468 = ~\pi079 & w1631 ;
  assign w3469 = w730 | w3467 ;
  assign w3470 = ( w1632 & w3467 ) | ( w1632 & w3469 ) | ( w3467 & w3469 ) ;
  assign w3471 = ( w1631 & ~w3468 ) | ( w1631 & w3470 ) | ( ~w3468 & w3470 ) ;
  assign w3472 = \pi026 ^ w3471 ;
  assign w3473 = ~\pi069 & w2712 ;
  assign w3474 = \pi068 & w2872 ;
  assign w3475 = ( w2712 & ~w3473 ) | ( w2712 & w3474 ) | ( ~w3473 & w3474 ) ;
  assign w3476 = ~\pi070 & w2714 ;
  assign w3477 = w271 | w3475 ;
  assign w3478 = ( w2715 & w3475 ) | ( w2715 & w3477 ) | ( w3475 & w3477 ) ;
  assign w3479 = ( w2714 & ~w3476 ) | ( w2714 & w3478 ) | ( ~w3476 & w3478 ) ;
  assign w3480 = \pi035 ^ w3479 ;
  assign w3481 = ~\pi066 & w3178 ;
  assign w3482 = \pi065 & w3340 ;
  assign w3483 = ( w3178 & ~w3481 ) | ( w3178 & w3482 ) | ( ~w3481 & w3482 ) ;
  assign w3484 = ~\pi067 & w3180 ;
  assign w3485 = w160 | w3483 ;
  assign w3486 = ( w3181 & w3483 ) | ( w3181 & w3485 ) | ( w3483 & w3485 ) ;
  assign w3487 = ( w3180 & ~w3484 ) | ( w3180 & w3486 ) | ( ~w3484 & w3486 ) ;
  assign w3488 = \pi038 ^ w3487 ;
  assign w3489 = w3349 ^ w3488 ;
  assign w3490 = \pi038 ^ \pi039 ;
  assign w3491 = \pi064 & w3490 ;
  assign w3492 = w3489 ^ w3491 ;
  assign w3493 = ( w3337 & w3350 ) | ( w3337 & w3358 ) | ( w3350 & w3358 ) ;
  assign w3494 = w3492 ^ w3493 ;
  assign w3495 = w3480 ^ w3494 ;
  assign w3496 = ~\pi072 & w2310 ;
  assign w3497 = \pi071 & w2443 ;
  assign w3498 = ( w2310 & ~w3496 ) | ( w2310 & w3497 ) | ( ~w3496 & w3497 ) ;
  assign w3499 = ~\pi073 & w2312 ;
  assign w3500 = w404 | w3498 ;
  assign w3501 = ( w2313 & w3498 ) | ( w2313 & w3500 ) | ( w3498 & w3500 ) ;
  assign w3502 = ( w2312 & ~w3499 ) | ( w2312 & w3501 ) | ( ~w3499 & w3501 ) ;
  assign w3503 = \pi032 ^ w3502 ;
  assign w3504 = ( w3336 & w3360 ) | ( w3336 & w3368 ) | ( w3360 & w3368 ) ;
  assign w3505 = w3495 ^ w3504 ;
  assign w3506 = w3503 ^ w3505 ;
  assign w3507 = ~\pi075 & w1944 ;
  assign w3508 = \pi074 & w2072 ;
  assign w3509 = ( w1944 & ~w3507 ) | ( w1944 & w3508 ) | ( ~w3507 & w3508 ) ;
  assign w3510 = ~\pi076 & w1946 ;
  assign w3511 = w538 | w3509 ;
  assign w3512 = ( w1947 & w3509 ) | ( w1947 & w3511 ) | ( w3509 & w3511 ) ;
  assign w3513 = ( w1946 & ~w3510 ) | ( w1946 & w3512 ) | ( ~w3510 & w3512 ) ;
  assign w3514 = \pi029 ^ w3513 ;
  assign w3515 = ( w3327 & w3335 ) | ( w3327 & w3370 ) | ( w3335 & w3370 ) ;
  assign w3516 = w3506 ^ w3515 ;
  assign w3517 = w3514 ^ w3516 ;
  assign w3518 = w3464 ^ w3517 ;
  assign w3519 = w3472 ^ w3518 ;
  assign w3520 = ~\pi081 & w1313 ;
  assign w3521 = \pi080 & w1417 ;
  assign w3522 = ( w1313 & ~w3520 ) | ( w1313 & w3521 ) | ( ~w3520 & w3521 ) ;
  assign w3523 = ~\pi082 & w1315 ;
  assign w3524 = w1008 | w3522 ;
  assign w3525 = ( w1316 & w3522 ) | ( w1316 & w3524 ) | ( w3522 & w3524 ) ;
  assign w3526 = ( w1315 & ~w3523 ) | ( w1315 & w3525 ) | ( ~w3523 & w3525 ) ;
  assign w3527 = \pi023 ^ w3526 ;
  assign w3528 = w3463 ^ w3519 ;
  assign w3529 = w3527 ^ w3528 ;
  assign w3530 = ~\pi084 & w1044 ;
  assign w3531 = \pi083 & w1138 ;
  assign w3532 = ( w1044 & ~w3530 ) | ( w1044 & w3531 ) | ( ~w3530 & w3531 ) ;
  assign w3533 = ~\pi085 & w1046 ;
  assign w3534 = w1274 | w3532 ;
  assign w3535 = ( w1047 & w3532 ) | ( w1047 & w3534 ) | ( w3532 & w3534 ) ;
  assign w3536 = ( w1046 & ~w3533 ) | ( w1046 & w3535 ) | ( ~w3533 & w3535 ) ;
  assign w3537 = \pi020 ^ w3536 ;
  assign w3538 = ( w3385 & w3393 ) | ( w3385 & w3394 ) | ( w3393 & w3394 ) ;
  assign w3539 = w3529 ^ w3538 ;
  assign w3540 = w3537 ^ w3539 ;
  assign w3541 = ~\pi087 & w837 ;
  assign w3542 = \pi086 & w902 ;
  assign w3543 = ( w837 & ~w3541 ) | ( w837 & w3542 ) | ( ~w3541 & w3542 ) ;
  assign w3544 = ~\pi088 & w839 ;
  assign w3545 = w1574 | w3543 ;
  assign w3546 = ( w840 & w3543 ) | ( w840 & w3545 ) | ( w3543 & w3545 ) ;
  assign w3547 = ( w839 & ~w3544 ) | ( w839 & w3546 ) | ( ~w3544 & w3546 ) ;
  assign w3548 = \pi017 ^ w3547 ;
  assign w3549 = w3405 ^ w3540 ;
  assign w3550 = w3548 ^ w3549 ;
  assign w3551 = w3454 ^ w3550 ;
  assign w3552 = w3462 ^ w3551 ;
  assign w3553 = ~\pi093 & w432 ;
  assign w3554 = \pi092 & w486 ;
  assign w3555 = ( w432 & ~w3553 ) | ( w432 & w3554 ) | ( ~w3553 & w3554 ) ;
  assign w3556 = ~\pi094 & w434 ;
  assign w3557 = w2274 | w3555 ;
  assign w3558 = ( w435 & w3555 ) | ( w435 & w3557 ) | ( w3555 & w3557 ) ;
  assign w3559 = ( w434 & ~w3556 ) | ( w434 & w3558 ) | ( ~w3556 & w3558 ) ;
  assign w3560 = \pi011 ^ w3559 ;
  assign w3561 = w3453 ^ w3552 ;
  assign w3562 = w3560 ^ w3561 ;
  assign w3563 = w3444 ^ w3562 ;
  assign w3564 = w3452 ^ w3563 ;
  assign w3565 = ~\pi099 & w189 ;
  assign w3566 = \pi098 & w229 ;
  assign w3567 = ( w189 & ~w3565 ) | ( w189 & w3566 ) | ( ~w3565 & w3566 ) ;
  assign w3568 = ~\pi100 & w191 ;
  assign w3569 = w3104 | w3567 ;
  assign w3570 = ( w192 & w3567 ) | ( w192 & w3569 ) | ( w3567 & w3569 ) ;
  assign w3571 = ( w191 & ~w3568 ) | ( w191 & w3570 ) | ( ~w3568 & w3570 ) ;
  assign w3572 = \pi005 ^ w3571 ;
  assign w3573 = w3443 ^ w3564 ;
  assign w3574 = w3572 ^ w3573 ;
  assign w3575 = ( w3289 & w3423 ) | ( w3289 & w3424 ) | ( w3423 & w3424 ) ;
  assign w3576 = w3574 ^ w3575 ;
  assign w3577 = w3442 ^ w3576 ;
  assign w3578 = ( w3442 & w3574 ) | ( w3442 & w3575 ) | ( w3574 & w3575 ) ;
  assign w3579 = ( w3443 & w3564 ) | ( w3443 & w3572 ) | ( w3564 & w3572 ) ;
  assign w3580 = ~\pi100 & w189 ;
  assign w3581 = \pi099 & w229 ;
  assign w3582 = ( w189 & ~w3580 ) | ( w189 & w3581 ) | ( ~w3580 & w3581 ) ;
  assign w3583 = ~\pi101 & w191 ;
  assign w3584 = w3264 | w3582 ;
  assign w3585 = ( w192 & w3582 ) | ( w192 & w3584 ) | ( w3582 & w3584 ) ;
  assign w3586 = ( w191 & ~w3583 ) | ( w191 & w3585 ) | ( ~w3583 & w3585 ) ;
  assign w3587 = \pi005 ^ w3586 ;
  assign w3588 = ( w3444 & w3452 ) | ( w3444 & w3562 ) | ( w3452 & w3562 ) ;
  assign w3589 = ~\pi097 & w305 ;
  assign w3590 = \pi096 & w328 ;
  assign w3591 = ( w305 & ~w3589 ) | ( w305 & w3590 ) | ( ~w3589 & w3590 ) ;
  assign w3592 = ~\pi098 & w307 ;
  assign w3593 = w2824 | w3591 ;
  assign w3594 = ( w308 & w3591 ) | ( w308 & w3593 ) | ( w3591 & w3593 ) ;
  assign w3595 = ( w307 & ~w3592 ) | ( w307 & w3594 ) | ( ~w3592 & w3594 ) ;
  assign w3596 = \pi008 ^ w3595 ;
  assign w3597 = ( w3453 & w3552 ) | ( w3453 & w3560 ) | ( w3552 & w3560 ) ;
  assign w3598 = ( w3454 & w3462 ) | ( w3454 & w3550 ) | ( w3462 & w3550 ) ;
  assign w3599 = ~\pi091 & w601 ;
  assign w3600 = \pi090 & w683 ;
  assign w3601 = ( w601 & ~w3599 ) | ( w601 & w3600 ) | ( ~w3599 & w3600 ) ;
  assign w3602 = ~\pi092 & w603 ;
  assign w3603 = w2033 | w3601 ;
  assign w3604 = ( w604 & w3601 ) | ( w604 & w3603 ) | ( w3601 & w3603 ) ;
  assign w3605 = ( w603 & ~w3602 ) | ( w603 & w3604 ) | ( ~w3602 & w3604 ) ;
  assign w3606 = \pi014 ^ w3605 ;
  assign w3607 = ~\pi079 & w1629 ;
  assign w3608 = \pi078 & w1722 ;
  assign w3609 = ( w1629 & ~w3607 ) | ( w1629 & w3608 ) | ( ~w3607 & w3608 ) ;
  assign w3610 = ~\pi080 & w1631 ;
  assign w3611 = w794 | w3609 ;
  assign w3612 = ( w1632 & w3609 ) | ( w1632 & w3611 ) | ( w3609 & w3611 ) ;
  assign w3613 = ( w1631 & ~w3610 ) | ( w1631 & w3612 ) | ( ~w3610 & w3612 ) ;
  assign w3614 = \pi026 ^ w3613 ;
  assign w3615 = ( w3506 & w3514 ) | ( w3506 & w3515 ) | ( w3514 & w3515 ) ;
  assign w3616 = ( w3495 & w3503 ) | ( w3495 & w3504 ) | ( w3503 & w3504 ) ;
  assign w3617 = ~\pi070 & w2712 ;
  assign w3618 = \pi069 & w2872 ;
  assign w3619 = ( w2712 & ~w3617 ) | ( w2712 & w3618 ) | ( ~w3617 & w3618 ) ;
  assign w3620 = ~\pi071 & w2714 ;
  assign w3621 = w290 | w3619 ;
  assign w3622 = ( w2715 & w3619 ) | ( w2715 & w3621 ) | ( w3619 & w3621 ) ;
  assign w3623 = ( w2714 & ~w3620 ) | ( w2714 & w3622 ) | ( ~w3620 & w3622 ) ;
  assign w3624 = \pi035 ^ w3623 ;
  assign w3625 = ( w3349 & w3488 ) | ( w3349 & w3491 ) | ( w3488 & w3491 ) ;
  assign w3626 = ~\pi067 & w3178 ;
  assign w3627 = \pi066 & w3340 ;
  assign w3628 = ( w3178 & ~w3626 ) | ( w3178 & w3627 ) | ( ~w3626 & w3627 ) ;
  assign w3629 = ~\pi068 & w3180 ;
  assign w3630 = w182 | w3628 ;
  assign w3631 = ( w3181 & w3628 ) | ( w3181 & w3630 ) | ( w3628 & w3630 ) ;
  assign w3632 = ( w3180 & ~w3629 ) | ( w3180 & w3631 ) | ( ~w3629 & w3631 ) ;
  assign w3633 = \pi038 ^ w3632 ;
  assign w3634 = ( \pi038 & \pi039 ) | ( \pi038 & \pi040 ) | ( \pi039 & \pi040 ) ;
  assign w3635 = \pi040 ^ w3634 ;
  assign w3636 = \pi040 ^ \pi041 ;
  assign w3637 = w3490 & ~w3636 ;
  assign w3638 = w3490 & w3636 ;
  assign w3639 = ( \pi038 & \pi039 ) | ( \pi038 & ~\pi041 ) | ( \pi039 & ~\pi041 ) ;
  assign w3640 = \pi041 & ~\pi064 ;
  assign w3641 = ~\pi065 & w3640 ;
  assign w3642 = ( \pi038 & \pi039 ) | ( \pi038 & ~w3641 ) | ( \pi039 & ~w3641 ) ;
  assign w3643 = ( \pi040 & \pi041 ) | ( \pi040 & ~w3642 ) | ( \pi041 & ~w3642 ) ;
  assign w3644 = ( \pi040 & ~w3640 ) | ( \pi040 & w3642 ) | ( ~w3640 & w3642 ) ;
  assign w3645 = ( w3639 & w3643 ) | ( w3639 & ~w3644 ) | ( w3643 & ~w3644 ) ;
  assign w3646 = ( \pi038 & \pi039 ) | ( \pi038 & \pi065 ) | ( \pi039 & \pi065 ) ;
  assign w3647 = \pi038 & \pi039 ;
  assign w3648 = \pi064 ^ w3647 ;
  assign w3649 = ( \pi040 & w3647 ) | ( \pi040 & w3648 ) | ( w3647 & w3648 ) ;
  assign w3650 = w3646 ^ w3649 ;
  assign w3651 = w3625 ^ w3633 ;
  assign w3652 = w3650 ^ w3651 ;
  assign w3653 = ( w3480 & w3492 ) | ( w3480 & w3493 ) | ( w3492 & w3493 ) ;
  assign w3654 = w3652 ^ w3653 ;
  assign w3655 = w3624 ^ w3654 ;
  assign w3656 = ~\pi073 & w2310 ;
  assign w3657 = \pi072 & w2443 ;
  assign w3658 = ( w2310 & ~w3656 ) | ( w2310 & w3657 ) | ( ~w3656 & w3657 ) ;
  assign w3659 = ~\pi074 & w2312 ;
  assign w3660 = w465 | w3658 ;
  assign w3661 = ( w2313 & w3658 ) | ( w2313 & w3660 ) | ( w3658 & w3660 ) ;
  assign w3662 = ( w2312 & ~w3659 ) | ( w2312 & w3661 ) | ( ~w3659 & w3661 ) ;
  assign w3663 = \pi032 ^ w3662 ;
  assign w3664 = ( w3616 & w3655 ) | ( w3616 & w3663 ) | ( w3655 & w3663 ) ;
  assign w3665 = w3616 ^ w3655 ;
  assign w3666 = w3663 ^ w3665 ;
  assign w3667 = ~\pi076 & w1944 ;
  assign w3668 = \pi075 & w2072 ;
  assign w3669 = ( w1944 & ~w3667 ) | ( w1944 & w3668 ) | ( ~w3667 & w3668 ) ;
  assign w3670 = ~\pi077 & w1946 ;
  assign w3671 = w644 | w3669 ;
  assign w3672 = ( w1947 & w3669 ) | ( w1947 & w3671 ) | ( w3669 & w3671 ) ;
  assign w3673 = ( w1946 & ~w3670 ) | ( w1946 & w3672 ) | ( ~w3670 & w3672 ) ;
  assign w3674 = \pi029 ^ w3673 ;
  assign w3675 = w3615 ^ w3666 ;
  assign w3676 = w3674 ^ w3675 ;
  assign w3677 = ( w3464 & w3472 ) | ( w3464 & w3517 ) | ( w3472 & w3517 ) ;
  assign w3678 = w3676 ^ w3677 ;
  assign w3679 = w3614 ^ w3678 ;
  assign w3680 = ~\pi082 & w1313 ;
  assign w3681 = \pi081 & w1417 ;
  assign w3682 = ( w1313 & ~w3680 ) | ( w1313 & w3681 ) | ( ~w3680 & w3681 ) ;
  assign w3683 = ~\pi083 & w1315 ;
  assign w3684 = w1099 | w3682 ;
  assign w3685 = ( w1316 & w3682 ) | ( w1316 & w3684 ) | ( w3682 & w3684 ) ;
  assign w3686 = ( w1315 & ~w3683 ) | ( w1315 & w3685 ) | ( ~w3683 & w3685 ) ;
  assign w3687 = \pi023 ^ w3686 ;
  assign w3688 = ( w3463 & w3519 ) | ( w3463 & w3527 ) | ( w3519 & w3527 ) ;
  assign w3689 = w3679 ^ w3688 ;
  assign w3690 = w3687 ^ w3689 ;
  assign w3691 = ~\pi085 & w1044 ;
  assign w3692 = \pi084 & w1138 ;
  assign w3693 = ( w1044 & ~w3691 ) | ( w1044 & w3692 ) | ( ~w3691 & w3692 ) ;
  assign w3694 = ~\pi086 & w1046 ;
  assign w3695 = w1379 | w3693 ;
  assign w3696 = ( w1047 & w3693 ) | ( w1047 & w3695 ) | ( w3693 & w3695 ) ;
  assign w3697 = ( w1046 & ~w3694 ) | ( w1046 & w3696 ) | ( ~w3694 & w3696 ) ;
  assign w3698 = \pi020 ^ w3697 ;
  assign w3699 = ( w3529 & w3537 ) | ( w3529 & w3538 ) | ( w3537 & w3538 ) ;
  assign w3700 = w3690 ^ w3699 ;
  assign w3701 = w3698 ^ w3700 ;
  assign w3702 = ~\pi088 & w837 ;
  assign w3703 = \pi087 & w902 ;
  assign w3704 = ( w837 & ~w3702 ) | ( w837 & w3703 ) | ( ~w3702 & w3703 ) ;
  assign w3705 = ~\pi089 & w839 ;
  assign w3706 = w1595 | w3704 ;
  assign w3707 = ( w840 & w3704 ) | ( w840 & w3706 ) | ( w3704 & w3706 ) ;
  assign w3708 = ( w839 & ~w3705 ) | ( w839 & w3707 ) | ( ~w3705 & w3707 ) ;
  assign w3709 = \pi017 ^ w3708 ;
  assign w3710 = ( w3405 & w3540 ) | ( w3405 & w3548 ) | ( w3540 & w3548 ) ;
  assign w3711 = w3701 ^ w3710 ;
  assign w3712 = w3709 ^ w3711 ;
  assign w3713 = w3598 ^ w3712 ;
  assign w3714 = w3606 ^ w3713 ;
  assign w3715 = ~\pi094 & w432 ;
  assign w3716 = \pi093 & w486 ;
  assign w3717 = ( w432 & ~w3715 ) | ( w432 & w3716 ) | ( ~w3715 & w3716 ) ;
  assign w3718 = ~\pi095 & w434 ;
  assign w3719 = w2409 | w3717 ;
  assign w3720 = ( w435 & w3717 ) | ( w435 & w3719 ) | ( w3717 & w3719 ) ;
  assign w3721 = ( w434 & ~w3718 ) | ( w434 & w3720 ) | ( ~w3718 & w3720 ) ;
  assign w3722 = \pi011 ^ w3721 ;
  assign w3723 = w3597 ^ w3714 ;
  assign w3724 = w3722 ^ w3723 ;
  assign w3725 = w3588 ^ w3724 ;
  assign w3726 = w3596 ^ w3725 ;
  assign w3727 = w3579 ^ w3726 ;
  assign w3728 = w3587 ^ w3727 ;
  assign w3729 = ( ~\pi002 & \pi103 ) | ( ~\pi002 & \pi104 ) | ( \pi103 & \pi104 ) ;
  assign w3730 = \pi000 ^ w3729 ;
  assign w3731 = ( \pi002 & \pi104 ) | ( \pi002 & ~w3730 ) | ( \pi104 & ~w3730 ) ;
  assign w3732 = ( \pi002 & \pi103 ) | ( \pi002 & w3730 ) | ( \pi103 & w3730 ) ;
  assign w3733 = \pi001 & w3732 ;
  assign w3734 = ( ~\pi000 & \pi102 ) | ( ~\pi000 & w3733 ) | ( \pi102 & w3733 ) ;
  assign w3735 = ( \pi001 & \pi002 ) | ( \pi001 & ~w3734 ) | ( \pi002 & ~w3734 ) ;
  assign w3736 = ( w3731 & w3733 ) | ( w3731 & ~w3735 ) | ( w3733 & ~w3735 ) ;
  assign w3737 = ( \pi101 & ~\pi103 ) | ( \pi101 & w3282 ) | ( ~\pi103 & w3282 ) ;
  assign w3738 = ( ~\pi102 & \pi103 ) | ( ~\pi102 & w3737 ) | ( \pi103 & w3737 ) ;
  assign w3739 = \pi104 ^ w3737 ;
  assign w3740 = w3738 ^ w3739 ;
  assign w3741 = \pi002 ^ w3736 ;
  assign w3742 = \pi000 & ~w3736 ;
  assign w3743 = w3740 & w3742 ;
  assign w3744 = \pi001 ^ w3743 ;
  assign w3745 = ( \pi001 & w3741 ) | ( \pi001 & ~w3744 ) | ( w3741 & ~w3744 ) ;
  assign w3746 = w3578 ^ w3728 ;
  assign w3747 = w3745 ^ w3746 ;
  assign w3748 = ( w3578 & w3728 ) | ( w3578 & w3745 ) | ( w3728 & w3745 ) ;
  assign w3749 = ( w3579 & w3587 ) | ( w3579 & w3726 ) | ( w3587 & w3726 ) ;
  assign w3750 = ( w3588 & w3596 ) | ( w3588 & w3724 ) | ( w3596 & w3724 ) ;
  assign w3751 = ~\pi098 & w305 ;
  assign w3752 = \pi097 & w328 ;
  assign w3753 = ( w305 & ~w3751 ) | ( w305 & w3752 ) | ( ~w3751 & w3752 ) ;
  assign w3754 = ~\pi099 & w307 ;
  assign w3755 = w2966 | w3753 ;
  assign w3756 = ( w308 & w3753 ) | ( w308 & w3755 ) | ( w3753 & w3755 ) ;
  assign w3757 = ( w307 & ~w3754 ) | ( w307 & w3756 ) | ( ~w3754 & w3756 ) ;
  assign w3758 = \pi008 ^ w3757 ;
  assign w3759 = ( w3597 & w3714 ) | ( w3597 & w3722 ) | ( w3714 & w3722 ) ;
  assign w3760 = ~\pi095 & w432 ;
  assign w3761 = \pi094 & w486 ;
  assign w3762 = ( w432 & ~w3760 ) | ( w432 & w3761 ) | ( ~w3760 & w3761 ) ;
  assign w3763 = ~\pi096 & w434 ;
  assign w3764 = w2546 | w3762 ;
  assign w3765 = ( w435 & w3762 ) | ( w435 & w3764 ) | ( w3762 & w3764 ) ;
  assign w3766 = ( w434 & ~w3763 ) | ( w434 & w3765 ) | ( ~w3763 & w3765 ) ;
  assign w3767 = \pi011 ^ w3766 ;
  assign w3768 = ( w3598 & w3606 ) | ( w3598 & w3712 ) | ( w3606 & w3712 ) ;
  assign w3769 = ~\pi092 & w601 ;
  assign w3770 = \pi091 & w683 ;
  assign w3771 = ( w601 & ~w3769 ) | ( w601 & w3770 ) | ( ~w3769 & w3770 ) ;
  assign w3772 = ~\pi093 & w603 ;
  assign w3773 = w2155 | w3771 ;
  assign w3774 = ( w604 & w3771 ) | ( w604 & w3773 ) | ( w3771 & w3773 ) ;
  assign w3775 = ( w603 & ~w3772 ) | ( w603 & w3774 ) | ( ~w3772 & w3774 ) ;
  assign w3776 = \pi014 ^ w3775 ;
  assign w3777 = ( w3701 & w3709 ) | ( w3701 & w3710 ) | ( w3709 & w3710 ) ;
  assign w3778 = ( w3690 & w3698 ) | ( w3690 & w3699 ) | ( w3698 & w3699 ) ;
  assign w3779 = ~\pi083 & w1313 ;
  assign w3780 = \pi082 & w1417 ;
  assign w3781 = ( w1313 & ~w3779 ) | ( w1313 & w3780 ) | ( ~w3779 & w3780 ) ;
  assign w3782 = ~\pi084 & w1315 ;
  assign w3783 = w1188 | w3781 ;
  assign w3784 = ( w1316 & w3781 ) | ( w1316 & w3783 ) | ( w3781 & w3783 ) ;
  assign w3785 = ( w1315 & ~w3782 ) | ( w1315 & w3784 ) | ( ~w3782 & w3784 ) ;
  assign w3786 = \pi023 ^ w3785 ;
  assign w3787 = ( w3614 & w3676 ) | ( w3614 & w3677 ) | ( w3676 & w3677 ) ;
  assign w3788 = ~\pi080 & w1629 ;
  assign w3789 = \pi079 & w1722 ;
  assign w3790 = ( w1629 & ~w3788 ) | ( w1629 & w3789 ) | ( ~w3788 & w3789 ) ;
  assign w3791 = ~\pi081 & w1631 ;
  assign w3792 = w874 | w3790 ;
  assign w3793 = ( w1632 & w3790 ) | ( w1632 & w3792 ) | ( w3790 & w3792 ) ;
  assign w3794 = ( w1631 & ~w3791 ) | ( w1631 & w3793 ) | ( ~w3791 & w3793 ) ;
  assign w3795 = \pi026 ^ w3794 ;
  assign w3796 = ( w3615 & w3666 ) | ( w3615 & w3674 ) | ( w3666 & w3674 ) ;
  assign w3797 = ~\pi077 & w1944 ;
  assign w3798 = \pi076 & w2072 ;
  assign w3799 = ( w1944 & ~w3797 ) | ( w1944 & w3798 ) | ( ~w3797 & w3798 ) ;
  assign w3800 = ~\pi078 & w1946 ;
  assign w3801 = w665 | w3799 ;
  assign w3802 = ( w1947 & w3799 ) | ( w1947 & w3801 ) | ( w3799 & w3801 ) ;
  assign w3803 = ( w1946 & ~w3800 ) | ( w1946 & w3802 ) | ( ~w3800 & w3802 ) ;
  assign w3804 = \pi029 ^ w3803 ;
  assign w3805 = ( w3624 & w3652 ) | ( w3624 & w3653 ) | ( w3652 & w3653 ) ;
  assign w3806 = ~\pi071 & w2712 ;
  assign w3807 = \pi070 & w2872 ;
  assign w3808 = ( w2712 & ~w3806 ) | ( w2712 & w3807 ) | ( ~w3806 & w3807 ) ;
  assign w3809 = ~\pi072 & w2714 ;
  assign w3810 = w361 | w3808 ;
  assign w3811 = ( w2715 & w3808 ) | ( w2715 & w3810 ) | ( w3808 & w3810 ) ;
  assign w3812 = ( w2714 & ~w3809 ) | ( w2714 & w3811 ) | ( ~w3809 & w3811 ) ;
  assign w3813 = \pi035 ^ w3812 ;
  assign w3814 = ( w3625 & w3633 ) | ( w3625 & w3650 ) | ( w3633 & w3650 ) ;
  assign w3815 = ( \pi039 & ~\pi040 ) | ( \pi039 & \pi041 ) | ( ~\pi040 & \pi041 ) ;
  assign w3816 = ( \pi038 & \pi039 ) | ( \pi038 & w3815 ) | ( \pi039 & w3815 ) ;
  assign w3817 = w3815 ^ w3816 ;
  assign w3818 = \pi064 & w3817 ;
  assign w3819 = ( \pi066 & w3637 ) | ( \pi066 & w3818 ) | ( w3637 & w3818 ) ;
  assign w3820 = \pi065 | w3819 ;
  assign w3821 = ( w3635 & w3819 ) | ( w3635 & w3820 ) | ( w3819 & w3820 ) ;
  assign w3822 = w3818 | w3821 ;
  assign w3823 = ~w134 & w3638 ;
  assign w3824 = ( w3638 & w3822 ) | ( w3638 & ~w3823 ) | ( w3822 & ~w3823 ) ;
  assign w3825 = \pi041 ^ w3824 ;
  assign w3826 = w3645 & w3825 ;
  assign w3827 = w3645 ^ w3825 ;
  assign w3828 = ~\pi068 & w3178 ;
  assign w3829 = \pi067 & w3340 ;
  assign w3830 = ( w3178 & ~w3828 ) | ( w3178 & w3829 ) | ( ~w3828 & w3829 ) ;
  assign w3831 = ~\pi069 & w3180 ;
  assign w3832 = w221 | w3830 ;
  assign w3833 = ( w3181 & w3830 ) | ( w3181 & w3832 ) | ( w3830 & w3832 ) ;
  assign w3834 = ( w3180 & ~w3831 ) | ( w3180 & w3833 ) | ( ~w3831 & w3833 ) ;
  assign w3835 = \pi038 ^ w3834 ;
  assign w3836 = w3814 ^ w3827 ;
  assign w3837 = w3835 ^ w3836 ;
  assign w3838 = w3805 ^ w3837 ;
  assign w3839 = w3813 ^ w3838 ;
  assign w3840 = ~\pi074 & w2310 ;
  assign w3841 = \pi073 & w2443 ;
  assign w3842 = ( w2310 & ~w3840 ) | ( w2310 & w3841 ) | ( ~w3840 & w3841 ) ;
  assign w3843 = ~\pi075 & w2312 ;
  assign w3844 = w519 | w3842 ;
  assign w3845 = ( w2313 & w3842 ) | ( w2313 & w3844 ) | ( w3842 & w3844 ) ;
  assign w3846 = ( w2312 & ~w3843 ) | ( w2312 & w3845 ) | ( ~w3843 & w3845 ) ;
  assign w3847 = \pi032 ^ w3846 ;
  assign w3848 = w3664 ^ w3839 ;
  assign w3849 = w3847 ^ w3848 ;
  assign w3850 = w3796 ^ w3849 ;
  assign w3851 = w3804 ^ w3850 ;
  assign w3852 = w3787 ^ w3851 ;
  assign w3853 = w3795 ^ w3852 ;
  assign w3854 = ( w3679 & w3687 ) | ( w3679 & w3688 ) | ( w3687 & w3688 ) ;
  assign w3855 = w3853 ^ w3854 ;
  assign w3856 = w3786 ^ w3855 ;
  assign w3857 = ~\pi086 & w1044 ;
  assign w3858 = \pi085 & w1138 ;
  assign w3859 = ( w1044 & ~w3857 ) | ( w1044 & w3858 ) | ( ~w3857 & w3858 ) ;
  assign w3860 = ~\pi087 & w1046 ;
  assign w3861 = w1477 | w3859 ;
  assign w3862 = ( w1047 & w3859 ) | ( w1047 & w3861 ) | ( w3859 & w3861 ) ;
  assign w3863 = ( w1046 & ~w3860 ) | ( w1046 & w3862 ) | ( ~w3860 & w3862 ) ;
  assign w3864 = \pi020 ^ w3863 ;
  assign w3865 = ( w3778 & w3856 ) | ( w3778 & w3864 ) | ( w3856 & w3864 ) ;
  assign w3866 = w3778 ^ w3856 ;
  assign w3867 = w3864 ^ w3866 ;
  assign w3868 = ~\pi089 & w837 ;
  assign w3869 = \pi088 & w902 ;
  assign w3870 = ( w837 & ~w3868 ) | ( w837 & w3869 ) | ( ~w3868 & w3869 ) ;
  assign w3871 = ~\pi090 & w839 ;
  assign w3872 = w1801 | w3870 ;
  assign w3873 = ( w840 & w3870 ) | ( w840 & w3872 ) | ( w3870 & w3872 ) ;
  assign w3874 = ( w839 & ~w3871 ) | ( w839 & w3873 ) | ( ~w3871 & w3873 ) ;
  assign w3875 = \pi017 ^ w3874 ;
  assign w3876 = w3777 ^ w3867 ;
  assign w3877 = w3875 ^ w3876 ;
  assign w3878 = w3768 ^ w3877 ;
  assign w3879 = w3776 ^ w3878 ;
  assign w3880 = w3759 ^ w3879 ;
  assign w3881 = w3767 ^ w3880 ;
  assign w3882 = w3750 ^ w3881 ;
  assign w3883 = w3758 ^ w3882 ;
  assign w3884 = ~\pi101 & w189 ;
  assign w3885 = \pi100 & w229 ;
  assign w3886 = ( w189 & ~w3884 ) | ( w189 & w3885 ) | ( ~w3884 & w3885 ) ;
  assign w3887 = ~\pi102 & w191 ;
  assign w3888 = w3284 | w3886 ;
  assign w3889 = ( w192 & w3886 ) | ( w192 & w3888 ) | ( w3886 & w3888 ) ;
  assign w3890 = ( w191 & ~w3887 ) | ( w191 & w3889 ) | ( ~w3887 & w3889 ) ;
  assign w3891 = \pi005 ^ w3890 ;
  assign w3892 = w3749 ^ w3883 ;
  assign w3893 = w3891 ^ w3892 ;
  assign w3894 = ( ~\pi002 & \pi104 ) | ( ~\pi002 & \pi105 ) | ( \pi104 & \pi105 ) ;
  assign w3895 = \pi000 ^ w3894 ;
  assign w3896 = ( \pi002 & \pi105 ) | ( \pi002 & ~w3895 ) | ( \pi105 & ~w3895 ) ;
  assign w3897 = ( \pi002 & \pi104 ) | ( \pi002 & w3895 ) | ( \pi104 & w3895 ) ;
  assign w3898 = \pi001 & w3897 ;
  assign w3899 = ( ~\pi000 & \pi103 ) | ( ~\pi000 & w3898 ) | ( \pi103 & w3898 ) ;
  assign w3900 = ( \pi001 & \pi002 ) | ( \pi001 & ~w3899 ) | ( \pi002 & ~w3899 ) ;
  assign w3901 = ( w3896 & w3898 ) | ( w3896 & ~w3900 ) | ( w3898 & ~w3900 ) ;
  assign w3902 = ( \pi102 & \pi103 ) | ( \pi102 & \pi104 ) | ( \pi103 & \pi104 ) ;
  assign w3903 = ( \pi103 & w3435 ) | ( \pi103 & w3902 ) | ( w3435 & w3902 ) ;
  assign w3904 = \pi104 ^ \pi105 ;
  assign w3905 = w3903 ^ w3904 ;
  assign w3906 = \pi002 ^ w3901 ;
  assign w3907 = \pi000 & ~w3901 ;
  assign w3908 = w3905 & w3907 ;
  assign w3909 = \pi001 ^ w3908 ;
  assign w3910 = ( \pi001 & w3906 ) | ( \pi001 & ~w3909 ) | ( w3906 & ~w3909 ) ;
  assign w3911 = w3748 ^ w3893 ;
  assign w3912 = w3910 ^ w3911 ;
  assign w3913 = ( w3749 & w3883 ) | ( w3749 & w3891 ) | ( w3883 & w3891 ) ;
  assign w3914 = ~\pi102 & w189 ;
  assign w3915 = \pi101 & w229 ;
  assign w3916 = ( w189 & ~w3914 ) | ( w189 & w3915 ) | ( ~w3914 & w3915 ) ;
  assign w3917 = ~\pi103 & w191 ;
  assign w3918 = w3437 | w3916 ;
  assign w3919 = ( w192 & w3916 ) | ( w192 & w3918 ) | ( w3916 & w3918 ) ;
  assign w3920 = ( w191 & ~w3917 ) | ( w191 & w3919 ) | ( ~w3917 & w3919 ) ;
  assign w3921 = \pi005 ^ w3920 ;
  assign w3922 = ( w3750 & w3758 ) | ( w3750 & w3881 ) | ( w3758 & w3881 ) ;
  assign w3923 = ( w3759 & w3767 ) | ( w3759 & w3879 ) | ( w3767 & w3879 ) ;
  assign w3924 = ~\pi096 & w432 ;
  assign w3925 = \pi095 & w486 ;
  assign w3926 = ( w432 & ~w3924 ) | ( w432 & w3925 ) | ( ~w3924 & w3925 ) ;
  assign w3927 = ~\pi097 & w434 ;
  assign w3928 = w2673 | w3926 ;
  assign w3929 = ( w435 & w3926 ) | ( w435 & w3928 ) | ( w3926 & w3928 ) ;
  assign w3930 = ( w434 & ~w3927 ) | ( w434 & w3929 ) | ( ~w3927 & w3929 ) ;
  assign w3931 = \pi011 ^ w3930 ;
  assign w3932 = ( w3768 & w3776 ) | ( w3768 & w3877 ) | ( w3776 & w3877 ) ;
  assign w3933 = ( w3777 & w3867 ) | ( w3777 & w3875 ) | ( w3867 & w3875 ) ;
  assign w3934 = ~\pi090 & w837 ;
  assign w3935 = \pi089 & w902 ;
  assign w3936 = ( w837 & ~w3934 ) | ( w837 & w3935 ) | ( ~w3934 & w3935 ) ;
  assign w3937 = ~\pi091 & w839 ;
  assign w3938 = w1908 | w3936 ;
  assign w3939 = ( w840 & w3936 ) | ( w840 & w3938 ) | ( w3936 & w3938 ) ;
  assign w3940 = ( w839 & ~w3937 ) | ( w839 & w3939 ) | ( ~w3937 & w3939 ) ;
  assign w3941 = \pi017 ^ w3940 ;
  assign w3942 = ~\pi084 & w1313 ;
  assign w3943 = \pi083 & w1417 ;
  assign w3944 = ( w1313 & ~w3942 ) | ( w1313 & w3943 ) | ( ~w3942 & w3943 ) ;
  assign w3945 = ~\pi085 & w1315 ;
  assign w3946 = w1274 | w3944 ;
  assign w3947 = ( w1316 & w3944 ) | ( w1316 & w3946 ) | ( w3944 & w3946 ) ;
  assign w3948 = ( w1315 & ~w3945 ) | ( w1315 & w3947 ) | ( ~w3945 & w3947 ) ;
  assign w3949 = \pi023 ^ w3948 ;
  assign w3950 = ( w3787 & w3795 ) | ( w3787 & w3851 ) | ( w3795 & w3851 ) ;
  assign w3951 = ( w3796 & w3804 ) | ( w3796 & w3849 ) | ( w3804 & w3849 ) ;
  assign w3952 = ( w3664 & w3839 ) | ( w3664 & w3847 ) | ( w3839 & w3847 ) ;
  assign w3953 = ~\pi075 & w2310 ;
  assign w3954 = \pi074 & w2443 ;
  assign w3955 = ( w2310 & ~w3953 ) | ( w2310 & w3954 ) | ( ~w3953 & w3954 ) ;
  assign w3956 = ~\pi076 & w2312 ;
  assign w3957 = w538 | w3955 ;
  assign w3958 = ( w2313 & w3955 ) | ( w2313 & w3957 ) | ( w3955 & w3957 ) ;
  assign w3959 = ( w2312 & ~w3956 ) | ( w2312 & w3958 ) | ( ~w3956 & w3958 ) ;
  assign w3960 = \pi032 ^ w3959 ;
  assign w3961 = ( w3805 & w3813 ) | ( w3805 & w3837 ) | ( w3813 & w3837 ) ;
  assign w3962 = ~\pi069 & w3178 ;
  assign w3963 = \pi068 & w3340 ;
  assign w3964 = ( w3178 & ~w3962 ) | ( w3178 & w3963 ) | ( ~w3962 & w3963 ) ;
  assign w3965 = ~\pi070 & w3180 ;
  assign w3966 = w271 | w3964 ;
  assign w3967 = ( w3181 & w3964 ) | ( w3181 & w3966 ) | ( w3964 & w3966 ) ;
  assign w3968 = ( w3180 & ~w3965 ) | ( w3180 & w3967 ) | ( ~w3965 & w3967 ) ;
  assign w3969 = \pi038 ^ w3968 ;
  assign w3970 = ~\pi066 & w3635 ;
  assign w3971 = \pi065 & w3817 ;
  assign w3972 = ( w3635 & ~w3970 ) | ( w3635 & w3971 ) | ( ~w3970 & w3971 ) ;
  assign w3973 = ~\pi067 & w3637 ;
  assign w3974 = w160 | w3972 ;
  assign w3975 = ( w3638 & w3972 ) | ( w3638 & w3974 ) | ( w3972 & w3974 ) ;
  assign w3976 = ( w3637 & ~w3973 ) | ( w3637 & w3975 ) | ( ~w3973 & w3975 ) ;
  assign w3977 = \pi041 ^ w3976 ;
  assign w3978 = w3826 ^ w3977 ;
  assign w3979 = \pi041 ^ \pi042 ;
  assign w3980 = \pi064 & w3979 ;
  assign w3981 = w3978 ^ w3980 ;
  assign w3982 = ( w3814 & w3827 ) | ( w3814 & w3835 ) | ( w3827 & w3835 ) ;
  assign w3983 = w3981 ^ w3982 ;
  assign w3984 = w3969 ^ w3983 ;
  assign w3985 = ~\pi072 & w2712 ;
  assign w3986 = \pi071 & w2872 ;
  assign w3987 = ( w2712 & ~w3985 ) | ( w2712 & w3986 ) | ( ~w3985 & w3986 ) ;
  assign w3988 = ~\pi073 & w2714 ;
  assign w3989 = w404 | w3987 ;
  assign w3990 = ( w2715 & w3987 ) | ( w2715 & w3989 ) | ( w3987 & w3989 ) ;
  assign w3991 = ( w2714 & ~w3988 ) | ( w2714 & w3990 ) | ( ~w3988 & w3990 ) ;
  assign w3992 = \pi035 ^ w3991 ;
  assign w3993 = w3961 ^ w3984 ;
  assign w3994 = w3992 ^ w3993 ;
  assign w3995 = w3952 ^ w3994 ;
  assign w3996 = w3960 ^ w3995 ;
  assign w3997 = ~\pi078 & w1944 ;
  assign w3998 = \pi077 & w2072 ;
  assign w3999 = ( w1944 & ~w3997 ) | ( w1944 & w3998 ) | ( ~w3997 & w3998 ) ;
  assign w4000 = ~\pi079 & w1946 ;
  assign w4001 = w730 | w3999 ;
  assign w4002 = ( w1947 & w3999 ) | ( w1947 & w4001 ) | ( w3999 & w4001 ) ;
  assign w4003 = ( w1946 & ~w4000 ) | ( w1946 & w4002 ) | ( ~w4000 & w4002 ) ;
  assign w4004 = \pi029 ^ w4003 ;
  assign w4005 = w3951 ^ w3996 ;
  assign w4006 = w4004 ^ w4005 ;
  assign w4007 = ~\pi081 & w1629 ;
  assign w4008 = \pi080 & w1722 ;
  assign w4009 = ( w1629 & ~w4007 ) | ( w1629 & w4008 ) | ( ~w4007 & w4008 ) ;
  assign w4010 = ~\pi082 & w1631 ;
  assign w4011 = w1008 | w4009 ;
  assign w4012 = ( w1632 & w4009 ) | ( w1632 & w4011 ) | ( w4009 & w4011 ) ;
  assign w4013 = ( w1631 & ~w4010 ) | ( w1631 & w4012 ) | ( ~w4010 & w4012 ) ;
  assign w4014 = \pi026 ^ w4013 ;
  assign w4015 = w3950 ^ w4006 ;
  assign w4016 = w4014 ^ w4015 ;
  assign w4017 = ( w3786 & w3853 ) | ( w3786 & w3854 ) | ( w3853 & w3854 ) ;
  assign w4018 = w4016 ^ w4017 ;
  assign w4019 = w3949 ^ w4018 ;
  assign w4020 = ~\pi087 & w1044 ;
  assign w4021 = \pi086 & w1138 ;
  assign w4022 = ( w1044 & ~w4020 ) | ( w1044 & w4021 ) | ( ~w4020 & w4021 ) ;
  assign w4023 = ~\pi088 & w1046 ;
  assign w4024 = w1574 | w4022 ;
  assign w4025 = ( w1047 & w4022 ) | ( w1047 & w4024 ) | ( w4022 & w4024 ) ;
  assign w4026 = ( w1046 & ~w4023 ) | ( w1046 & w4025 ) | ( ~w4023 & w4025 ) ;
  assign w4027 = \pi020 ^ w4026 ;
  assign w4028 = w3865 ^ w4019 ;
  assign w4029 = w4027 ^ w4028 ;
  assign w4030 = w3933 ^ w4029 ;
  assign w4031 = w3941 ^ w4030 ;
  assign w4032 = ~\pi093 & w601 ;
  assign w4033 = \pi092 & w683 ;
  assign w4034 = ( w601 & ~w4032 ) | ( w601 & w4033 ) | ( ~w4032 & w4033 ) ;
  assign w4035 = ~\pi094 & w603 ;
  assign w4036 = w2274 | w4034 ;
  assign w4037 = ( w604 & w4034 ) | ( w604 & w4036 ) | ( w4034 & w4036 ) ;
  assign w4038 = ( w603 & ~w4035 ) | ( w603 & w4037 ) | ( ~w4035 & w4037 ) ;
  assign w4039 = \pi014 ^ w4038 ;
  assign w4040 = w3932 ^ w4031 ;
  assign w4041 = w4039 ^ w4040 ;
  assign w4042 = w3923 ^ w4041 ;
  assign w4043 = w3931 ^ w4042 ;
  assign w4044 = ~\pi099 & w305 ;
  assign w4045 = \pi098 & w328 ;
  assign w4046 = ( w305 & ~w4044 ) | ( w305 & w4045 ) | ( ~w4044 & w4045 ) ;
  assign w4047 = ~\pi100 & w307 ;
  assign w4048 = w3104 | w4046 ;
  assign w4049 = ( w308 & w4046 ) | ( w308 & w4048 ) | ( w4046 & w4048 ) ;
  assign w4050 = ( w307 & ~w4047 ) | ( w307 & w4049 ) | ( ~w4047 & w4049 ) ;
  assign w4051 = \pi008 ^ w4050 ;
  assign w4052 = w3922 ^ w4043 ;
  assign w4053 = w4051 ^ w4052 ;
  assign w4054 = w3913 ^ w4053 ;
  assign w4055 = w3921 ^ w4054 ;
  assign w4056 = ( ~\pi002 & \pi105 ) | ( ~\pi002 & \pi106 ) | ( \pi105 & \pi106 ) ;
  assign w4057 = \pi000 ^ w4056 ;
  assign w4058 = ( \pi002 & \pi106 ) | ( \pi002 & ~w4057 ) | ( \pi106 & ~w4057 ) ;
  assign w4059 = ( \pi002 & \pi105 ) | ( \pi002 & w4057 ) | ( \pi105 & w4057 ) ;
  assign w4060 = \pi001 & w4059 ;
  assign w4061 = ( ~\pi000 & \pi104 ) | ( ~\pi000 & w4060 ) | ( \pi104 & w4060 ) ;
  assign w4062 = ( \pi001 & \pi002 ) | ( \pi001 & ~w4061 ) | ( \pi002 & ~w4061 ) ;
  assign w4063 = ( w4058 & w4060 ) | ( w4058 & ~w4062 ) | ( w4060 & ~w4062 ) ;
  assign w4064 = ( \pi102 & \pi103 ) | ( \pi102 & ~\pi105 ) | ( \pi103 & ~\pi105 ) ;
  assign w4065 = ( \pi103 & w3435 ) | ( \pi103 & w4064 ) | ( w3435 & w4064 ) ;
  assign w4066 = ( \pi104 & \pi105 ) | ( \pi104 & w4065 ) | ( \pi105 & w4065 ) ;
  assign w4067 = \pi105 ^ w4066 ;
  assign w4068 = \pi106 ^ w4067 ;
  assign w4069 = \pi002 ^ w4063 ;
  assign w4070 = \pi000 & ~w4063 ;
  assign w4071 = w4068 & w4070 ;
  assign w4072 = \pi001 ^ w4071 ;
  assign w4073 = ( \pi001 & w4069 ) | ( \pi001 & ~w4072 ) | ( w4069 & ~w4072 ) ;
  assign w4074 = ( w3748 & w3893 ) | ( w3748 & w3910 ) | ( w3893 & w3910 ) ;
  assign w4075 = w4055 ^ w4074 ;
  assign w4076 = w4073 ^ w4075 ;
  assign w4077 = ( ~\pi002 & \pi106 ) | ( ~\pi002 & \pi107 ) | ( \pi106 & \pi107 ) ;
  assign w4078 = \pi000 ^ w4077 ;
  assign w4079 = ( \pi002 & \pi107 ) | ( \pi002 & ~w4078 ) | ( \pi107 & ~w4078 ) ;
  assign w4080 = ( \pi002 & \pi106 ) | ( \pi002 & w4078 ) | ( \pi106 & w4078 ) ;
  assign w4081 = \pi001 & w4080 ;
  assign w4082 = ( ~\pi000 & \pi105 ) | ( ~\pi000 & w4081 ) | ( \pi105 & w4081 ) ;
  assign w4083 = ( \pi001 & \pi002 ) | ( \pi001 & ~w4082 ) | ( \pi002 & ~w4082 ) ;
  assign w4084 = ( w4079 & w4081 ) | ( w4079 & ~w4083 ) | ( w4081 & ~w4083 ) ;
  assign w4085 = ( \pi105 & \pi106 ) | ( \pi105 & w4066 ) | ( \pi106 & w4066 ) ;
  assign w4086 = \pi106 ^ w4085 ;
  assign w4087 = \pi107 ^ w4086 ;
  assign w4088 = \pi002 ^ w4084 ;
  assign w4089 = \pi000 & ~w4084 ;
  assign w4090 = w4087 & w4089 ;
  assign w4091 = \pi001 ^ w4090 ;
  assign w4092 = ( \pi001 & w4088 ) | ( \pi001 & ~w4091 ) | ( w4088 & ~w4091 ) ;
  assign w4093 = ( w3913 & w3921 ) | ( w3913 & w4053 ) | ( w3921 & w4053 ) ;
  assign w4094 = ( w3922 & w4043 ) | ( w3922 & w4051 ) | ( w4043 & w4051 ) ;
  assign w4095 = ~\pi097 & w432 ;
  assign w4096 = \pi096 & w486 ;
  assign w4097 = ( w432 & ~w4095 ) | ( w432 & w4096 ) | ( ~w4095 & w4096 ) ;
  assign w4098 = ~\pi098 & w434 ;
  assign w4099 = w2824 | w4097 ;
  assign w4100 = ( w435 & w4097 ) | ( w435 & w4099 ) | ( w4097 & w4099 ) ;
  assign w4101 = ( w434 & ~w4098 ) | ( w434 & w4100 ) | ( ~w4098 & w4100 ) ;
  assign w4102 = \pi011 ^ w4101 ;
  assign w4103 = ( w3932 & w4031 ) | ( w3932 & w4039 ) | ( w4031 & w4039 ) ;
  assign w4104 = ( w3933 & w3941 ) | ( w3933 & w4029 ) | ( w3941 & w4029 ) ;
  assign w4105 = ~\pi091 & w837 ;
  assign w4106 = \pi090 & w902 ;
  assign w4107 = ( w837 & ~w4105 ) | ( w837 & w4106 ) | ( ~w4105 & w4106 ) ;
  assign w4108 = ~\pi092 & w839 ;
  assign w4109 = w2033 | w4107 ;
  assign w4110 = ( w840 & w4107 ) | ( w840 & w4109 ) | ( w4107 & w4109 ) ;
  assign w4111 = ( w839 & ~w4108 ) | ( w839 & w4110 ) | ( ~w4108 & w4110 ) ;
  assign w4112 = \pi017 ^ w4111 ;
  assign w4113 = ~\pi079 & w1944 ;
  assign w4114 = \pi078 & w2072 ;
  assign w4115 = ( w1944 & ~w4113 ) | ( w1944 & w4114 ) | ( ~w4113 & w4114 ) ;
  assign w4116 = ~\pi080 & w1946 ;
  assign w4117 = w794 | w4115 ;
  assign w4118 = ( w1947 & w4115 ) | ( w1947 & w4117 ) | ( w4115 & w4117 ) ;
  assign w4119 = ( w1946 & ~w4116 ) | ( w1946 & w4118 ) | ( ~w4116 & w4118 ) ;
  assign w4120 = \pi029 ^ w4119 ;
  assign w4121 = ( w3952 & w3960 ) | ( w3952 & w3994 ) | ( w3960 & w3994 ) ;
  assign w4122 = ( w3961 & w3984 ) | ( w3961 & w3992 ) | ( w3984 & w3992 ) ;
  assign w4123 = ~\pi070 & w3178 ;
  assign w4124 = \pi069 & w3340 ;
  assign w4125 = ( w3178 & ~w4123 ) | ( w3178 & w4124 ) | ( ~w4123 & w4124 ) ;
  assign w4126 = ~\pi071 & w3180 ;
  assign w4127 = w290 | w4125 ;
  assign w4128 = ( w3181 & w4125 ) | ( w3181 & w4127 ) | ( w4125 & w4127 ) ;
  assign w4129 = ( w3180 & ~w4126 ) | ( w3180 & w4128 ) | ( ~w4126 & w4128 ) ;
  assign w4130 = \pi038 ^ w4129 ;
  assign w4131 = ( w3826 & w3977 ) | ( w3826 & w3980 ) | ( w3977 & w3980 ) ;
  assign w4132 = ~\pi067 & w3635 ;
  assign w4133 = \pi066 & w3817 ;
  assign w4134 = ( w3635 & ~w4132 ) | ( w3635 & w4133 ) | ( ~w4132 & w4133 ) ;
  assign w4135 = ~\pi068 & w3637 ;
  assign w4136 = w182 | w4134 ;
  assign w4137 = ( w3638 & w4134 ) | ( w3638 & w4136 ) | ( w4134 & w4136 ) ;
  assign w4138 = ( w3637 & ~w4135 ) | ( w3637 & w4137 ) | ( ~w4135 & w4137 ) ;
  assign w4139 = \pi041 ^ w4138 ;
  assign w4140 = ( \pi041 & \pi042 ) | ( \pi041 & \pi043 ) | ( \pi042 & \pi043 ) ;
  assign w4141 = \pi043 ^ w4140 ;
  assign w4142 = \pi043 ^ \pi044 ;
  assign w4143 = w3979 & ~w4142 ;
  assign w4144 = w3979 & w4142 ;
  assign w4145 = ( \pi041 & \pi042 ) | ( \pi041 & ~\pi044 ) | ( \pi042 & ~\pi044 ) ;
  assign w4146 = \pi044 & ~\pi064 ;
  assign w4147 = ~\pi065 & w4146 ;
  assign w4148 = ( \pi041 & \pi042 ) | ( \pi041 & ~w4147 ) | ( \pi042 & ~w4147 ) ;
  assign w4149 = ( \pi043 & \pi044 ) | ( \pi043 & ~w4148 ) | ( \pi044 & ~w4148 ) ;
  assign w4150 = ( \pi043 & ~w4146 ) | ( \pi043 & w4148 ) | ( ~w4146 & w4148 ) ;
  assign w4151 = ( w4145 & w4149 ) | ( w4145 & ~w4150 ) | ( w4149 & ~w4150 ) ;
  assign w4152 = ( \pi041 & \pi042 ) | ( \pi041 & \pi065 ) | ( \pi042 & \pi065 ) ;
  assign w4153 = \pi041 & \pi042 ;
  assign w4154 = \pi064 ^ w4153 ;
  assign w4155 = ( \pi043 & w4153 ) | ( \pi043 & w4154 ) | ( w4153 & w4154 ) ;
  assign w4156 = w4152 ^ w4155 ;
  assign w4157 = w4131 ^ w4139 ;
  assign w4158 = w4156 ^ w4157 ;
  assign w4159 = ( w3969 & w3981 ) | ( w3969 & w3982 ) | ( w3981 & w3982 ) ;
  assign w4160 = w4158 ^ w4159 ;
  assign w4161 = w4130 ^ w4160 ;
  assign w4162 = ~\pi073 & w2712 ;
  assign w4163 = \pi072 & w2872 ;
  assign w4164 = ( w2712 & ~w4162 ) | ( w2712 & w4163 ) | ( ~w4162 & w4163 ) ;
  assign w4165 = ~\pi074 & w2714 ;
  assign w4166 = w465 | w4164 ;
  assign w4167 = ( w2715 & w4164 ) | ( w2715 & w4166 ) | ( w4164 & w4166 ) ;
  assign w4168 = ( w2714 & ~w4165 ) | ( w2714 & w4167 ) | ( ~w4165 & w4167 ) ;
  assign w4169 = \pi035 ^ w4168 ;
  assign w4170 = ( w4122 & w4161 ) | ( w4122 & w4169 ) | ( w4161 & w4169 ) ;
  assign w4171 = w4122 ^ w4161 ;
  assign w4172 = w4169 ^ w4171 ;
  assign w4173 = ~\pi076 & w2310 ;
  assign w4174 = \pi075 & w2443 ;
  assign w4175 = ( w2310 & ~w4173 ) | ( w2310 & w4174 ) | ( ~w4173 & w4174 ) ;
  assign w4176 = ~\pi077 & w2312 ;
  assign w4177 = w644 | w4175 ;
  assign w4178 = ( w2313 & w4175 ) | ( w2313 & w4177 ) | ( w4175 & w4177 ) ;
  assign w4179 = ( w2312 & ~w4176 ) | ( w2312 & w4178 ) | ( ~w4176 & w4178 ) ;
  assign w4180 = \pi032 ^ w4179 ;
  assign w4181 = w4121 ^ w4172 ;
  assign w4182 = w4180 ^ w4181 ;
  assign w4183 = ( w3951 & w3996 ) | ( w3951 & w4004 ) | ( w3996 & w4004 ) ;
  assign w4184 = w4182 ^ w4183 ;
  assign w4185 = w4120 ^ w4184 ;
  assign w4186 = ~\pi082 & w1629 ;
  assign w4187 = \pi081 & w1722 ;
  assign w4188 = ( w1629 & ~w4186 ) | ( w1629 & w4187 ) | ( ~w4186 & w4187 ) ;
  assign w4189 = ~\pi083 & w1631 ;
  assign w4190 = w1099 | w4188 ;
  assign w4191 = ( w1632 & w4188 ) | ( w1632 & w4190 ) | ( w4188 & w4190 ) ;
  assign w4192 = ( w1631 & ~w4189 ) | ( w1631 & w4191 ) | ( ~w4189 & w4191 ) ;
  assign w4193 = \pi026 ^ w4192 ;
  assign w4194 = ( w3950 & w4006 ) | ( w3950 & w4014 ) | ( w4006 & w4014 ) ;
  assign w4195 = w4185 ^ w4194 ;
  assign w4196 = w4193 ^ w4195 ;
  assign w4197 = ~\pi085 & w1313 ;
  assign w4198 = \pi084 & w1417 ;
  assign w4199 = ( w1313 & ~w4197 ) | ( w1313 & w4198 ) | ( ~w4197 & w4198 ) ;
  assign w4200 = ~\pi086 & w1315 ;
  assign w4201 = w1379 | w4199 ;
  assign w4202 = ( w1316 & w4199 ) | ( w1316 & w4201 ) | ( w4199 & w4201 ) ;
  assign w4203 = ( w1315 & ~w4200 ) | ( w1315 & w4202 ) | ( ~w4200 & w4202 ) ;
  assign w4204 = \pi023 ^ w4203 ;
  assign w4205 = ( w3949 & w4016 ) | ( w3949 & w4017 ) | ( w4016 & w4017 ) ;
  assign w4206 = w4196 ^ w4205 ;
  assign w4207 = w4204 ^ w4206 ;
  assign w4208 = ~\pi088 & w1044 ;
  assign w4209 = \pi087 & w1138 ;
  assign w4210 = ( w1044 & ~w4208 ) | ( w1044 & w4209 ) | ( ~w4208 & w4209 ) ;
  assign w4211 = ~\pi089 & w1046 ;
  assign w4212 = w1595 | w4210 ;
  assign w4213 = ( w1047 & w4210 ) | ( w1047 & w4212 ) | ( w4210 & w4212 ) ;
  assign w4214 = ( w1046 & ~w4211 ) | ( w1046 & w4213 ) | ( ~w4211 & w4213 ) ;
  assign w4215 = \pi020 ^ w4214 ;
  assign w4216 = ( w3865 & w4019 ) | ( w3865 & w4027 ) | ( w4019 & w4027 ) ;
  assign w4217 = w4207 ^ w4216 ;
  assign w4218 = w4215 ^ w4217 ;
  assign w4219 = w4104 ^ w4218 ;
  assign w4220 = w4112 ^ w4219 ;
  assign w4221 = ~\pi094 & w601 ;
  assign w4222 = \pi093 & w683 ;
  assign w4223 = ( w601 & ~w4221 ) | ( w601 & w4222 ) | ( ~w4221 & w4222 ) ;
  assign w4224 = ~\pi095 & w603 ;
  assign w4225 = w2409 | w4223 ;
  assign w4226 = ( w604 & w4223 ) | ( w604 & w4225 ) | ( w4223 & w4225 ) ;
  assign w4227 = ( w603 & ~w4224 ) | ( w603 & w4226 ) | ( ~w4224 & w4226 ) ;
  assign w4228 = \pi014 ^ w4227 ;
  assign w4229 = w4103 ^ w4220 ;
  assign w4230 = w4228 ^ w4229 ;
  assign w4231 = ( w3923 & w3931 ) | ( w3923 & w4041 ) | ( w3931 & w4041 ) ;
  assign w4232 = w4230 ^ w4231 ;
  assign w4233 = w4102 ^ w4232 ;
  assign w4234 = ~\pi100 & w305 ;
  assign w4235 = \pi099 & w328 ;
  assign w4236 = ( w305 & ~w4234 ) | ( w305 & w4235 ) | ( ~w4234 & w4235 ) ;
  assign w4237 = ~\pi101 & w307 ;
  assign w4238 = w3264 | w4236 ;
  assign w4239 = ( w308 & w4236 ) | ( w308 & w4238 ) | ( w4236 & w4238 ) ;
  assign w4240 = ( w307 & ~w4237 ) | ( w307 & w4239 ) | ( ~w4237 & w4239 ) ;
  assign w4241 = \pi008 ^ w4240 ;
  assign w4242 = ( w4094 & w4233 ) | ( w4094 & w4241 ) | ( w4233 & w4241 ) ;
  assign w4243 = w4094 ^ w4233 ;
  assign w4244 = w4241 ^ w4243 ;
  assign w4245 = ~\pi103 & w189 ;
  assign w4246 = \pi102 & w229 ;
  assign w4247 = ( w189 & ~w4245 ) | ( w189 & w4246 ) | ( ~w4245 & w4246 ) ;
  assign w4248 = ~\pi104 & w191 ;
  assign w4249 = w3740 | w4247 ;
  assign w4250 = ( w192 & w4247 ) | ( w192 & w4249 ) | ( w4247 & w4249 ) ;
  assign w4251 = ( w191 & ~w4248 ) | ( w191 & w4250 ) | ( ~w4248 & w4250 ) ;
  assign w4252 = \pi005 ^ w4251 ;
  assign w4253 = w4093 ^ w4244 ;
  assign w4254 = w4252 ^ w4253 ;
  assign w4255 = ( w4055 & w4073 ) | ( w4055 & w4074 ) | ( w4073 & w4074 ) ;
  assign w4256 = w4254 ^ w4255 ;
  assign w4257 = w4092 ^ w4256 ;
  assign w4258 = ( w4092 & w4254 ) | ( w4092 & w4255 ) | ( w4254 & w4255 ) ;
  assign w4259 = ( w4093 & w4244 ) | ( w4093 & w4252 ) | ( w4244 & w4252 ) ;
  assign w4260 = ~\pi104 & w189 ;
  assign w4261 = \pi103 & w229 ;
  assign w4262 = ( w189 & ~w4260 ) | ( w189 & w4261 ) | ( ~w4260 & w4261 ) ;
  assign w4263 = ~\pi105 & w191 ;
  assign w4264 = w3905 | w4262 ;
  assign w4265 = ( w192 & w4262 ) | ( w192 & w4264 ) | ( w4262 & w4264 ) ;
  assign w4266 = ( w191 & ~w4263 ) | ( w191 & w4265 ) | ( ~w4263 & w4265 ) ;
  assign w4267 = \pi005 ^ w4266 ;
  assign w4268 = ~\pi098 & w432 ;
  assign w4269 = \pi097 & w486 ;
  assign w4270 = ( w432 & ~w4268 ) | ( w432 & w4269 ) | ( ~w4268 & w4269 ) ;
  assign w4271 = ~\pi099 & w434 ;
  assign w4272 = w2966 | w4270 ;
  assign w4273 = ( w435 & w4270 ) | ( w435 & w4272 ) | ( w4270 & w4272 ) ;
  assign w4274 = ( w434 & ~w4271 ) | ( w434 & w4273 ) | ( ~w4271 & w4273 ) ;
  assign w4275 = \pi011 ^ w4274 ;
  assign w4276 = ( w4103 & w4220 ) | ( w4103 & w4228 ) | ( w4220 & w4228 ) ;
  assign w4277 = ~\pi095 & w601 ;
  assign w4278 = \pi094 & w683 ;
  assign w4279 = ( w601 & ~w4277 ) | ( w601 & w4278 ) | ( ~w4277 & w4278 ) ;
  assign w4280 = ~\pi096 & w603 ;
  assign w4281 = w2546 | w4279 ;
  assign w4282 = ( w604 & w4279 ) | ( w604 & w4281 ) | ( w4279 & w4281 ) ;
  assign w4283 = ( w603 & ~w4280 ) | ( w603 & w4282 ) | ( ~w4280 & w4282 ) ;
  assign w4284 = \pi014 ^ w4283 ;
  assign w4285 = ( w4104 & w4112 ) | ( w4104 & w4218 ) | ( w4112 & w4218 ) ;
  assign w4286 = ~\pi092 & w837 ;
  assign w4287 = \pi091 & w902 ;
  assign w4288 = ( w837 & ~w4286 ) | ( w837 & w4287 ) | ( ~w4286 & w4287 ) ;
  assign w4289 = ~\pi093 & w839 ;
  assign w4290 = w2155 | w4288 ;
  assign w4291 = ( w840 & w4288 ) | ( w840 & w4290 ) | ( w4288 & w4290 ) ;
  assign w4292 = ( w839 & ~w4289 ) | ( w839 & w4291 ) | ( ~w4289 & w4291 ) ;
  assign w4293 = \pi017 ^ w4292 ;
  assign w4294 = ( w4207 & w4215 ) | ( w4207 & w4216 ) | ( w4215 & w4216 ) ;
  assign w4295 = ( w4196 & w4204 ) | ( w4196 & w4205 ) | ( w4204 & w4205 ) ;
  assign w4296 = ~\pi083 & w1629 ;
  assign w4297 = \pi082 & w1722 ;
  assign w4298 = ( w1629 & ~w4296 ) | ( w1629 & w4297 ) | ( ~w4296 & w4297 ) ;
  assign w4299 = ~\pi084 & w1631 ;
  assign w4300 = w1188 | w4298 ;
  assign w4301 = ( w1632 & w4298 ) | ( w1632 & w4300 ) | ( w4298 & w4300 ) ;
  assign w4302 = ( w1631 & ~w4299 ) | ( w1631 & w4301 ) | ( ~w4299 & w4301 ) ;
  assign w4303 = \pi026 ^ w4302 ;
  assign w4304 = ( w4120 & w4182 ) | ( w4120 & w4183 ) | ( w4182 & w4183 ) ;
  assign w4305 = ~\pi080 & w1944 ;
  assign w4306 = \pi079 & w2072 ;
  assign w4307 = ( w1944 & ~w4305 ) | ( w1944 & w4306 ) | ( ~w4305 & w4306 ) ;
  assign w4308 = ~\pi081 & w1946 ;
  assign w4309 = w874 | w4307 ;
  assign w4310 = ( w1947 & w4307 ) | ( w1947 & w4309 ) | ( w4307 & w4309 ) ;
  assign w4311 = ( w1946 & ~w4308 ) | ( w1946 & w4310 ) | ( ~w4308 & w4310 ) ;
  assign w4312 = \pi029 ^ w4311 ;
  assign w4313 = ( w4121 & w4172 ) | ( w4121 & w4180 ) | ( w4172 & w4180 ) ;
  assign w4314 = ~\pi077 & w2310 ;
  assign w4315 = \pi076 & w2443 ;
  assign w4316 = ( w2310 & ~w4314 ) | ( w2310 & w4315 ) | ( ~w4314 & w4315 ) ;
  assign w4317 = ~\pi078 & w2312 ;
  assign w4318 = w665 | w4316 ;
  assign w4319 = ( w2313 & w4316 ) | ( w2313 & w4318 ) | ( w4316 & w4318 ) ;
  assign w4320 = ( w2312 & ~w4317 ) | ( w2312 & w4319 ) | ( ~w4317 & w4319 ) ;
  assign w4321 = \pi032 ^ w4320 ;
  assign w4322 = ( w4130 & w4158 ) | ( w4130 & w4159 ) | ( w4158 & w4159 ) ;
  assign w4323 = ~\pi071 & w3178 ;
  assign w4324 = \pi070 & w3340 ;
  assign w4325 = ( w3178 & ~w4323 ) | ( w3178 & w4324 ) | ( ~w4323 & w4324 ) ;
  assign w4326 = ~\pi072 & w3180 ;
  assign w4327 = w361 | w4325 ;
  assign w4328 = ( w3181 & w4325 ) | ( w3181 & w4327 ) | ( w4325 & w4327 ) ;
  assign w4329 = ( w3180 & ~w4326 ) | ( w3180 & w4328 ) | ( ~w4326 & w4328 ) ;
  assign w4330 = \pi038 ^ w4329 ;
  assign w4331 = ( w4131 & w4139 ) | ( w4131 & w4156 ) | ( w4139 & w4156 ) ;
  assign w4332 = ( \pi042 & ~\pi043 ) | ( \pi042 & \pi044 ) | ( ~\pi043 & \pi044 ) ;
  assign w4333 = ( \pi041 & \pi042 ) | ( \pi041 & w4332 ) | ( \pi042 & w4332 ) ;
  assign w4334 = w4332 ^ w4333 ;
  assign w4335 = \pi064 & w4334 ;
  assign w4336 = ( \pi066 & w4143 ) | ( \pi066 & w4335 ) | ( w4143 & w4335 ) ;
  assign w4337 = \pi065 | w4336 ;
  assign w4338 = ( w4141 & w4336 ) | ( w4141 & w4337 ) | ( w4336 & w4337 ) ;
  assign w4339 = w4335 | w4338 ;
  assign w4340 = ~w134 & w4144 ;
  assign w4341 = ( w4144 & w4339 ) | ( w4144 & ~w4340 ) | ( w4339 & ~w4340 ) ;
  assign w4342 = \pi044 ^ w4341 ;
  assign w4343 = w4151 & w4342 ;
  assign w4344 = w4151 ^ w4342 ;
  assign w4345 = ~\pi068 & w3635 ;
  assign w4346 = \pi067 & w3817 ;
  assign w4347 = ( w3635 & ~w4345 ) | ( w3635 & w4346 ) | ( ~w4345 & w4346 ) ;
  assign w4348 = ~\pi069 & w3637 ;
  assign w4349 = w221 | w4347 ;
  assign w4350 = ( w3638 & w4347 ) | ( w3638 & w4349 ) | ( w4347 & w4349 ) ;
  assign w4351 = ( w3637 & ~w4348 ) | ( w3637 & w4350 ) | ( ~w4348 & w4350 ) ;
  assign w4352 = \pi041 ^ w4351 ;
  assign w4353 = w4331 ^ w4344 ;
  assign w4354 = w4352 ^ w4353 ;
  assign w4355 = w4322 ^ w4354 ;
  assign w4356 = w4330 ^ w4355 ;
  assign w4357 = ~\pi074 & w2712 ;
  assign w4358 = \pi073 & w2872 ;
  assign w4359 = ( w2712 & ~w4357 ) | ( w2712 & w4358 ) | ( ~w4357 & w4358 ) ;
  assign w4360 = ~\pi075 & w2714 ;
  assign w4361 = w519 | w4359 ;
  assign w4362 = ( w2715 & w4359 ) | ( w2715 & w4361 ) | ( w4359 & w4361 ) ;
  assign w4363 = ( w2714 & ~w4360 ) | ( w2714 & w4362 ) | ( ~w4360 & w4362 ) ;
  assign w4364 = \pi035 ^ w4363 ;
  assign w4365 = w4170 ^ w4356 ;
  assign w4366 = w4364 ^ w4365 ;
  assign w4367 = w4313 ^ w4366 ;
  assign w4368 = w4321 ^ w4367 ;
  assign w4369 = w4304 ^ w4368 ;
  assign w4370 = w4312 ^ w4369 ;
  assign w4371 = ( w4185 & w4193 ) | ( w4185 & w4194 ) | ( w4193 & w4194 ) ;
  assign w4372 = w4370 ^ w4371 ;
  assign w4373 = w4303 ^ w4372 ;
  assign w4374 = ~\pi086 & w1313 ;
  assign w4375 = \pi085 & w1417 ;
  assign w4376 = ( w1313 & ~w4374 ) | ( w1313 & w4375 ) | ( ~w4374 & w4375 ) ;
  assign w4377 = ~\pi087 & w1315 ;
  assign w4378 = w1477 | w4376 ;
  assign w4379 = ( w1316 & w4376 ) | ( w1316 & w4378 ) | ( w4376 & w4378 ) ;
  assign w4380 = ( w1315 & ~w4377 ) | ( w1315 & w4379 ) | ( ~w4377 & w4379 ) ;
  assign w4381 = \pi023 ^ w4380 ;
  assign w4382 = ( w4295 & w4373 ) | ( w4295 & w4381 ) | ( w4373 & w4381 ) ;
  assign w4383 = w4295 ^ w4373 ;
  assign w4384 = w4381 ^ w4383 ;
  assign w4385 = ~\pi089 & w1044 ;
  assign w4386 = \pi088 & w1138 ;
  assign w4387 = ( w1044 & ~w4385 ) | ( w1044 & w4386 ) | ( ~w4385 & w4386 ) ;
  assign w4388 = ~\pi090 & w1046 ;
  assign w4389 = w1801 | w4387 ;
  assign w4390 = ( w1047 & w4387 ) | ( w1047 & w4389 ) | ( w4387 & w4389 ) ;
  assign w4391 = ( w1046 & ~w4388 ) | ( w1046 & w4390 ) | ( ~w4388 & w4390 ) ;
  assign w4392 = \pi020 ^ w4391 ;
  assign w4393 = w4294 ^ w4384 ;
  assign w4394 = w4392 ^ w4393 ;
  assign w4395 = w4285 ^ w4394 ;
  assign w4396 = w4293 ^ w4395 ;
  assign w4397 = w4276 ^ w4396 ;
  assign w4398 = w4284 ^ w4397 ;
  assign w4399 = ( w4102 & w4230 ) | ( w4102 & w4231 ) | ( w4230 & w4231 ) ;
  assign w4400 = w4398 ^ w4399 ;
  assign w4401 = w4275 ^ w4400 ;
  assign w4402 = ~\pi101 & w305 ;
  assign w4403 = \pi100 & w328 ;
  assign w4404 = ( w305 & ~w4402 ) | ( w305 & w4403 ) | ( ~w4402 & w4403 ) ;
  assign w4405 = ~\pi102 & w307 ;
  assign w4406 = w3284 | w4404 ;
  assign w4407 = ( w308 & w4404 ) | ( w308 & w4406 ) | ( w4404 & w4406 ) ;
  assign w4408 = ( w307 & ~w4405 ) | ( w307 & w4407 ) | ( ~w4405 & w4407 ) ;
  assign w4409 = \pi008 ^ w4408 ;
  assign w4410 = w4242 ^ w4401 ;
  assign w4411 = w4409 ^ w4410 ;
  assign w4412 = w4259 ^ w4411 ;
  assign w4413 = w4267 ^ w4412 ;
  assign w4414 = ( ~\pi002 & \pi107 ) | ( ~\pi002 & \pi108 ) | ( \pi107 & \pi108 ) ;
  assign w4415 = \pi000 ^ w4414 ;
  assign w4416 = ( \pi002 & \pi108 ) | ( \pi002 & ~w4415 ) | ( \pi108 & ~w4415 ) ;
  assign w4417 = ( \pi002 & \pi107 ) | ( \pi002 & w4415 ) | ( \pi107 & w4415 ) ;
  assign w4418 = \pi001 & w4417 ;
  assign w4419 = ( ~\pi000 & \pi106 ) | ( ~\pi000 & w4418 ) | ( \pi106 & w4418 ) ;
  assign w4420 = ( \pi001 & \pi002 ) | ( \pi001 & ~w4419 ) | ( \pi002 & ~w4419 ) ;
  assign w4421 = ( w4416 & w4418 ) | ( w4416 & ~w4420 ) | ( w4418 & ~w4420 ) ;
  assign w4422 = ( \pi105 & ~\pi107 ) | ( \pi105 & w4066 ) | ( ~\pi107 & w4066 ) ;
  assign w4423 = ( ~\pi106 & \pi107 ) | ( ~\pi106 & w4422 ) | ( \pi107 & w4422 ) ;
  assign w4424 = \pi108 ^ w4422 ;
  assign w4425 = w4423 ^ w4424 ;
  assign w4426 = \pi002 ^ w4421 ;
  assign w4427 = \pi000 & ~w4421 ;
  assign w4428 = w4425 & w4427 ;
  assign w4429 = \pi001 ^ w4428 ;
  assign w4430 = ( \pi001 & w4426 ) | ( \pi001 & ~w4429 ) | ( w4426 & ~w4429 ) ;
  assign w4431 = w4258 ^ w4413 ;
  assign w4432 = w4430 ^ w4431 ;
  assign w4433 = ( w4258 & w4413 ) | ( w4258 & w4430 ) | ( w4413 & w4430 ) ;
  assign w4434 = ( w4275 & w4398 ) | ( w4275 & w4399 ) | ( w4398 & w4399 ) ;
  assign w4435 = ( w4276 & w4284 ) | ( w4276 & w4396 ) | ( w4284 & w4396 ) ;
  assign w4436 = ~\pi096 & w601 ;
  assign w4437 = \pi095 & w683 ;
  assign w4438 = ( w601 & ~w4436 ) | ( w601 & w4437 ) | ( ~w4436 & w4437 ) ;
  assign w4439 = ~\pi097 & w603 ;
  assign w4440 = w2673 | w4438 ;
  assign w4441 = ( w604 & w4438 ) | ( w604 & w4440 ) | ( w4438 & w4440 ) ;
  assign w4442 = ( w603 & ~w4439 ) | ( w603 & w4441 ) | ( ~w4439 & w4441 ) ;
  assign w4443 = \pi014 ^ w4442 ;
  assign w4444 = ( w4285 & w4293 ) | ( w4285 & w4394 ) | ( w4293 & w4394 ) ;
  assign w4445 = ( w4294 & w4384 ) | ( w4294 & w4392 ) | ( w4384 & w4392 ) ;
  assign w4446 = ~\pi090 & w1044 ;
  assign w4447 = \pi089 & w1138 ;
  assign w4448 = ( w1044 & ~w4446 ) | ( w1044 & w4447 ) | ( ~w4446 & w4447 ) ;
  assign w4449 = ~\pi091 & w1046 ;
  assign w4450 = w1908 | w4448 ;
  assign w4451 = ( w1047 & w4448 ) | ( w1047 & w4450 ) | ( w4448 & w4450 ) ;
  assign w4452 = ( w1046 & ~w4449 ) | ( w1046 & w4451 ) | ( ~w4449 & w4451 ) ;
  assign w4453 = \pi020 ^ w4452 ;
  assign w4454 = ~\pi084 & w1629 ;
  assign w4455 = \pi083 & w1722 ;
  assign w4456 = ( w1629 & ~w4454 ) | ( w1629 & w4455 ) | ( ~w4454 & w4455 ) ;
  assign w4457 = ~\pi085 & w1631 ;
  assign w4458 = w1274 | w4456 ;
  assign w4459 = ( w1632 & w4456 ) | ( w1632 & w4458 ) | ( w4456 & w4458 ) ;
  assign w4460 = ( w1631 & ~w4457 ) | ( w1631 & w4459 ) | ( ~w4457 & w4459 ) ;
  assign w4461 = \pi026 ^ w4460 ;
  assign w4462 = ( w4304 & w4312 ) | ( w4304 & w4368 ) | ( w4312 & w4368 ) ;
  assign w4463 = ( w4313 & w4321 ) | ( w4313 & w4366 ) | ( w4321 & w4366 ) ;
  assign w4464 = ( w4170 & w4356 ) | ( w4170 & w4364 ) | ( w4356 & w4364 ) ;
  assign w4465 = ~\pi075 & w2712 ;
  assign w4466 = \pi074 & w2872 ;
  assign w4467 = ( w2712 & ~w4465 ) | ( w2712 & w4466 ) | ( ~w4465 & w4466 ) ;
  assign w4468 = ~\pi076 & w2714 ;
  assign w4469 = w538 | w4467 ;
  assign w4470 = ( w2715 & w4467 ) | ( w2715 & w4469 ) | ( w4467 & w4469 ) ;
  assign w4471 = ( w2714 & ~w4468 ) | ( w2714 & w4470 ) | ( ~w4468 & w4470 ) ;
  assign w4472 = \pi035 ^ w4471 ;
  assign w4473 = ( w4322 & w4330 ) | ( w4322 & w4354 ) | ( w4330 & w4354 ) ;
  assign w4474 = ~\pi069 & w3635 ;
  assign w4475 = \pi068 & w3817 ;
  assign w4476 = ( w3635 & ~w4474 ) | ( w3635 & w4475 ) | ( ~w4474 & w4475 ) ;
  assign w4477 = ~\pi070 & w3637 ;
  assign w4478 = w271 | w4476 ;
  assign w4479 = ( w3638 & w4476 ) | ( w3638 & w4478 ) | ( w4476 & w4478 ) ;
  assign w4480 = ( w3637 & ~w4477 ) | ( w3637 & w4479 ) | ( ~w4477 & w4479 ) ;
  assign w4481 = \pi041 ^ w4480 ;
  assign w4482 = ~\pi066 & w4141 ;
  assign w4483 = \pi065 & w4334 ;
  assign w4484 = ( w4141 & ~w4482 ) | ( w4141 & w4483 ) | ( ~w4482 & w4483 ) ;
  assign w4485 = ~\pi067 & w4143 ;
  assign w4486 = w160 | w4484 ;
  assign w4487 = ( w4144 & w4484 ) | ( w4144 & w4486 ) | ( w4484 & w4486 ) ;
  assign w4488 = ( w4143 & ~w4485 ) | ( w4143 & w4487 ) | ( ~w4485 & w4487 ) ;
  assign w4489 = \pi044 ^ w4488 ;
  assign w4490 = w4343 ^ w4489 ;
  assign w4491 = \pi044 ^ \pi045 ;
  assign w4492 = \pi064 & w4491 ;
  assign w4493 = w4490 ^ w4492 ;
  assign w4494 = ( w4331 & w4344 ) | ( w4331 & w4352 ) | ( w4344 & w4352 ) ;
  assign w4495 = w4493 ^ w4494 ;
  assign w4496 = w4481 ^ w4495 ;
  assign w4497 = ~\pi072 & w3178 ;
  assign w4498 = \pi071 & w3340 ;
  assign w4499 = ( w3178 & ~w4497 ) | ( w3178 & w4498 ) | ( ~w4497 & w4498 ) ;
  assign w4500 = ~\pi073 & w3180 ;
  assign w4501 = w404 | w4499 ;
  assign w4502 = ( w3181 & w4499 ) | ( w3181 & w4501 ) | ( w4499 & w4501 ) ;
  assign w4503 = ( w3180 & ~w4500 ) | ( w3180 & w4502 ) | ( ~w4500 & w4502 ) ;
  assign w4504 = \pi038 ^ w4503 ;
  assign w4505 = w4473 ^ w4496 ;
  assign w4506 = w4504 ^ w4505 ;
  assign w4507 = w4464 ^ w4506 ;
  assign w4508 = w4472 ^ w4507 ;
  assign w4509 = ~\pi078 & w2310 ;
  assign w4510 = \pi077 & w2443 ;
  assign w4511 = ( w2310 & ~w4509 ) | ( w2310 & w4510 ) | ( ~w4509 & w4510 ) ;
  assign w4512 = ~\pi079 & w2312 ;
  assign w4513 = w730 | w4511 ;
  assign w4514 = ( w2313 & w4511 ) | ( w2313 & w4513 ) | ( w4511 & w4513 ) ;
  assign w4515 = ( w2312 & ~w4512 ) | ( w2312 & w4514 ) | ( ~w4512 & w4514 ) ;
  assign w4516 = \pi032 ^ w4515 ;
  assign w4517 = w4463 ^ w4508 ;
  assign w4518 = w4516 ^ w4517 ;
  assign w4519 = ~\pi081 & w1944 ;
  assign w4520 = \pi080 & w2072 ;
  assign w4521 = ( w1944 & ~w4519 ) | ( w1944 & w4520 ) | ( ~w4519 & w4520 ) ;
  assign w4522 = ~\pi082 & w1946 ;
  assign w4523 = w1008 | w4521 ;
  assign w4524 = ( w1947 & w4521 ) | ( w1947 & w4523 ) | ( w4521 & w4523 ) ;
  assign w4525 = ( w1946 & ~w4522 ) | ( w1946 & w4524 ) | ( ~w4522 & w4524 ) ;
  assign w4526 = \pi029 ^ w4525 ;
  assign w4527 = w4462 ^ w4518 ;
  assign w4528 = w4526 ^ w4527 ;
  assign w4529 = ( w4303 & w4370 ) | ( w4303 & w4371 ) | ( w4370 & w4371 ) ;
  assign w4530 = w4528 ^ w4529 ;
  assign w4531 = w4461 ^ w4530 ;
  assign w4532 = ~\pi087 & w1313 ;
  assign w4533 = \pi086 & w1417 ;
  assign w4534 = ( w1313 & ~w4532 ) | ( w1313 & w4533 ) | ( ~w4532 & w4533 ) ;
  assign w4535 = ~\pi088 & w1315 ;
  assign w4536 = w1574 | w4534 ;
  assign w4537 = ( w1316 & w4534 ) | ( w1316 & w4536 ) | ( w4534 & w4536 ) ;
  assign w4538 = ( w1315 & ~w4535 ) | ( w1315 & w4537 ) | ( ~w4535 & w4537 ) ;
  assign w4539 = \pi023 ^ w4538 ;
  assign w4540 = w4382 ^ w4531 ;
  assign w4541 = w4539 ^ w4540 ;
  assign w4542 = w4445 ^ w4541 ;
  assign w4543 = w4453 ^ w4542 ;
  assign w4544 = ~\pi093 & w837 ;
  assign w4545 = \pi092 & w902 ;
  assign w4546 = ( w837 & ~w4544 ) | ( w837 & w4545 ) | ( ~w4544 & w4545 ) ;
  assign w4547 = ~\pi094 & w839 ;
  assign w4548 = w2274 | w4546 ;
  assign w4549 = ( w840 & w4546 ) | ( w840 & w4548 ) | ( w4546 & w4548 ) ;
  assign w4550 = ( w839 & ~w4547 ) | ( w839 & w4549 ) | ( ~w4547 & w4549 ) ;
  assign w4551 = \pi017 ^ w4550 ;
  assign w4552 = w4444 ^ w4543 ;
  assign w4553 = w4551 ^ w4552 ;
  assign w4554 = w4435 ^ w4553 ;
  assign w4555 = w4443 ^ w4554 ;
  assign w4556 = ~\pi099 & w432 ;
  assign w4557 = \pi098 & w486 ;
  assign w4558 = ( w432 & ~w4556 ) | ( w432 & w4557 ) | ( ~w4556 & w4557 ) ;
  assign w4559 = ~\pi100 & w434 ;
  assign w4560 = w3104 | w4558 ;
  assign w4561 = ( w435 & w4558 ) | ( w435 & w4560 ) | ( w4558 & w4560 ) ;
  assign w4562 = ( w434 & ~w4559 ) | ( w434 & w4561 ) | ( ~w4559 & w4561 ) ;
  assign w4563 = \pi011 ^ w4562 ;
  assign w4564 = w4434 ^ w4555 ;
  assign w4565 = w4563 ^ w4564 ;
  assign w4566 = ~\pi102 & w305 ;
  assign w4567 = \pi101 & w328 ;
  assign w4568 = ( w305 & ~w4566 ) | ( w305 & w4567 ) | ( ~w4566 & w4567 ) ;
  assign w4569 = ~\pi103 & w307 ;
  assign w4570 = w3437 | w4568 ;
  assign w4571 = ( w308 & w4568 ) | ( w308 & w4570 ) | ( w4568 & w4570 ) ;
  assign w4572 = ( w307 & ~w4569 ) | ( w307 & w4571 ) | ( ~w4569 & w4571 ) ;
  assign w4573 = \pi008 ^ w4572 ;
  assign w4574 = ( w4242 & w4401 ) | ( w4242 & w4409 ) | ( w4401 & w4409 ) ;
  assign w4575 = w4565 ^ w4574 ;
  assign w4576 = w4573 ^ w4575 ;
  assign w4577 = ~\pi105 & w189 ;
  assign w4578 = \pi104 & w229 ;
  assign w4579 = ( w189 & ~w4577 ) | ( w189 & w4578 ) | ( ~w4577 & w4578 ) ;
  assign w4580 = ~\pi106 & w191 ;
  assign w4581 = w4068 | w4579 ;
  assign w4582 = ( w192 & w4579 ) | ( w192 & w4581 ) | ( w4579 & w4581 ) ;
  assign w4583 = ( w191 & ~w4580 ) | ( w191 & w4582 ) | ( ~w4580 & w4582 ) ;
  assign w4584 = \pi005 ^ w4583 ;
  assign w4585 = ( w4259 & w4267 ) | ( w4259 & w4411 ) | ( w4267 & w4411 ) ;
  assign w4586 = w4576 ^ w4585 ;
  assign w4587 = w4584 ^ w4586 ;
  assign w4588 = ( ~\pi002 & \pi108 ) | ( ~\pi002 & \pi109 ) | ( \pi108 & \pi109 ) ;
  assign w4589 = \pi000 ^ w4588 ;
  assign w4590 = ( \pi002 & \pi109 ) | ( \pi002 & ~w4589 ) | ( \pi109 & ~w4589 ) ;
  assign w4591 = ( \pi002 & \pi108 ) | ( \pi002 & w4589 ) | ( \pi108 & w4589 ) ;
  assign w4592 = \pi001 & w4591 ;
  assign w4593 = ( ~\pi000 & \pi107 ) | ( ~\pi000 & w4592 ) | ( \pi107 & w4592 ) ;
  assign w4594 = ( \pi001 & \pi002 ) | ( \pi001 & ~w4593 ) | ( \pi002 & ~w4593 ) ;
  assign w4595 = ( w4590 & w4592 ) | ( w4590 & ~w4594 ) | ( w4592 & ~w4594 ) ;
  assign w4596 = ( \pi106 & \pi107 ) | ( \pi106 & \pi108 ) | ( \pi107 & \pi108 ) ;
  assign w4597 = ( \pi107 & w4085 ) | ( \pi107 & w4596 ) | ( w4085 & w4596 ) ;
  assign w4598 = \pi108 ^ \pi109 ;
  assign w4599 = w4597 ^ w4598 ;
  assign w4600 = \pi002 ^ w4595 ;
  assign w4601 = \pi000 & ~w4595 ;
  assign w4602 = w4599 & w4601 ;
  assign w4603 = \pi001 ^ w4602 ;
  assign w4604 = ( \pi001 & w4600 ) | ( \pi001 & ~w4603 ) | ( w4600 & ~w4603 ) ;
  assign w4605 = w4433 ^ w4587 ;
  assign w4606 = w4604 ^ w4605 ;
  assign w4607 = ( w4565 & w4573 ) | ( w4565 & w4574 ) | ( w4573 & w4574 ) ;
  assign w4608 = ~\pi097 & w601 ;
  assign w4609 = \pi096 & w683 ;
  assign w4610 = ( w601 & ~w4608 ) | ( w601 & w4609 ) | ( ~w4608 & w4609 ) ;
  assign w4611 = ~\pi098 & w603 ;
  assign w4612 = w2824 | w4610 ;
  assign w4613 = ( w604 & w4610 ) | ( w604 & w4612 ) | ( w4610 & w4612 ) ;
  assign w4614 = ( w603 & ~w4611 ) | ( w603 & w4613 ) | ( ~w4611 & w4613 ) ;
  assign w4615 = \pi014 ^ w4614 ;
  assign w4616 = ( w4444 & w4543 ) | ( w4444 & w4551 ) | ( w4543 & w4551 ) ;
  assign w4617 = ( w4445 & w4453 ) | ( w4445 & w4541 ) | ( w4453 & w4541 ) ;
  assign w4618 = ~\pi091 & w1044 ;
  assign w4619 = \pi090 & w1138 ;
  assign w4620 = ( w1044 & ~w4618 ) | ( w1044 & w4619 ) | ( ~w4618 & w4619 ) ;
  assign w4621 = ~\pi092 & w1046 ;
  assign w4622 = w2033 | w4620 ;
  assign w4623 = ( w1047 & w4620 ) | ( w1047 & w4622 ) | ( w4620 & w4622 ) ;
  assign w4624 = ( w1046 & ~w4621 ) | ( w1046 & w4623 ) | ( ~w4621 & w4623 ) ;
  assign w4625 = \pi020 ^ w4624 ;
  assign w4626 = ~\pi079 & w2310 ;
  assign w4627 = \pi078 & w2443 ;
  assign w4628 = ( w2310 & ~w4626 ) | ( w2310 & w4627 ) | ( ~w4626 & w4627 ) ;
  assign w4629 = ~\pi080 & w2312 ;
  assign w4630 = w794 | w4628 ;
  assign w4631 = ( w2313 & w4628 ) | ( w2313 & w4630 ) | ( w4628 & w4630 ) ;
  assign w4632 = ( w2312 & ~w4629 ) | ( w2312 & w4631 ) | ( ~w4629 & w4631 ) ;
  assign w4633 = \pi032 ^ w4632 ;
  assign w4634 = ( w4464 & w4472 ) | ( w4464 & w4506 ) | ( w4472 & w4506 ) ;
  assign w4635 = ( w4473 & w4496 ) | ( w4473 & w4504 ) | ( w4496 & w4504 ) ;
  assign w4636 = ~\pi070 & w3635 ;
  assign w4637 = \pi069 & w3817 ;
  assign w4638 = ( w3635 & ~w4636 ) | ( w3635 & w4637 ) | ( ~w4636 & w4637 ) ;
  assign w4639 = ~\pi071 & w3637 ;
  assign w4640 = w290 | w4638 ;
  assign w4641 = ( w3638 & w4638 ) | ( w3638 & w4640 ) | ( w4638 & w4640 ) ;
  assign w4642 = ( w3637 & ~w4639 ) | ( w3637 & w4641 ) | ( ~w4639 & w4641 ) ;
  assign w4643 = \pi041 ^ w4642 ;
  assign w4644 = ( w4343 & w4489 ) | ( w4343 & w4492 ) | ( w4489 & w4492 ) ;
  assign w4645 = ~\pi067 & w4141 ;
  assign w4646 = \pi066 & w4334 ;
  assign w4647 = ( w4141 & ~w4645 ) | ( w4141 & w4646 ) | ( ~w4645 & w4646 ) ;
  assign w4648 = ~\pi068 & w4143 ;
  assign w4649 = w182 | w4647 ;
  assign w4650 = ( w4144 & w4647 ) | ( w4144 & w4649 ) | ( w4647 & w4649 ) ;
  assign w4651 = ( w4143 & ~w4648 ) | ( w4143 & w4650 ) | ( ~w4648 & w4650 ) ;
  assign w4652 = \pi044 ^ w4651 ;
  assign w4653 = ( \pi044 & \pi045 ) | ( \pi044 & \pi046 ) | ( \pi045 & \pi046 ) ;
  assign w4654 = \pi046 ^ w4653 ;
  assign w4655 = \pi046 ^ \pi047 ;
  assign w4656 = w4491 & ~w4655 ;
  assign w4657 = w4491 & w4655 ;
  assign w4658 = ( \pi044 & \pi045 ) | ( \pi044 & ~\pi047 ) | ( \pi045 & ~\pi047 ) ;
  assign w4659 = \pi047 & ~\pi064 ;
  assign w4660 = ~\pi065 & w4659 ;
  assign w4661 = ( \pi044 & \pi045 ) | ( \pi044 & ~w4660 ) | ( \pi045 & ~w4660 ) ;
  assign w4662 = ( \pi046 & \pi047 ) | ( \pi046 & ~w4661 ) | ( \pi047 & ~w4661 ) ;
  assign w4663 = ( \pi046 & ~w4659 ) | ( \pi046 & w4661 ) | ( ~w4659 & w4661 ) ;
  assign w4664 = ( w4658 & w4662 ) | ( w4658 & ~w4663 ) | ( w4662 & ~w4663 ) ;
  assign w4665 = ( \pi044 & \pi045 ) | ( \pi044 & \pi065 ) | ( \pi045 & \pi065 ) ;
  assign w4666 = \pi044 & \pi045 ;
  assign w4667 = \pi064 ^ w4666 ;
  assign w4668 = ( \pi046 & w4666 ) | ( \pi046 & w4667 ) | ( w4666 & w4667 ) ;
  assign w4669 = w4665 ^ w4668 ;
  assign w4670 = w4644 ^ w4652 ;
  assign w4671 = w4669 ^ w4670 ;
  assign w4672 = ( w4481 & w4493 ) | ( w4481 & w4494 ) | ( w4493 & w4494 ) ;
  assign w4673 = w4671 ^ w4672 ;
  assign w4674 = w4643 ^ w4673 ;
  assign w4675 = ~\pi073 & w3178 ;
  assign w4676 = \pi072 & w3340 ;
  assign w4677 = ( w3178 & ~w4675 ) | ( w3178 & w4676 ) | ( ~w4675 & w4676 ) ;
  assign w4678 = ~\pi074 & w3180 ;
  assign w4679 = w465 | w4677 ;
  assign w4680 = ( w3181 & w4677 ) | ( w3181 & w4679 ) | ( w4677 & w4679 ) ;
  assign w4681 = ( w3180 & ~w4678 ) | ( w3180 & w4680 ) | ( ~w4678 & w4680 ) ;
  assign w4682 = \pi038 ^ w4681 ;
  assign w4683 = ( w4635 & w4674 ) | ( w4635 & w4682 ) | ( w4674 & w4682 ) ;
  assign w4684 = w4635 ^ w4674 ;
  assign w4685 = w4682 ^ w4684 ;
  assign w4686 = ~\pi076 & w2712 ;
  assign w4687 = \pi075 & w2872 ;
  assign w4688 = ( w2712 & ~w4686 ) | ( w2712 & w4687 ) | ( ~w4686 & w4687 ) ;
  assign w4689 = ~\pi077 & w2714 ;
  assign w4690 = w644 | w4688 ;
  assign w4691 = ( w2715 & w4688 ) | ( w2715 & w4690 ) | ( w4688 & w4690 ) ;
  assign w4692 = ( w2714 & ~w4689 ) | ( w2714 & w4691 ) | ( ~w4689 & w4691 ) ;
  assign w4693 = \pi035 ^ w4692 ;
  assign w4694 = w4634 ^ w4685 ;
  assign w4695 = w4693 ^ w4694 ;
  assign w4696 = ( w4463 & w4508 ) | ( w4463 & w4516 ) | ( w4508 & w4516 ) ;
  assign w4697 = w4695 ^ w4696 ;
  assign w4698 = w4633 ^ w4697 ;
  assign w4699 = ~\pi082 & w1944 ;
  assign w4700 = \pi081 & w2072 ;
  assign w4701 = ( w1944 & ~w4699 ) | ( w1944 & w4700 ) | ( ~w4699 & w4700 ) ;
  assign w4702 = ~\pi083 & w1946 ;
  assign w4703 = w1099 | w4701 ;
  assign w4704 = ( w1947 & w4701 ) | ( w1947 & w4703 ) | ( w4701 & w4703 ) ;
  assign w4705 = ( w1946 & ~w4702 ) | ( w1946 & w4704 ) | ( ~w4702 & w4704 ) ;
  assign w4706 = \pi029 ^ w4705 ;
  assign w4707 = ( w4462 & w4518 ) | ( w4462 & w4526 ) | ( w4518 & w4526 ) ;
  assign w4708 = w4698 ^ w4707 ;
  assign w4709 = w4706 ^ w4708 ;
  assign w4710 = ~\pi085 & w1629 ;
  assign w4711 = \pi084 & w1722 ;
  assign w4712 = ( w1629 & ~w4710 ) | ( w1629 & w4711 ) | ( ~w4710 & w4711 ) ;
  assign w4713 = ~\pi086 & w1631 ;
  assign w4714 = w1379 | w4712 ;
  assign w4715 = ( w1632 & w4712 ) | ( w1632 & w4714 ) | ( w4712 & w4714 ) ;
  assign w4716 = ( w1631 & ~w4713 ) | ( w1631 & w4715 ) | ( ~w4713 & w4715 ) ;
  assign w4717 = \pi026 ^ w4716 ;
  assign w4718 = ( w4461 & w4528 ) | ( w4461 & w4529 ) | ( w4528 & w4529 ) ;
  assign w4719 = w4709 ^ w4718 ;
  assign w4720 = w4717 ^ w4719 ;
  assign w4721 = ~\pi088 & w1313 ;
  assign w4722 = \pi087 & w1417 ;
  assign w4723 = ( w1313 & ~w4721 ) | ( w1313 & w4722 ) | ( ~w4721 & w4722 ) ;
  assign w4724 = ~\pi089 & w1315 ;
  assign w4725 = w1595 | w4723 ;
  assign w4726 = ( w1316 & w4723 ) | ( w1316 & w4725 ) | ( w4723 & w4725 ) ;
  assign w4727 = ( w1315 & ~w4724 ) | ( w1315 & w4726 ) | ( ~w4724 & w4726 ) ;
  assign w4728 = \pi023 ^ w4727 ;
  assign w4729 = ( w4382 & w4531 ) | ( w4382 & w4539 ) | ( w4531 & w4539 ) ;
  assign w4730 = w4720 ^ w4729 ;
  assign w4731 = w4728 ^ w4730 ;
  assign w4732 = w4617 ^ w4731 ;
  assign w4733 = w4625 ^ w4732 ;
  assign w4734 = ~\pi094 & w837 ;
  assign w4735 = \pi093 & w902 ;
  assign w4736 = ( w837 & ~w4734 ) | ( w837 & w4735 ) | ( ~w4734 & w4735 ) ;
  assign w4737 = ~\pi095 & w839 ;
  assign w4738 = w2409 | w4736 ;
  assign w4739 = ( w840 & w4736 ) | ( w840 & w4738 ) | ( w4736 & w4738 ) ;
  assign w4740 = ( w839 & ~w4737 ) | ( w839 & w4739 ) | ( ~w4737 & w4739 ) ;
  assign w4741 = \pi017 ^ w4740 ;
  assign w4742 = w4616 ^ w4733 ;
  assign w4743 = w4741 ^ w4742 ;
  assign w4744 = ( w4435 & w4443 ) | ( w4435 & w4553 ) | ( w4443 & w4553 ) ;
  assign w4745 = w4743 ^ w4744 ;
  assign w4746 = w4615 ^ w4745 ;
  assign w4747 = ~\pi100 & w432 ;
  assign w4748 = \pi099 & w486 ;
  assign w4749 = ( w432 & ~w4747 ) | ( w432 & w4748 ) | ( ~w4747 & w4748 ) ;
  assign w4750 = ~\pi101 & w434 ;
  assign w4751 = w3264 | w4749 ;
  assign w4752 = ( w435 & w4749 ) | ( w435 & w4751 ) | ( w4749 & w4751 ) ;
  assign w4753 = ( w434 & ~w4750 ) | ( w434 & w4752 ) | ( ~w4750 & w4752 ) ;
  assign w4754 = \pi011 ^ w4753 ;
  assign w4755 = ( w4434 & w4555 ) | ( w4434 & w4563 ) | ( w4555 & w4563 ) ;
  assign w4756 = w4746 ^ w4755 ;
  assign w4757 = w4754 ^ w4756 ;
  assign w4758 = ~\pi103 & w305 ;
  assign w4759 = \pi102 & w328 ;
  assign w4760 = ( w305 & ~w4758 ) | ( w305 & w4759 ) | ( ~w4758 & w4759 ) ;
  assign w4761 = ~\pi104 & w307 ;
  assign w4762 = w3740 | w4760 ;
  assign w4763 = ( w308 & w4760 ) | ( w308 & w4762 ) | ( w4760 & w4762 ) ;
  assign w4764 = ( w307 & ~w4761 ) | ( w307 & w4763 ) | ( ~w4761 & w4763 ) ;
  assign w4765 = \pi008 ^ w4764 ;
  assign w4766 = ( w4607 & w4757 ) | ( w4607 & w4765 ) | ( w4757 & w4765 ) ;
  assign w4767 = w4607 ^ w4757 ;
  assign w4768 = w4765 ^ w4767 ;
  assign w4769 = ~\pi106 & w189 ;
  assign w4770 = \pi105 & w229 ;
  assign w4771 = ( w189 & ~w4769 ) | ( w189 & w4770 ) | ( ~w4769 & w4770 ) ;
  assign w4772 = ~\pi107 & w191 ;
  assign w4773 = w4087 | w4771 ;
  assign w4774 = ( w192 & w4771 ) | ( w192 & w4773 ) | ( w4771 & w4773 ) ;
  assign w4775 = ( w191 & ~w4772 ) | ( w191 & w4774 ) | ( ~w4772 & w4774 ) ;
  assign w4776 = \pi005 ^ w4775 ;
  assign w4777 = ( w4576 & w4584 ) | ( w4576 & w4585 ) | ( w4584 & w4585 ) ;
  assign w4778 = w4768 ^ w4777 ;
  assign w4779 = w4776 ^ w4778 ;
  assign w4780 = ( ~\pi002 & \pi109 ) | ( ~\pi002 & \pi110 ) | ( \pi109 & \pi110 ) ;
  assign w4781 = \pi000 ^ w4780 ;
  assign w4782 = ( \pi002 & \pi110 ) | ( \pi002 & ~w4781 ) | ( \pi110 & ~w4781 ) ;
  assign w4783 = ( \pi002 & \pi109 ) | ( \pi002 & w4781 ) | ( \pi109 & w4781 ) ;
  assign w4784 = \pi001 & w4783 ;
  assign w4785 = ( ~\pi000 & \pi108 ) | ( ~\pi000 & w4784 ) | ( \pi108 & w4784 ) ;
  assign w4786 = ( \pi001 & \pi002 ) | ( \pi001 & ~w4785 ) | ( \pi002 & ~w4785 ) ;
  assign w4787 = ( w4782 & w4784 ) | ( w4782 & ~w4786 ) | ( w4784 & ~w4786 ) ;
  assign w4788 = ( \pi106 & \pi107 ) | ( \pi106 & ~\pi109 ) | ( \pi107 & ~\pi109 ) ;
  assign w4789 = ( \pi107 & w4085 ) | ( \pi107 & w4788 ) | ( w4085 & w4788 ) ;
  assign w4790 = ( \pi108 & \pi109 ) | ( \pi108 & w4789 ) | ( \pi109 & w4789 ) ;
  assign w4791 = \pi109 ^ w4790 ;
  assign w4792 = \pi110 ^ w4791 ;
  assign w4793 = \pi002 ^ w4787 ;
  assign w4794 = \pi000 & ~w4787 ;
  assign w4795 = w4792 & w4794 ;
  assign w4796 = \pi001 ^ w4795 ;
  assign w4797 = ( \pi001 & w4793 ) | ( \pi001 & ~w4796 ) | ( w4793 & ~w4796 ) ;
  assign w4798 = ( w4433 & w4587 ) | ( w4433 & w4604 ) | ( w4587 & w4604 ) ;
  assign w4799 = w4779 ^ w4798 ;
  assign w4800 = w4797 ^ w4799 ;
  assign w4801 = ( ~\pi002 & \pi110 ) | ( ~\pi002 & \pi111 ) | ( \pi110 & \pi111 ) ;
  assign w4802 = \pi000 ^ w4801 ;
  assign w4803 = ( \pi002 & \pi111 ) | ( \pi002 & ~w4802 ) | ( \pi111 & ~w4802 ) ;
  assign w4804 = ( \pi002 & \pi110 ) | ( \pi002 & w4802 ) | ( \pi110 & w4802 ) ;
  assign w4805 = \pi001 & w4804 ;
  assign w4806 = ( ~\pi000 & \pi109 ) | ( ~\pi000 & w4805 ) | ( \pi109 & w4805 ) ;
  assign w4807 = ( \pi001 & \pi002 ) | ( \pi001 & ~w4806 ) | ( \pi002 & ~w4806 ) ;
  assign w4808 = ( w4803 & w4805 ) | ( w4803 & ~w4807 ) | ( w4805 & ~w4807 ) ;
  assign w4809 = ( \pi109 & \pi110 ) | ( \pi109 & w4790 ) | ( \pi110 & w4790 ) ;
  assign w4810 = \pi110 ^ w4809 ;
  assign w4811 = \pi111 ^ w4810 ;
  assign w4812 = \pi002 ^ w4808 ;
  assign w4813 = \pi000 & ~w4808 ;
  assign w4814 = w4811 & w4813 ;
  assign w4815 = \pi001 ^ w4814 ;
  assign w4816 = ( \pi001 & w4812 ) | ( \pi001 & ~w4815 ) | ( w4812 & ~w4815 ) ;
  assign w4817 = ( w4768 & w4776 ) | ( w4768 & w4777 ) | ( w4776 & w4777 ) ;
  assign w4818 = ~\pi098 & w601 ;
  assign w4819 = \pi097 & w683 ;
  assign w4820 = ( w601 & ~w4818 ) | ( w601 & w4819 ) | ( ~w4818 & w4819 ) ;
  assign w4821 = ~\pi099 & w603 ;
  assign w4822 = w2966 | w4820 ;
  assign w4823 = ( w604 & w4820 ) | ( w604 & w4822 ) | ( w4820 & w4822 ) ;
  assign w4824 = ( w603 & ~w4821 ) | ( w603 & w4823 ) | ( ~w4821 & w4823 ) ;
  assign w4825 = \pi014 ^ w4824 ;
  assign w4826 = ( w4616 & w4733 ) | ( w4616 & w4741 ) | ( w4733 & w4741 ) ;
  assign w4827 = ~\pi095 & w837 ;
  assign w4828 = \pi094 & w902 ;
  assign w4829 = ( w837 & ~w4827 ) | ( w837 & w4828 ) | ( ~w4827 & w4828 ) ;
  assign w4830 = ~\pi096 & w839 ;
  assign w4831 = w2546 | w4829 ;
  assign w4832 = ( w840 & w4829 ) | ( w840 & w4831 ) | ( w4829 & w4831 ) ;
  assign w4833 = ( w839 & ~w4830 ) | ( w839 & w4832 ) | ( ~w4830 & w4832 ) ;
  assign w4834 = \pi017 ^ w4833 ;
  assign w4835 = ( w4617 & w4625 ) | ( w4617 & w4731 ) | ( w4625 & w4731 ) ;
  assign w4836 = ~\pi092 & w1044 ;
  assign w4837 = \pi091 & w1138 ;
  assign w4838 = ( w1044 & ~w4836 ) | ( w1044 & w4837 ) | ( ~w4836 & w4837 ) ;
  assign w4839 = ~\pi093 & w1046 ;
  assign w4840 = w2155 | w4838 ;
  assign w4841 = ( w1047 & w4838 ) | ( w1047 & w4840 ) | ( w4838 & w4840 ) ;
  assign w4842 = ( w1046 & ~w4839 ) | ( w1046 & w4841 ) | ( ~w4839 & w4841 ) ;
  assign w4843 = \pi020 ^ w4842 ;
  assign w4844 = ( w4720 & w4728 ) | ( w4720 & w4729 ) | ( w4728 & w4729 ) ;
  assign w4845 = ( w4709 & w4717 ) | ( w4709 & w4718 ) | ( w4717 & w4718 ) ;
  assign w4846 = ( w4633 & w4695 ) | ( w4633 & w4696 ) | ( w4695 & w4696 ) ;
  assign w4847 = ~\pi080 & w2310 ;
  assign w4848 = \pi079 & w2443 ;
  assign w4849 = ( w2310 & ~w4847 ) | ( w2310 & w4848 ) | ( ~w4847 & w4848 ) ;
  assign w4850 = ~\pi081 & w2312 ;
  assign w4851 = w874 | w4849 ;
  assign w4852 = ( w2313 & w4849 ) | ( w2313 & w4851 ) | ( w4849 & w4851 ) ;
  assign w4853 = ( w2312 & ~w4850 ) | ( w2312 & w4852 ) | ( ~w4850 & w4852 ) ;
  assign w4854 = \pi032 ^ w4853 ;
  assign w4855 = ( w4634 & w4685 ) | ( w4634 & w4693 ) | ( w4685 & w4693 ) ;
  assign w4856 = ~\pi077 & w2712 ;
  assign w4857 = \pi076 & w2872 ;
  assign w4858 = ( w2712 & ~w4856 ) | ( w2712 & w4857 ) | ( ~w4856 & w4857 ) ;
  assign w4859 = ~\pi078 & w2714 ;
  assign w4860 = w665 | w4858 ;
  assign w4861 = ( w2715 & w4858 ) | ( w2715 & w4860 ) | ( w4858 & w4860 ) ;
  assign w4862 = ( w2714 & ~w4859 ) | ( w2714 & w4861 ) | ( ~w4859 & w4861 ) ;
  assign w4863 = \pi035 ^ w4862 ;
  assign w4864 = ( w4643 & w4671 ) | ( w4643 & w4672 ) | ( w4671 & w4672 ) ;
  assign w4865 = ~\pi071 & w3635 ;
  assign w4866 = \pi070 & w3817 ;
  assign w4867 = ( w3635 & ~w4865 ) | ( w3635 & w4866 ) | ( ~w4865 & w4866 ) ;
  assign w4868 = ~\pi072 & w3637 ;
  assign w4869 = w361 | w4867 ;
  assign w4870 = ( w3638 & w4867 ) | ( w3638 & w4869 ) | ( w4867 & w4869 ) ;
  assign w4871 = ( w3637 & ~w4868 ) | ( w3637 & w4870 ) | ( ~w4868 & w4870 ) ;
  assign w4872 = \pi041 ^ w4871 ;
  assign w4873 = ( w4644 & w4652 ) | ( w4644 & w4669 ) | ( w4652 & w4669 ) ;
  assign w4874 = ( \pi045 & ~\pi046 ) | ( \pi045 & \pi047 ) | ( ~\pi046 & \pi047 ) ;
  assign w4875 = ( \pi044 & \pi045 ) | ( \pi044 & w4874 ) | ( \pi045 & w4874 ) ;
  assign w4876 = w4874 ^ w4875 ;
  assign w4877 = \pi064 & w4876 ;
  assign w4878 = ( \pi066 & w4656 ) | ( \pi066 & w4877 ) | ( w4656 & w4877 ) ;
  assign w4879 = \pi065 | w4878 ;
  assign w4880 = ( w4654 & w4878 ) | ( w4654 & w4879 ) | ( w4878 & w4879 ) ;
  assign w4881 = w4877 | w4880 ;
  assign w4882 = ~w134 & w4657 ;
  assign w4883 = ( w4657 & w4881 ) | ( w4657 & ~w4882 ) | ( w4881 & ~w4882 ) ;
  assign w4884 = \pi047 ^ w4883 ;
  assign w4885 = w4664 & w4884 ;
  assign w4886 = w4664 ^ w4884 ;
  assign w4887 = ~\pi068 & w4141 ;
  assign w4888 = \pi067 & w4334 ;
  assign w4889 = ( w4141 & ~w4887 ) | ( w4141 & w4888 ) | ( ~w4887 & w4888 ) ;
  assign w4890 = ~\pi069 & w4143 ;
  assign w4891 = w221 | w4889 ;
  assign w4892 = ( w4144 & w4889 ) | ( w4144 & w4891 ) | ( w4889 & w4891 ) ;
  assign w4893 = ( w4143 & ~w4890 ) | ( w4143 & w4892 ) | ( ~w4890 & w4892 ) ;
  assign w4894 = \pi044 ^ w4893 ;
  assign w4895 = w4873 ^ w4886 ;
  assign w4896 = w4894 ^ w4895 ;
  assign w4897 = w4864 ^ w4896 ;
  assign w4898 = w4872 ^ w4897 ;
  assign w4899 = ~\pi074 & w3178 ;
  assign w4900 = \pi073 & w3340 ;
  assign w4901 = ( w3178 & ~w4899 ) | ( w3178 & w4900 ) | ( ~w4899 & w4900 ) ;
  assign w4902 = ~\pi075 & w3180 ;
  assign w4903 = w519 | w4901 ;
  assign w4904 = ( w3181 & w4901 ) | ( w3181 & w4903 ) | ( w4901 & w4903 ) ;
  assign w4905 = ( w3180 & ~w4902 ) | ( w3180 & w4904 ) | ( ~w4902 & w4904 ) ;
  assign w4906 = \pi038 ^ w4905 ;
  assign w4907 = w4683 ^ w4898 ;
  assign w4908 = w4906 ^ w4907 ;
  assign w4909 = w4855 ^ w4908 ;
  assign w4910 = w4863 ^ w4909 ;
  assign w4911 = w4846 ^ w4910 ;
  assign w4912 = w4854 ^ w4911 ;
  assign w4913 = ~\pi083 & w1944 ;
  assign w4914 = \pi082 & w2072 ;
  assign w4915 = ( w1944 & ~w4913 ) | ( w1944 & w4914 ) | ( ~w4913 & w4914 ) ;
  assign w4916 = ~\pi084 & w1946 ;
  assign w4917 = w1188 | w4915 ;
  assign w4918 = ( w1947 & w4915 ) | ( w1947 & w4917 ) | ( w4915 & w4917 ) ;
  assign w4919 = ( w1946 & ~w4916 ) | ( w1946 & w4918 ) | ( ~w4916 & w4918 ) ;
  assign w4920 = \pi029 ^ w4919 ;
  assign w4921 = ( w4698 & w4706 ) | ( w4698 & w4707 ) | ( w4706 & w4707 ) ;
  assign w4922 = w4912 ^ w4921 ;
  assign w4923 = w4920 ^ w4922 ;
  assign w4924 = ~\pi086 & w1629 ;
  assign w4925 = \pi085 & w1722 ;
  assign w4926 = ( w1629 & ~w4924 ) | ( w1629 & w4925 ) | ( ~w4924 & w4925 ) ;
  assign w4927 = ~\pi087 & w1631 ;
  assign w4928 = w1477 | w4926 ;
  assign w4929 = ( w1632 & w4926 ) | ( w1632 & w4928 ) | ( w4926 & w4928 ) ;
  assign w4930 = ( w1631 & ~w4927 ) | ( w1631 & w4929 ) | ( ~w4927 & w4929 ) ;
  assign w4931 = \pi026 ^ w4930 ;
  assign w4932 = ( w4845 & w4923 ) | ( w4845 & w4931 ) | ( w4923 & w4931 ) ;
  assign w4933 = w4845 ^ w4923 ;
  assign w4934 = w4931 ^ w4933 ;
  assign w4935 = ~\pi089 & w1313 ;
  assign w4936 = \pi088 & w1417 ;
  assign w4937 = ( w1313 & ~w4935 ) | ( w1313 & w4936 ) | ( ~w4935 & w4936 ) ;
  assign w4938 = ~\pi090 & w1315 ;
  assign w4939 = w1801 | w4937 ;
  assign w4940 = ( w1316 & w4937 ) | ( w1316 & w4939 ) | ( w4937 & w4939 ) ;
  assign w4941 = ( w1315 & ~w4938 ) | ( w1315 & w4940 ) | ( ~w4938 & w4940 ) ;
  assign w4942 = \pi023 ^ w4941 ;
  assign w4943 = w4844 ^ w4934 ;
  assign w4944 = w4942 ^ w4943 ;
  assign w4945 = w4835 ^ w4944 ;
  assign w4946 = w4843 ^ w4945 ;
  assign w4947 = w4826 ^ w4946 ;
  assign w4948 = w4834 ^ w4947 ;
  assign w4949 = ( w4615 & w4743 ) | ( w4615 & w4744 ) | ( w4743 & w4744 ) ;
  assign w4950 = w4948 ^ w4949 ;
  assign w4951 = w4825 ^ w4950 ;
  assign w4952 = ~\pi101 & w432 ;
  assign w4953 = \pi100 & w486 ;
  assign w4954 = ( w432 & ~w4952 ) | ( w432 & w4953 ) | ( ~w4952 & w4953 ) ;
  assign w4955 = ~\pi102 & w434 ;
  assign w4956 = w3284 | w4954 ;
  assign w4957 = ( w435 & w4954 ) | ( w435 & w4956 ) | ( w4954 & w4956 ) ;
  assign w4958 = ( w434 & ~w4955 ) | ( w434 & w4957 ) | ( ~w4955 & w4957 ) ;
  assign w4959 = \pi011 ^ w4958 ;
  assign w4960 = ( w4746 & w4754 ) | ( w4746 & w4755 ) | ( w4754 & w4755 ) ;
  assign w4961 = w4951 ^ w4960 ;
  assign w4962 = w4959 ^ w4961 ;
  assign w4963 = ~\pi104 & w305 ;
  assign w4964 = \pi103 & w328 ;
  assign w4965 = ( w305 & ~w4963 ) | ( w305 & w4964 ) | ( ~w4963 & w4964 ) ;
  assign w4966 = ~\pi105 & w307 ;
  assign w4967 = w3905 | w4965 ;
  assign w4968 = ( w308 & w4965 ) | ( w308 & w4967 ) | ( w4965 & w4967 ) ;
  assign w4969 = ( w307 & ~w4966 ) | ( w307 & w4968 ) | ( ~w4966 & w4968 ) ;
  assign w4970 = \pi008 ^ w4969 ;
  assign w4971 = ( w4766 & w4962 ) | ( w4766 & w4970 ) | ( w4962 & w4970 ) ;
  assign w4972 = w4766 ^ w4962 ;
  assign w4973 = w4970 ^ w4972 ;
  assign w4974 = ~\pi107 & w189 ;
  assign w4975 = \pi106 & w229 ;
  assign w4976 = ( w189 & ~w4974 ) | ( w189 & w4975 ) | ( ~w4974 & w4975 ) ;
  assign w4977 = ~\pi108 & w191 ;
  assign w4978 = w4425 | w4976 ;
  assign w4979 = ( w192 & w4976 ) | ( w192 & w4978 ) | ( w4976 & w4978 ) ;
  assign w4980 = ( w191 & ~w4977 ) | ( w191 & w4979 ) | ( ~w4977 & w4979 ) ;
  assign w4981 = \pi005 ^ w4980 ;
  assign w4982 = w4817 ^ w4973 ;
  assign w4983 = w4981 ^ w4982 ;
  assign w4984 = ( w4779 & w4797 ) | ( w4779 & w4798 ) | ( w4797 & w4798 ) ;
  assign w4985 = w4983 ^ w4984 ;
  assign w4986 = w4816 ^ w4985 ;
  assign w4987 = ( w4816 & w4983 ) | ( w4816 & w4984 ) | ( w4983 & w4984 ) ;
  assign w4988 = ( ~\pi002 & \pi111 ) | ( ~\pi002 & \pi112 ) | ( \pi111 & \pi112 ) ;
  assign w4989 = \pi000 ^ w4988 ;
  assign w4990 = ( \pi002 & \pi112 ) | ( \pi002 & ~w4989 ) | ( \pi112 & ~w4989 ) ;
  assign w4991 = ( \pi002 & \pi111 ) | ( \pi002 & w4989 ) | ( \pi111 & w4989 ) ;
  assign w4992 = \pi001 & w4991 ;
  assign w4993 = ( ~\pi000 & \pi110 ) | ( ~\pi000 & w4992 ) | ( \pi110 & w4992 ) ;
  assign w4994 = ( \pi001 & \pi002 ) | ( \pi001 & ~w4993 ) | ( \pi002 & ~w4993 ) ;
  assign w4995 = ( w4990 & w4992 ) | ( w4990 & ~w4994 ) | ( w4992 & ~w4994 ) ;
  assign w4996 = ( \pi109 & ~\pi111 ) | ( \pi109 & w4790 ) | ( ~\pi111 & w4790 ) ;
  assign w4997 = ( ~\pi110 & \pi111 ) | ( ~\pi110 & w4996 ) | ( \pi111 & w4996 ) ;
  assign w4998 = \pi112 ^ w4996 ;
  assign w4999 = w4997 ^ w4998 ;
  assign w5000 = \pi002 ^ w4995 ;
  assign w5001 = \pi000 & ~w4995 ;
  assign w5002 = w4999 & w5001 ;
  assign w5003 = \pi001 ^ w5002 ;
  assign w5004 = ( \pi001 & w5000 ) | ( \pi001 & ~w5003 ) | ( w5000 & ~w5003 ) ;
  assign w5005 = ( w4817 & w4973 ) | ( w4817 & w4981 ) | ( w4973 & w4981 ) ;
  assign w5006 = ( w4825 & w4948 ) | ( w4825 & w4949 ) | ( w4948 & w4949 ) ;
  assign w5007 = ( w4826 & w4834 ) | ( w4826 & w4946 ) | ( w4834 & w4946 ) ;
  assign w5008 = ~\pi096 & w837 ;
  assign w5009 = \pi095 & w902 ;
  assign w5010 = ( w837 & ~w5008 ) | ( w837 & w5009 ) | ( ~w5008 & w5009 ) ;
  assign w5011 = ~\pi097 & w839 ;
  assign w5012 = w2673 | w5010 ;
  assign w5013 = ( w840 & w5010 ) | ( w840 & w5012 ) | ( w5010 & w5012 ) ;
  assign w5014 = ( w839 & ~w5011 ) | ( w839 & w5013 ) | ( ~w5011 & w5013 ) ;
  assign w5015 = \pi017 ^ w5014 ;
  assign w5016 = ( w4835 & w4843 ) | ( w4835 & w4944 ) | ( w4843 & w4944 ) ;
  assign w5017 = ( w4844 & w4934 ) | ( w4844 & w4942 ) | ( w4934 & w4942 ) ;
  assign w5018 = ~\pi090 & w1313 ;
  assign w5019 = \pi089 & w1417 ;
  assign w5020 = ( w1313 & ~w5018 ) | ( w1313 & w5019 ) | ( ~w5018 & w5019 ) ;
  assign w5021 = ~\pi091 & w1315 ;
  assign w5022 = w1908 | w5020 ;
  assign w5023 = ( w1316 & w5020 ) | ( w1316 & w5022 ) | ( w5020 & w5022 ) ;
  assign w5024 = ( w1315 & ~w5021 ) | ( w1315 & w5023 ) | ( ~w5021 & w5023 ) ;
  assign w5025 = \pi023 ^ w5024 ;
  assign w5026 = ( w4855 & w4863 ) | ( w4855 & w4908 ) | ( w4863 & w4908 ) ;
  assign w5027 = ~\pi078 & w2712 ;
  assign w5028 = \pi077 & w2872 ;
  assign w5029 = ( w2712 & ~w5027 ) | ( w2712 & w5028 ) | ( ~w5027 & w5028 ) ;
  assign w5030 = ~\pi079 & w2714 ;
  assign w5031 = w730 | w5029 ;
  assign w5032 = ( w2715 & w5029 ) | ( w2715 & w5031 ) | ( w5029 & w5031 ) ;
  assign w5033 = ( w2714 & ~w5030 ) | ( w2714 & w5032 ) | ( ~w5030 & w5032 ) ;
  assign w5034 = \pi035 ^ w5033 ;
  assign w5035 = ( w4683 & w4898 ) | ( w4683 & w4906 ) | ( w4898 & w4906 ) ;
  assign w5036 = ~\pi075 & w3178 ;
  assign w5037 = \pi074 & w3340 ;
  assign w5038 = ( w3178 & ~w5036 ) | ( w3178 & w5037 ) | ( ~w5036 & w5037 ) ;
  assign w5039 = ~\pi076 & w3180 ;
  assign w5040 = w538 | w5038 ;
  assign w5041 = ( w3181 & w5038 ) | ( w3181 & w5040 ) | ( w5038 & w5040 ) ;
  assign w5042 = ( w3180 & ~w5039 ) | ( w3180 & w5041 ) | ( ~w5039 & w5041 ) ;
  assign w5043 = \pi038 ^ w5042 ;
  assign w5044 = ( w4864 & w4872 ) | ( w4864 & w4896 ) | ( w4872 & w4896 ) ;
  assign w5045 = ~\pi069 & w4141 ;
  assign w5046 = \pi068 & w4334 ;
  assign w5047 = ( w4141 & ~w5045 ) | ( w4141 & w5046 ) | ( ~w5045 & w5046 ) ;
  assign w5048 = ~\pi070 & w4143 ;
  assign w5049 = w271 | w5047 ;
  assign w5050 = ( w4144 & w5047 ) | ( w4144 & w5049 ) | ( w5047 & w5049 ) ;
  assign w5051 = ( w4143 & ~w5048 ) | ( w4143 & w5050 ) | ( ~w5048 & w5050 ) ;
  assign w5052 = \pi044 ^ w5051 ;
  assign w5053 = ~\pi066 & w4654 ;
  assign w5054 = \pi065 & w4876 ;
  assign w5055 = ( w4654 & ~w5053 ) | ( w4654 & w5054 ) | ( ~w5053 & w5054 ) ;
  assign w5056 = ~\pi067 & w4656 ;
  assign w5057 = w160 | w5055 ;
  assign w5058 = ( w4657 & w5055 ) | ( w4657 & w5057 ) | ( w5055 & w5057 ) ;
  assign w5059 = ( w4656 & ~w5056 ) | ( w4656 & w5058 ) | ( ~w5056 & w5058 ) ;
  assign w5060 = \pi047 ^ w5059 ;
  assign w5061 = w4885 ^ w5060 ;
  assign w5062 = \pi047 ^ \pi048 ;
  assign w5063 = \pi064 & w5062 ;
  assign w5064 = w5061 ^ w5063 ;
  assign w5065 = ( w4873 & w4886 ) | ( w4873 & w4894 ) | ( w4886 & w4894 ) ;
  assign w5066 = w5064 ^ w5065 ;
  assign w5067 = w5052 ^ w5066 ;
  assign w5068 = ~\pi072 & w3635 ;
  assign w5069 = \pi071 & w3817 ;
  assign w5070 = ( w3635 & ~w5068 ) | ( w3635 & w5069 ) | ( ~w5068 & w5069 ) ;
  assign w5071 = ~\pi073 & w3637 ;
  assign w5072 = w404 | w5070 ;
  assign w5073 = ( w3638 & w5070 ) | ( w3638 & w5072 ) | ( w5070 & w5072 ) ;
  assign w5074 = ( w3637 & ~w5071 ) | ( w3637 & w5073 ) | ( ~w5071 & w5073 ) ;
  assign w5075 = \pi041 ^ w5074 ;
  assign w5076 = w5044 ^ w5067 ;
  assign w5077 = w5075 ^ w5076 ;
  assign w5078 = w5035 ^ w5077 ;
  assign w5079 = w5043 ^ w5078 ;
  assign w5080 = w5026 ^ w5079 ;
  assign w5081 = w5034 ^ w5080 ;
  assign w5082 = ~\pi081 & w2310 ;
  assign w5083 = \pi080 & w2443 ;
  assign w5084 = ( w2310 & ~w5082 ) | ( w2310 & w5083 ) | ( ~w5082 & w5083 ) ;
  assign w5085 = ~\pi082 & w2312 ;
  assign w5086 = w1008 | w5084 ;
  assign w5087 = ( w2313 & w5084 ) | ( w2313 & w5086 ) | ( w5084 & w5086 ) ;
  assign w5088 = ( w2312 & ~w5085 ) | ( w2312 & w5087 ) | ( ~w5085 & w5087 ) ;
  assign w5089 = \pi032 ^ w5088 ;
  assign w5090 = ( w4846 & w4854 ) | ( w4846 & w4910 ) | ( w4854 & w4910 ) ;
  assign w5091 = w5081 ^ w5090 ;
  assign w5092 = w5089 ^ w5091 ;
  assign w5093 = ~\pi084 & w1944 ;
  assign w5094 = \pi083 & w2072 ;
  assign w5095 = ( w1944 & ~w5093 ) | ( w1944 & w5094 ) | ( ~w5093 & w5094 ) ;
  assign w5096 = ~\pi085 & w1946 ;
  assign w5097 = w1274 | w5095 ;
  assign w5098 = ( w1947 & w5095 ) | ( w1947 & w5097 ) | ( w5095 & w5097 ) ;
  assign w5099 = ( w1946 & ~w5096 ) | ( w1946 & w5098 ) | ( ~w5096 & w5098 ) ;
  assign w5100 = \pi029 ^ w5099 ;
  assign w5101 = ( w4912 & w4920 ) | ( w4912 & w4921 ) | ( w4920 & w4921 ) ;
  assign w5102 = w5092 ^ w5101 ;
  assign w5103 = w5100 ^ w5102 ;
  assign w5104 = ~\pi087 & w1629 ;
  assign w5105 = \pi086 & w1722 ;
  assign w5106 = ( w1629 & ~w5104 ) | ( w1629 & w5105 ) | ( ~w5104 & w5105 ) ;
  assign w5107 = ~\pi088 & w1631 ;
  assign w5108 = w1574 | w5106 ;
  assign w5109 = ( w1632 & w5106 ) | ( w1632 & w5108 ) | ( w5106 & w5108 ) ;
  assign w5110 = ( w1631 & ~w5107 ) | ( w1631 & w5109 ) | ( ~w5107 & w5109 ) ;
  assign w5111 = \pi026 ^ w5110 ;
  assign w5112 = w4932 ^ w5103 ;
  assign w5113 = w5111 ^ w5112 ;
  assign w5114 = w5017 ^ w5113 ;
  assign w5115 = w5025 ^ w5114 ;
  assign w5116 = ~\pi093 & w1044 ;
  assign w5117 = \pi092 & w1138 ;
  assign w5118 = ( w1044 & ~w5116 ) | ( w1044 & w5117 ) | ( ~w5116 & w5117 ) ;
  assign w5119 = ~\pi094 & w1046 ;
  assign w5120 = w2274 | w5118 ;
  assign w5121 = ( w1047 & w5118 ) | ( w1047 & w5120 ) | ( w5118 & w5120 ) ;
  assign w5122 = ( w1046 & ~w5119 ) | ( w1046 & w5121 ) | ( ~w5119 & w5121 ) ;
  assign w5123 = \pi020 ^ w5122 ;
  assign w5124 = w5016 ^ w5115 ;
  assign w5125 = w5123 ^ w5124 ;
  assign w5126 = w5007 ^ w5125 ;
  assign w5127 = w5015 ^ w5126 ;
  assign w5128 = ~\pi099 & w601 ;
  assign w5129 = \pi098 & w683 ;
  assign w5130 = ( w601 & ~w5128 ) | ( w601 & w5129 ) | ( ~w5128 & w5129 ) ;
  assign w5131 = ~\pi100 & w603 ;
  assign w5132 = w3104 | w5130 ;
  assign w5133 = ( w604 & w5130 ) | ( w604 & w5132 ) | ( w5130 & w5132 ) ;
  assign w5134 = ( w603 & ~w5131 ) | ( w603 & w5133 ) | ( ~w5131 & w5133 ) ;
  assign w5135 = \pi014 ^ w5134 ;
  assign w5136 = w5006 ^ w5127 ;
  assign w5137 = w5135 ^ w5136 ;
  assign w5138 = ~\pi102 & w432 ;
  assign w5139 = \pi101 & w486 ;
  assign w5140 = ( w432 & ~w5138 ) | ( w432 & w5139 ) | ( ~w5138 & w5139 ) ;
  assign w5141 = ~\pi103 & w434 ;
  assign w5142 = w3437 | w5140 ;
  assign w5143 = ( w435 & w5140 ) | ( w435 & w5142 ) | ( w5140 & w5142 ) ;
  assign w5144 = ( w434 & ~w5141 ) | ( w434 & w5143 ) | ( ~w5141 & w5143 ) ;
  assign w5145 = \pi011 ^ w5144 ;
  assign w5146 = ( w4951 & w4959 ) | ( w4951 & w4960 ) | ( w4959 & w4960 ) ;
  assign w5147 = w5137 ^ w5146 ;
  assign w5148 = w5145 ^ w5147 ;
  assign w5149 = ~\pi105 & w305 ;
  assign w5150 = \pi104 & w328 ;
  assign w5151 = ( w305 & ~w5149 ) | ( w305 & w5150 ) | ( ~w5149 & w5150 ) ;
  assign w5152 = ~\pi106 & w307 ;
  assign w5153 = w4068 | w5151 ;
  assign w5154 = ( w308 & w5151 ) | ( w308 & w5153 ) | ( w5151 & w5153 ) ;
  assign w5155 = ( w307 & ~w5152 ) | ( w307 & w5154 ) | ( ~w5152 & w5154 ) ;
  assign w5156 = \pi008 ^ w5155 ;
  assign w5157 = w4971 ^ w5148 ;
  assign w5158 = w5156 ^ w5157 ;
  assign w5159 = ~\pi108 & w189 ;
  assign w5160 = \pi107 & w229 ;
  assign w5161 = ( w189 & ~w5159 ) | ( w189 & w5160 ) | ( ~w5159 & w5160 ) ;
  assign w5162 = ~\pi109 & w191 ;
  assign w5163 = w4599 | w5161 ;
  assign w5164 = ( w192 & w5161 ) | ( w192 & w5163 ) | ( w5161 & w5163 ) ;
  assign w5165 = ( w191 & ~w5162 ) | ( w191 & w5164 ) | ( ~w5162 & w5164 ) ;
  assign w5166 = \pi005 ^ w5165 ;
  assign w5167 = w5005 ^ w5158 ;
  assign w5168 = w5166 ^ w5167 ;
  assign w5169 = w4987 ^ w5168 ;
  assign w5170 = w5004 ^ w5169 ;
  assign w5171 = ( w4987 & w5004 ) | ( w4987 & w5168 ) | ( w5004 & w5168 ) ;
  assign w5172 = ( w5017 & w5025 ) | ( w5017 & w5113 ) | ( w5025 & w5113 ) ;
  assign w5173 = ~\pi091 & w1313 ;
  assign w5174 = \pi090 & w1417 ;
  assign w5175 = ( w1313 & ~w5173 ) | ( w1313 & w5174 ) | ( ~w5173 & w5174 ) ;
  assign w5176 = ~\pi092 & w1315 ;
  assign w5177 = w2033 | w5175 ;
  assign w5178 = ( w1316 & w5175 ) | ( w1316 & w5177 ) | ( w5175 & w5177 ) ;
  assign w5179 = ( w1315 & ~w5176 ) | ( w1315 & w5178 ) | ( ~w5176 & w5178 ) ;
  assign w5180 = \pi023 ^ w5179 ;
  assign w5181 = ~\pi079 & w2712 ;
  assign w5182 = \pi078 & w2872 ;
  assign w5183 = ( w2712 & ~w5181 ) | ( w2712 & w5182 ) | ( ~w5181 & w5182 ) ;
  assign w5184 = ~\pi080 & w2714 ;
  assign w5185 = w794 | w5183 ;
  assign w5186 = ( w2715 & w5183 ) | ( w2715 & w5185 ) | ( w5183 & w5185 ) ;
  assign w5187 = ( w2714 & ~w5184 ) | ( w2714 & w5186 ) | ( ~w5184 & w5186 ) ;
  assign w5188 = \pi035 ^ w5187 ;
  assign w5189 = ( w5035 & w5043 ) | ( w5035 & w5077 ) | ( w5043 & w5077 ) ;
  assign w5190 = ( w5044 & w5067 ) | ( w5044 & w5075 ) | ( w5067 & w5075 ) ;
  assign w5191 = ~\pi070 & w4141 ;
  assign w5192 = \pi069 & w4334 ;
  assign w5193 = ( w4141 & ~w5191 ) | ( w4141 & w5192 ) | ( ~w5191 & w5192 ) ;
  assign w5194 = ~\pi071 & w4143 ;
  assign w5195 = w290 | w5193 ;
  assign w5196 = ( w4144 & w5193 ) | ( w4144 & w5195 ) | ( w5193 & w5195 ) ;
  assign w5197 = ( w4143 & ~w5194 ) | ( w4143 & w5196 ) | ( ~w5194 & w5196 ) ;
  assign w5198 = \pi044 ^ w5197 ;
  assign w5199 = ( w4885 & w5060 ) | ( w4885 & w5063 ) | ( w5060 & w5063 ) ;
  assign w5200 = ~\pi067 & w4654 ;
  assign w5201 = \pi066 & w4876 ;
  assign w5202 = ( w4654 & ~w5200 ) | ( w4654 & w5201 ) | ( ~w5200 & w5201 ) ;
  assign w5203 = ~\pi068 & w4656 ;
  assign w5204 = w182 | w5202 ;
  assign w5205 = ( w4657 & w5202 ) | ( w4657 & w5204 ) | ( w5202 & w5204 ) ;
  assign w5206 = ( w4656 & ~w5203 ) | ( w4656 & w5205 ) | ( ~w5203 & w5205 ) ;
  assign w5207 = \pi047 ^ w5206 ;
  assign w5208 = ( \pi047 & \pi048 ) | ( \pi047 & \pi049 ) | ( \pi048 & \pi049 ) ;
  assign w5209 = \pi049 ^ w5208 ;
  assign w5210 = \pi049 ^ \pi050 ;
  assign w5211 = w5062 & ~w5210 ;
  assign w5212 = w5062 & w5210 ;
  assign w5213 = ( \pi047 & \pi048 ) | ( \pi047 & ~\pi050 ) | ( \pi048 & ~\pi050 ) ;
  assign w5214 = \pi050 & ~\pi064 ;
  assign w5215 = ~\pi065 & w5214 ;
  assign w5216 = ( \pi047 & \pi048 ) | ( \pi047 & ~w5215 ) | ( \pi048 & ~w5215 ) ;
  assign w5217 = ( \pi049 & \pi050 ) | ( \pi049 & ~w5216 ) | ( \pi050 & ~w5216 ) ;
  assign w5218 = ( \pi049 & ~w5214 ) | ( \pi049 & w5216 ) | ( ~w5214 & w5216 ) ;
  assign w5219 = ( w5213 & w5217 ) | ( w5213 & ~w5218 ) | ( w5217 & ~w5218 ) ;
  assign w5220 = ( \pi047 & \pi048 ) | ( \pi047 & \pi065 ) | ( \pi048 & \pi065 ) ;
  assign w5221 = \pi047 & \pi048 ;
  assign w5222 = \pi064 ^ w5221 ;
  assign w5223 = ( \pi049 & w5221 ) | ( \pi049 & w5222 ) | ( w5221 & w5222 ) ;
  assign w5224 = w5220 ^ w5223 ;
  assign w5225 = w5199 ^ w5207 ;
  assign w5226 = w5224 ^ w5225 ;
  assign w5227 = ( w5052 & w5064 ) | ( w5052 & w5065 ) | ( w5064 & w5065 ) ;
  assign w5228 = w5226 ^ w5227 ;
  assign w5229 = w5198 ^ w5228 ;
  assign w5230 = ~\pi073 & w3635 ;
  assign w5231 = \pi072 & w3817 ;
  assign w5232 = ( w3635 & ~w5230 ) | ( w3635 & w5231 ) | ( ~w5230 & w5231 ) ;
  assign w5233 = ~\pi074 & w3637 ;
  assign w5234 = w465 | w5232 ;
  assign w5235 = ( w3638 & w5232 ) | ( w3638 & w5234 ) | ( w5232 & w5234 ) ;
  assign w5236 = ( w3637 & ~w5233 ) | ( w3637 & w5235 ) | ( ~w5233 & w5235 ) ;
  assign w5237 = \pi041 ^ w5236 ;
  assign w5238 = ( w5190 & w5229 ) | ( w5190 & w5237 ) | ( w5229 & w5237 ) ;
  assign w5239 = w5190 ^ w5229 ;
  assign w5240 = w5237 ^ w5239 ;
  assign w5241 = ~\pi076 & w3178 ;
  assign w5242 = \pi075 & w3340 ;
  assign w5243 = ( w3178 & ~w5241 ) | ( w3178 & w5242 ) | ( ~w5241 & w5242 ) ;
  assign w5244 = ~\pi077 & w3180 ;
  assign w5245 = w644 | w5243 ;
  assign w5246 = ( w3181 & w5243 ) | ( w3181 & w5245 ) | ( w5243 & w5245 ) ;
  assign w5247 = ( w3180 & ~w5244 ) | ( w3180 & w5246 ) | ( ~w5244 & w5246 ) ;
  assign w5248 = \pi038 ^ w5247 ;
  assign w5249 = w5189 ^ w5240 ;
  assign w5250 = w5248 ^ w5249 ;
  assign w5251 = ( w5026 & w5034 ) | ( w5026 & w5079 ) | ( w5034 & w5079 ) ;
  assign w5252 = w5250 ^ w5251 ;
  assign w5253 = w5188 ^ w5252 ;
  assign w5254 = ~\pi082 & w2310 ;
  assign w5255 = \pi081 & w2443 ;
  assign w5256 = ( w2310 & ~w5254 ) | ( w2310 & w5255 ) | ( ~w5254 & w5255 ) ;
  assign w5257 = ~\pi083 & w2312 ;
  assign w5258 = w1099 | w5256 ;
  assign w5259 = ( w2313 & w5256 ) | ( w2313 & w5258 ) | ( w5256 & w5258 ) ;
  assign w5260 = ( w2312 & ~w5257 ) | ( w2312 & w5259 ) | ( ~w5257 & w5259 ) ;
  assign w5261 = \pi032 ^ w5260 ;
  assign w5262 = ( w5081 & w5089 ) | ( w5081 & w5090 ) | ( w5089 & w5090 ) ;
  assign w5263 = w5253 ^ w5262 ;
  assign w5264 = w5261 ^ w5263 ;
  assign w5265 = ~\pi085 & w1944 ;
  assign w5266 = \pi084 & w2072 ;
  assign w5267 = ( w1944 & ~w5265 ) | ( w1944 & w5266 ) | ( ~w5265 & w5266 ) ;
  assign w5268 = ~\pi086 & w1946 ;
  assign w5269 = w1379 | w5267 ;
  assign w5270 = ( w1947 & w5267 ) | ( w1947 & w5269 ) | ( w5267 & w5269 ) ;
  assign w5271 = ( w1946 & ~w5268 ) | ( w1946 & w5270 ) | ( ~w5268 & w5270 ) ;
  assign w5272 = \pi029 ^ w5271 ;
  assign w5273 = ( w5092 & w5100 ) | ( w5092 & w5101 ) | ( w5100 & w5101 ) ;
  assign w5274 = w5264 ^ w5273 ;
  assign w5275 = w5272 ^ w5274 ;
  assign w5276 = ~\pi088 & w1629 ;
  assign w5277 = \pi087 & w1722 ;
  assign w5278 = ( w1629 & ~w5276 ) | ( w1629 & w5277 ) | ( ~w5276 & w5277 ) ;
  assign w5279 = ~\pi089 & w1631 ;
  assign w5280 = w1595 | w5278 ;
  assign w5281 = ( w1632 & w5278 ) | ( w1632 & w5280 ) | ( w5278 & w5280 ) ;
  assign w5282 = ( w1631 & ~w5279 ) | ( w1631 & w5281 ) | ( ~w5279 & w5281 ) ;
  assign w5283 = \pi026 ^ w5282 ;
  assign w5284 = ( w4932 & w5103 ) | ( w4932 & w5111 ) | ( w5103 & w5111 ) ;
  assign w5285 = w5275 ^ w5284 ;
  assign w5286 = w5283 ^ w5285 ;
  assign w5287 = w5172 ^ w5286 ;
  assign w5288 = w5180 ^ w5287 ;
  assign w5289 = ~\pi094 & w1044 ;
  assign w5290 = \pi093 & w1138 ;
  assign w5291 = ( w1044 & ~w5289 ) | ( w1044 & w5290 ) | ( ~w5289 & w5290 ) ;
  assign w5292 = ~\pi095 & w1046 ;
  assign w5293 = w2409 | w5291 ;
  assign w5294 = ( w1047 & w5291 ) | ( w1047 & w5293 ) | ( w5291 & w5293 ) ;
  assign w5295 = ( w1046 & ~w5292 ) | ( w1046 & w5294 ) | ( ~w5292 & w5294 ) ;
  assign w5296 = \pi020 ^ w5295 ;
  assign w5297 = ( w5016 & w5115 ) | ( w5016 & w5123 ) | ( w5115 & w5123 ) ;
  assign w5298 = w5288 ^ w5297 ;
  assign w5299 = w5296 ^ w5298 ;
  assign w5300 = ~\pi097 & w837 ;
  assign w5301 = \pi096 & w902 ;
  assign w5302 = ( w837 & ~w5300 ) | ( w837 & w5301 ) | ( ~w5300 & w5301 ) ;
  assign w5303 = ~\pi098 & w839 ;
  assign w5304 = w2824 | w5302 ;
  assign w5305 = ( w840 & w5302 ) | ( w840 & w5304 ) | ( w5302 & w5304 ) ;
  assign w5306 = ( w839 & ~w5303 ) | ( w839 & w5305 ) | ( ~w5303 & w5305 ) ;
  assign w5307 = \pi017 ^ w5306 ;
  assign w5308 = ( w5007 & w5015 ) | ( w5007 & w5125 ) | ( w5015 & w5125 ) ;
  assign w5309 = w5299 ^ w5308 ;
  assign w5310 = w5307 ^ w5309 ;
  assign w5311 = ~\pi100 & w601 ;
  assign w5312 = \pi099 & w683 ;
  assign w5313 = ( w601 & ~w5311 ) | ( w601 & w5312 ) | ( ~w5311 & w5312 ) ;
  assign w5314 = ~\pi101 & w603 ;
  assign w5315 = w3264 | w5313 ;
  assign w5316 = ( w604 & w5313 ) | ( w604 & w5315 ) | ( w5313 & w5315 ) ;
  assign w5317 = ( w603 & ~w5314 ) | ( w603 & w5316 ) | ( ~w5314 & w5316 ) ;
  assign w5318 = \pi014 ^ w5317 ;
  assign w5319 = ( w5006 & w5127 ) | ( w5006 & w5135 ) | ( w5127 & w5135 ) ;
  assign w5320 = w5310 ^ w5319 ;
  assign w5321 = w5318 ^ w5320 ;
  assign w5322 = ~\pi103 & w432 ;
  assign w5323 = \pi102 & w486 ;
  assign w5324 = ( w432 & ~w5322 ) | ( w432 & w5323 ) | ( ~w5322 & w5323 ) ;
  assign w5325 = ~\pi104 & w434 ;
  assign w5326 = w3740 | w5324 ;
  assign w5327 = ( w435 & w5324 ) | ( w435 & w5326 ) | ( w5324 & w5326 ) ;
  assign w5328 = ( w434 & ~w5325 ) | ( w434 & w5327 ) | ( ~w5325 & w5327 ) ;
  assign w5329 = \pi011 ^ w5328 ;
  assign w5330 = ( w5137 & w5145 ) | ( w5137 & w5146 ) | ( w5145 & w5146 ) ;
  assign w5331 = w5321 ^ w5330 ;
  assign w5332 = w5329 ^ w5331 ;
  assign w5333 = ~\pi106 & w305 ;
  assign w5334 = \pi105 & w328 ;
  assign w5335 = ( w305 & ~w5333 ) | ( w305 & w5334 ) | ( ~w5333 & w5334 ) ;
  assign w5336 = ~\pi107 & w307 ;
  assign w5337 = w4087 | w5335 ;
  assign w5338 = ( w308 & w5335 ) | ( w308 & w5337 ) | ( w5335 & w5337 ) ;
  assign w5339 = ( w307 & ~w5336 ) | ( w307 & w5338 ) | ( ~w5336 & w5338 ) ;
  assign w5340 = \pi008 ^ w5339 ;
  assign w5341 = ( w4971 & w5148 ) | ( w4971 & w5156 ) | ( w5148 & w5156 ) ;
  assign w5342 = w5332 ^ w5341 ;
  assign w5343 = w5340 ^ w5342 ;
  assign w5344 = ~\pi109 & w189 ;
  assign w5345 = \pi108 & w229 ;
  assign w5346 = ( w189 & ~w5344 ) | ( w189 & w5345 ) | ( ~w5344 & w5345 ) ;
  assign w5347 = ~\pi110 & w191 ;
  assign w5348 = w4792 | w5346 ;
  assign w5349 = ( w192 & w5346 ) | ( w192 & w5348 ) | ( w5346 & w5348 ) ;
  assign w5350 = ( w191 & ~w5347 ) | ( w191 & w5349 ) | ( ~w5347 & w5349 ) ;
  assign w5351 = \pi005 ^ w5350 ;
  assign w5352 = ( w5005 & w5158 ) | ( w5005 & w5166 ) | ( w5158 & w5166 ) ;
  assign w5353 = w5343 ^ w5352 ;
  assign w5354 = w5351 ^ w5353 ;
  assign w5355 = ( ~\pi002 & \pi112 ) | ( ~\pi002 & \pi113 ) | ( \pi112 & \pi113 ) ;
  assign w5356 = \pi000 ^ w5355 ;
  assign w5357 = ( \pi002 & \pi113 ) | ( \pi002 & ~w5356 ) | ( \pi113 & ~w5356 ) ;
  assign w5358 = ( \pi002 & \pi112 ) | ( \pi002 & w5356 ) | ( \pi112 & w5356 ) ;
  assign w5359 = \pi001 & w5358 ;
  assign w5360 = ( ~\pi000 & \pi111 ) | ( ~\pi000 & w5359 ) | ( \pi111 & w5359 ) ;
  assign w5361 = ( \pi001 & \pi002 ) | ( \pi001 & ~w5360 ) | ( \pi002 & ~w5360 ) ;
  assign w5362 = ( w5357 & w5359 ) | ( w5357 & ~w5361 ) | ( w5359 & ~w5361 ) ;
  assign w5363 = ( \pi110 & \pi111 ) | ( \pi110 & \pi112 ) | ( \pi111 & \pi112 ) ;
  assign w5364 = ( \pi111 & w4809 ) | ( \pi111 & w5363 ) | ( w4809 & w5363 ) ;
  assign w5365 = \pi112 ^ \pi113 ;
  assign w5366 = w5364 ^ w5365 ;
  assign w5367 = \pi002 ^ w5362 ;
  assign w5368 = \pi000 & ~w5362 ;
  assign w5369 = w5366 & w5368 ;
  assign w5370 = \pi001 ^ w5369 ;
  assign w5371 = ( \pi001 & w5367 ) | ( \pi001 & ~w5370 ) | ( w5367 & ~w5370 ) ;
  assign w5372 = w5171 ^ w5354 ;
  assign w5373 = w5371 ^ w5372 ;
  assign w5374 = ( w5332 & w5340 ) | ( w5332 & w5341 ) | ( w5340 & w5341 ) ;
  assign w5375 = ~\pi098 & w837 ;
  assign w5376 = \pi097 & w902 ;
  assign w5377 = ( w837 & ~w5375 ) | ( w837 & w5376 ) | ( ~w5375 & w5376 ) ;
  assign w5378 = ~\pi099 & w839 ;
  assign w5379 = w2966 | w5377 ;
  assign w5380 = ( w840 & w5377 ) | ( w840 & w5379 ) | ( w5377 & w5379 ) ;
  assign w5381 = ( w839 & ~w5378 ) | ( w839 & w5380 ) | ( ~w5378 & w5380 ) ;
  assign w5382 = \pi017 ^ w5381 ;
  assign w5383 = ( w5288 & w5296 ) | ( w5288 & w5297 ) | ( w5296 & w5297 ) ;
  assign w5384 = ~\pi095 & w1044 ;
  assign w5385 = \pi094 & w1138 ;
  assign w5386 = ( w1044 & ~w5384 ) | ( w1044 & w5385 ) | ( ~w5384 & w5385 ) ;
  assign w5387 = ~\pi096 & w1046 ;
  assign w5388 = w2546 | w5386 ;
  assign w5389 = ( w1047 & w5386 ) | ( w1047 & w5388 ) | ( w5386 & w5388 ) ;
  assign w5390 = ( w1046 & ~w5387 ) | ( w1046 & w5389 ) | ( ~w5387 & w5389 ) ;
  assign w5391 = \pi020 ^ w5390 ;
  assign w5392 = ( w5172 & w5180 ) | ( w5172 & w5286 ) | ( w5180 & w5286 ) ;
  assign w5393 = ~\pi092 & w1313 ;
  assign w5394 = \pi091 & w1417 ;
  assign w5395 = ( w1313 & ~w5393 ) | ( w1313 & w5394 ) | ( ~w5393 & w5394 ) ;
  assign w5396 = ~\pi093 & w1315 ;
  assign w5397 = w2155 | w5395 ;
  assign w5398 = ( w1316 & w5395 ) | ( w1316 & w5397 ) | ( w5395 & w5397 ) ;
  assign w5399 = ( w1315 & ~w5396 ) | ( w1315 & w5398 ) | ( ~w5396 & w5398 ) ;
  assign w5400 = \pi023 ^ w5399 ;
  assign w5401 = ( w5275 & w5283 ) | ( w5275 & w5284 ) | ( w5283 & w5284 ) ;
  assign w5402 = ( w5264 & w5272 ) | ( w5264 & w5273 ) | ( w5272 & w5273 ) ;
  assign w5403 = ( w5188 & w5250 ) | ( w5188 & w5251 ) | ( w5250 & w5251 ) ;
  assign w5404 = ~\pi080 & w2712 ;
  assign w5405 = \pi079 & w2872 ;
  assign w5406 = ( w2712 & ~w5404 ) | ( w2712 & w5405 ) | ( ~w5404 & w5405 ) ;
  assign w5407 = ~\pi081 & w2714 ;
  assign w5408 = w874 | w5406 ;
  assign w5409 = ( w2715 & w5406 ) | ( w2715 & w5408 ) | ( w5406 & w5408 ) ;
  assign w5410 = ( w2714 & ~w5407 ) | ( w2714 & w5409 ) | ( ~w5407 & w5409 ) ;
  assign w5411 = \pi035 ^ w5410 ;
  assign w5412 = ( w5189 & w5240 ) | ( w5189 & w5248 ) | ( w5240 & w5248 ) ;
  assign w5413 = ~\pi077 & w3178 ;
  assign w5414 = \pi076 & w3340 ;
  assign w5415 = ( w3178 & ~w5413 ) | ( w3178 & w5414 ) | ( ~w5413 & w5414 ) ;
  assign w5416 = ~\pi078 & w3180 ;
  assign w5417 = w665 | w5415 ;
  assign w5418 = ( w3181 & w5415 ) | ( w3181 & w5417 ) | ( w5415 & w5417 ) ;
  assign w5419 = ( w3180 & ~w5416 ) | ( w3180 & w5418 ) | ( ~w5416 & w5418 ) ;
  assign w5420 = \pi038 ^ w5419 ;
  assign w5421 = ( w5198 & w5226 ) | ( w5198 & w5227 ) | ( w5226 & w5227 ) ;
  assign w5422 = ~\pi071 & w4141 ;
  assign w5423 = \pi070 & w4334 ;
  assign w5424 = ( w4141 & ~w5422 ) | ( w4141 & w5423 ) | ( ~w5422 & w5423 ) ;
  assign w5425 = ~\pi072 & w4143 ;
  assign w5426 = w361 | w5424 ;
  assign w5427 = ( w4144 & w5424 ) | ( w4144 & w5426 ) | ( w5424 & w5426 ) ;
  assign w5428 = ( w4143 & ~w5425 ) | ( w4143 & w5427 ) | ( ~w5425 & w5427 ) ;
  assign w5429 = \pi044 ^ w5428 ;
  assign w5430 = ( w5199 & w5207 ) | ( w5199 & w5224 ) | ( w5207 & w5224 ) ;
  assign w5431 = ( \pi048 & ~\pi049 ) | ( \pi048 & \pi050 ) | ( ~\pi049 & \pi050 ) ;
  assign w5432 = ( \pi047 & \pi048 ) | ( \pi047 & w5431 ) | ( \pi048 & w5431 ) ;
  assign w5433 = w5431 ^ w5432 ;
  assign w5434 = \pi064 & w5433 ;
  assign w5435 = ( \pi066 & w5211 ) | ( \pi066 & w5434 ) | ( w5211 & w5434 ) ;
  assign w5436 = \pi065 | w5435 ;
  assign w5437 = ( w5209 & w5435 ) | ( w5209 & w5436 ) | ( w5435 & w5436 ) ;
  assign w5438 = w5434 | w5437 ;
  assign w5439 = ~w134 & w5212 ;
  assign w5440 = ( w5212 & w5438 ) | ( w5212 & ~w5439 ) | ( w5438 & ~w5439 ) ;
  assign w5441 = \pi050 ^ w5440 ;
  assign w5442 = w5219 & w5441 ;
  assign w5443 = w5219 ^ w5441 ;
  assign w5444 = ~\pi068 & w4654 ;
  assign w5445 = \pi067 & w4876 ;
  assign w5446 = ( w4654 & ~w5444 ) | ( w4654 & w5445 ) | ( ~w5444 & w5445 ) ;
  assign w5447 = ~\pi069 & w4656 ;
  assign w5448 = w221 | w5446 ;
  assign w5449 = ( w4657 & w5446 ) | ( w4657 & w5448 ) | ( w5446 & w5448 ) ;
  assign w5450 = ( w4656 & ~w5447 ) | ( w4656 & w5449 ) | ( ~w5447 & w5449 ) ;
  assign w5451 = \pi047 ^ w5450 ;
  assign w5452 = w5430 ^ w5443 ;
  assign w5453 = w5451 ^ w5452 ;
  assign w5454 = w5421 ^ w5453 ;
  assign w5455 = w5429 ^ w5454 ;
  assign w5456 = ~\pi074 & w3635 ;
  assign w5457 = \pi073 & w3817 ;
  assign w5458 = ( w3635 & ~w5456 ) | ( w3635 & w5457 ) | ( ~w5456 & w5457 ) ;
  assign w5459 = ~\pi075 & w3637 ;
  assign w5460 = w519 | w5458 ;
  assign w5461 = ( w3638 & w5458 ) | ( w3638 & w5460 ) | ( w5458 & w5460 ) ;
  assign w5462 = ( w3637 & ~w5459 ) | ( w3637 & w5461 ) | ( ~w5459 & w5461 ) ;
  assign w5463 = \pi041 ^ w5462 ;
  assign w5464 = w5238 ^ w5455 ;
  assign w5465 = w5463 ^ w5464 ;
  assign w5466 = w5412 ^ w5465 ;
  assign w5467 = w5420 ^ w5466 ;
  assign w5468 = w5403 ^ w5467 ;
  assign w5469 = w5411 ^ w5468 ;
  assign w5470 = ~\pi083 & w2310 ;
  assign w5471 = \pi082 & w2443 ;
  assign w5472 = ( w2310 & ~w5470 ) | ( w2310 & w5471 ) | ( ~w5470 & w5471 ) ;
  assign w5473 = ~\pi084 & w2312 ;
  assign w5474 = w1188 | w5472 ;
  assign w5475 = ( w2313 & w5472 ) | ( w2313 & w5474 ) | ( w5472 & w5474 ) ;
  assign w5476 = ( w2312 & ~w5473 ) | ( w2312 & w5475 ) | ( ~w5473 & w5475 ) ;
  assign w5477 = \pi032 ^ w5476 ;
  assign w5478 = ( w5253 & w5261 ) | ( w5253 & w5262 ) | ( w5261 & w5262 ) ;
  assign w5479 = w5469 ^ w5478 ;
  assign w5480 = w5477 ^ w5479 ;
  assign w5481 = ~\pi086 & w1944 ;
  assign w5482 = \pi085 & w2072 ;
  assign w5483 = ( w1944 & ~w5481 ) | ( w1944 & w5482 ) | ( ~w5481 & w5482 ) ;
  assign w5484 = ~\pi087 & w1946 ;
  assign w5485 = w1477 | w5483 ;
  assign w5486 = ( w1947 & w5483 ) | ( w1947 & w5485 ) | ( w5483 & w5485 ) ;
  assign w5487 = ( w1946 & ~w5484 ) | ( w1946 & w5486 ) | ( ~w5484 & w5486 ) ;
  assign w5488 = \pi029 ^ w5487 ;
  assign w5489 = ( w5402 & w5480 ) | ( w5402 & w5488 ) | ( w5480 & w5488 ) ;
  assign w5490 = w5402 ^ w5480 ;
  assign w5491 = w5488 ^ w5490 ;
  assign w5492 = ~\pi089 & w1629 ;
  assign w5493 = \pi088 & w1722 ;
  assign w5494 = ( w1629 & ~w5492 ) | ( w1629 & w5493 ) | ( ~w5492 & w5493 ) ;
  assign w5495 = ~\pi090 & w1631 ;
  assign w5496 = w1801 | w5494 ;
  assign w5497 = ( w1632 & w5494 ) | ( w1632 & w5496 ) | ( w5494 & w5496 ) ;
  assign w5498 = ( w1631 & ~w5495 ) | ( w1631 & w5497 ) | ( ~w5495 & w5497 ) ;
  assign w5499 = \pi026 ^ w5498 ;
  assign w5500 = w5401 ^ w5491 ;
  assign w5501 = w5499 ^ w5500 ;
  assign w5502 = w5392 ^ w5501 ;
  assign w5503 = w5400 ^ w5502 ;
  assign w5504 = w5383 ^ w5503 ;
  assign w5505 = w5391 ^ w5504 ;
  assign w5506 = ( w5299 & w5307 ) | ( w5299 & w5308 ) | ( w5307 & w5308 ) ;
  assign w5507 = w5505 ^ w5506 ;
  assign w5508 = w5382 ^ w5507 ;
  assign w5509 = ~\pi101 & w601 ;
  assign w5510 = \pi100 & w683 ;
  assign w5511 = ( w601 & ~w5509 ) | ( w601 & w5510 ) | ( ~w5509 & w5510 ) ;
  assign w5512 = ~\pi102 & w603 ;
  assign w5513 = w3284 | w5511 ;
  assign w5514 = ( w604 & w5511 ) | ( w604 & w5513 ) | ( w5511 & w5513 ) ;
  assign w5515 = ( w603 & ~w5512 ) | ( w603 & w5514 ) | ( ~w5512 & w5514 ) ;
  assign w5516 = \pi014 ^ w5515 ;
  assign w5517 = ( w5310 & w5318 ) | ( w5310 & w5319 ) | ( w5318 & w5319 ) ;
  assign w5518 = w5508 ^ w5517 ;
  assign w5519 = w5516 ^ w5518 ;
  assign w5520 = ~\pi104 & w432 ;
  assign w5521 = \pi103 & w486 ;
  assign w5522 = ( w432 & ~w5520 ) | ( w432 & w5521 ) | ( ~w5520 & w5521 ) ;
  assign w5523 = ~\pi105 & w434 ;
  assign w5524 = w3905 | w5522 ;
  assign w5525 = ( w435 & w5522 ) | ( w435 & w5524 ) | ( w5522 & w5524 ) ;
  assign w5526 = ( w434 & ~w5523 ) | ( w434 & w5525 ) | ( ~w5523 & w5525 ) ;
  assign w5527 = \pi011 ^ w5526 ;
  assign w5528 = ( w5321 & w5329 ) | ( w5321 & w5330 ) | ( w5329 & w5330 ) ;
  assign w5529 = w5519 ^ w5528 ;
  assign w5530 = w5527 ^ w5529 ;
  assign w5531 = ~\pi107 & w305 ;
  assign w5532 = \pi106 & w328 ;
  assign w5533 = ( w305 & ~w5531 ) | ( w305 & w5532 ) | ( ~w5531 & w5532 ) ;
  assign w5534 = ~\pi108 & w307 ;
  assign w5535 = w4425 | w5533 ;
  assign w5536 = ( w308 & w5533 ) | ( w308 & w5535 ) | ( w5533 & w5535 ) ;
  assign w5537 = ( w307 & ~w5534 ) | ( w307 & w5536 ) | ( ~w5534 & w5536 ) ;
  assign w5538 = \pi008 ^ w5537 ;
  assign w5539 = ( w5374 & w5530 ) | ( w5374 & w5538 ) | ( w5530 & w5538 ) ;
  assign w5540 = w5374 ^ w5530 ;
  assign w5541 = w5538 ^ w5540 ;
  assign w5542 = ~\pi110 & w189 ;
  assign w5543 = \pi109 & w229 ;
  assign w5544 = ( w189 & ~w5542 ) | ( w189 & w5543 ) | ( ~w5542 & w5543 ) ;
  assign w5545 = ~\pi111 & w191 ;
  assign w5546 = w4811 | w5544 ;
  assign w5547 = ( w192 & w5544 ) | ( w192 & w5546 ) | ( w5544 & w5546 ) ;
  assign w5548 = ( w191 & ~w5545 ) | ( w191 & w5547 ) | ( ~w5545 & w5547 ) ;
  assign w5549 = \pi005 ^ w5548 ;
  assign w5550 = ( w5343 & w5351 ) | ( w5343 & w5352 ) | ( w5351 & w5352 ) ;
  assign w5551 = w5541 ^ w5550 ;
  assign w5552 = w5549 ^ w5551 ;
  assign w5553 = ( ~\pi002 & \pi113 ) | ( ~\pi002 & \pi114 ) | ( \pi113 & \pi114 ) ;
  assign w5554 = \pi000 ^ w5553 ;
  assign w5555 = ( \pi002 & \pi114 ) | ( \pi002 & ~w5554 ) | ( \pi114 & ~w5554 ) ;
  assign w5556 = ( \pi002 & \pi113 ) | ( \pi002 & w5554 ) | ( \pi113 & w5554 ) ;
  assign w5557 = \pi001 & w5556 ;
  assign w5558 = ( ~\pi000 & \pi112 ) | ( ~\pi000 & w5557 ) | ( \pi112 & w5557 ) ;
  assign w5559 = ( \pi001 & \pi002 ) | ( \pi001 & ~w5558 ) | ( \pi002 & ~w5558 ) ;
  assign w5560 = ( w5555 & w5557 ) | ( w5555 & ~w5559 ) | ( w5557 & ~w5559 ) ;
  assign w5561 = ( \pi110 & \pi111 ) | ( \pi110 & ~\pi113 ) | ( \pi111 & ~\pi113 ) ;
  assign w5562 = ( \pi111 & w4809 ) | ( \pi111 & w5561 ) | ( w4809 & w5561 ) ;
  assign w5563 = ( \pi112 & \pi113 ) | ( \pi112 & w5562 ) | ( \pi113 & w5562 ) ;
  assign w5564 = \pi113 ^ w5563 ;
  assign w5565 = \pi114 ^ w5564 ;
  assign w5566 = \pi002 ^ w5560 ;
  assign w5567 = \pi000 & ~w5560 ;
  assign w5568 = w5565 & w5567 ;
  assign w5569 = \pi001 ^ w5568 ;
  assign w5570 = ( \pi001 & w5566 ) | ( \pi001 & ~w5569 ) | ( w5566 & ~w5569 ) ;
  assign w5571 = ( w5171 & w5354 ) | ( w5171 & w5371 ) | ( w5354 & w5371 ) ;
  assign w5572 = w5552 ^ w5571 ;
  assign w5573 = w5570 ^ w5572 ;
  assign w5574 = ( w5552 & w5570 ) | ( w5552 & w5571 ) | ( w5570 & w5571 ) ;
  assign w5575 = ( ~\pi002 & \pi114 ) | ( ~\pi002 & \pi115 ) | ( \pi114 & \pi115 ) ;
  assign w5576 = \pi000 ^ w5575 ;
  assign w5577 = ( \pi002 & \pi115 ) | ( \pi002 & ~w5576 ) | ( \pi115 & ~w5576 ) ;
  assign w5578 = ( \pi002 & \pi114 ) | ( \pi002 & w5576 ) | ( \pi114 & w5576 ) ;
  assign w5579 = \pi001 & w5578 ;
  assign w5580 = ( ~\pi000 & \pi113 ) | ( ~\pi000 & w5579 ) | ( \pi113 & w5579 ) ;
  assign w5581 = ( \pi001 & \pi002 ) | ( \pi001 & ~w5580 ) | ( \pi002 & ~w5580 ) ;
  assign w5582 = ( w5577 & w5579 ) | ( w5577 & ~w5581 ) | ( w5579 & ~w5581 ) ;
  assign w5583 = ( \pi113 & \pi114 ) | ( \pi113 & w5563 ) | ( \pi114 & w5563 ) ;
  assign w5584 = \pi114 ^ w5583 ;
  assign w5585 = \pi115 ^ w5584 ;
  assign w5586 = \pi002 ^ w5582 ;
  assign w5587 = \pi000 & ~w5582 ;
  assign w5588 = w5585 & w5587 ;
  assign w5589 = \pi001 ^ w5588 ;
  assign w5590 = ( \pi001 & w5586 ) | ( \pi001 & ~w5589 ) | ( w5586 & ~w5589 ) ;
  assign w5591 = ( w5541 & w5549 ) | ( w5541 & w5550 ) | ( w5549 & w5550 ) ;
  assign w5592 = ~\pi108 & w305 ;
  assign w5593 = \pi107 & w328 ;
  assign w5594 = ( w305 & ~w5592 ) | ( w305 & w5593 ) | ( ~w5592 & w5593 ) ;
  assign w5595 = ~\pi109 & w307 ;
  assign w5596 = w4599 | w5594 ;
  assign w5597 = ( w308 & w5594 ) | ( w308 & w5596 ) | ( w5594 & w5596 ) ;
  assign w5598 = ( w307 & ~w5595 ) | ( w307 & w5597 ) | ( ~w5595 & w5597 ) ;
  assign w5599 = \pi008 ^ w5598 ;
  assign w5600 = ( w5382 & w5505 ) | ( w5382 & w5506 ) | ( w5505 & w5506 ) ;
  assign w5601 = ( w5383 & w5391 ) | ( w5383 & w5503 ) | ( w5391 & w5503 ) ;
  assign w5602 = ~\pi096 & w1044 ;
  assign w5603 = \pi095 & w1138 ;
  assign w5604 = ( w1044 & ~w5602 ) | ( w1044 & w5603 ) | ( ~w5602 & w5603 ) ;
  assign w5605 = ~\pi097 & w1046 ;
  assign w5606 = w2673 | w5604 ;
  assign w5607 = ( w1047 & w5604 ) | ( w1047 & w5606 ) | ( w5604 & w5606 ) ;
  assign w5608 = ( w1046 & ~w5605 ) | ( w1046 & w5607 ) | ( ~w5605 & w5607 ) ;
  assign w5609 = \pi020 ^ w5608 ;
  assign w5610 = ( w5392 & w5400 ) | ( w5392 & w5501 ) | ( w5400 & w5501 ) ;
  assign w5611 = ( w5401 & w5491 ) | ( w5401 & w5499 ) | ( w5491 & w5499 ) ;
  assign w5612 = ~\pi090 & w1629 ;
  assign w5613 = \pi089 & w1722 ;
  assign w5614 = ( w1629 & ~w5612 ) | ( w1629 & w5613 ) | ( ~w5612 & w5613 ) ;
  assign w5615 = ~\pi091 & w1631 ;
  assign w5616 = w1908 | w5614 ;
  assign w5617 = ( w1632 & w5614 ) | ( w1632 & w5616 ) | ( w5614 & w5616 ) ;
  assign w5618 = ( w1631 & ~w5615 ) | ( w1631 & w5617 ) | ( ~w5615 & w5617 ) ;
  assign w5619 = \pi026 ^ w5618 ;
  assign w5620 = ( w5403 & w5411 ) | ( w5403 & w5467 ) | ( w5411 & w5467 ) ;
  assign w5621 = ~\pi081 & w2712 ;
  assign w5622 = \pi080 & w2872 ;
  assign w5623 = ( w2712 & ~w5621 ) | ( w2712 & w5622 ) | ( ~w5621 & w5622 ) ;
  assign w5624 = ~\pi082 & w2714 ;
  assign w5625 = w1008 | w5623 ;
  assign w5626 = ( w2715 & w5623 ) | ( w2715 & w5625 ) | ( w5623 & w5625 ) ;
  assign w5627 = ( w2714 & ~w5624 ) | ( w2714 & w5626 ) | ( ~w5624 & w5626 ) ;
  assign w5628 = \pi035 ^ w5627 ;
  assign w5629 = ( w5412 & w5420 ) | ( w5412 & w5465 ) | ( w5420 & w5465 ) ;
  assign w5630 = ~\pi078 & w3178 ;
  assign w5631 = \pi077 & w3340 ;
  assign w5632 = ( w3178 & ~w5630 ) | ( w3178 & w5631 ) | ( ~w5630 & w5631 ) ;
  assign w5633 = ~\pi079 & w3180 ;
  assign w5634 = w730 | w5632 ;
  assign w5635 = ( w3181 & w5632 ) | ( w3181 & w5634 ) | ( w5632 & w5634 ) ;
  assign w5636 = ( w3180 & ~w5633 ) | ( w3180 & w5635 ) | ( ~w5633 & w5635 ) ;
  assign w5637 = \pi038 ^ w5636 ;
  assign w5638 = ( w5238 & w5455 ) | ( w5238 & w5463 ) | ( w5455 & w5463 ) ;
  assign w5639 = ~\pi075 & w3635 ;
  assign w5640 = \pi074 & w3817 ;
  assign w5641 = ( w3635 & ~w5639 ) | ( w3635 & w5640 ) | ( ~w5639 & w5640 ) ;
  assign w5642 = ~\pi076 & w3637 ;
  assign w5643 = w538 | w5641 ;
  assign w5644 = ( w3638 & w5641 ) | ( w3638 & w5643 ) | ( w5641 & w5643 ) ;
  assign w5645 = ( w3637 & ~w5642 ) | ( w3637 & w5644 ) | ( ~w5642 & w5644 ) ;
  assign w5646 = \pi041 ^ w5645 ;
  assign w5647 = ( w5421 & w5429 ) | ( w5421 & w5453 ) | ( w5429 & w5453 ) ;
  assign w5648 = ~\pi069 & w4654 ;
  assign w5649 = \pi068 & w4876 ;
  assign w5650 = ( w4654 & ~w5648 ) | ( w4654 & w5649 ) | ( ~w5648 & w5649 ) ;
  assign w5651 = ~\pi070 & w4656 ;
  assign w5652 = w271 | w5650 ;
  assign w5653 = ( w4657 & w5650 ) | ( w4657 & w5652 ) | ( w5650 & w5652 ) ;
  assign w5654 = ( w4656 & ~w5651 ) | ( w4656 & w5653 ) | ( ~w5651 & w5653 ) ;
  assign w5655 = \pi047 ^ w5654 ;
  assign w5656 = ~\pi066 & w5209 ;
  assign w5657 = \pi065 & w5433 ;
  assign w5658 = ( w5209 & ~w5656 ) | ( w5209 & w5657 ) | ( ~w5656 & w5657 ) ;
  assign w5659 = ~\pi067 & w5211 ;
  assign w5660 = w160 | w5658 ;
  assign w5661 = ( w5212 & w5658 ) | ( w5212 & w5660 ) | ( w5658 & w5660 ) ;
  assign w5662 = ( w5211 & ~w5659 ) | ( w5211 & w5661 ) | ( ~w5659 & w5661 ) ;
  assign w5663 = \pi050 ^ w5662 ;
  assign w5664 = w5442 ^ w5663 ;
  assign w5665 = \pi050 ^ \pi051 ;
  assign w5666 = \pi064 & w5665 ;
  assign w5667 = w5664 ^ w5666 ;
  assign w5668 = ( w5430 & w5443 ) | ( w5430 & w5451 ) | ( w5443 & w5451 ) ;
  assign w5669 = w5667 ^ w5668 ;
  assign w5670 = w5655 ^ w5669 ;
  assign w5671 = ~\pi072 & w4141 ;
  assign w5672 = \pi071 & w4334 ;
  assign w5673 = ( w4141 & ~w5671 ) | ( w4141 & w5672 ) | ( ~w5671 & w5672 ) ;
  assign w5674 = ~\pi073 & w4143 ;
  assign w5675 = w404 | w5673 ;
  assign w5676 = ( w4144 & w5673 ) | ( w4144 & w5675 ) | ( w5673 & w5675 ) ;
  assign w5677 = ( w4143 & ~w5674 ) | ( w4143 & w5676 ) | ( ~w5674 & w5676 ) ;
  assign w5678 = \pi044 ^ w5677 ;
  assign w5679 = w5647 ^ w5670 ;
  assign w5680 = w5678 ^ w5679 ;
  assign w5681 = w5638 ^ w5680 ;
  assign w5682 = w5646 ^ w5681 ;
  assign w5683 = w5629 ^ w5682 ;
  assign w5684 = w5637 ^ w5683 ;
  assign w5685 = w5620 ^ w5684 ;
  assign w5686 = w5628 ^ w5685 ;
  assign w5687 = ~\pi084 & w2310 ;
  assign w5688 = \pi083 & w2443 ;
  assign w5689 = ( w2310 & ~w5687 ) | ( w2310 & w5688 ) | ( ~w5687 & w5688 ) ;
  assign w5690 = ~\pi085 & w2312 ;
  assign w5691 = w1274 | w5689 ;
  assign w5692 = ( w2313 & w5689 ) | ( w2313 & w5691 ) | ( w5689 & w5691 ) ;
  assign w5693 = ( w2312 & ~w5690 ) | ( w2312 & w5692 ) | ( ~w5690 & w5692 ) ;
  assign w5694 = \pi032 ^ w5693 ;
  assign w5695 = ( w5469 & w5477 ) | ( w5469 & w5478 ) | ( w5477 & w5478 ) ;
  assign w5696 = w5686 ^ w5695 ;
  assign w5697 = w5694 ^ w5696 ;
  assign w5698 = ~\pi087 & w1944 ;
  assign w5699 = \pi086 & w2072 ;
  assign w5700 = ( w1944 & ~w5698 ) | ( w1944 & w5699 ) | ( ~w5698 & w5699 ) ;
  assign w5701 = ~\pi088 & w1946 ;
  assign w5702 = w1574 | w5700 ;
  assign w5703 = ( w1947 & w5700 ) | ( w1947 & w5702 ) | ( w5700 & w5702 ) ;
  assign w5704 = ( w1946 & ~w5701 ) | ( w1946 & w5703 ) | ( ~w5701 & w5703 ) ;
  assign w5705 = \pi029 ^ w5704 ;
  assign w5706 = w5489 ^ w5697 ;
  assign w5707 = w5705 ^ w5706 ;
  assign w5708 = w5611 ^ w5707 ;
  assign w5709 = w5619 ^ w5708 ;
  assign w5710 = ~\pi093 & w1313 ;
  assign w5711 = \pi092 & w1417 ;
  assign w5712 = ( w1313 & ~w5710 ) | ( w1313 & w5711 ) | ( ~w5710 & w5711 ) ;
  assign w5713 = ~\pi094 & w1315 ;
  assign w5714 = w2274 | w5712 ;
  assign w5715 = ( w1316 & w5712 ) | ( w1316 & w5714 ) | ( w5712 & w5714 ) ;
  assign w5716 = ( w1315 & ~w5713 ) | ( w1315 & w5715 ) | ( ~w5713 & w5715 ) ;
  assign w5717 = \pi023 ^ w5716 ;
  assign w5718 = w5610 ^ w5709 ;
  assign w5719 = w5717 ^ w5718 ;
  assign w5720 = w5601 ^ w5719 ;
  assign w5721 = w5609 ^ w5720 ;
  assign w5722 = ~\pi099 & w837 ;
  assign w5723 = \pi098 & w902 ;
  assign w5724 = ( w837 & ~w5722 ) | ( w837 & w5723 ) | ( ~w5722 & w5723 ) ;
  assign w5725 = ~\pi100 & w839 ;
  assign w5726 = w3104 | w5724 ;
  assign w5727 = ( w840 & w5724 ) | ( w840 & w5726 ) | ( w5724 & w5726 ) ;
  assign w5728 = ( w839 & ~w5725 ) | ( w839 & w5727 ) | ( ~w5725 & w5727 ) ;
  assign w5729 = \pi017 ^ w5728 ;
  assign w5730 = w5600 ^ w5721 ;
  assign w5731 = w5729 ^ w5730 ;
  assign w5732 = ~\pi102 & w601 ;
  assign w5733 = \pi101 & w683 ;
  assign w5734 = ( w601 & ~w5732 ) | ( w601 & w5733 ) | ( ~w5732 & w5733 ) ;
  assign w5735 = ~\pi103 & w603 ;
  assign w5736 = w3437 | w5734 ;
  assign w5737 = ( w604 & w5734 ) | ( w604 & w5736 ) | ( w5734 & w5736 ) ;
  assign w5738 = ( w603 & ~w5735 ) | ( w603 & w5737 ) | ( ~w5735 & w5737 ) ;
  assign w5739 = \pi014 ^ w5738 ;
  assign w5740 = ( w5508 & w5516 ) | ( w5508 & w5517 ) | ( w5516 & w5517 ) ;
  assign w5741 = w5731 ^ w5740 ;
  assign w5742 = w5739 ^ w5741 ;
  assign w5743 = ~\pi105 & w432 ;
  assign w5744 = \pi104 & w486 ;
  assign w5745 = ( w432 & ~w5743 ) | ( w432 & w5744 ) | ( ~w5743 & w5744 ) ;
  assign w5746 = ~\pi106 & w434 ;
  assign w5747 = w4068 | w5745 ;
  assign w5748 = ( w435 & w5745 ) | ( w435 & w5747 ) | ( w5745 & w5747 ) ;
  assign w5749 = ( w434 & ~w5746 ) | ( w434 & w5748 ) | ( ~w5746 & w5748 ) ;
  assign w5750 = \pi011 ^ w5749 ;
  assign w5751 = ( w5519 & w5527 ) | ( w5519 & w5528 ) | ( w5527 & w5528 ) ;
  assign w5752 = w5742 ^ w5751 ;
  assign w5753 = w5750 ^ w5752 ;
  assign w5754 = w5539 ^ w5753 ;
  assign w5755 = w5599 ^ w5754 ;
  assign w5756 = ~\pi111 & w189 ;
  assign w5757 = \pi110 & w229 ;
  assign w5758 = ( w189 & ~w5756 ) | ( w189 & w5757 ) | ( ~w5756 & w5757 ) ;
  assign w5759 = ~\pi112 & w191 ;
  assign w5760 = w4999 | w5758 ;
  assign w5761 = ( w192 & w5758 ) | ( w192 & w5760 ) | ( w5758 & w5760 ) ;
  assign w5762 = ( w191 & ~w5759 ) | ( w191 & w5761 ) | ( ~w5759 & w5761 ) ;
  assign w5763 = \pi005 ^ w5762 ;
  assign w5764 = w5591 ^ w5755 ;
  assign w5765 = w5763 ^ w5764 ;
  assign w5766 = w5574 ^ w5765 ;
  assign w5767 = w5590 ^ w5766 ;
  assign w5768 = ( w5574 & w5590 ) | ( w5574 & w5765 ) | ( w5590 & w5765 ) ;
  assign w5769 = ( w5591 & w5755 ) | ( w5591 & w5763 ) | ( w5755 & w5763 ) ;
  assign w5770 = ( w5742 & w5750 ) | ( w5742 & w5751 ) | ( w5750 & w5751 ) ;
  assign w5771 = ( w5611 & w5619 ) | ( w5611 & w5707 ) | ( w5619 & w5707 ) ;
  assign w5772 = ( w5489 & w5697 ) | ( w5489 & w5705 ) | ( w5697 & w5705 ) ;
  assign w5773 = ( w5620 & w5628 ) | ( w5620 & w5684 ) | ( w5628 & w5684 ) ;
  assign w5774 = ~\pi079 & w3178 ;
  assign w5775 = \pi078 & w3340 ;
  assign w5776 = ( w3178 & ~w5774 ) | ( w3178 & w5775 ) | ( ~w5774 & w5775 ) ;
  assign w5777 = ~\pi080 & w3180 ;
  assign w5778 = w794 | w5776 ;
  assign w5779 = ( w3181 & w5776 ) | ( w3181 & w5778 ) | ( w5776 & w5778 ) ;
  assign w5780 = ( w3180 & ~w5777 ) | ( w3180 & w5779 ) | ( ~w5777 & w5779 ) ;
  assign w5781 = \pi038 ^ w5780 ;
  assign w5782 = ( w5638 & w5646 ) | ( w5638 & w5680 ) | ( w5646 & w5680 ) ;
  assign w5783 = ( w5647 & w5670 ) | ( w5647 & w5678 ) | ( w5670 & w5678 ) ;
  assign w5784 = ~\pi070 & w4654 ;
  assign w5785 = \pi069 & w4876 ;
  assign w5786 = ( w4654 & ~w5784 ) | ( w4654 & w5785 ) | ( ~w5784 & w5785 ) ;
  assign w5787 = ~\pi071 & w4656 ;
  assign w5788 = w290 | w5786 ;
  assign w5789 = ( w4657 & w5786 ) | ( w4657 & w5788 ) | ( w5786 & w5788 ) ;
  assign w5790 = ( w4656 & ~w5787 ) | ( w4656 & w5789 ) | ( ~w5787 & w5789 ) ;
  assign w5791 = \pi047 ^ w5790 ;
  assign w5792 = ( w5442 & w5663 ) | ( w5442 & w5666 ) | ( w5663 & w5666 ) ;
  assign w5793 = ~\pi067 & w5209 ;
  assign w5794 = \pi066 & w5433 ;
  assign w5795 = ( w5209 & ~w5793 ) | ( w5209 & w5794 ) | ( ~w5793 & w5794 ) ;
  assign w5796 = ~\pi068 & w5211 ;
  assign w5797 = w182 | w5795 ;
  assign w5798 = ( w5212 & w5795 ) | ( w5212 & w5797 ) | ( w5795 & w5797 ) ;
  assign w5799 = ( w5211 & ~w5796 ) | ( w5211 & w5798 ) | ( ~w5796 & w5798 ) ;
  assign w5800 = \pi050 ^ w5799 ;
  assign w5801 = ( \pi050 & \pi051 ) | ( \pi050 & \pi052 ) | ( \pi051 & \pi052 ) ;
  assign w5802 = \pi052 ^ w5801 ;
  assign w5803 = \pi052 ^ \pi053 ;
  assign w5804 = w5665 & ~w5803 ;
  assign w5805 = w5665 & w5803 ;
  assign w5806 = ( \pi050 & \pi051 ) | ( \pi050 & ~\pi053 ) | ( \pi051 & ~\pi053 ) ;
  assign w5807 = \pi053 & ~\pi064 ;
  assign w5808 = ~\pi065 & w5807 ;
  assign w5809 = ( \pi050 & \pi051 ) | ( \pi050 & ~w5808 ) | ( \pi051 & ~w5808 ) ;
  assign w5810 = ( \pi052 & \pi053 ) | ( \pi052 & ~w5809 ) | ( \pi053 & ~w5809 ) ;
  assign w5811 = ( \pi052 & ~w5807 ) | ( \pi052 & w5809 ) | ( ~w5807 & w5809 ) ;
  assign w5812 = ( w5806 & w5810 ) | ( w5806 & ~w5811 ) | ( w5810 & ~w5811 ) ;
  assign w5813 = ( \pi050 & \pi051 ) | ( \pi050 & \pi065 ) | ( \pi051 & \pi065 ) ;
  assign w5814 = \pi050 & \pi051 ;
  assign w5815 = \pi064 ^ w5814 ;
  assign w5816 = ( \pi052 & w5814 ) | ( \pi052 & w5815 ) | ( w5814 & w5815 ) ;
  assign w5817 = w5813 ^ w5816 ;
  assign w5818 = w5792 ^ w5800 ;
  assign w5819 = w5817 ^ w5818 ;
  assign w5820 = ( w5655 & w5667 ) | ( w5655 & w5668 ) | ( w5667 & w5668 ) ;
  assign w5821 = w5819 ^ w5820 ;
  assign w5822 = w5791 ^ w5821 ;
  assign w5823 = ~\pi073 & w4141 ;
  assign w5824 = \pi072 & w4334 ;
  assign w5825 = ( w4141 & ~w5823 ) | ( w4141 & w5824 ) | ( ~w5823 & w5824 ) ;
  assign w5826 = ~\pi074 & w4143 ;
  assign w5827 = w465 | w5825 ;
  assign w5828 = ( w4144 & w5825 ) | ( w4144 & w5827 ) | ( w5825 & w5827 ) ;
  assign w5829 = ( w4143 & ~w5826 ) | ( w4143 & w5828 ) | ( ~w5826 & w5828 ) ;
  assign w5830 = \pi044 ^ w5829 ;
  assign w5831 = ( w5783 & w5822 ) | ( w5783 & w5830 ) | ( w5822 & w5830 ) ;
  assign w5832 = w5783 ^ w5822 ;
  assign w5833 = w5830 ^ w5832 ;
  assign w5834 = ~\pi076 & w3635 ;
  assign w5835 = \pi075 & w3817 ;
  assign w5836 = ( w3635 & ~w5834 ) | ( w3635 & w5835 ) | ( ~w5834 & w5835 ) ;
  assign w5837 = ~\pi077 & w3637 ;
  assign w5838 = w644 | w5836 ;
  assign w5839 = ( w3638 & w5836 ) | ( w3638 & w5838 ) | ( w5836 & w5838 ) ;
  assign w5840 = ( w3637 & ~w5837 ) | ( w3637 & w5839 ) | ( ~w5837 & w5839 ) ;
  assign w5841 = \pi041 ^ w5840 ;
  assign w5842 = w5782 ^ w5833 ;
  assign w5843 = w5841 ^ w5842 ;
  assign w5844 = ( w5629 & w5637 ) | ( w5629 & w5682 ) | ( w5637 & w5682 ) ;
  assign w5845 = w5843 ^ w5844 ;
  assign w5846 = w5781 ^ w5845 ;
  assign w5847 = ~\pi082 & w2712 ;
  assign w5848 = \pi081 & w2872 ;
  assign w5849 = ( w2712 & ~w5847 ) | ( w2712 & w5848 ) | ( ~w5847 & w5848 ) ;
  assign w5850 = ~\pi083 & w2714 ;
  assign w5851 = w1099 | w5849 ;
  assign w5852 = ( w2715 & w5849 ) | ( w2715 & w5851 ) | ( w5849 & w5851 ) ;
  assign w5853 = ( w2714 & ~w5850 ) | ( w2714 & w5852 ) | ( ~w5850 & w5852 ) ;
  assign w5854 = \pi035 ^ w5853 ;
  assign w5855 = ( w5773 & w5846 ) | ( w5773 & w5854 ) | ( w5846 & w5854 ) ;
  assign w5856 = w5773 ^ w5846 ;
  assign w5857 = w5854 ^ w5856 ;
  assign w5858 = ~\pi085 & w2310 ;
  assign w5859 = \pi084 & w2443 ;
  assign w5860 = ( w2310 & ~w5858 ) | ( w2310 & w5859 ) | ( ~w5858 & w5859 ) ;
  assign w5861 = ~\pi086 & w2312 ;
  assign w5862 = w1379 | w5860 ;
  assign w5863 = ( w2313 & w5860 ) | ( w2313 & w5862 ) | ( w5860 & w5862 ) ;
  assign w5864 = ( w2312 & ~w5861 ) | ( w2312 & w5863 ) | ( ~w5861 & w5863 ) ;
  assign w5865 = \pi032 ^ w5864 ;
  assign w5866 = ( w5686 & w5694 ) | ( w5686 & w5695 ) | ( w5694 & w5695 ) ;
  assign w5867 = w5857 ^ w5866 ;
  assign w5868 = w5865 ^ w5867 ;
  assign w5869 = ~\pi088 & w1944 ;
  assign w5870 = \pi087 & w2072 ;
  assign w5871 = ( w1944 & ~w5869 ) | ( w1944 & w5870 ) | ( ~w5869 & w5870 ) ;
  assign w5872 = ~\pi089 & w1946 ;
  assign w5873 = w1595 | w5871 ;
  assign w5874 = ( w1947 & w5871 ) | ( w1947 & w5873 ) | ( w5871 & w5873 ) ;
  assign w5875 = ( w1946 & ~w5872 ) | ( w1946 & w5874 ) | ( ~w5872 & w5874 ) ;
  assign w5876 = \pi029 ^ w5875 ;
  assign w5877 = w5772 ^ w5868 ;
  assign w5878 = w5876 ^ w5877 ;
  assign w5879 = ~\pi091 & w1629 ;
  assign w5880 = \pi090 & w1722 ;
  assign w5881 = ( w1629 & ~w5879 ) | ( w1629 & w5880 ) | ( ~w5879 & w5880 ) ;
  assign w5882 = ~\pi092 & w1631 ;
  assign w5883 = w2033 | w5881 ;
  assign w5884 = ( w1632 & w5881 ) | ( w1632 & w5883 ) | ( w5881 & w5883 ) ;
  assign w5885 = ( w1631 & ~w5882 ) | ( w1631 & w5884 ) | ( ~w5882 & w5884 ) ;
  assign w5886 = \pi026 ^ w5885 ;
  assign w5887 = w5771 ^ w5878 ;
  assign w5888 = w5886 ^ w5887 ;
  assign w5889 = ~\pi094 & w1313 ;
  assign w5890 = \pi093 & w1417 ;
  assign w5891 = ( w1313 & ~w5889 ) | ( w1313 & w5890 ) | ( ~w5889 & w5890 ) ;
  assign w5892 = ~\pi095 & w1315 ;
  assign w5893 = w2409 | w5891 ;
  assign w5894 = ( w1316 & w5891 ) | ( w1316 & w5893 ) | ( w5891 & w5893 ) ;
  assign w5895 = ( w1315 & ~w5892 ) | ( w1315 & w5894 ) | ( ~w5892 & w5894 ) ;
  assign w5896 = \pi023 ^ w5895 ;
  assign w5897 = ( w5610 & w5709 ) | ( w5610 & w5717 ) | ( w5709 & w5717 ) ;
  assign w5898 = w5888 ^ w5897 ;
  assign w5899 = w5896 ^ w5898 ;
  assign w5900 = ~\pi097 & w1044 ;
  assign w5901 = \pi096 & w1138 ;
  assign w5902 = ( w1044 & ~w5900 ) | ( w1044 & w5901 ) | ( ~w5900 & w5901 ) ;
  assign w5903 = ~\pi098 & w1046 ;
  assign w5904 = w2824 | w5902 ;
  assign w5905 = ( w1047 & w5902 ) | ( w1047 & w5904 ) | ( w5902 & w5904 ) ;
  assign w5906 = ( w1046 & ~w5903 ) | ( w1046 & w5905 ) | ( ~w5903 & w5905 ) ;
  assign w5907 = \pi020 ^ w5906 ;
  assign w5908 = ( w5601 & w5609 ) | ( w5601 & w5719 ) | ( w5609 & w5719 ) ;
  assign w5909 = w5899 ^ w5908 ;
  assign w5910 = w5907 ^ w5909 ;
  assign w5911 = ~\pi100 & w837 ;
  assign w5912 = \pi099 & w902 ;
  assign w5913 = ( w837 & ~w5911 ) | ( w837 & w5912 ) | ( ~w5911 & w5912 ) ;
  assign w5914 = ~\pi101 & w839 ;
  assign w5915 = w3264 | w5913 ;
  assign w5916 = ( w840 & w5913 ) | ( w840 & w5915 ) | ( w5913 & w5915 ) ;
  assign w5917 = ( w839 & ~w5914 ) | ( w839 & w5916 ) | ( ~w5914 & w5916 ) ;
  assign w5918 = \pi017 ^ w5917 ;
  assign w5919 = ( w5600 & w5721 ) | ( w5600 & w5729 ) | ( w5721 & w5729 ) ;
  assign w5920 = w5910 ^ w5919 ;
  assign w5921 = w5918 ^ w5920 ;
  assign w5922 = ~\pi103 & w601 ;
  assign w5923 = \pi102 & w683 ;
  assign w5924 = ( w601 & ~w5922 ) | ( w601 & w5923 ) | ( ~w5922 & w5923 ) ;
  assign w5925 = ~\pi104 & w603 ;
  assign w5926 = w3740 | w5924 ;
  assign w5927 = ( w604 & w5924 ) | ( w604 & w5926 ) | ( w5924 & w5926 ) ;
  assign w5928 = ( w603 & ~w5925 ) | ( w603 & w5927 ) | ( ~w5925 & w5927 ) ;
  assign w5929 = \pi014 ^ w5928 ;
  assign w5930 = ( w5731 & w5739 ) | ( w5731 & w5740 ) | ( w5739 & w5740 ) ;
  assign w5931 = w5921 ^ w5930 ;
  assign w5932 = w5929 ^ w5931 ;
  assign w5933 = ~\pi106 & w432 ;
  assign w5934 = \pi105 & w486 ;
  assign w5935 = ( w432 & ~w5933 ) | ( w432 & w5934 ) | ( ~w5933 & w5934 ) ;
  assign w5936 = ~\pi107 & w434 ;
  assign w5937 = w4087 | w5935 ;
  assign w5938 = ( w435 & w5935 ) | ( w435 & w5937 ) | ( w5935 & w5937 ) ;
  assign w5939 = ( w434 & ~w5936 ) | ( w434 & w5938 ) | ( ~w5936 & w5938 ) ;
  assign w5940 = \pi011 ^ w5939 ;
  assign w5941 = ( w5770 & w5932 ) | ( w5770 & w5940 ) | ( w5932 & w5940 ) ;
  assign w5942 = w5770 ^ w5932 ;
  assign w5943 = w5940 ^ w5942 ;
  assign w5944 = ~\pi109 & w305 ;
  assign w5945 = \pi108 & w328 ;
  assign w5946 = ( w305 & ~w5944 ) | ( w305 & w5945 ) | ( ~w5944 & w5945 ) ;
  assign w5947 = ~\pi110 & w307 ;
  assign w5948 = w4792 | w5946 ;
  assign w5949 = ( w308 & w5946 ) | ( w308 & w5948 ) | ( w5946 & w5948 ) ;
  assign w5950 = ( w307 & ~w5947 ) | ( w307 & w5949 ) | ( ~w5947 & w5949 ) ;
  assign w5951 = \pi008 ^ w5950 ;
  assign w5952 = ( w5539 & w5599 ) | ( w5539 & w5753 ) | ( w5599 & w5753 ) ;
  assign w5953 = w5943 ^ w5952 ;
  assign w5954 = w5951 ^ w5953 ;
  assign w5955 = ~\pi112 & w189 ;
  assign w5956 = \pi111 & w229 ;
  assign w5957 = ( w189 & ~w5955 ) | ( w189 & w5956 ) | ( ~w5955 & w5956 ) ;
  assign w5958 = ~\pi113 & w191 ;
  assign w5959 = w5366 | w5957 ;
  assign w5960 = ( w192 & w5957 ) | ( w192 & w5959 ) | ( w5957 & w5959 ) ;
  assign w5961 = ( w191 & ~w5958 ) | ( w191 & w5960 ) | ( ~w5958 & w5960 ) ;
  assign w5962 = \pi005 ^ w5961 ;
  assign w5963 = w5769 ^ w5954 ;
  assign w5964 = w5962 ^ w5963 ;
  assign w5965 = ( ~\pi002 & \pi115 ) | ( ~\pi002 & \pi116 ) | ( \pi115 & \pi116 ) ;
  assign w5966 = \pi000 ^ w5965 ;
  assign w5967 = ( \pi002 & \pi116 ) | ( \pi002 & ~w5966 ) | ( \pi116 & ~w5966 ) ;
  assign w5968 = ( \pi002 & \pi115 ) | ( \pi002 & w5966 ) | ( \pi115 & w5966 ) ;
  assign w5969 = \pi001 & w5968 ;
  assign w5970 = ( ~\pi000 & \pi114 ) | ( ~\pi000 & w5969 ) | ( \pi114 & w5969 ) ;
  assign w5971 = ( \pi001 & \pi002 ) | ( \pi001 & ~w5970 ) | ( \pi002 & ~w5970 ) ;
  assign w5972 = ( w5967 & w5969 ) | ( w5967 & ~w5971 ) | ( w5969 & ~w5971 ) ;
  assign w5973 = ( \pi113 & ~\pi115 ) | ( \pi113 & w5563 ) | ( ~\pi115 & w5563 ) ;
  assign w5974 = ( ~\pi114 & \pi115 ) | ( ~\pi114 & w5973 ) | ( \pi115 & w5973 ) ;
  assign w5975 = \pi116 ^ w5973 ;
  assign w5976 = w5974 ^ w5975 ;
  assign w5977 = \pi002 ^ w5972 ;
  assign w5978 = \pi000 & ~w5972 ;
  assign w5979 = w5976 & w5978 ;
  assign w5980 = \pi001 ^ w5979 ;
  assign w5981 = ( \pi001 & w5977 ) | ( \pi001 & ~w5980 ) | ( w5977 & ~w5980 ) ;
  assign w5982 = w5768 ^ w5964 ;
  assign w5983 = w5981 ^ w5982 ;
  assign w5984 = ( w5768 & w5964 ) | ( w5768 & w5981 ) | ( w5964 & w5981 ) ;
  assign w5985 = ( w5769 & w5954 ) | ( w5769 & w5962 ) | ( w5954 & w5962 ) ;
  assign w5986 = ~\pi098 & w1044 ;
  assign w5987 = \pi097 & w1138 ;
  assign w5988 = ( w1044 & ~w5986 ) | ( w1044 & w5987 ) | ( ~w5986 & w5987 ) ;
  assign w5989 = ~\pi099 & w1046 ;
  assign w5990 = w2966 | w5988 ;
  assign w5991 = ( w1047 & w5988 ) | ( w1047 & w5990 ) | ( w5988 & w5990 ) ;
  assign w5992 = ( w1046 & ~w5989 ) | ( w1046 & w5991 ) | ( ~w5989 & w5991 ) ;
  assign w5993 = \pi020 ^ w5992 ;
  assign w5994 = ( w5888 & w5896 ) | ( w5888 & w5897 ) | ( w5896 & w5897 ) ;
  assign w5995 = ~\pi095 & w1313 ;
  assign w5996 = \pi094 & w1417 ;
  assign w5997 = ( w1313 & ~w5995 ) | ( w1313 & w5996 ) | ( ~w5995 & w5996 ) ;
  assign w5998 = ~\pi096 & w1315 ;
  assign w5999 = w2546 | w5997 ;
  assign w6000 = ( w1316 & w5997 ) | ( w1316 & w5999 ) | ( w5997 & w5999 ) ;
  assign w6001 = ( w1315 & ~w5998 ) | ( w1315 & w6000 ) | ( ~w5998 & w6000 ) ;
  assign w6002 = \pi023 ^ w6001 ;
  assign w6003 = ( w5771 & w5878 ) | ( w5771 & w5886 ) | ( w5878 & w5886 ) ;
  assign w6004 = ~\pi092 & w1629 ;
  assign w6005 = \pi091 & w1722 ;
  assign w6006 = ( w1629 & ~w6004 ) | ( w1629 & w6005 ) | ( ~w6004 & w6005 ) ;
  assign w6007 = ~\pi093 & w1631 ;
  assign w6008 = w2155 | w6006 ;
  assign w6009 = ( w1632 & w6006 ) | ( w1632 & w6008 ) | ( w6006 & w6008 ) ;
  assign w6010 = ( w1631 & ~w6007 ) | ( w1631 & w6009 ) | ( ~w6007 & w6009 ) ;
  assign w6011 = \pi026 ^ w6010 ;
  assign w6012 = ( w5772 & w5868 ) | ( w5772 & w5876 ) | ( w5868 & w5876 ) ;
  assign w6013 = ( w5857 & w5865 ) | ( w5857 & w5866 ) | ( w5865 & w5866 ) ;
  assign w6014 = ~\pi086 & w2310 ;
  assign w6015 = \pi085 & w2443 ;
  assign w6016 = ( w2310 & ~w6014 ) | ( w2310 & w6015 ) | ( ~w6014 & w6015 ) ;
  assign w6017 = ~\pi087 & w2312 ;
  assign w6018 = w1477 | w6016 ;
  assign w6019 = ( w2313 & w6016 ) | ( w2313 & w6018 ) | ( w6016 & w6018 ) ;
  assign w6020 = ( w2312 & ~w6017 ) | ( w2312 & w6019 ) | ( ~w6017 & w6019 ) ;
  assign w6021 = \pi032 ^ w6020 ;
  assign w6022 = ( w5781 & w5843 ) | ( w5781 & w5844 ) | ( w5843 & w5844 ) ;
  assign w6023 = ~\pi080 & w3178 ;
  assign w6024 = \pi079 & w3340 ;
  assign w6025 = ( w3178 & ~w6023 ) | ( w3178 & w6024 ) | ( ~w6023 & w6024 ) ;
  assign w6026 = ~\pi081 & w3180 ;
  assign w6027 = w874 | w6025 ;
  assign w6028 = ( w3181 & w6025 ) | ( w3181 & w6027 ) | ( w6025 & w6027 ) ;
  assign w6029 = ( w3180 & ~w6026 ) | ( w3180 & w6028 ) | ( ~w6026 & w6028 ) ;
  assign w6030 = \pi038 ^ w6029 ;
  assign w6031 = ( w5782 & w5833 ) | ( w5782 & w5841 ) | ( w5833 & w5841 ) ;
  assign w6032 = ~\pi077 & w3635 ;
  assign w6033 = \pi076 & w3817 ;
  assign w6034 = ( w3635 & ~w6032 ) | ( w3635 & w6033 ) | ( ~w6032 & w6033 ) ;
  assign w6035 = ~\pi078 & w3637 ;
  assign w6036 = w665 | w6034 ;
  assign w6037 = ( w3638 & w6034 ) | ( w3638 & w6036 ) | ( w6034 & w6036 ) ;
  assign w6038 = ( w3637 & ~w6035 ) | ( w3637 & w6037 ) | ( ~w6035 & w6037 ) ;
  assign w6039 = \pi041 ^ w6038 ;
  assign w6040 = ~\pi074 & w4141 ;
  assign w6041 = \pi073 & w4334 ;
  assign w6042 = ( w4141 & ~w6040 ) | ( w4141 & w6041 ) | ( ~w6040 & w6041 ) ;
  assign w6043 = ~\pi075 & w4143 ;
  assign w6044 = w519 | w6042 ;
  assign w6045 = ( w4144 & w6042 ) | ( w4144 & w6044 ) | ( w6042 & w6044 ) ;
  assign w6046 = ( w4143 & ~w6043 ) | ( w4143 & w6045 ) | ( ~w6043 & w6045 ) ;
  assign w6047 = \pi044 ^ w6046 ;
  assign w6048 = ( w5791 & w5819 ) | ( w5791 & w5820 ) | ( w5819 & w5820 ) ;
  assign w6049 = ( w5792 & w5800 ) | ( w5792 & w5817 ) | ( w5800 & w5817 ) ;
  assign w6050 = ( \pi051 & ~\pi052 ) | ( \pi051 & \pi053 ) | ( ~\pi052 & \pi053 ) ;
  assign w6051 = ( \pi050 & \pi051 ) | ( \pi050 & w6050 ) | ( \pi051 & w6050 ) ;
  assign w6052 = w6050 ^ w6051 ;
  assign w6053 = \pi064 & w6052 ;
  assign w6054 = ( \pi066 & w5804 ) | ( \pi066 & w6053 ) | ( w5804 & w6053 ) ;
  assign w6055 = \pi065 | w6054 ;
  assign w6056 = ( w5802 & w6054 ) | ( w5802 & w6055 ) | ( w6054 & w6055 ) ;
  assign w6057 = w6053 | w6056 ;
  assign w6058 = ~w134 & w5805 ;
  assign w6059 = ( w5805 & w6057 ) | ( w5805 & ~w6058 ) | ( w6057 & ~w6058 ) ;
  assign w6060 = \pi053 ^ w6059 ;
  assign w6061 = w5812 & w6060 ;
  assign w6062 = w5812 ^ w6060 ;
  assign w6063 = ~\pi068 & w5209 ;
  assign w6064 = \pi067 & w5433 ;
  assign w6065 = ( w5209 & ~w6063 ) | ( w5209 & w6064 ) | ( ~w6063 & w6064 ) ;
  assign w6066 = ~\pi069 & w5211 ;
  assign w6067 = w221 | w6065 ;
  assign w6068 = ( w5212 & w6065 ) | ( w5212 & w6067 ) | ( w6065 & w6067 ) ;
  assign w6069 = ( w5211 & ~w6066 ) | ( w5211 & w6068 ) | ( ~w6066 & w6068 ) ;
  assign w6070 = \pi050 ^ w6069 ;
  assign w6071 = ( w6049 & w6062 ) | ( w6049 & w6070 ) | ( w6062 & w6070 ) ;
  assign w6072 = w6049 ^ w6062 ;
  assign w6073 = w6070 ^ w6072 ;
  assign w6074 = ~\pi071 & w4654 ;
  assign w6075 = \pi070 & w4876 ;
  assign w6076 = ( w4654 & ~w6074 ) | ( w4654 & w6075 ) | ( ~w6074 & w6075 ) ;
  assign w6077 = ~\pi072 & w4656 ;
  assign w6078 = w361 | w6076 ;
  assign w6079 = ( w4657 & w6076 ) | ( w4657 & w6078 ) | ( w6076 & w6078 ) ;
  assign w6080 = ( w4656 & ~w6077 ) | ( w4656 & w6079 ) | ( ~w6077 & w6079 ) ;
  assign w6081 = \pi047 ^ w6080 ;
  assign w6082 = w6048 ^ w6073 ;
  assign w6083 = w6081 ^ w6082 ;
  assign w6084 = w5831 ^ w6083 ;
  assign w6085 = w6047 ^ w6084 ;
  assign w6086 = w6031 ^ w6085 ;
  assign w6087 = w6039 ^ w6086 ;
  assign w6088 = w6022 ^ w6087 ;
  assign w6089 = w6030 ^ w6088 ;
  assign w6090 = ~\pi083 & w2712 ;
  assign w6091 = \pi082 & w2872 ;
  assign w6092 = ( w2712 & ~w6090 ) | ( w2712 & w6091 ) | ( ~w6090 & w6091 ) ;
  assign w6093 = ~\pi084 & w2714 ;
  assign w6094 = w1188 | w6092 ;
  assign w6095 = ( w2715 & w6092 ) | ( w2715 & w6094 ) | ( w6092 & w6094 ) ;
  assign w6096 = ( w2714 & ~w6093 ) | ( w2714 & w6095 ) | ( ~w6093 & w6095 ) ;
  assign w6097 = \pi035 ^ w6096 ;
  assign w6098 = w5855 ^ w6089 ;
  assign w6099 = w6097 ^ w6098 ;
  assign w6100 = w6013 ^ w6099 ;
  assign w6101 = w6021 ^ w6100 ;
  assign w6102 = ~\pi089 & w1944 ;
  assign w6103 = \pi088 & w2072 ;
  assign w6104 = ( w1944 & ~w6102 ) | ( w1944 & w6103 ) | ( ~w6102 & w6103 ) ;
  assign w6105 = ~\pi090 & w1946 ;
  assign w6106 = w1801 | w6104 ;
  assign w6107 = ( w1947 & w6104 ) | ( w1947 & w6106 ) | ( w6104 & w6106 ) ;
  assign w6108 = ( w1946 & ~w6105 ) | ( w1946 & w6107 ) | ( ~w6105 & w6107 ) ;
  assign w6109 = \pi029 ^ w6108 ;
  assign w6110 = w6012 ^ w6101 ;
  assign w6111 = w6109 ^ w6110 ;
  assign w6112 = w6003 ^ w6111 ;
  assign w6113 = w6011 ^ w6112 ;
  assign w6114 = w5994 ^ w6113 ;
  assign w6115 = w6002 ^ w6114 ;
  assign w6116 = ( w5899 & w5907 ) | ( w5899 & w5908 ) | ( w5907 & w5908 ) ;
  assign w6117 = w6115 ^ w6116 ;
  assign w6118 = w5993 ^ w6117 ;
  assign w6119 = ~\pi101 & w837 ;
  assign w6120 = \pi100 & w902 ;
  assign w6121 = ( w837 & ~w6119 ) | ( w837 & w6120 ) | ( ~w6119 & w6120 ) ;
  assign w6122 = ~\pi102 & w839 ;
  assign w6123 = w3284 | w6121 ;
  assign w6124 = ( w840 & w6121 ) | ( w840 & w6123 ) | ( w6121 & w6123 ) ;
  assign w6125 = ( w839 & ~w6122 ) | ( w839 & w6124 ) | ( ~w6122 & w6124 ) ;
  assign w6126 = \pi017 ^ w6125 ;
  assign w6127 = ( w5910 & w5918 ) | ( w5910 & w5919 ) | ( w5918 & w5919 ) ;
  assign w6128 = w6118 ^ w6127 ;
  assign w6129 = w6126 ^ w6128 ;
  assign w6130 = ~\pi104 & w601 ;
  assign w6131 = \pi103 & w683 ;
  assign w6132 = ( w601 & ~w6130 ) | ( w601 & w6131 ) | ( ~w6130 & w6131 ) ;
  assign w6133 = ~\pi105 & w603 ;
  assign w6134 = w3905 | w6132 ;
  assign w6135 = ( w604 & w6132 ) | ( w604 & w6134 ) | ( w6132 & w6134 ) ;
  assign w6136 = ( w603 & ~w6133 ) | ( w603 & w6135 ) | ( ~w6133 & w6135 ) ;
  assign w6137 = \pi014 ^ w6136 ;
  assign w6138 = ( w5921 & w5929 ) | ( w5921 & w5930 ) | ( w5929 & w5930 ) ;
  assign w6139 = w6129 ^ w6138 ;
  assign w6140 = w6137 ^ w6139 ;
  assign w6141 = ~\pi107 & w432 ;
  assign w6142 = \pi106 & w486 ;
  assign w6143 = ( w432 & ~w6141 ) | ( w432 & w6142 ) | ( ~w6141 & w6142 ) ;
  assign w6144 = ~\pi108 & w434 ;
  assign w6145 = w4425 | w6143 ;
  assign w6146 = ( w435 & w6143 ) | ( w435 & w6145 ) | ( w6143 & w6145 ) ;
  assign w6147 = ( w434 & ~w6144 ) | ( w434 & w6146 ) | ( ~w6144 & w6146 ) ;
  assign w6148 = \pi011 ^ w6147 ;
  assign w6149 = ( w5941 & w6140 ) | ( w5941 & w6148 ) | ( w6140 & w6148 ) ;
  assign w6150 = w5941 ^ w6140 ;
  assign w6151 = w6148 ^ w6150 ;
  assign w6152 = ~\pi110 & w305 ;
  assign w6153 = \pi109 & w328 ;
  assign w6154 = ( w305 & ~w6152 ) | ( w305 & w6153 ) | ( ~w6152 & w6153 ) ;
  assign w6155 = ~\pi111 & w307 ;
  assign w6156 = w4811 | w6154 ;
  assign w6157 = ( w308 & w6154 ) | ( w308 & w6156 ) | ( w6154 & w6156 ) ;
  assign w6158 = ( w307 & ~w6155 ) | ( w307 & w6157 ) | ( ~w6155 & w6157 ) ;
  assign w6159 = \pi008 ^ w6158 ;
  assign w6160 = ( w5943 & w5951 ) | ( w5943 & w5952 ) | ( w5951 & w5952 ) ;
  assign w6161 = w6151 ^ w6160 ;
  assign w6162 = w6159 ^ w6161 ;
  assign w6163 = ~\pi113 & w189 ;
  assign w6164 = \pi112 & w229 ;
  assign w6165 = ( w189 & ~w6163 ) | ( w189 & w6164 ) | ( ~w6163 & w6164 ) ;
  assign w6166 = ~\pi114 & w191 ;
  assign w6167 = w5565 | w6165 ;
  assign w6168 = ( w192 & w6165 ) | ( w192 & w6167 ) | ( w6165 & w6167 ) ;
  assign w6169 = ( w191 & ~w6166 ) | ( w191 & w6168 ) | ( ~w6166 & w6168 ) ;
  assign w6170 = \pi005 ^ w6169 ;
  assign w6171 = ( w5985 & w6162 ) | ( w5985 & w6170 ) | ( w6162 & w6170 ) ;
  assign w6172 = w5985 ^ w6162 ;
  assign w6173 = w6170 ^ w6172 ;
  assign w6174 = ( ~\pi002 & \pi116 ) | ( ~\pi002 & \pi117 ) | ( \pi116 & \pi117 ) ;
  assign w6175 = \pi000 ^ w6174 ;
  assign w6176 = ( \pi002 & \pi117 ) | ( \pi002 & ~w6175 ) | ( \pi117 & ~w6175 ) ;
  assign w6177 = ( \pi002 & \pi116 ) | ( \pi002 & w6175 ) | ( \pi116 & w6175 ) ;
  assign w6178 = \pi001 & w6177 ;
  assign w6179 = ( ~\pi000 & \pi115 ) | ( ~\pi000 & w6178 ) | ( \pi115 & w6178 ) ;
  assign w6180 = ( \pi001 & \pi002 ) | ( \pi001 & ~w6179 ) | ( \pi002 & ~w6179 ) ;
  assign w6181 = ( w6176 & w6178 ) | ( w6176 & ~w6180 ) | ( w6178 & ~w6180 ) ;
  assign w6182 = ( \pi114 & \pi115 ) | ( \pi114 & \pi116 ) | ( \pi115 & \pi116 ) ;
  assign w6183 = ( \pi115 & w5583 ) | ( \pi115 & w6182 ) | ( w5583 & w6182 ) ;
  assign w6184 = \pi116 ^ \pi117 ;
  assign w6185 = w6183 ^ w6184 ;
  assign w6186 = \pi002 ^ w6181 ;
  assign w6187 = \pi000 & ~w6181 ;
  assign w6188 = w6185 & w6187 ;
  assign w6189 = \pi001 ^ w6188 ;
  assign w6190 = ( \pi001 & w6186 ) | ( \pi001 & ~w6189 ) | ( w6186 & ~w6189 ) ;
  assign w6191 = w5984 ^ w6173 ;
  assign w6192 = w6190 ^ w6191 ;
  assign w6193 = ( w5984 & w6173 ) | ( w5984 & w6190 ) | ( w6173 & w6190 ) ;
  assign w6194 = ( ~\pi002 & \pi117 ) | ( ~\pi002 & \pi118 ) | ( \pi117 & \pi118 ) ;
  assign w6195 = \pi000 ^ w6194 ;
  assign w6196 = ( \pi002 & \pi118 ) | ( \pi002 & ~w6195 ) | ( \pi118 & ~w6195 ) ;
  assign w6197 = ( \pi002 & \pi117 ) | ( \pi002 & w6195 ) | ( \pi117 & w6195 ) ;
  assign w6198 = \pi001 & w6197 ;
  assign w6199 = ( ~\pi000 & \pi116 ) | ( ~\pi000 & w6198 ) | ( \pi116 & w6198 ) ;
  assign w6200 = ( \pi001 & \pi002 ) | ( \pi001 & ~w6199 ) | ( \pi002 & ~w6199 ) ;
  assign w6201 = ( w6196 & w6198 ) | ( w6196 & ~w6200 ) | ( w6198 & ~w6200 ) ;
  assign w6202 = ( \pi114 & \pi115 ) | ( \pi114 & ~\pi117 ) | ( \pi115 & ~\pi117 ) ;
  assign w6203 = ( \pi115 & w5583 ) | ( \pi115 & w6202 ) | ( w5583 & w6202 ) ;
  assign w6204 = ( \pi116 & \pi117 ) | ( \pi116 & w6203 ) | ( \pi117 & w6203 ) ;
  assign w6205 = \pi117 ^ w6204 ;
  assign w6206 = \pi118 ^ w6205 ;
  assign w6207 = \pi002 ^ w6201 ;
  assign w6208 = \pi000 & ~w6201 ;
  assign w6209 = w6206 & w6208 ;
  assign w6210 = \pi001 ^ w6209 ;
  assign w6211 = ( \pi001 & w6207 ) | ( \pi001 & ~w6210 ) | ( w6207 & ~w6210 ) ;
  assign w6212 = ~\pi108 & w432 ;
  assign w6213 = \pi107 & w486 ;
  assign w6214 = ( w432 & ~w6212 ) | ( w432 & w6213 ) | ( ~w6212 & w6213 ) ;
  assign w6215 = ~\pi109 & w434 ;
  assign w6216 = w4599 | w6214 ;
  assign w6217 = ( w435 & w6214 ) | ( w435 & w6216 ) | ( w6214 & w6216 ) ;
  assign w6218 = ( w434 & ~w6215 ) | ( w434 & w6217 ) | ( ~w6215 & w6217 ) ;
  assign w6219 = \pi011 ^ w6218 ;
  assign w6220 = ( w6129 & w6137 ) | ( w6129 & w6138 ) | ( w6137 & w6138 ) ;
  assign w6221 = ( w5993 & w6115 ) | ( w5993 & w6116 ) | ( w6115 & w6116 ) ;
  assign w6222 = ( w5994 & w6002 ) | ( w5994 & w6113 ) | ( w6002 & w6113 ) ;
  assign w6223 = ( w6003 & w6011 ) | ( w6003 & w6111 ) | ( w6011 & w6111 ) ;
  assign w6224 = ~\pi093 & w1629 ;
  assign w6225 = \pi092 & w1722 ;
  assign w6226 = ( w1629 & ~w6224 ) | ( w1629 & w6225 ) | ( ~w6224 & w6225 ) ;
  assign w6227 = ~\pi094 & w1631 ;
  assign w6228 = w2274 | w6226 ;
  assign w6229 = ( w1632 & w6226 ) | ( w1632 & w6228 ) | ( w6226 & w6228 ) ;
  assign w6230 = ( w1631 & ~w6227 ) | ( w1631 & w6229 ) | ( ~w6227 & w6229 ) ;
  assign w6231 = \pi026 ^ w6230 ;
  assign w6232 = ( w6012 & w6101 ) | ( w6012 & w6109 ) | ( w6101 & w6109 ) ;
  assign w6233 = ~\pi090 & w1944 ;
  assign w6234 = \pi089 & w2072 ;
  assign w6235 = ( w1944 & ~w6233 ) | ( w1944 & w6234 ) | ( ~w6233 & w6234 ) ;
  assign w6236 = ~\pi091 & w1946 ;
  assign w6237 = w1908 | w6235 ;
  assign w6238 = ( w1947 & w6235 ) | ( w1947 & w6237 ) | ( w6235 & w6237 ) ;
  assign w6239 = ( w1946 & ~w6236 ) | ( w1946 & w6238 ) | ( ~w6236 & w6238 ) ;
  assign w6240 = \pi029 ^ w6239 ;
  assign w6241 = ( w6013 & w6021 ) | ( w6013 & w6099 ) | ( w6021 & w6099 ) ;
  assign w6242 = ~\pi087 & w2310 ;
  assign w6243 = \pi086 & w2443 ;
  assign w6244 = ( w2310 & ~w6242 ) | ( w2310 & w6243 ) | ( ~w6242 & w6243 ) ;
  assign w6245 = ~\pi088 & w2312 ;
  assign w6246 = w1574 | w6244 ;
  assign w6247 = ( w2313 & w6244 ) | ( w2313 & w6246 ) | ( w6244 & w6246 ) ;
  assign w6248 = ( w2312 & ~w6245 ) | ( w2312 & w6247 ) | ( ~w6245 & w6247 ) ;
  assign w6249 = \pi032 ^ w6248 ;
  assign w6250 = ( w5855 & w6089 ) | ( w5855 & w6097 ) | ( w6089 & w6097 ) ;
  assign w6251 = ~\pi084 & w2712 ;
  assign w6252 = \pi083 & w2872 ;
  assign w6253 = ( w2712 & ~w6251 ) | ( w2712 & w6252 ) | ( ~w6251 & w6252 ) ;
  assign w6254 = ~\pi085 & w2714 ;
  assign w6255 = w1274 | w6253 ;
  assign w6256 = ( w2715 & w6253 ) | ( w2715 & w6255 ) | ( w6253 & w6255 ) ;
  assign w6257 = ( w2714 & ~w6254 ) | ( w2714 & w6256 ) | ( ~w6254 & w6256 ) ;
  assign w6258 = \pi035 ^ w6257 ;
  assign w6259 = ( w6022 & w6030 ) | ( w6022 & w6087 ) | ( w6030 & w6087 ) ;
  assign w6260 = ~\pi081 & w3178 ;
  assign w6261 = \pi080 & w3340 ;
  assign w6262 = ( w3178 & ~w6260 ) | ( w3178 & w6261 ) | ( ~w6260 & w6261 ) ;
  assign w6263 = ~\pi082 & w3180 ;
  assign w6264 = w1008 | w6262 ;
  assign w6265 = ( w3181 & w6262 ) | ( w3181 & w6264 ) | ( w6262 & w6264 ) ;
  assign w6266 = ( w3180 & ~w6263 ) | ( w3180 & w6265 ) | ( ~w6263 & w6265 ) ;
  assign w6267 = \pi038 ^ w6266 ;
  assign w6268 = ( w6031 & w6039 ) | ( w6031 & w6085 ) | ( w6039 & w6085 ) ;
  assign w6269 = ~\pi078 & w3635 ;
  assign w6270 = \pi077 & w3817 ;
  assign w6271 = ( w3635 & ~w6269 ) | ( w3635 & w6270 ) | ( ~w6269 & w6270 ) ;
  assign w6272 = ~\pi079 & w3637 ;
  assign w6273 = w730 | w6271 ;
  assign w6274 = ( w3638 & w6271 ) | ( w3638 & w6273 ) | ( w6271 & w6273 ) ;
  assign w6275 = ( w3637 & ~w6272 ) | ( w3637 & w6274 ) | ( ~w6272 & w6274 ) ;
  assign w6276 = \pi041 ^ w6275 ;
  assign w6277 = ( w5831 & w6047 ) | ( w5831 & w6083 ) | ( w6047 & w6083 ) ;
  assign w6278 = ~\pi075 & w4141 ;
  assign w6279 = \pi074 & w4334 ;
  assign w6280 = ( w4141 & ~w6278 ) | ( w4141 & w6279 ) | ( ~w6278 & w6279 ) ;
  assign w6281 = ~\pi076 & w4143 ;
  assign w6282 = w538 | w6280 ;
  assign w6283 = ( w4144 & w6280 ) | ( w4144 & w6282 ) | ( w6280 & w6282 ) ;
  assign w6284 = ( w4143 & ~w6281 ) | ( w4143 & w6283 ) | ( ~w6281 & w6283 ) ;
  assign w6285 = \pi044 ^ w6284 ;
  assign w6286 = ( w6048 & w6073 ) | ( w6048 & w6081 ) | ( w6073 & w6081 ) ;
  assign w6287 = ~\pi072 & w4654 ;
  assign w6288 = \pi071 & w4876 ;
  assign w6289 = ( w4654 & ~w6287 ) | ( w4654 & w6288 ) | ( ~w6287 & w6288 ) ;
  assign w6290 = ~\pi073 & w4656 ;
  assign w6291 = w404 | w6289 ;
  assign w6292 = ( w4657 & w6289 ) | ( w4657 & w6291 ) | ( w6289 & w6291 ) ;
  assign w6293 = ( w4656 & ~w6290 ) | ( w4656 & w6292 ) | ( ~w6290 & w6292 ) ;
  assign w6294 = \pi047 ^ w6293 ;
  assign w6295 = ~\pi069 & w5209 ;
  assign w6296 = \pi068 & w5433 ;
  assign w6297 = ( w5209 & ~w6295 ) | ( w5209 & w6296 ) | ( ~w6295 & w6296 ) ;
  assign w6298 = ~\pi070 & w5211 ;
  assign w6299 = w271 | w6297 ;
  assign w6300 = ( w5212 & w6297 ) | ( w5212 & w6299 ) | ( w6297 & w6299 ) ;
  assign w6301 = ( w5211 & ~w6298 ) | ( w5211 & w6300 ) | ( ~w6298 & w6300 ) ;
  assign w6302 = \pi050 ^ w6301 ;
  assign w6303 = ~\pi066 & w5802 ;
  assign w6304 = \pi065 & w6052 ;
  assign w6305 = ( w5802 & ~w6303 ) | ( w5802 & w6304 ) | ( ~w6303 & w6304 ) ;
  assign w6306 = ~\pi067 & w5804 ;
  assign w6307 = w160 | w6305 ;
  assign w6308 = ( w5805 & w6305 ) | ( w5805 & w6307 ) | ( w6305 & w6307 ) ;
  assign w6309 = ( w5804 & ~w6306 ) | ( w5804 & w6308 ) | ( ~w6306 & w6308 ) ;
  assign w6310 = \pi053 ^ w6309 ;
  assign w6311 = w6061 ^ w6310 ;
  assign w6312 = \pi053 ^ \pi054 ;
  assign w6313 = \pi064 & w6312 ;
  assign w6314 = w6311 ^ w6313 ;
  assign w6315 = w6071 ^ w6314 ;
  assign w6316 = w6302 ^ w6315 ;
  assign w6317 = w6286 ^ w6316 ;
  assign w6318 = w6294 ^ w6317 ;
  assign w6319 = w6277 ^ w6318 ;
  assign w6320 = w6285 ^ w6319 ;
  assign w6321 = w6268 ^ w6320 ;
  assign w6322 = w6276 ^ w6321 ;
  assign w6323 = w6259 ^ w6322 ;
  assign w6324 = w6267 ^ w6323 ;
  assign w6325 = w6250 ^ w6324 ;
  assign w6326 = w6258 ^ w6325 ;
  assign w6327 = w6241 ^ w6326 ;
  assign w6328 = w6249 ^ w6327 ;
  assign w6329 = w6232 ^ w6328 ;
  assign w6330 = w6240 ^ w6329 ;
  assign w6331 = w6223 ^ w6330 ;
  assign w6332 = w6231 ^ w6331 ;
  assign w6333 = ~\pi096 & w1313 ;
  assign w6334 = \pi095 & w1417 ;
  assign w6335 = ( w1313 & ~w6333 ) | ( w1313 & w6334 ) | ( ~w6333 & w6334 ) ;
  assign w6336 = ~\pi097 & w1315 ;
  assign w6337 = w2673 | w6335 ;
  assign w6338 = ( w1316 & w6335 ) | ( w1316 & w6337 ) | ( w6335 & w6337 ) ;
  assign w6339 = ( w1315 & ~w6336 ) | ( w1315 & w6338 ) | ( ~w6336 & w6338 ) ;
  assign w6340 = \pi023 ^ w6339 ;
  assign w6341 = w6222 ^ w6332 ;
  assign w6342 = w6340 ^ w6341 ;
  assign w6343 = ~\pi099 & w1044 ;
  assign w6344 = \pi098 & w1138 ;
  assign w6345 = ( w1044 & ~w6343 ) | ( w1044 & w6344 ) | ( ~w6343 & w6344 ) ;
  assign w6346 = ~\pi100 & w1046 ;
  assign w6347 = w3104 | w6345 ;
  assign w6348 = ( w1047 & w6345 ) | ( w1047 & w6347 ) | ( w6345 & w6347 ) ;
  assign w6349 = ( w1046 & ~w6346 ) | ( w1046 & w6348 ) | ( ~w6346 & w6348 ) ;
  assign w6350 = \pi020 ^ w6349 ;
  assign w6351 = w6221 ^ w6342 ;
  assign w6352 = w6350 ^ w6351 ;
  assign w6353 = ~\pi102 & w837 ;
  assign w6354 = \pi101 & w902 ;
  assign w6355 = ( w837 & ~w6353 ) | ( w837 & w6354 ) | ( ~w6353 & w6354 ) ;
  assign w6356 = ~\pi103 & w839 ;
  assign w6357 = w3437 | w6355 ;
  assign w6358 = ( w840 & w6355 ) | ( w840 & w6357 ) | ( w6355 & w6357 ) ;
  assign w6359 = ( w839 & ~w6356 ) | ( w839 & w6358 ) | ( ~w6356 & w6358 ) ;
  assign w6360 = \pi017 ^ w6359 ;
  assign w6361 = ( w6118 & w6126 ) | ( w6118 & w6127 ) | ( w6126 & w6127 ) ;
  assign w6362 = w6352 ^ w6361 ;
  assign w6363 = w6360 ^ w6362 ;
  assign w6364 = ~\pi105 & w601 ;
  assign w6365 = \pi104 & w683 ;
  assign w6366 = ( w601 & ~w6364 ) | ( w601 & w6365 ) | ( ~w6364 & w6365 ) ;
  assign w6367 = ~\pi106 & w603 ;
  assign w6368 = w4068 | w6366 ;
  assign w6369 = ( w604 & w6366 ) | ( w604 & w6368 ) | ( w6366 & w6368 ) ;
  assign w6370 = ( w603 & ~w6367 ) | ( w603 & w6369 ) | ( ~w6367 & w6369 ) ;
  assign w6371 = \pi014 ^ w6370 ;
  assign w6372 = w6220 ^ w6363 ;
  assign w6373 = w6371 ^ w6372 ;
  assign w6374 = w6149 ^ w6373 ;
  assign w6375 = w6219 ^ w6374 ;
  assign w6376 = ~\pi111 & w305 ;
  assign w6377 = \pi110 & w328 ;
  assign w6378 = ( w305 & ~w6376 ) | ( w305 & w6377 ) | ( ~w6376 & w6377 ) ;
  assign w6379 = ~\pi112 & w307 ;
  assign w6380 = w4999 | w6378 ;
  assign w6381 = ( w308 & w6378 ) | ( w308 & w6380 ) | ( w6378 & w6380 ) ;
  assign w6382 = ( w307 & ~w6379 ) | ( w307 & w6381 ) | ( ~w6379 & w6381 ) ;
  assign w6383 = \pi008 ^ w6382 ;
  assign w6384 = ( w6151 & w6159 ) | ( w6151 & w6160 ) | ( w6159 & w6160 ) ;
  assign w6385 = w6375 ^ w6384 ;
  assign w6386 = w6383 ^ w6385 ;
  assign w6387 = ~\pi114 & w189 ;
  assign w6388 = \pi113 & w229 ;
  assign w6389 = ( w189 & ~w6387 ) | ( w189 & w6388 ) | ( ~w6387 & w6388 ) ;
  assign w6390 = ~\pi115 & w191 ;
  assign w6391 = w5585 | w6389 ;
  assign w6392 = ( w192 & w6389 ) | ( w192 & w6391 ) | ( w6389 & w6391 ) ;
  assign w6393 = ( w191 & ~w6390 ) | ( w191 & w6392 ) | ( ~w6390 & w6392 ) ;
  assign w6394 = \pi005 ^ w6393 ;
  assign w6395 = w6171 ^ w6386 ;
  assign w6396 = w6394 ^ w6395 ;
  assign w6397 = w6193 ^ w6396 ;
  assign w6398 = w6211 ^ w6397 ;
  assign w6399 = ( w6193 & w6211 ) | ( w6193 & w6396 ) | ( w6211 & w6396 ) ;
  assign w6400 = ( w6171 & w6386 ) | ( w6171 & w6394 ) | ( w6386 & w6394 ) ;
  assign w6401 = ~\pi115 & w189 ;
  assign w6402 = \pi114 & w229 ;
  assign w6403 = ( w189 & ~w6401 ) | ( w189 & w6402 ) | ( ~w6401 & w6402 ) ;
  assign w6404 = ~\pi116 & w191 ;
  assign w6405 = w5976 | w6403 ;
  assign w6406 = ( w192 & w6403 ) | ( w192 & w6405 ) | ( w6403 & w6405 ) ;
  assign w6407 = ( w191 & ~w6404 ) | ( w191 & w6406 ) | ( ~w6404 & w6406 ) ;
  assign w6408 = \pi005 ^ w6407 ;
  assign w6409 = ( w6375 & w6383 ) | ( w6375 & w6384 ) | ( w6383 & w6384 ) ;
  assign w6410 = ~\pi112 & w305 ;
  assign w6411 = \pi111 & w328 ;
  assign w6412 = ( w305 & ~w6410 ) | ( w305 & w6411 ) | ( ~w6410 & w6411 ) ;
  assign w6413 = ~\pi113 & w307 ;
  assign w6414 = w5366 | w6412 ;
  assign w6415 = ( w308 & w6412 ) | ( w308 & w6414 ) | ( w6412 & w6414 ) ;
  assign w6416 = ( w307 & ~w6413 ) | ( w307 & w6415 ) | ( ~w6413 & w6415 ) ;
  assign w6417 = \pi008 ^ w6416 ;
  assign w6418 = ( w6149 & w6219 ) | ( w6149 & w6373 ) | ( w6219 & w6373 ) ;
  assign w6419 = ( w6220 & w6363 ) | ( w6220 & w6371 ) | ( w6363 & w6371 ) ;
  assign w6420 = ( w6259 & w6267 ) | ( w6259 & w6322 ) | ( w6267 & w6322 ) ;
  assign w6421 = ~\pi079 & w3635 ;
  assign w6422 = \pi078 & w3817 ;
  assign w6423 = ( w3635 & ~w6421 ) | ( w3635 & w6422 ) | ( ~w6421 & w6422 ) ;
  assign w6424 = ~\pi080 & w3637 ;
  assign w6425 = w794 | w6423 ;
  assign w6426 = ( w3638 & w6423 ) | ( w3638 & w6425 ) | ( w6423 & w6425 ) ;
  assign w6427 = ( w3637 & ~w6424 ) | ( w3637 & w6426 ) | ( ~w6424 & w6426 ) ;
  assign w6428 = \pi041 ^ w6427 ;
  assign w6429 = ( w6277 & w6285 ) | ( w6277 & w6318 ) | ( w6285 & w6318 ) ;
  assign w6430 = ~\pi076 & w4141 ;
  assign w6431 = \pi075 & w4334 ;
  assign w6432 = ( w4141 & ~w6430 ) | ( w4141 & w6431 ) | ( ~w6430 & w6431 ) ;
  assign w6433 = ~\pi077 & w4143 ;
  assign w6434 = w644 | w6432 ;
  assign w6435 = ( w4144 & w6432 ) | ( w4144 & w6434 ) | ( w6432 & w6434 ) ;
  assign w6436 = ( w4143 & ~w6433 ) | ( w4143 & w6435 ) | ( ~w6433 & w6435 ) ;
  assign w6437 = \pi044 ^ w6436 ;
  assign w6438 = ( w6286 & w6294 ) | ( w6286 & w6316 ) | ( w6294 & w6316 ) ;
  assign w6439 = ~\pi073 & w4654 ;
  assign w6440 = \pi072 & w4876 ;
  assign w6441 = ( w4654 & ~w6439 ) | ( w4654 & w6440 ) | ( ~w6439 & w6440 ) ;
  assign w6442 = ~\pi074 & w4656 ;
  assign w6443 = w465 | w6441 ;
  assign w6444 = ( w4657 & w6441 ) | ( w4657 & w6443 ) | ( w6441 & w6443 ) ;
  assign w6445 = ( w4656 & ~w6442 ) | ( w4656 & w6444 ) | ( ~w6442 & w6444 ) ;
  assign w6446 = \pi047 ^ w6445 ;
  assign w6447 = ( w6071 & w6302 ) | ( w6071 & w6314 ) | ( w6302 & w6314 ) ;
  assign w6448 = ~\pi070 & w5209 ;
  assign w6449 = \pi069 & w5433 ;
  assign w6450 = ( w5209 & ~w6448 ) | ( w5209 & w6449 ) | ( ~w6448 & w6449 ) ;
  assign w6451 = ~\pi071 & w5211 ;
  assign w6452 = w290 | w6450 ;
  assign w6453 = ( w5212 & w6450 ) | ( w5212 & w6452 ) | ( w6450 & w6452 ) ;
  assign w6454 = ( w5211 & ~w6451 ) | ( w5211 & w6453 ) | ( ~w6451 & w6453 ) ;
  assign w6455 = \pi050 ^ w6454 ;
  assign w6456 = ( w6061 & w6310 ) | ( w6061 & w6313 ) | ( w6310 & w6313 ) ;
  assign w6457 = ~\pi067 & w5802 ;
  assign w6458 = \pi066 & w6052 ;
  assign w6459 = ( w5802 & ~w6457 ) | ( w5802 & w6458 ) | ( ~w6457 & w6458 ) ;
  assign w6460 = ~\pi068 & w5804 ;
  assign w6461 = w182 | w6459 ;
  assign w6462 = ( w5805 & w6459 ) | ( w5805 & w6461 ) | ( w6459 & w6461 ) ;
  assign w6463 = ( w5804 & ~w6460 ) | ( w5804 & w6462 ) | ( ~w6460 & w6462 ) ;
  assign w6464 = \pi053 ^ w6463 ;
  assign w6465 = ( \pi053 & \pi054 ) | ( \pi053 & \pi055 ) | ( \pi054 & \pi055 ) ;
  assign w6466 = \pi055 ^ w6465 ;
  assign w6467 = \pi055 ^ \pi056 ;
  assign w6468 = w6312 & ~w6467 ;
  assign w6469 = w6312 & w6467 ;
  assign w6470 = ( \pi053 & \pi054 ) | ( \pi053 & ~\pi056 ) | ( \pi054 & ~\pi056 ) ;
  assign w6471 = \pi056 & ~\pi064 ;
  assign w6472 = ~\pi065 & w6471 ;
  assign w6473 = ( \pi053 & \pi054 ) | ( \pi053 & ~w6472 ) | ( \pi054 & ~w6472 ) ;
  assign w6474 = ( \pi055 & \pi056 ) | ( \pi055 & ~w6473 ) | ( \pi056 & ~w6473 ) ;
  assign w6475 = ( \pi055 & ~w6471 ) | ( \pi055 & w6473 ) | ( ~w6471 & w6473 ) ;
  assign w6476 = ( w6470 & w6474 ) | ( w6470 & ~w6475 ) | ( w6474 & ~w6475 ) ;
  assign w6477 = ( \pi053 & \pi054 ) | ( \pi053 & \pi065 ) | ( \pi054 & \pi065 ) ;
  assign w6478 = \pi053 & \pi054 ;
  assign w6479 = \pi064 ^ w6478 ;
  assign w6480 = ( \pi055 & w6478 ) | ( \pi055 & w6479 ) | ( w6478 & w6479 ) ;
  assign w6481 = w6477 ^ w6480 ;
  assign w6482 = w6456 ^ w6464 ;
  assign w6483 = w6481 ^ w6482 ;
  assign w6484 = w6447 ^ w6483 ;
  assign w6485 = w6455 ^ w6484 ;
  assign w6486 = w6438 ^ w6485 ;
  assign w6487 = w6446 ^ w6486 ;
  assign w6488 = w6429 ^ w6487 ;
  assign w6489 = w6437 ^ w6488 ;
  assign w6490 = ( w6268 & w6276 ) | ( w6268 & w6320 ) | ( w6276 & w6320 ) ;
  assign w6491 = w6489 ^ w6490 ;
  assign w6492 = w6428 ^ w6491 ;
  assign w6493 = ~\pi082 & w3178 ;
  assign w6494 = \pi081 & w3340 ;
  assign w6495 = ( w3178 & ~w6493 ) | ( w3178 & w6494 ) | ( ~w6493 & w6494 ) ;
  assign w6496 = ~\pi083 & w3180 ;
  assign w6497 = w1099 | w6495 ;
  assign w6498 = ( w3181 & w6495 ) | ( w3181 & w6497 ) | ( w6495 & w6497 ) ;
  assign w6499 = ( w3180 & ~w6496 ) | ( w3180 & w6498 ) | ( ~w6496 & w6498 ) ;
  assign w6500 = \pi038 ^ w6499 ;
  assign w6501 = ( w6420 & w6492 ) | ( w6420 & w6500 ) | ( w6492 & w6500 ) ;
  assign w6502 = w6420 ^ w6492 ;
  assign w6503 = w6500 ^ w6502 ;
  assign w6504 = ~\pi085 & w2712 ;
  assign w6505 = \pi084 & w2872 ;
  assign w6506 = ( w2712 & ~w6504 ) | ( w2712 & w6505 ) | ( ~w6504 & w6505 ) ;
  assign w6507 = ~\pi086 & w2714 ;
  assign w6508 = w1379 | w6506 ;
  assign w6509 = ( w2715 & w6506 ) | ( w2715 & w6508 ) | ( w6506 & w6508 ) ;
  assign w6510 = ( w2714 & ~w6507 ) | ( w2714 & w6509 ) | ( ~w6507 & w6509 ) ;
  assign w6511 = \pi035 ^ w6510 ;
  assign w6512 = ( w6250 & w6258 ) | ( w6250 & w6324 ) | ( w6258 & w6324 ) ;
  assign w6513 = w6503 ^ w6512 ;
  assign w6514 = w6511 ^ w6513 ;
  assign w6515 = ~\pi088 & w2310 ;
  assign w6516 = \pi087 & w2443 ;
  assign w6517 = ( w2310 & ~w6515 ) | ( w2310 & w6516 ) | ( ~w6515 & w6516 ) ;
  assign w6518 = ~\pi089 & w2312 ;
  assign w6519 = w1595 | w6517 ;
  assign w6520 = ( w2313 & w6517 ) | ( w2313 & w6519 ) | ( w6517 & w6519 ) ;
  assign w6521 = ( w2312 & ~w6518 ) | ( w2312 & w6520 ) | ( ~w6518 & w6520 ) ;
  assign w6522 = \pi032 ^ w6521 ;
  assign w6523 = ( w6241 & w6249 ) | ( w6241 & w6326 ) | ( w6249 & w6326 ) ;
  assign w6524 = w6514 ^ w6523 ;
  assign w6525 = w6522 ^ w6524 ;
  assign w6526 = ~\pi091 & w1944 ;
  assign w6527 = \pi090 & w2072 ;
  assign w6528 = ( w1944 & ~w6526 ) | ( w1944 & w6527 ) | ( ~w6526 & w6527 ) ;
  assign w6529 = ~\pi092 & w1946 ;
  assign w6530 = w2033 | w6528 ;
  assign w6531 = ( w1947 & w6528 ) | ( w1947 & w6530 ) | ( w6528 & w6530 ) ;
  assign w6532 = ( w1946 & ~w6529 ) | ( w1946 & w6531 ) | ( ~w6529 & w6531 ) ;
  assign w6533 = \pi029 ^ w6532 ;
  assign w6534 = ( w6232 & w6240 ) | ( w6232 & w6328 ) | ( w6240 & w6328 ) ;
  assign w6535 = w6525 ^ w6534 ;
  assign w6536 = w6533 ^ w6535 ;
  assign w6537 = ~\pi094 & w1629 ;
  assign w6538 = \pi093 & w1722 ;
  assign w6539 = ( w1629 & ~w6537 ) | ( w1629 & w6538 ) | ( ~w6537 & w6538 ) ;
  assign w6540 = ~\pi095 & w1631 ;
  assign w6541 = w2409 | w6539 ;
  assign w6542 = ( w1632 & w6539 ) | ( w1632 & w6541 ) | ( w6539 & w6541 ) ;
  assign w6543 = ( w1631 & ~w6540 ) | ( w1631 & w6542 ) | ( ~w6540 & w6542 ) ;
  assign w6544 = \pi026 ^ w6543 ;
  assign w6545 = ( w6223 & w6231 ) | ( w6223 & w6330 ) | ( w6231 & w6330 ) ;
  assign w6546 = w6536 ^ w6545 ;
  assign w6547 = w6544 ^ w6546 ;
  assign w6548 = ~\pi097 & w1313 ;
  assign w6549 = \pi096 & w1417 ;
  assign w6550 = ( w1313 & ~w6548 ) | ( w1313 & w6549 ) | ( ~w6548 & w6549 ) ;
  assign w6551 = ~\pi098 & w1315 ;
  assign w6552 = w2824 | w6550 ;
  assign w6553 = ( w1316 & w6550 ) | ( w1316 & w6552 ) | ( w6550 & w6552 ) ;
  assign w6554 = ( w1315 & ~w6551 ) | ( w1315 & w6553 ) | ( ~w6551 & w6553 ) ;
  assign w6555 = \pi023 ^ w6554 ;
  assign w6556 = ( w6222 & w6332 ) | ( w6222 & w6340 ) | ( w6332 & w6340 ) ;
  assign w6557 = w6547 ^ w6556 ;
  assign w6558 = w6555 ^ w6557 ;
  assign w6559 = ~\pi100 & w1044 ;
  assign w6560 = \pi099 & w1138 ;
  assign w6561 = ( w1044 & ~w6559 ) | ( w1044 & w6560 ) | ( ~w6559 & w6560 ) ;
  assign w6562 = ~\pi101 & w1046 ;
  assign w6563 = w3264 | w6561 ;
  assign w6564 = ( w1047 & w6561 ) | ( w1047 & w6563 ) | ( w6561 & w6563 ) ;
  assign w6565 = ( w1046 & ~w6562 ) | ( w1046 & w6564 ) | ( ~w6562 & w6564 ) ;
  assign w6566 = \pi020 ^ w6565 ;
  assign w6567 = ( w6221 & w6342 ) | ( w6221 & w6350 ) | ( w6342 & w6350 ) ;
  assign w6568 = w6558 ^ w6567 ;
  assign w6569 = w6566 ^ w6568 ;
  assign w6570 = ~\pi103 & w837 ;
  assign w6571 = \pi102 & w902 ;
  assign w6572 = ( w837 & ~w6570 ) | ( w837 & w6571 ) | ( ~w6570 & w6571 ) ;
  assign w6573 = ~\pi104 & w839 ;
  assign w6574 = w3740 | w6572 ;
  assign w6575 = ( w840 & w6572 ) | ( w840 & w6574 ) | ( w6572 & w6574 ) ;
  assign w6576 = ( w839 & ~w6573 ) | ( w839 & w6575 ) | ( ~w6573 & w6575 ) ;
  assign w6577 = \pi017 ^ w6576 ;
  assign w6578 = ( w6352 & w6360 ) | ( w6352 & w6361 ) | ( w6360 & w6361 ) ;
  assign w6579 = w6569 ^ w6578 ;
  assign w6580 = w6577 ^ w6579 ;
  assign w6581 = ~\pi106 & w601 ;
  assign w6582 = \pi105 & w683 ;
  assign w6583 = ( w601 & ~w6581 ) | ( w601 & w6582 ) | ( ~w6581 & w6582 ) ;
  assign w6584 = ~\pi107 & w603 ;
  assign w6585 = w4087 | w6583 ;
  assign w6586 = ( w604 & w6583 ) | ( w604 & w6585 ) | ( w6583 & w6585 ) ;
  assign w6587 = ( w603 & ~w6584 ) | ( w603 & w6586 ) | ( ~w6584 & w6586 ) ;
  assign w6588 = \pi014 ^ w6587 ;
  assign w6589 = ( w6419 & w6580 ) | ( w6419 & w6588 ) | ( w6580 & w6588 ) ;
  assign w6590 = w6419 ^ w6580 ;
  assign w6591 = w6588 ^ w6590 ;
  assign w6592 = ~\pi109 & w432 ;
  assign w6593 = \pi108 & w486 ;
  assign w6594 = ( w432 & ~w6592 ) | ( w432 & w6593 ) | ( ~w6592 & w6593 ) ;
  assign w6595 = ~\pi110 & w434 ;
  assign w6596 = w4792 | w6594 ;
  assign w6597 = ( w435 & w6594 ) | ( w435 & w6596 ) | ( w6594 & w6596 ) ;
  assign w6598 = ( w434 & ~w6595 ) | ( w434 & w6597 ) | ( ~w6595 & w6597 ) ;
  assign w6599 = \pi011 ^ w6598 ;
  assign w6600 = w6418 ^ w6591 ;
  assign w6601 = w6599 ^ w6600 ;
  assign w6602 = w6409 ^ w6601 ;
  assign w6603 = w6417 ^ w6602 ;
  assign w6604 = w6400 ^ w6603 ;
  assign w6605 = w6408 ^ w6604 ;
  assign w6606 = ( ~\pi002 & \pi118 ) | ( ~\pi002 & \pi119 ) | ( \pi118 & \pi119 ) ;
  assign w6607 = \pi000 ^ w6606 ;
  assign w6608 = ( \pi002 & \pi119 ) | ( \pi002 & ~w6607 ) | ( \pi119 & ~w6607 ) ;
  assign w6609 = ( \pi002 & \pi118 ) | ( \pi002 & w6607 ) | ( \pi118 & w6607 ) ;
  assign w6610 = \pi001 & w6609 ;
  assign w6611 = ( ~\pi000 & \pi117 ) | ( ~\pi000 & w6610 ) | ( \pi117 & w6610 ) ;
  assign w6612 = ( \pi001 & \pi002 ) | ( \pi001 & ~w6611 ) | ( \pi002 & ~w6611 ) ;
  assign w6613 = ( w6608 & w6610 ) | ( w6608 & ~w6612 ) | ( w6610 & ~w6612 ) ;
  assign w6614 = ( \pi117 & \pi118 ) | ( \pi117 & w6204 ) | ( \pi118 & w6204 ) ;
  assign w6615 = \pi118 ^ w6614 ;
  assign w6616 = \pi119 ^ w6615 ;
  assign w6617 = \pi002 ^ w6613 ;
  assign w6618 = \pi000 & ~w6613 ;
  assign w6619 = w6616 & w6618 ;
  assign w6620 = \pi001 ^ w6619 ;
  assign w6621 = ( \pi001 & w6617 ) | ( \pi001 & ~w6620 ) | ( w6617 & ~w6620 ) ;
  assign w6622 = w6399 ^ w6605 ;
  assign w6623 = w6621 ^ w6622 ;
  assign w6624 = ( ~\pi002 & \pi119 ) | ( ~\pi002 & \pi120 ) | ( \pi119 & \pi120 ) ;
  assign w6625 = \pi000 ^ w6624 ;
  assign w6626 = ( \pi002 & \pi120 ) | ( \pi002 & ~w6625 ) | ( \pi120 & ~w6625 ) ;
  assign w6627 = ( \pi002 & \pi119 ) | ( \pi002 & w6625 ) | ( \pi119 & w6625 ) ;
  assign w6628 = \pi001 & w6627 ;
  assign w6629 = ( ~\pi000 & \pi118 ) | ( ~\pi000 & w6628 ) | ( \pi118 & w6628 ) ;
  assign w6630 = ( \pi001 & \pi002 ) | ( \pi001 & ~w6629 ) | ( \pi002 & ~w6629 ) ;
  assign w6631 = ( w6626 & w6628 ) | ( w6626 & ~w6630 ) | ( w6628 & ~w6630 ) ;
  assign w6632 = ( \pi118 & \pi119 ) | ( \pi118 & w6614 ) | ( \pi119 & w6614 ) ;
  assign w6633 = \pi119 ^ w6632 ;
  assign w6634 = \pi120 ^ w6633 ;
  assign w6635 = \pi002 ^ w6631 ;
  assign w6636 = \pi000 & ~w6631 ;
  assign w6637 = w6634 & w6636 ;
  assign w6638 = \pi001 ^ w6637 ;
  assign w6639 = ( \pi001 & w6635 ) | ( \pi001 & ~w6638 ) | ( w6635 & ~w6638 ) ;
  assign w6640 = ( w6400 & w6408 ) | ( w6400 & w6603 ) | ( w6408 & w6603 ) ;
  assign w6641 = ( w6409 & w6417 ) | ( w6409 & w6601 ) | ( w6417 & w6601 ) ;
  assign w6642 = ~\pi113 & w305 ;
  assign w6643 = \pi112 & w328 ;
  assign w6644 = ( w305 & ~w6642 ) | ( w305 & w6643 ) | ( ~w6642 & w6643 ) ;
  assign w6645 = ~\pi114 & w307 ;
  assign w6646 = w5565 | w6644 ;
  assign w6647 = ( w308 & w6644 ) | ( w308 & w6646 ) | ( w6644 & w6646 ) ;
  assign w6648 = ( w307 & ~w6645 ) | ( w307 & w6647 ) | ( ~w6645 & w6647 ) ;
  assign w6649 = \pi008 ^ w6648 ;
  assign w6650 = ( w6418 & w6591 ) | ( w6418 & w6599 ) | ( w6591 & w6599 ) ;
  assign w6651 = ~\pi098 & w1313 ;
  assign w6652 = \pi097 & w1417 ;
  assign w6653 = ( w1313 & ~w6651 ) | ( w1313 & w6652 ) | ( ~w6651 & w6652 ) ;
  assign w6654 = ~\pi099 & w1315 ;
  assign w6655 = w2966 | w6653 ;
  assign w6656 = ( w1316 & w6653 ) | ( w1316 & w6655 ) | ( w6653 & w6655 ) ;
  assign w6657 = ( w1315 & ~w6654 ) | ( w1315 & w6656 ) | ( ~w6654 & w6656 ) ;
  assign w6658 = \pi023 ^ w6657 ;
  assign w6659 = ( w6536 & w6544 ) | ( w6536 & w6545 ) | ( w6544 & w6545 ) ;
  assign w6660 = ~\pi095 & w1629 ;
  assign w6661 = \pi094 & w1722 ;
  assign w6662 = ( w1629 & ~w6660 ) | ( w1629 & w6661 ) | ( ~w6660 & w6661 ) ;
  assign w6663 = ~\pi096 & w1631 ;
  assign w6664 = w2546 | w6662 ;
  assign w6665 = ( w1632 & w6662 ) | ( w1632 & w6664 ) | ( w6662 & w6664 ) ;
  assign w6666 = ( w1631 & ~w6663 ) | ( w1631 & w6665 ) | ( ~w6663 & w6665 ) ;
  assign w6667 = \pi026 ^ w6666 ;
  assign w6668 = ( w6525 & w6533 ) | ( w6525 & w6534 ) | ( w6533 & w6534 ) ;
  assign w6669 = ( w6514 & w6522 ) | ( w6514 & w6523 ) | ( w6522 & w6523 ) ;
  assign w6670 = ( w6503 & w6511 ) | ( w6503 & w6512 ) | ( w6511 & w6512 ) ;
  assign w6671 = ( w6428 & w6489 ) | ( w6428 & w6490 ) | ( w6489 & w6490 ) ;
  assign w6672 = ~\pi080 & w3635 ;
  assign w6673 = \pi079 & w3817 ;
  assign w6674 = ( w3635 & ~w6672 ) | ( w3635 & w6673 ) | ( ~w6672 & w6673 ) ;
  assign w6675 = ~\pi081 & w3637 ;
  assign w6676 = w874 | w6674 ;
  assign w6677 = ( w3638 & w6674 ) | ( w3638 & w6676 ) | ( w6674 & w6676 ) ;
  assign w6678 = ( w3637 & ~w6675 ) | ( w3637 & w6677 ) | ( ~w6675 & w6677 ) ;
  assign w6679 = \pi041 ^ w6678 ;
  assign w6680 = ( w6429 & w6437 ) | ( w6429 & w6487 ) | ( w6437 & w6487 ) ;
  assign w6681 = ~\pi077 & w4141 ;
  assign w6682 = \pi076 & w4334 ;
  assign w6683 = ( w4141 & ~w6681 ) | ( w4141 & w6682 ) | ( ~w6681 & w6682 ) ;
  assign w6684 = ~\pi078 & w4143 ;
  assign w6685 = w665 | w6683 ;
  assign w6686 = ( w4144 & w6683 ) | ( w4144 & w6685 ) | ( w6683 & w6685 ) ;
  assign w6687 = ( w4143 & ~w6684 ) | ( w4143 & w6686 ) | ( ~w6684 & w6686 ) ;
  assign w6688 = \pi044 ^ w6687 ;
  assign w6689 = ( w6438 & w6446 ) | ( w6438 & w6485 ) | ( w6446 & w6485 ) ;
  assign w6690 = ~\pi074 & w4654 ;
  assign w6691 = \pi073 & w4876 ;
  assign w6692 = ( w4654 & ~w6690 ) | ( w4654 & w6691 ) | ( ~w6690 & w6691 ) ;
  assign w6693 = ~\pi075 & w4656 ;
  assign w6694 = w519 | w6692 ;
  assign w6695 = ( w4657 & w6692 ) | ( w4657 & w6694 ) | ( w6692 & w6694 ) ;
  assign w6696 = ( w4656 & ~w6693 ) | ( w4656 & w6695 ) | ( ~w6693 & w6695 ) ;
  assign w6697 = \pi047 ^ w6696 ;
  assign w6698 = ( w6447 & w6455 ) | ( w6447 & w6483 ) | ( w6455 & w6483 ) ;
  assign w6699 = ( w6456 & w6464 ) | ( w6456 & w6481 ) | ( w6464 & w6481 ) ;
  assign w6700 = ( \pi054 & ~\pi055 ) | ( \pi054 & \pi056 ) | ( ~\pi055 & \pi056 ) ;
  assign w6701 = ( \pi053 & \pi054 ) | ( \pi053 & w6700 ) | ( \pi054 & w6700 ) ;
  assign w6702 = w6700 ^ w6701 ;
  assign w6703 = \pi064 & w6702 ;
  assign w6704 = ( \pi066 & w6468 ) | ( \pi066 & w6703 ) | ( w6468 & w6703 ) ;
  assign w6705 = \pi065 | w6704 ;
  assign w6706 = ( w6466 & w6704 ) | ( w6466 & w6705 ) | ( w6704 & w6705 ) ;
  assign w6707 = w6703 | w6706 ;
  assign w6708 = ~w134 & w6469 ;
  assign w6709 = ( w6469 & w6707 ) | ( w6469 & ~w6708 ) | ( w6707 & ~w6708 ) ;
  assign w6710 = \pi056 ^ w6709 ;
  assign w6711 = w6476 & w6710 ;
  assign w6712 = w6476 ^ w6710 ;
  assign w6713 = ~\pi068 & w5802 ;
  assign w6714 = \pi067 & w6052 ;
  assign w6715 = ( w5802 & ~w6713 ) | ( w5802 & w6714 ) | ( ~w6713 & w6714 ) ;
  assign w6716 = ~\pi069 & w5804 ;
  assign w6717 = w221 | w6715 ;
  assign w6718 = ( w5805 & w6715 ) | ( w5805 & w6717 ) | ( w6715 & w6717 ) ;
  assign w6719 = ( w5804 & ~w6716 ) | ( w5804 & w6718 ) | ( ~w6716 & w6718 ) ;
  assign w6720 = \pi053 ^ w6719 ;
  assign w6721 = ( w6699 & w6712 ) | ( w6699 & w6720 ) | ( w6712 & w6720 ) ;
  assign w6722 = w6699 ^ w6712 ;
  assign w6723 = w6720 ^ w6722 ;
  assign w6724 = ~\pi071 & w5209 ;
  assign w6725 = \pi070 & w5433 ;
  assign w6726 = ( w5209 & ~w6724 ) | ( w5209 & w6725 ) | ( ~w6724 & w6725 ) ;
  assign w6727 = ~\pi072 & w5211 ;
  assign w6728 = w361 | w6726 ;
  assign w6729 = ( w5212 & w6726 ) | ( w5212 & w6728 ) | ( w6726 & w6728 ) ;
  assign w6730 = ( w5211 & ~w6727 ) | ( w5211 & w6729 ) | ( ~w6727 & w6729 ) ;
  assign w6731 = \pi050 ^ w6730 ;
  assign w6732 = w6698 ^ w6723 ;
  assign w6733 = w6731 ^ w6732 ;
  assign w6734 = w6689 ^ w6733 ;
  assign w6735 = w6697 ^ w6734 ;
  assign w6736 = w6680 ^ w6735 ;
  assign w6737 = w6688 ^ w6736 ;
  assign w6738 = w6671 ^ w6737 ;
  assign w6739 = w6679 ^ w6738 ;
  assign w6740 = ~\pi083 & w3178 ;
  assign w6741 = \pi082 & w3340 ;
  assign w6742 = ( w3178 & ~w6740 ) | ( w3178 & w6741 ) | ( ~w6740 & w6741 ) ;
  assign w6743 = ~\pi084 & w3180 ;
  assign w6744 = w1188 | w6742 ;
  assign w6745 = ( w3181 & w6742 ) | ( w3181 & w6744 ) | ( w6742 & w6744 ) ;
  assign w6746 = ( w3180 & ~w6743 ) | ( w3180 & w6745 ) | ( ~w6743 & w6745 ) ;
  assign w6747 = \pi038 ^ w6746 ;
  assign w6748 = w6501 ^ w6739 ;
  assign w6749 = w6747 ^ w6748 ;
  assign w6750 = ~\pi086 & w2712 ;
  assign w6751 = \pi085 & w2872 ;
  assign w6752 = ( w2712 & ~w6750 ) | ( w2712 & w6751 ) | ( ~w6750 & w6751 ) ;
  assign w6753 = ~\pi087 & w2714 ;
  assign w6754 = w1477 | w6752 ;
  assign w6755 = ( w2715 & w6752 ) | ( w2715 & w6754 ) | ( w6752 & w6754 ) ;
  assign w6756 = ( w2714 & ~w6753 ) | ( w2714 & w6755 ) | ( ~w6753 & w6755 ) ;
  assign w6757 = \pi035 ^ w6756 ;
  assign w6758 = w6670 ^ w6749 ;
  assign w6759 = w6757 ^ w6758 ;
  assign w6760 = ~\pi089 & w2310 ;
  assign w6761 = \pi088 & w2443 ;
  assign w6762 = ( w2310 & ~w6760 ) | ( w2310 & w6761 ) | ( ~w6760 & w6761 ) ;
  assign w6763 = ~\pi090 & w2312 ;
  assign w6764 = w1801 | w6762 ;
  assign w6765 = ( w2313 & w6762 ) | ( w2313 & w6764 ) | ( w6762 & w6764 ) ;
  assign w6766 = ( w2312 & ~w6763 ) | ( w2312 & w6765 ) | ( ~w6763 & w6765 ) ;
  assign w6767 = \pi032 ^ w6766 ;
  assign w6768 = ( w6669 & w6759 ) | ( w6669 & w6767 ) | ( w6759 & w6767 ) ;
  assign w6769 = w6669 ^ w6759 ;
  assign w6770 = w6767 ^ w6769 ;
  assign w6771 = ~\pi092 & w1944 ;
  assign w6772 = \pi091 & w2072 ;
  assign w6773 = ( w1944 & ~w6771 ) | ( w1944 & w6772 ) | ( ~w6771 & w6772 ) ;
  assign w6774 = ~\pi093 & w1946 ;
  assign w6775 = w2155 | w6773 ;
  assign w6776 = ( w1947 & w6773 ) | ( w1947 & w6775 ) | ( w6773 & w6775 ) ;
  assign w6777 = ( w1946 & ~w6774 ) | ( w1946 & w6776 ) | ( ~w6774 & w6776 ) ;
  assign w6778 = \pi029 ^ w6777 ;
  assign w6779 = w6668 ^ w6770 ;
  assign w6780 = w6778 ^ w6779 ;
  assign w6781 = w6659 ^ w6780 ;
  assign w6782 = w6667 ^ w6781 ;
  assign w6783 = ( w6547 & w6555 ) | ( w6547 & w6556 ) | ( w6555 & w6556 ) ;
  assign w6784 = w6782 ^ w6783 ;
  assign w6785 = w6658 ^ w6784 ;
  assign w6786 = ~\pi101 & w1044 ;
  assign w6787 = \pi100 & w1138 ;
  assign w6788 = ( w1044 & ~w6786 ) | ( w1044 & w6787 ) | ( ~w6786 & w6787 ) ;
  assign w6789 = ~\pi102 & w1046 ;
  assign w6790 = w3284 | w6788 ;
  assign w6791 = ( w1047 & w6788 ) | ( w1047 & w6790 ) | ( w6788 & w6790 ) ;
  assign w6792 = ( w1046 & ~w6789 ) | ( w1046 & w6791 ) | ( ~w6789 & w6791 ) ;
  assign w6793 = \pi020 ^ w6792 ;
  assign w6794 = ( w6558 & w6566 ) | ( w6558 & w6567 ) | ( w6566 & w6567 ) ;
  assign w6795 = w6785 ^ w6794 ;
  assign w6796 = w6793 ^ w6795 ;
  assign w6797 = ~\pi104 & w837 ;
  assign w6798 = \pi103 & w902 ;
  assign w6799 = ( w837 & ~w6797 ) | ( w837 & w6798 ) | ( ~w6797 & w6798 ) ;
  assign w6800 = ~\pi105 & w839 ;
  assign w6801 = w3905 | w6799 ;
  assign w6802 = ( w840 & w6799 ) | ( w840 & w6801 ) | ( w6799 & w6801 ) ;
  assign w6803 = ( w839 & ~w6800 ) | ( w839 & w6802 ) | ( ~w6800 & w6802 ) ;
  assign w6804 = \pi017 ^ w6803 ;
  assign w6805 = ( w6569 & w6577 ) | ( w6569 & w6578 ) | ( w6577 & w6578 ) ;
  assign w6806 = w6796 ^ w6805 ;
  assign w6807 = w6804 ^ w6806 ;
  assign w6808 = ~\pi107 & w601 ;
  assign w6809 = \pi106 & w683 ;
  assign w6810 = ( w601 & ~w6808 ) | ( w601 & w6809 ) | ( ~w6808 & w6809 ) ;
  assign w6811 = ~\pi108 & w603 ;
  assign w6812 = w4425 | w6810 ;
  assign w6813 = ( w604 & w6810 ) | ( w604 & w6812 ) | ( w6810 & w6812 ) ;
  assign w6814 = ( w603 & ~w6811 ) | ( w603 & w6813 ) | ( ~w6811 & w6813 ) ;
  assign w6815 = \pi014 ^ w6814 ;
  assign w6816 = ( w6589 & w6807 ) | ( w6589 & w6815 ) | ( w6807 & w6815 ) ;
  assign w6817 = w6589 ^ w6807 ;
  assign w6818 = w6815 ^ w6817 ;
  assign w6819 = ~\pi110 & w432 ;
  assign w6820 = \pi109 & w486 ;
  assign w6821 = ( w432 & ~w6819 ) | ( w432 & w6820 ) | ( ~w6819 & w6820 ) ;
  assign w6822 = ~\pi111 & w434 ;
  assign w6823 = w4811 | w6821 ;
  assign w6824 = ( w435 & w6821 ) | ( w435 & w6823 ) | ( w6821 & w6823 ) ;
  assign w6825 = ( w434 & ~w6822 ) | ( w434 & w6824 ) | ( ~w6822 & w6824 ) ;
  assign w6826 = \pi011 ^ w6825 ;
  assign w6827 = w6650 ^ w6818 ;
  assign w6828 = w6826 ^ w6827 ;
  assign w6829 = w6641 ^ w6828 ;
  assign w6830 = w6649 ^ w6829 ;
  assign w6831 = ~\pi116 & w189 ;
  assign w6832 = \pi115 & w229 ;
  assign w6833 = ( w189 & ~w6831 ) | ( w189 & w6832 ) | ( ~w6831 & w6832 ) ;
  assign w6834 = ~\pi117 & w191 ;
  assign w6835 = w6185 | w6833 ;
  assign w6836 = ( w192 & w6833 ) | ( w192 & w6835 ) | ( w6833 & w6835 ) ;
  assign w6837 = ( w191 & ~w6834 ) | ( w191 & w6836 ) | ( ~w6834 & w6836 ) ;
  assign w6838 = \pi005 ^ w6837 ;
  assign w6839 = w6640 ^ w6830 ;
  assign w6840 = w6838 ^ w6839 ;
  assign w6841 = ( w6399 & w6605 ) | ( w6399 & w6621 ) | ( w6605 & w6621 ) ;
  assign w6842 = w6840 ^ w6841 ;
  assign w6843 = w6639 ^ w6842 ;
  assign w6844 = ( w6640 & w6830 ) | ( w6640 & w6838 ) | ( w6830 & w6838 ) ;
  assign w6845 = ~\pi117 & w189 ;
  assign w6846 = \pi116 & w229 ;
  assign w6847 = ( w189 & ~w6845 ) | ( w189 & w6846 ) | ( ~w6845 & w6846 ) ;
  assign w6848 = ~\pi118 & w191 ;
  assign w6849 = w6206 | w6847 ;
  assign w6850 = ( w192 & w6847 ) | ( w192 & w6849 ) | ( w6847 & w6849 ) ;
  assign w6851 = ( w191 & ~w6848 ) | ( w191 & w6850 ) | ( ~w6848 & w6850 ) ;
  assign w6852 = \pi005 ^ w6851 ;
  assign w6853 = ( w6641 & w6649 ) | ( w6641 & w6828 ) | ( w6649 & w6828 ) ;
  assign w6854 = ~\pi114 & w305 ;
  assign w6855 = \pi113 & w328 ;
  assign w6856 = ( w305 & ~w6854 ) | ( w305 & w6855 ) | ( ~w6854 & w6855 ) ;
  assign w6857 = ~\pi115 & w307 ;
  assign w6858 = w5585 | w6856 ;
  assign w6859 = ( w308 & w6856 ) | ( w308 & w6858 ) | ( w6856 & w6858 ) ;
  assign w6860 = ( w307 & ~w6857 ) | ( w307 & w6859 ) | ( ~w6857 & w6859 ) ;
  assign w6861 = \pi008 ^ w6860 ;
  assign w6862 = ( w6650 & w6818 ) | ( w6650 & w6826 ) | ( w6818 & w6826 ) ;
  assign w6863 = ~\pi111 & w432 ;
  assign w6864 = \pi110 & w486 ;
  assign w6865 = ( w432 & ~w6863 ) | ( w432 & w6864 ) | ( ~w6863 & w6864 ) ;
  assign w6866 = ~\pi112 & w434 ;
  assign w6867 = w4999 | w6865 ;
  assign w6868 = ( w435 & w6865 ) | ( w435 & w6867 ) | ( w6865 & w6867 ) ;
  assign w6869 = ( w434 & ~w6866 ) | ( w434 & w6868 ) | ( ~w6866 & w6868 ) ;
  assign w6870 = \pi011 ^ w6869 ;
  assign w6871 = ~\pi108 & w601 ;
  assign w6872 = \pi107 & w683 ;
  assign w6873 = ( w601 & ~w6871 ) | ( w601 & w6872 ) | ( ~w6871 & w6872 ) ;
  assign w6874 = ~\pi109 & w603 ;
  assign w6875 = w4599 | w6873 ;
  assign w6876 = ( w604 & w6873 ) | ( w604 & w6875 ) | ( w6873 & w6875 ) ;
  assign w6877 = ( w603 & ~w6874 ) | ( w603 & w6876 ) | ( ~w6874 & w6876 ) ;
  assign w6878 = \pi014 ^ w6877 ;
  assign w6879 = ( w6796 & w6804 ) | ( w6796 & w6805 ) | ( w6804 & w6805 ) ;
  assign w6880 = ( w6658 & w6782 ) | ( w6658 & w6783 ) | ( w6782 & w6783 ) ;
  assign w6881 = ( w6659 & w6667 ) | ( w6659 & w6780 ) | ( w6667 & w6780 ) ;
  assign w6882 = ( w6668 & w6770 ) | ( w6668 & w6778 ) | ( w6770 & w6778 ) ;
  assign w6883 = ~\pi093 & w1944 ;
  assign w6884 = \pi092 & w2072 ;
  assign w6885 = ( w1944 & ~w6883 ) | ( w1944 & w6884 ) | ( ~w6883 & w6884 ) ;
  assign w6886 = ~\pi094 & w1946 ;
  assign w6887 = w2274 | w6885 ;
  assign w6888 = ( w1947 & w6885 ) | ( w1947 & w6887 ) | ( w6885 & w6887 ) ;
  assign w6889 = ( w1946 & ~w6886 ) | ( w1946 & w6888 ) | ( ~w6886 & w6888 ) ;
  assign w6890 = \pi029 ^ w6889 ;
  assign w6891 = ( w6501 & w6739 ) | ( w6501 & w6747 ) | ( w6739 & w6747 ) ;
  assign w6892 = ~\pi084 & w3178 ;
  assign w6893 = \pi083 & w3340 ;
  assign w6894 = ( w3178 & ~w6892 ) | ( w3178 & w6893 ) | ( ~w6892 & w6893 ) ;
  assign w6895 = ~\pi085 & w3180 ;
  assign w6896 = w1274 | w6894 ;
  assign w6897 = ( w3181 & w6894 ) | ( w3181 & w6896 ) | ( w6894 & w6896 ) ;
  assign w6898 = ( w3180 & ~w6895 ) | ( w3180 & w6897 ) | ( ~w6895 & w6897 ) ;
  assign w6899 = \pi038 ^ w6898 ;
  assign w6900 = ( w6671 & w6679 ) | ( w6671 & w6737 ) | ( w6679 & w6737 ) ;
  assign w6901 = ~\pi081 & w3635 ;
  assign w6902 = \pi080 & w3817 ;
  assign w6903 = ( w3635 & ~w6901 ) | ( w3635 & w6902 ) | ( ~w6901 & w6902 ) ;
  assign w6904 = ~\pi082 & w3637 ;
  assign w6905 = w1008 | w6903 ;
  assign w6906 = ( w3638 & w6903 ) | ( w3638 & w6905 ) | ( w6903 & w6905 ) ;
  assign w6907 = ( w3637 & ~w6904 ) | ( w3637 & w6906 ) | ( ~w6904 & w6906 ) ;
  assign w6908 = \pi041 ^ w6907 ;
  assign w6909 = ( w6680 & w6688 ) | ( w6680 & w6735 ) | ( w6688 & w6735 ) ;
  assign w6910 = ~\pi078 & w4141 ;
  assign w6911 = \pi077 & w4334 ;
  assign w6912 = ( w4141 & ~w6910 ) | ( w4141 & w6911 ) | ( ~w6910 & w6911 ) ;
  assign w6913 = ~\pi079 & w4143 ;
  assign w6914 = w730 | w6912 ;
  assign w6915 = ( w4144 & w6912 ) | ( w4144 & w6914 ) | ( w6912 & w6914 ) ;
  assign w6916 = ( w4143 & ~w6913 ) | ( w4143 & w6915 ) | ( ~w6913 & w6915 ) ;
  assign w6917 = \pi044 ^ w6916 ;
  assign w6918 = ( w6689 & w6697 ) | ( w6689 & w6733 ) | ( w6697 & w6733 ) ;
  assign w6919 = ~\pi075 & w4654 ;
  assign w6920 = \pi074 & w4876 ;
  assign w6921 = ( w4654 & ~w6919 ) | ( w4654 & w6920 ) | ( ~w6919 & w6920 ) ;
  assign w6922 = ~\pi076 & w4656 ;
  assign w6923 = w538 | w6921 ;
  assign w6924 = ( w4657 & w6921 ) | ( w4657 & w6923 ) | ( w6921 & w6923 ) ;
  assign w6925 = ( w4656 & ~w6922 ) | ( w4656 & w6924 ) | ( ~w6922 & w6924 ) ;
  assign w6926 = \pi047 ^ w6925 ;
  assign w6927 = ( w6698 & w6723 ) | ( w6698 & w6731 ) | ( w6723 & w6731 ) ;
  assign w6928 = ~\pi069 & w5802 ;
  assign w6929 = \pi068 & w6052 ;
  assign w6930 = ( w5802 & ~w6928 ) | ( w5802 & w6929 ) | ( ~w6928 & w6929 ) ;
  assign w6931 = ~\pi070 & w5804 ;
  assign w6932 = w271 | w6930 ;
  assign w6933 = ( w5805 & w6930 ) | ( w5805 & w6932 ) | ( w6930 & w6932 ) ;
  assign w6934 = ( w5804 & ~w6931 ) | ( w5804 & w6933 ) | ( ~w6931 & w6933 ) ;
  assign w6935 = \pi053 ^ w6934 ;
  assign w6936 = ~\pi066 & w6466 ;
  assign w6937 = \pi065 & w6702 ;
  assign w6938 = ( w6466 & ~w6936 ) | ( w6466 & w6937 ) | ( ~w6936 & w6937 ) ;
  assign w6939 = ~\pi067 & w6468 ;
  assign w6940 = w160 | w6938 ;
  assign w6941 = ( w6469 & w6938 ) | ( w6469 & w6940 ) | ( w6938 & w6940 ) ;
  assign w6942 = ( w6468 & ~w6939 ) | ( w6468 & w6941 ) | ( ~w6939 & w6941 ) ;
  assign w6943 = \pi056 ^ w6942 ;
  assign w6944 = w6711 ^ w6943 ;
  assign w6945 = \pi056 ^ \pi057 ;
  assign w6946 = \pi064 & w6945 ;
  assign w6947 = w6944 ^ w6946 ;
  assign w6948 = w6721 ^ w6947 ;
  assign w6949 = w6935 ^ w6948 ;
  assign w6950 = ~\pi072 & w5209 ;
  assign w6951 = \pi071 & w5433 ;
  assign w6952 = ( w5209 & ~w6950 ) | ( w5209 & w6951 ) | ( ~w6950 & w6951 ) ;
  assign w6953 = ~\pi073 & w5211 ;
  assign w6954 = w404 | w6952 ;
  assign w6955 = ( w5212 & w6952 ) | ( w5212 & w6954 ) | ( w6952 & w6954 ) ;
  assign w6956 = ( w5211 & ~w6953 ) | ( w5211 & w6955 ) | ( ~w6953 & w6955 ) ;
  assign w6957 = \pi050 ^ w6956 ;
  assign w6958 = w6927 ^ w6949 ;
  assign w6959 = w6957 ^ w6958 ;
  assign w6960 = w6918 ^ w6959 ;
  assign w6961 = w6926 ^ w6960 ;
  assign w6962 = w6909 ^ w6961 ;
  assign w6963 = w6917 ^ w6962 ;
  assign w6964 = w6900 ^ w6963 ;
  assign w6965 = w6908 ^ w6964 ;
  assign w6966 = w6891 ^ w6965 ;
  assign w6967 = w6899 ^ w6966 ;
  assign w6968 = ~\pi087 & w2712 ;
  assign w6969 = \pi086 & w2872 ;
  assign w6970 = ( w2712 & ~w6968 ) | ( w2712 & w6969 ) | ( ~w6968 & w6969 ) ;
  assign w6971 = ~\pi088 & w2714 ;
  assign w6972 = w1574 | w6970 ;
  assign w6973 = ( w2715 & w6970 ) | ( w2715 & w6972 ) | ( w6970 & w6972 ) ;
  assign w6974 = ( w2714 & ~w6971 ) | ( w2714 & w6973 ) | ( ~w6971 & w6973 ) ;
  assign w6975 = \pi035 ^ w6974 ;
  assign w6976 = ( w6670 & w6749 ) | ( w6670 & w6757 ) | ( w6749 & w6757 ) ;
  assign w6977 = w6967 ^ w6976 ;
  assign w6978 = w6975 ^ w6977 ;
  assign w6979 = ~\pi090 & w2310 ;
  assign w6980 = \pi089 & w2443 ;
  assign w6981 = ( w2310 & ~w6979 ) | ( w2310 & w6980 ) | ( ~w6979 & w6980 ) ;
  assign w6982 = ~\pi091 & w2312 ;
  assign w6983 = w1908 | w6981 ;
  assign w6984 = ( w2313 & w6981 ) | ( w2313 & w6983 ) | ( w6981 & w6983 ) ;
  assign w6985 = ( w2312 & ~w6982 ) | ( w2312 & w6984 ) | ( ~w6982 & w6984 ) ;
  assign w6986 = \pi032 ^ w6985 ;
  assign w6987 = w6768 ^ w6978 ;
  assign w6988 = w6986 ^ w6987 ;
  assign w6989 = w6882 ^ w6988 ;
  assign w6990 = w6890 ^ w6989 ;
  assign w6991 = ~\pi096 & w1629 ;
  assign w6992 = \pi095 & w1722 ;
  assign w6993 = ( w1629 & ~w6991 ) | ( w1629 & w6992 ) | ( ~w6991 & w6992 ) ;
  assign w6994 = ~\pi097 & w1631 ;
  assign w6995 = w2673 | w6993 ;
  assign w6996 = ( w1632 & w6993 ) | ( w1632 & w6995 ) | ( w6993 & w6995 ) ;
  assign w6997 = ( w1631 & ~w6994 ) | ( w1631 & w6996 ) | ( ~w6994 & w6996 ) ;
  assign w6998 = \pi026 ^ w6997 ;
  assign w6999 = w6881 ^ w6990 ;
  assign w7000 = w6998 ^ w6999 ;
  assign w7001 = ~\pi099 & w1313 ;
  assign w7002 = \pi098 & w1417 ;
  assign w7003 = ( w1313 & ~w7001 ) | ( w1313 & w7002 ) | ( ~w7001 & w7002 ) ;
  assign w7004 = ~\pi100 & w1315 ;
  assign w7005 = w3104 | w7003 ;
  assign w7006 = ( w1316 & w7003 ) | ( w1316 & w7005 ) | ( w7003 & w7005 ) ;
  assign w7007 = ( w1315 & ~w7004 ) | ( w1315 & w7006 ) | ( ~w7004 & w7006 ) ;
  assign w7008 = \pi023 ^ w7007 ;
  assign w7009 = w6880 ^ w7000 ;
  assign w7010 = w7008 ^ w7009 ;
  assign w7011 = ~\pi102 & w1044 ;
  assign w7012 = \pi101 & w1138 ;
  assign w7013 = ( w1044 & ~w7011 ) | ( w1044 & w7012 ) | ( ~w7011 & w7012 ) ;
  assign w7014 = ~\pi103 & w1046 ;
  assign w7015 = w3437 | w7013 ;
  assign w7016 = ( w1047 & w7013 ) | ( w1047 & w7015 ) | ( w7013 & w7015 ) ;
  assign w7017 = ( w1046 & ~w7014 ) | ( w1046 & w7016 ) | ( ~w7014 & w7016 ) ;
  assign w7018 = \pi020 ^ w7017 ;
  assign w7019 = ( w6785 & w6793 ) | ( w6785 & w6794 ) | ( w6793 & w6794 ) ;
  assign w7020 = w7010 ^ w7019 ;
  assign w7021 = w7018 ^ w7020 ;
  assign w7022 = ~\pi105 & w837 ;
  assign w7023 = \pi104 & w902 ;
  assign w7024 = ( w837 & ~w7022 ) | ( w837 & w7023 ) | ( ~w7022 & w7023 ) ;
  assign w7025 = ~\pi106 & w839 ;
  assign w7026 = w4068 | w7024 ;
  assign w7027 = ( w840 & w7024 ) | ( w840 & w7026 ) | ( w7024 & w7026 ) ;
  assign w7028 = ( w839 & ~w7025 ) | ( w839 & w7027 ) | ( ~w7025 & w7027 ) ;
  assign w7029 = \pi017 ^ w7028 ;
  assign w7030 = w6879 ^ w7021 ;
  assign w7031 = w7029 ^ w7030 ;
  assign w7032 = w6816 ^ w7031 ;
  assign w7033 = w6878 ^ w7032 ;
  assign w7034 = w6862 ^ w7033 ;
  assign w7035 = w6870 ^ w7034 ;
  assign w7036 = w6853 ^ w7035 ;
  assign w7037 = w6861 ^ w7036 ;
  assign w7038 = w6844 ^ w7037 ;
  assign w7039 = w6852 ^ w7038 ;
  assign w7040 = ( ~\pi002 & \pi120 ) | ( ~\pi002 & \pi121 ) | ( \pi120 & \pi121 ) ;
  assign w7041 = \pi000 ^ w7040 ;
  assign w7042 = ( \pi002 & \pi121 ) | ( \pi002 & ~w7041 ) | ( \pi121 & ~w7041 ) ;
  assign w7043 = ( \pi002 & \pi120 ) | ( \pi002 & w7041 ) | ( \pi120 & w7041 ) ;
  assign w7044 = \pi001 & w7043 ;
  assign w7045 = ( ~\pi000 & \pi119 ) | ( ~\pi000 & w7044 ) | ( \pi119 & w7044 ) ;
  assign w7046 = ( \pi001 & \pi002 ) | ( \pi001 & ~w7045 ) | ( \pi002 & ~w7045 ) ;
  assign w7047 = ( w7042 & w7044 ) | ( w7042 & ~w7046 ) | ( w7044 & ~w7046 ) ;
  assign w7048 = ( \pi119 & \pi120 ) | ( \pi119 & w6632 ) | ( \pi120 & w6632 ) ;
  assign w7049 = \pi120 ^ w7048 ;
  assign w7050 = \pi121 ^ w7049 ;
  assign w7051 = \pi002 ^ w7047 ;
  assign w7052 = \pi000 & ~w7047 ;
  assign w7053 = w7050 & w7052 ;
  assign w7054 = \pi001 ^ w7053 ;
  assign w7055 = ( \pi001 & w7051 ) | ( \pi001 & ~w7054 ) | ( w7051 & ~w7054 ) ;
  assign w7056 = ( w6639 & w6840 ) | ( w6639 & w6841 ) | ( w6840 & w6841 ) ;
  assign w7057 = w7039 ^ w7056 ;
  assign w7058 = w7055 ^ w7057 ;
  assign w7059 = ( ~\pi002 & \pi121 ) | ( ~\pi002 & \pi122 ) | ( \pi121 & \pi122 ) ;
  assign w7060 = \pi000 ^ w7059 ;
  assign w7061 = ( \pi002 & \pi122 ) | ( \pi002 & ~w7060 ) | ( \pi122 & ~w7060 ) ;
  assign w7062 = ( \pi002 & \pi121 ) | ( \pi002 & w7060 ) | ( \pi121 & w7060 ) ;
  assign w7063 = \pi001 & w7062 ;
  assign w7064 = ( ~\pi000 & \pi120 ) | ( ~\pi000 & w7063 ) | ( \pi120 & w7063 ) ;
  assign w7065 = ( \pi001 & \pi002 ) | ( \pi001 & ~w7064 ) | ( \pi002 & ~w7064 ) ;
  assign w7066 = ( w7061 & w7063 ) | ( w7061 & ~w7065 ) | ( w7063 & ~w7065 ) ;
  assign w7067 = ( \pi120 & \pi121 ) | ( \pi120 & w7048 ) | ( \pi121 & w7048 ) ;
  assign w7068 = \pi121 ^ w7067 ;
  assign w7069 = \pi122 ^ w7068 ;
  assign w7070 = \pi002 ^ w7066 ;
  assign w7071 = \pi000 & ~w7066 ;
  assign w7072 = w7069 & w7071 ;
  assign w7073 = \pi001 ^ w7072 ;
  assign w7074 = ( \pi001 & w7070 ) | ( \pi001 & ~w7073 ) | ( w7070 & ~w7073 ) ;
  assign w7075 = ( w6844 & w6852 ) | ( w6844 & w7037 ) | ( w6852 & w7037 ) ;
  assign w7076 = ~\pi118 & w189 ;
  assign w7077 = \pi117 & w229 ;
  assign w7078 = ( w189 & ~w7076 ) | ( w189 & w7077 ) | ( ~w7076 & w7077 ) ;
  assign w7079 = ~\pi119 & w191 ;
  assign w7080 = w6616 | w7078 ;
  assign w7081 = ( w192 & w7078 ) | ( w192 & w7080 ) | ( w7078 & w7080 ) ;
  assign w7082 = ( w191 & ~w7079 ) | ( w191 & w7081 ) | ( ~w7079 & w7081 ) ;
  assign w7083 = \pi005 ^ w7082 ;
  assign w7084 = ( w6853 & w6861 ) | ( w6853 & w7035 ) | ( w6861 & w7035 ) ;
  assign w7085 = ~\pi115 & w305 ;
  assign w7086 = \pi114 & w328 ;
  assign w7087 = ( w305 & ~w7085 ) | ( w305 & w7086 ) | ( ~w7085 & w7086 ) ;
  assign w7088 = ~\pi116 & w307 ;
  assign w7089 = w5976 | w7087 ;
  assign w7090 = ( w308 & w7087 ) | ( w308 & w7089 ) | ( w7087 & w7089 ) ;
  assign w7091 = ( w307 & ~w7088 ) | ( w307 & w7090 ) | ( ~w7088 & w7090 ) ;
  assign w7092 = \pi008 ^ w7091 ;
  assign w7093 = ( w6862 & w6870 ) | ( w6862 & w7033 ) | ( w6870 & w7033 ) ;
  assign w7094 = ~\pi112 & w432 ;
  assign w7095 = \pi111 & w486 ;
  assign w7096 = ( w432 & ~w7094 ) | ( w432 & w7095 ) | ( ~w7094 & w7095 ) ;
  assign w7097 = ~\pi113 & w434 ;
  assign w7098 = w5366 | w7096 ;
  assign w7099 = ( w435 & w7096 ) | ( w435 & w7098 ) | ( w7096 & w7098 ) ;
  assign w7100 = ( w434 & ~w7097 ) | ( w434 & w7099 ) | ( ~w7097 & w7099 ) ;
  assign w7101 = \pi011 ^ w7100 ;
  assign w7102 = ( w6816 & w6878 ) | ( w6816 & w7031 ) | ( w6878 & w7031 ) ;
  assign w7103 = ( w6879 & w7021 ) | ( w6879 & w7029 ) | ( w7021 & w7029 ) ;
  assign w7104 = ( w6882 & w6890 ) | ( w6882 & w6988 ) | ( w6890 & w6988 ) ;
  assign w7105 = ( w6768 & w6978 ) | ( w6768 & w6986 ) | ( w6978 & w6986 ) ;
  assign w7106 = ( w6900 & w6908 ) | ( w6900 & w6963 ) | ( w6908 & w6963 ) ;
  assign w7107 = ( w6918 & w6926 ) | ( w6918 & w6959 ) | ( w6926 & w6959 ) ;
  assign w7108 = ~\pi073 & w5209 ;
  assign w7109 = \pi072 & w5433 ;
  assign w7110 = ( w5209 & ~w7108 ) | ( w5209 & w7109 ) | ( ~w7108 & w7109 ) ;
  assign w7111 = ~\pi074 & w5211 ;
  assign w7112 = w465 | w7110 ;
  assign w7113 = ( w5212 & w7110 ) | ( w5212 & w7112 ) | ( w7110 & w7112 ) ;
  assign w7114 = ( w5211 & ~w7111 ) | ( w5211 & w7113 ) | ( ~w7111 & w7113 ) ;
  assign w7115 = \pi050 ^ w7114 ;
  assign w7116 = ( w6721 & w6935 ) | ( w6721 & w6947 ) | ( w6935 & w6947 ) ;
  assign w7117 = ~\pi070 & w5802 ;
  assign w7118 = \pi069 & w6052 ;
  assign w7119 = ( w5802 & ~w7117 ) | ( w5802 & w7118 ) | ( ~w7117 & w7118 ) ;
  assign w7120 = ~\pi071 & w5804 ;
  assign w7121 = w290 | w7119 ;
  assign w7122 = ( w5805 & w7119 ) | ( w5805 & w7121 ) | ( w7119 & w7121 ) ;
  assign w7123 = ( w5804 & ~w7120 ) | ( w5804 & w7122 ) | ( ~w7120 & w7122 ) ;
  assign w7124 = \pi053 ^ w7123 ;
  assign w7125 = ( w6711 & w6943 ) | ( w6711 & w6946 ) | ( w6943 & w6946 ) ;
  assign w7126 = ~\pi067 & w6466 ;
  assign w7127 = \pi066 & w6702 ;
  assign w7128 = ( w6466 & ~w7126 ) | ( w6466 & w7127 ) | ( ~w7126 & w7127 ) ;
  assign w7129 = ~\pi068 & w6468 ;
  assign w7130 = w182 | w7128 ;
  assign w7131 = ( w6469 & w7128 ) | ( w6469 & w7130 ) | ( w7128 & w7130 ) ;
  assign w7132 = ( w6468 & ~w7129 ) | ( w6468 & w7131 ) | ( ~w7129 & w7131 ) ;
  assign w7133 = \pi056 ^ w7132 ;
  assign w7134 = ( \pi056 & \pi057 ) | ( \pi056 & \pi058 ) | ( \pi057 & \pi058 ) ;
  assign w7135 = \pi058 ^ w7134 ;
  assign w7136 = \pi058 ^ \pi059 ;
  assign w7137 = w6945 & ~w7136 ;
  assign w7138 = w6945 & w7136 ;
  assign w7139 = ( \pi056 & \pi057 ) | ( \pi056 & ~\pi059 ) | ( \pi057 & ~\pi059 ) ;
  assign w7140 = \pi059 & ~\pi064 ;
  assign w7141 = ~\pi065 & w7140 ;
  assign w7142 = ( \pi056 & \pi057 ) | ( \pi056 & ~w7141 ) | ( \pi057 & ~w7141 ) ;
  assign w7143 = ( \pi058 & \pi059 ) | ( \pi058 & ~w7142 ) | ( \pi059 & ~w7142 ) ;
  assign w7144 = ( \pi058 & ~w7140 ) | ( \pi058 & w7142 ) | ( ~w7140 & w7142 ) ;
  assign w7145 = ( w7139 & w7143 ) | ( w7139 & ~w7144 ) | ( w7143 & ~w7144 ) ;
  assign w7146 = ( \pi056 & \pi057 ) | ( \pi056 & \pi065 ) | ( \pi057 & \pi065 ) ;
  assign w7147 = \pi056 & \pi057 ;
  assign w7148 = \pi064 ^ w7147 ;
  assign w7149 = ( \pi058 & w7147 ) | ( \pi058 & w7148 ) | ( w7147 & w7148 ) ;
  assign w7150 = w7146 ^ w7149 ;
  assign w7151 = w7125 ^ w7133 ;
  assign w7152 = w7150 ^ w7151 ;
  assign w7153 = w7116 ^ w7152 ;
  assign w7154 = w7124 ^ w7153 ;
  assign w7155 = ( w6927 & w6949 ) | ( w6927 & w6957 ) | ( w6949 & w6957 ) ;
  assign w7156 = w7154 ^ w7155 ;
  assign w7157 = w7115 ^ w7156 ;
  assign w7158 = ~\pi076 & w4654 ;
  assign w7159 = \pi075 & w4876 ;
  assign w7160 = ( w4654 & ~w7158 ) | ( w4654 & w7159 ) | ( ~w7158 & w7159 ) ;
  assign w7161 = ~\pi077 & w4656 ;
  assign w7162 = w644 | w7160 ;
  assign w7163 = ( w4657 & w7160 ) | ( w4657 & w7162 ) | ( w7160 & w7162 ) ;
  assign w7164 = ( w4656 & ~w7161 ) | ( w4656 & w7163 ) | ( ~w7161 & w7163 ) ;
  assign w7165 = \pi047 ^ w7164 ;
  assign w7166 = ( w7107 & w7157 ) | ( w7107 & w7165 ) | ( w7157 & w7165 ) ;
  assign w7167 = w7107 ^ w7157 ;
  assign w7168 = w7165 ^ w7167 ;
  assign w7169 = ~\pi079 & w4141 ;
  assign w7170 = \pi078 & w4334 ;
  assign w7171 = ( w4141 & ~w7169 ) | ( w4141 & w7170 ) | ( ~w7169 & w7170 ) ;
  assign w7172 = ~\pi080 & w4143 ;
  assign w7173 = w794 | w7171 ;
  assign w7174 = ( w4144 & w7171 ) | ( w4144 & w7173 ) | ( w7171 & w7173 ) ;
  assign w7175 = ( w4143 & ~w7172 ) | ( w4143 & w7174 ) | ( ~w7172 & w7174 ) ;
  assign w7176 = \pi044 ^ w7175 ;
  assign w7177 = ( w6909 & w6917 ) | ( w6909 & w6961 ) | ( w6917 & w6961 ) ;
  assign w7178 = w7168 ^ w7177 ;
  assign w7179 = w7176 ^ w7178 ;
  assign w7180 = ~\pi082 & w3635 ;
  assign w7181 = \pi081 & w3817 ;
  assign w7182 = ( w3635 & ~w7180 ) | ( w3635 & w7181 ) | ( ~w7180 & w7181 ) ;
  assign w7183 = ~\pi083 & w3637 ;
  assign w7184 = w1099 | w7182 ;
  assign w7185 = ( w3638 & w7182 ) | ( w3638 & w7184 ) | ( w7182 & w7184 ) ;
  assign w7186 = ( w3637 & ~w7183 ) | ( w3637 & w7185 ) | ( ~w7183 & w7185 ) ;
  assign w7187 = \pi041 ^ w7186 ;
  assign w7188 = ( w7106 & w7179 ) | ( w7106 & w7187 ) | ( w7179 & w7187 ) ;
  assign w7189 = w7106 ^ w7179 ;
  assign w7190 = w7187 ^ w7189 ;
  assign w7191 = ~\pi085 & w3178 ;
  assign w7192 = \pi084 & w3340 ;
  assign w7193 = ( w3178 & ~w7191 ) | ( w3178 & w7192 ) | ( ~w7191 & w7192 ) ;
  assign w7194 = ~\pi086 & w3180 ;
  assign w7195 = w1379 | w7193 ;
  assign w7196 = ( w3181 & w7193 ) | ( w3181 & w7195 ) | ( w7193 & w7195 ) ;
  assign w7197 = ( w3180 & ~w7194 ) | ( w3180 & w7196 ) | ( ~w7194 & w7196 ) ;
  assign w7198 = \pi038 ^ w7197 ;
  assign w7199 = ( w6891 & w6899 ) | ( w6891 & w6965 ) | ( w6899 & w6965 ) ;
  assign w7200 = w7190 ^ w7199 ;
  assign w7201 = w7198 ^ w7200 ;
  assign w7202 = ~\pi088 & w2712 ;
  assign w7203 = \pi087 & w2872 ;
  assign w7204 = ( w2712 & ~w7202 ) | ( w2712 & w7203 ) | ( ~w7202 & w7203 ) ;
  assign w7205 = ~\pi089 & w2714 ;
  assign w7206 = w1595 | w7204 ;
  assign w7207 = ( w2715 & w7204 ) | ( w2715 & w7206 ) | ( w7204 & w7206 ) ;
  assign w7208 = ( w2714 & ~w7205 ) | ( w2714 & w7207 ) | ( ~w7205 & w7207 ) ;
  assign w7209 = \pi035 ^ w7208 ;
  assign w7210 = ( w6967 & w6975 ) | ( w6967 & w6976 ) | ( w6975 & w6976 ) ;
  assign w7211 = w7201 ^ w7210 ;
  assign w7212 = w7209 ^ w7211 ;
  assign w7213 = ~\pi091 & w2310 ;
  assign w7214 = \pi090 & w2443 ;
  assign w7215 = ( w2310 & ~w7213 ) | ( w2310 & w7214 ) | ( ~w7213 & w7214 ) ;
  assign w7216 = ~\pi092 & w2312 ;
  assign w7217 = w2033 | w7215 ;
  assign w7218 = ( w2313 & w7215 ) | ( w2313 & w7217 ) | ( w7215 & w7217 ) ;
  assign w7219 = ( w2312 & ~w7216 ) | ( w2312 & w7218 ) | ( ~w7216 & w7218 ) ;
  assign w7220 = \pi032 ^ w7219 ;
  assign w7221 = w7105 ^ w7212 ;
  assign w7222 = w7220 ^ w7221 ;
  assign w7223 = ~\pi094 & w1944 ;
  assign w7224 = \pi093 & w2072 ;
  assign w7225 = ( w1944 & ~w7223 ) | ( w1944 & w7224 ) | ( ~w7223 & w7224 ) ;
  assign w7226 = ~\pi095 & w1946 ;
  assign w7227 = w2409 | w7225 ;
  assign w7228 = ( w1947 & w7225 ) | ( w1947 & w7227 ) | ( w7225 & w7227 ) ;
  assign w7229 = ( w1946 & ~w7226 ) | ( w1946 & w7228 ) | ( ~w7226 & w7228 ) ;
  assign w7230 = \pi029 ^ w7229 ;
  assign w7231 = w7104 ^ w7222 ;
  assign w7232 = w7230 ^ w7231 ;
  assign w7233 = ~\pi097 & w1629 ;
  assign w7234 = \pi096 & w1722 ;
  assign w7235 = ( w1629 & ~w7233 ) | ( w1629 & w7234 ) | ( ~w7233 & w7234 ) ;
  assign w7236 = ~\pi098 & w1631 ;
  assign w7237 = w2824 | w7235 ;
  assign w7238 = ( w1632 & w7235 ) | ( w1632 & w7237 ) | ( w7235 & w7237 ) ;
  assign w7239 = ( w1631 & ~w7236 ) | ( w1631 & w7238 ) | ( ~w7236 & w7238 ) ;
  assign w7240 = \pi026 ^ w7239 ;
  assign w7241 = ( w6881 & w6990 ) | ( w6881 & w6998 ) | ( w6990 & w6998 ) ;
  assign w7242 = w7232 ^ w7241 ;
  assign w7243 = w7240 ^ w7242 ;
  assign w7244 = ~\pi100 & w1313 ;
  assign w7245 = \pi099 & w1417 ;
  assign w7246 = ( w1313 & ~w7244 ) | ( w1313 & w7245 ) | ( ~w7244 & w7245 ) ;
  assign w7247 = ~\pi101 & w1315 ;
  assign w7248 = w3264 | w7246 ;
  assign w7249 = ( w1316 & w7246 ) | ( w1316 & w7248 ) | ( w7246 & w7248 ) ;
  assign w7250 = ( w1315 & ~w7247 ) | ( w1315 & w7249 ) | ( ~w7247 & w7249 ) ;
  assign w7251 = \pi023 ^ w7250 ;
  assign w7252 = ( w6880 & w7000 ) | ( w6880 & w7008 ) | ( w7000 & w7008 ) ;
  assign w7253 = w7243 ^ w7252 ;
  assign w7254 = w7251 ^ w7253 ;
  assign w7255 = ~\pi103 & w1044 ;
  assign w7256 = \pi102 & w1138 ;
  assign w7257 = ( w1044 & ~w7255 ) | ( w1044 & w7256 ) | ( ~w7255 & w7256 ) ;
  assign w7258 = ~\pi104 & w1046 ;
  assign w7259 = w3740 | w7257 ;
  assign w7260 = ( w1047 & w7257 ) | ( w1047 & w7259 ) | ( w7257 & w7259 ) ;
  assign w7261 = ( w1046 & ~w7258 ) | ( w1046 & w7260 ) | ( ~w7258 & w7260 ) ;
  assign w7262 = \pi020 ^ w7261 ;
  assign w7263 = ( w7010 & w7018 ) | ( w7010 & w7019 ) | ( w7018 & w7019 ) ;
  assign w7264 = w7254 ^ w7263 ;
  assign w7265 = w7262 ^ w7264 ;
  assign w7266 = ~\pi106 & w837 ;
  assign w7267 = \pi105 & w902 ;
  assign w7268 = ( w837 & ~w7266 ) | ( w837 & w7267 ) | ( ~w7266 & w7267 ) ;
  assign w7269 = ~\pi107 & w839 ;
  assign w7270 = w4087 | w7268 ;
  assign w7271 = ( w840 & w7268 ) | ( w840 & w7270 ) | ( w7268 & w7270 ) ;
  assign w7272 = ( w839 & ~w7269 ) | ( w839 & w7271 ) | ( ~w7269 & w7271 ) ;
  assign w7273 = \pi017 ^ w7272 ;
  assign w7274 = ( w7103 & w7265 ) | ( w7103 & w7273 ) | ( w7265 & w7273 ) ;
  assign w7275 = w7103 ^ w7265 ;
  assign w7276 = w7273 ^ w7275 ;
  assign w7277 = ~\pi109 & w601 ;
  assign w7278 = \pi108 & w683 ;
  assign w7279 = ( w601 & ~w7277 ) | ( w601 & w7278 ) | ( ~w7277 & w7278 ) ;
  assign w7280 = ~\pi110 & w603 ;
  assign w7281 = w4792 | w7279 ;
  assign w7282 = ( w604 & w7279 ) | ( w604 & w7281 ) | ( w7279 & w7281 ) ;
  assign w7283 = ( w603 & ~w7280 ) | ( w603 & w7282 ) | ( ~w7280 & w7282 ) ;
  assign w7284 = \pi014 ^ w7283 ;
  assign w7285 = w7102 ^ w7276 ;
  assign w7286 = w7284 ^ w7285 ;
  assign w7287 = w7093 ^ w7286 ;
  assign w7288 = w7101 ^ w7287 ;
  assign w7289 = w7084 ^ w7288 ;
  assign w7290 = w7092 ^ w7289 ;
  assign w7291 = w7075 ^ w7290 ;
  assign w7292 = w7083 ^ w7291 ;
  assign w7293 = ( w7039 & w7055 ) | ( w7039 & w7056 ) | ( w7055 & w7056 ) ;
  assign w7294 = w7292 ^ w7293 ;
  assign w7295 = w7074 ^ w7294 ;
  assign w7296 = ( w7074 & w7292 ) | ( w7074 & w7293 ) | ( w7292 & w7293 ) ;
  assign w7297 = ( w7075 & w7083 ) | ( w7075 & w7290 ) | ( w7083 & w7290 ) ;
  assign w7298 = ( w7084 & w7092 ) | ( w7084 & w7288 ) | ( w7092 & w7288 ) ;
  assign w7299 = ~\pi116 & w305 ;
  assign w7300 = \pi115 & w328 ;
  assign w7301 = ( w305 & ~w7299 ) | ( w305 & w7300 ) | ( ~w7299 & w7300 ) ;
  assign w7302 = ~\pi117 & w307 ;
  assign w7303 = w6185 | w7301 ;
  assign w7304 = ( w308 & w7301 ) | ( w308 & w7303 ) | ( w7301 & w7303 ) ;
  assign w7305 = ( w307 & ~w7302 ) | ( w307 & w7304 ) | ( ~w7302 & w7304 ) ;
  assign w7306 = \pi008 ^ w7305 ;
  assign w7307 = ( w7093 & w7101 ) | ( w7093 & w7286 ) | ( w7101 & w7286 ) ;
  assign w7308 = ~\pi113 & w432 ;
  assign w7309 = \pi112 & w486 ;
  assign w7310 = ( w432 & ~w7308 ) | ( w432 & w7309 ) | ( ~w7308 & w7309 ) ;
  assign w7311 = ~\pi114 & w434 ;
  assign w7312 = w5565 | w7310 ;
  assign w7313 = ( w435 & w7310 ) | ( w435 & w7312 ) | ( w7310 & w7312 ) ;
  assign w7314 = ( w434 & ~w7311 ) | ( w434 & w7313 ) | ( ~w7311 & w7313 ) ;
  assign w7315 = \pi011 ^ w7314 ;
  assign w7316 = ( w7102 & w7276 ) | ( w7102 & w7284 ) | ( w7276 & w7284 ) ;
  assign w7317 = ( w7254 & w7262 ) | ( w7254 & w7263 ) | ( w7262 & w7263 ) ;
  assign w7318 = ~\pi098 & w1629 ;
  assign w7319 = \pi097 & w1722 ;
  assign w7320 = ( w1629 & ~w7318 ) | ( w1629 & w7319 ) | ( ~w7318 & w7319 ) ;
  assign w7321 = ~\pi099 & w1631 ;
  assign w7322 = w2966 | w7320 ;
  assign w7323 = ( w1632 & w7320 ) | ( w1632 & w7322 ) | ( w7320 & w7322 ) ;
  assign w7324 = ( w1631 & ~w7321 ) | ( w1631 & w7323 ) | ( ~w7321 & w7323 ) ;
  assign w7325 = \pi026 ^ w7324 ;
  assign w7326 = ( w7104 & w7222 ) | ( w7104 & w7230 ) | ( w7222 & w7230 ) ;
  assign w7327 = ( w7105 & w7212 ) | ( w7105 & w7220 ) | ( w7212 & w7220 ) ;
  assign w7328 = ( w7190 & w7198 ) | ( w7190 & w7199 ) | ( w7198 & w7199 ) ;
  assign w7329 = ( w7168 & w7176 ) | ( w7168 & w7177 ) | ( w7176 & w7177 ) ;
  assign w7330 = ~\pi080 & w4141 ;
  assign w7331 = \pi079 & w4334 ;
  assign w7332 = ( w4141 & ~w7330 ) | ( w4141 & w7331 ) | ( ~w7330 & w7331 ) ;
  assign w7333 = ~\pi081 & w4143 ;
  assign w7334 = w874 | w7332 ;
  assign w7335 = ( w4144 & w7332 ) | ( w4144 & w7334 ) | ( w7332 & w7334 ) ;
  assign w7336 = ( w4143 & ~w7333 ) | ( w4143 & w7335 ) | ( ~w7333 & w7335 ) ;
  assign w7337 = \pi044 ^ w7336 ;
  assign w7338 = ~\pi077 & w4654 ;
  assign w7339 = \pi076 & w4876 ;
  assign w7340 = ( w4654 & ~w7338 ) | ( w4654 & w7339 ) | ( ~w7338 & w7339 ) ;
  assign w7341 = ~\pi078 & w4656 ;
  assign w7342 = w665 | w7340 ;
  assign w7343 = ( w4657 & w7340 ) | ( w4657 & w7342 ) | ( w7340 & w7342 ) ;
  assign w7344 = ( w4656 & ~w7341 ) | ( w4656 & w7343 ) | ( ~w7341 & w7343 ) ;
  assign w7345 = \pi047 ^ w7344 ;
  assign w7346 = ( w7115 & w7154 ) | ( w7115 & w7155 ) | ( w7154 & w7155 ) ;
  assign w7347 = ~\pi074 & w5209 ;
  assign w7348 = \pi073 & w5433 ;
  assign w7349 = ( w5209 & ~w7347 ) | ( w5209 & w7348 ) | ( ~w7347 & w7348 ) ;
  assign w7350 = ~\pi075 & w5211 ;
  assign w7351 = w519 | w7349 ;
  assign w7352 = ( w5212 & w7349 ) | ( w5212 & w7351 ) | ( w7349 & w7351 ) ;
  assign w7353 = ( w5211 & ~w7350 ) | ( w5211 & w7352 ) | ( ~w7350 & w7352 ) ;
  assign w7354 = \pi050 ^ w7353 ;
  assign w7355 = ( w7116 & w7124 ) | ( w7116 & w7152 ) | ( w7124 & w7152 ) ;
  assign w7356 = ( w7125 & w7133 ) | ( w7125 & w7150 ) | ( w7133 & w7150 ) ;
  assign w7357 = ( \pi057 & ~\pi058 ) | ( \pi057 & \pi059 ) | ( ~\pi058 & \pi059 ) ;
  assign w7358 = ( \pi056 & \pi057 ) | ( \pi056 & w7357 ) | ( \pi057 & w7357 ) ;
  assign w7359 = w7357 ^ w7358 ;
  assign w7360 = \pi064 & w7359 ;
  assign w7361 = ( \pi066 & w7137 ) | ( \pi066 & w7360 ) | ( w7137 & w7360 ) ;
  assign w7362 = \pi065 | w7361 ;
  assign w7363 = ( w7135 & w7361 ) | ( w7135 & w7362 ) | ( w7361 & w7362 ) ;
  assign w7364 = w7360 | w7363 ;
  assign w7365 = ~w134 & w7138 ;
  assign w7366 = ( w7138 & w7364 ) | ( w7138 & ~w7365 ) | ( w7364 & ~w7365 ) ;
  assign w7367 = \pi059 ^ w7366 ;
  assign w7368 = w7145 & w7367 ;
  assign w7369 = w7145 ^ w7367 ;
  assign w7370 = ~\pi068 & w6466 ;
  assign w7371 = \pi067 & w6702 ;
  assign w7372 = ( w6466 & ~w7370 ) | ( w6466 & w7371 ) | ( ~w7370 & w7371 ) ;
  assign w7373 = ~\pi069 & w6468 ;
  assign w7374 = w221 | w7372 ;
  assign w7375 = ( w6469 & w7372 ) | ( w6469 & w7374 ) | ( w7372 & w7374 ) ;
  assign w7376 = ( w6468 & ~w7373 ) | ( w6468 & w7375 ) | ( ~w7373 & w7375 ) ;
  assign w7377 = \pi056 ^ w7376 ;
  assign w7378 = ( w7356 & w7369 ) | ( w7356 & w7377 ) | ( w7369 & w7377 ) ;
  assign w7379 = w7356 ^ w7369 ;
  assign w7380 = w7377 ^ w7379 ;
  assign w7381 = ~\pi071 & w5802 ;
  assign w7382 = \pi070 & w6052 ;
  assign w7383 = ( w5802 & ~w7381 ) | ( w5802 & w7382 ) | ( ~w7381 & w7382 ) ;
  assign w7384 = ~\pi072 & w5804 ;
  assign w7385 = w361 | w7383 ;
  assign w7386 = ( w5805 & w7383 ) | ( w5805 & w7385 ) | ( w7383 & w7385 ) ;
  assign w7387 = ( w5804 & ~w7384 ) | ( w5804 & w7386 ) | ( ~w7384 & w7386 ) ;
  assign w7388 = \pi053 ^ w7387 ;
  assign w7389 = w7355 ^ w7380 ;
  assign w7390 = w7388 ^ w7389 ;
  assign w7391 = w7346 ^ w7390 ;
  assign w7392 = w7354 ^ w7391 ;
  assign w7393 = w7166 ^ w7392 ;
  assign w7394 = w7345 ^ w7393 ;
  assign w7395 = w7329 ^ w7394 ;
  assign w7396 = w7337 ^ w7395 ;
  assign w7397 = ~\pi083 & w3635 ;
  assign w7398 = \pi082 & w3817 ;
  assign w7399 = ( w3635 & ~w7397 ) | ( w3635 & w7398 ) | ( ~w7397 & w7398 ) ;
  assign w7400 = ~\pi084 & w3637 ;
  assign w7401 = w1188 | w7399 ;
  assign w7402 = ( w3638 & w7399 ) | ( w3638 & w7401 ) | ( w7399 & w7401 ) ;
  assign w7403 = ( w3637 & ~w7400 ) | ( w3637 & w7402 ) | ( ~w7400 & w7402 ) ;
  assign w7404 = \pi041 ^ w7403 ;
  assign w7405 = w7188 ^ w7396 ;
  assign w7406 = w7404 ^ w7405 ;
  assign w7407 = ~\pi086 & w3178 ;
  assign w7408 = \pi085 & w3340 ;
  assign w7409 = ( w3178 & ~w7407 ) | ( w3178 & w7408 ) | ( ~w7407 & w7408 ) ;
  assign w7410 = ~\pi087 & w3180 ;
  assign w7411 = w1477 | w7409 ;
  assign w7412 = ( w3181 & w7409 ) | ( w3181 & w7411 ) | ( w7409 & w7411 ) ;
  assign w7413 = ( w3180 & ~w7410 ) | ( w3180 & w7412 ) | ( ~w7410 & w7412 ) ;
  assign w7414 = \pi038 ^ w7413 ;
  assign w7415 = w7328 ^ w7406 ;
  assign w7416 = w7414 ^ w7415 ;
  assign w7417 = ~\pi089 & w2712 ;
  assign w7418 = \pi088 & w2872 ;
  assign w7419 = ( w2712 & ~w7417 ) | ( w2712 & w7418 ) | ( ~w7417 & w7418 ) ;
  assign w7420 = ~\pi090 & w2714 ;
  assign w7421 = w1801 | w7419 ;
  assign w7422 = ( w2715 & w7419 ) | ( w2715 & w7421 ) | ( w7419 & w7421 ) ;
  assign w7423 = ( w2714 & ~w7420 ) | ( w2714 & w7422 ) | ( ~w7420 & w7422 ) ;
  assign w7424 = \pi035 ^ w7423 ;
  assign w7425 = ( w7201 & w7209 ) | ( w7201 & w7210 ) | ( w7209 & w7210 ) ;
  assign w7426 = w7416 ^ w7425 ;
  assign w7427 = w7424 ^ w7426 ;
  assign w7428 = ~\pi092 & w2310 ;
  assign w7429 = \pi091 & w2443 ;
  assign w7430 = ( w2310 & ~w7428 ) | ( w2310 & w7429 ) | ( ~w7428 & w7429 ) ;
  assign w7431 = ~\pi093 & w2312 ;
  assign w7432 = w2155 | w7430 ;
  assign w7433 = ( w2313 & w7430 ) | ( w2313 & w7432 ) | ( w7430 & w7432 ) ;
  assign w7434 = ( w2312 & ~w7431 ) | ( w2312 & w7433 ) | ( ~w7431 & w7433 ) ;
  assign w7435 = \pi032 ^ w7434 ;
  assign w7436 = ( w7327 & w7427 ) | ( w7327 & w7435 ) | ( w7427 & w7435 ) ;
  assign w7437 = w7327 ^ w7427 ;
  assign w7438 = w7435 ^ w7437 ;
  assign w7439 = ~\pi095 & w1944 ;
  assign w7440 = \pi094 & w2072 ;
  assign w7441 = ( w1944 & ~w7439 ) | ( w1944 & w7440 ) | ( ~w7439 & w7440 ) ;
  assign w7442 = ~\pi096 & w1946 ;
  assign w7443 = w2546 | w7441 ;
  assign w7444 = ( w1947 & w7441 ) | ( w1947 & w7443 ) | ( w7441 & w7443 ) ;
  assign w7445 = ( w1946 & ~w7442 ) | ( w1946 & w7444 ) | ( ~w7442 & w7444 ) ;
  assign w7446 = \pi029 ^ w7445 ;
  assign w7447 = w7326 ^ w7438 ;
  assign w7448 = w7446 ^ w7447 ;
  assign w7449 = ( w7232 & w7240 ) | ( w7232 & w7241 ) | ( w7240 & w7241 ) ;
  assign w7450 = w7448 ^ w7449 ;
  assign w7451 = w7325 ^ w7450 ;
  assign w7452 = ~\pi101 & w1313 ;
  assign w7453 = \pi100 & w1417 ;
  assign w7454 = ( w1313 & ~w7452 ) | ( w1313 & w7453 ) | ( ~w7452 & w7453 ) ;
  assign w7455 = ~\pi102 & w1315 ;
  assign w7456 = w3284 | w7454 ;
  assign w7457 = ( w1316 & w7454 ) | ( w1316 & w7456 ) | ( w7454 & w7456 ) ;
  assign w7458 = ( w1315 & ~w7455 ) | ( w1315 & w7457 ) | ( ~w7455 & w7457 ) ;
  assign w7459 = \pi023 ^ w7458 ;
  assign w7460 = ( w7243 & w7251 ) | ( w7243 & w7252 ) | ( w7251 & w7252 ) ;
  assign w7461 = w7451 ^ w7460 ;
  assign w7462 = w7459 ^ w7461 ;
  assign w7463 = ~\pi104 & w1044 ;
  assign w7464 = \pi103 & w1138 ;
  assign w7465 = ( w1044 & ~w7463 ) | ( w1044 & w7464 ) | ( ~w7463 & w7464 ) ;
  assign w7466 = ~\pi105 & w1046 ;
  assign w7467 = w3905 | w7465 ;
  assign w7468 = ( w1047 & w7465 ) | ( w1047 & w7467 ) | ( w7465 & w7467 ) ;
  assign w7469 = ( w1046 & ~w7466 ) | ( w1046 & w7468 ) | ( ~w7466 & w7468 ) ;
  assign w7470 = \pi020 ^ w7469 ;
  assign w7471 = ( w7317 & w7462 ) | ( w7317 & w7470 ) | ( w7462 & w7470 ) ;
  assign w7472 = w7317 ^ w7462 ;
  assign w7473 = w7470 ^ w7472 ;
  assign w7474 = ~\pi107 & w837 ;
  assign w7475 = \pi106 & w902 ;
  assign w7476 = ( w837 & ~w7474 ) | ( w837 & w7475 ) | ( ~w7474 & w7475 ) ;
  assign w7477 = ~\pi108 & w839 ;
  assign w7478 = w4425 | w7476 ;
  assign w7479 = ( w840 & w7476 ) | ( w840 & w7478 ) | ( w7476 & w7478 ) ;
  assign w7480 = ( w839 & ~w7477 ) | ( w839 & w7479 ) | ( ~w7477 & w7479 ) ;
  assign w7481 = \pi017 ^ w7480 ;
  assign w7482 = w7274 ^ w7473 ;
  assign w7483 = w7481 ^ w7482 ;
  assign w7484 = ~\pi110 & w601 ;
  assign w7485 = \pi109 & w683 ;
  assign w7486 = ( w601 & ~w7484 ) | ( w601 & w7485 ) | ( ~w7484 & w7485 ) ;
  assign w7487 = ~\pi111 & w603 ;
  assign w7488 = w4811 | w7486 ;
  assign w7489 = ( w604 & w7486 ) | ( w604 & w7488 ) | ( w7486 & w7488 ) ;
  assign w7490 = ( w603 & ~w7487 ) | ( w603 & w7489 ) | ( ~w7487 & w7489 ) ;
  assign w7491 = \pi014 ^ w7490 ;
  assign w7492 = w7316 ^ w7483 ;
  assign w7493 = w7491 ^ w7492 ;
  assign w7494 = w7307 ^ w7493 ;
  assign w7495 = w7315 ^ w7494 ;
  assign w7496 = w7298 ^ w7495 ;
  assign w7497 = w7306 ^ w7496 ;
  assign w7498 = ~\pi119 & w189 ;
  assign w7499 = \pi118 & w229 ;
  assign w7500 = ( w189 & ~w7498 ) | ( w189 & w7499 ) | ( ~w7498 & w7499 ) ;
  assign w7501 = ~\pi120 & w191 ;
  assign w7502 = w6634 | w7500 ;
  assign w7503 = ( w192 & w7500 ) | ( w192 & w7502 ) | ( w7500 & w7502 ) ;
  assign w7504 = ( w191 & ~w7501 ) | ( w191 & w7503 ) | ( ~w7501 & w7503 ) ;
  assign w7505 = \pi005 ^ w7504 ;
  assign w7506 = ( ~\pi002 & \pi122 ) | ( ~\pi002 & \pi123 ) | ( \pi122 & \pi123 ) ;
  assign w7507 = \pi000 ^ w7506 ;
  assign w7508 = ( \pi002 & \pi123 ) | ( \pi002 & ~w7507 ) | ( \pi123 & ~w7507 ) ;
  assign w7509 = ( \pi002 & \pi122 ) | ( \pi002 & w7507 ) | ( \pi122 & w7507 ) ;
  assign w7510 = \pi001 & w7509 ;
  assign w7511 = ( ~\pi000 & \pi121 ) | ( ~\pi000 & w7510 ) | ( \pi121 & w7510 ) ;
  assign w7512 = ( \pi001 & \pi002 ) | ( \pi001 & ~w7511 ) | ( \pi002 & ~w7511 ) ;
  assign w7513 = ( w7508 & w7510 ) | ( w7508 & ~w7512 ) | ( w7510 & ~w7512 ) ;
  assign w7514 = ( \pi121 & \pi122 ) | ( \pi121 & w7067 ) | ( \pi122 & w7067 ) ;
  assign w7515 = \pi122 ^ w7514 ;
  assign w7516 = \pi123 ^ w7515 ;
  assign w7517 = \pi002 ^ w7513 ;
  assign w7518 = \pi000 & ~w7513 ;
  assign w7519 = w7516 & w7518 ;
  assign w7520 = \pi001 ^ w7519 ;
  assign w7521 = ( \pi001 & w7517 ) | ( \pi001 & ~w7520 ) | ( w7517 & ~w7520 ) ;
  assign w7522 = w7497 ^ w7521 ;
  assign w7523 = w7505 ^ w7522 ;
  assign w7524 = w7296 ^ w7297 ;
  assign w7525 = w7523 ^ w7524 ;
  assign w7526 = ( w7296 & w7297 ) | ( w7296 & w7523 ) | ( w7297 & w7523 ) ;
  assign w7527 = ( w7497 & w7505 ) | ( w7497 & w7521 ) | ( w7505 & w7521 ) ;
  assign w7528 = ( ~\pi002 & \pi123 ) | ( ~\pi002 & \pi124 ) | ( \pi123 & \pi124 ) ;
  assign w7529 = \pi000 ^ w7528 ;
  assign w7530 = ( \pi002 & \pi124 ) | ( \pi002 & ~w7529 ) | ( \pi124 & ~w7529 ) ;
  assign w7531 = ( \pi002 & \pi123 ) | ( \pi002 & w7529 ) | ( \pi123 & w7529 ) ;
  assign w7532 = \pi001 & w7531 ;
  assign w7533 = ( ~\pi000 & \pi122 ) | ( ~\pi000 & w7532 ) | ( \pi122 & w7532 ) ;
  assign w7534 = ( \pi001 & \pi002 ) | ( \pi001 & ~w7533 ) | ( \pi002 & ~w7533 ) ;
  assign w7535 = ( w7530 & w7532 ) | ( w7530 & ~w7534 ) | ( w7532 & ~w7534 ) ;
  assign w7536 = ( \pi122 & \pi123 ) | ( \pi122 & w7514 ) | ( \pi123 & w7514 ) ;
  assign w7537 = \pi123 ^ w7536 ;
  assign w7538 = \pi124 ^ w7537 ;
  assign w7539 = \pi002 ^ w7535 ;
  assign w7540 = \pi000 & ~w7535 ;
  assign w7541 = w7538 & w7540 ;
  assign w7542 = \pi001 ^ w7541 ;
  assign w7543 = ( \pi001 & w7539 ) | ( \pi001 & ~w7542 ) | ( w7539 & ~w7542 ) ;
  assign w7544 = ~\pi120 & w189 ;
  assign w7545 = \pi119 & w229 ;
  assign w7546 = ( w189 & ~w7544 ) | ( w189 & w7545 ) | ( ~w7544 & w7545 ) ;
  assign w7547 = ~\pi121 & w191 ;
  assign w7548 = w7050 | w7546 ;
  assign w7549 = ( w192 & w7546 ) | ( w192 & w7548 ) | ( w7546 & w7548 ) ;
  assign w7550 = ( w191 & ~w7547 ) | ( w191 & w7549 ) | ( ~w7547 & w7549 ) ;
  assign w7551 = \pi005 ^ w7550 ;
  assign w7552 = ( w7298 & w7306 ) | ( w7298 & w7495 ) | ( w7306 & w7495 ) ;
  assign w7553 = ~\pi117 & w305 ;
  assign w7554 = \pi116 & w328 ;
  assign w7555 = ( w305 & ~w7553 ) | ( w305 & w7554 ) | ( ~w7553 & w7554 ) ;
  assign w7556 = ~\pi118 & w307 ;
  assign w7557 = w6206 | w7555 ;
  assign w7558 = ( w308 & w7555 ) | ( w308 & w7557 ) | ( w7555 & w7557 ) ;
  assign w7559 = ( w307 & ~w7556 ) | ( w307 & w7558 ) | ( ~w7556 & w7558 ) ;
  assign w7560 = \pi008 ^ w7559 ;
  assign w7561 = ( w7307 & w7315 ) | ( w7307 & w7493 ) | ( w7315 & w7493 ) ;
  assign w7562 = ~\pi114 & w432 ;
  assign w7563 = \pi113 & w486 ;
  assign w7564 = ( w432 & ~w7562 ) | ( w432 & w7563 ) | ( ~w7562 & w7563 ) ;
  assign w7565 = ~\pi115 & w434 ;
  assign w7566 = w5585 | w7564 ;
  assign w7567 = ( w435 & w7564 ) | ( w435 & w7566 ) | ( w7564 & w7566 ) ;
  assign w7568 = ( w434 & ~w7565 ) | ( w434 & w7567 ) | ( ~w7565 & w7567 ) ;
  assign w7569 = \pi011 ^ w7568 ;
  assign w7570 = ( w7316 & w7483 ) | ( w7316 & w7491 ) | ( w7483 & w7491 ) ;
  assign w7571 = ~\pi111 & w601 ;
  assign w7572 = \pi110 & w683 ;
  assign w7573 = ( w601 & ~w7571 ) | ( w601 & w7572 ) | ( ~w7571 & w7572 ) ;
  assign w7574 = ~\pi112 & w603 ;
  assign w7575 = w4999 | w7573 ;
  assign w7576 = ( w604 & w7573 ) | ( w604 & w7575 ) | ( w7573 & w7575 ) ;
  assign w7577 = ( w603 & ~w7574 ) | ( w603 & w7576 ) | ( ~w7574 & w7576 ) ;
  assign w7578 = \pi014 ^ w7577 ;
  assign w7579 = ( w7274 & w7473 ) | ( w7274 & w7481 ) | ( w7473 & w7481 ) ;
  assign w7580 = ~\pi108 & w837 ;
  assign w7581 = \pi107 & w902 ;
  assign w7582 = ( w837 & ~w7580 ) | ( w837 & w7581 ) | ( ~w7580 & w7581 ) ;
  assign w7583 = ~\pi109 & w839 ;
  assign w7584 = w4599 | w7582 ;
  assign w7585 = ( w840 & w7582 ) | ( w840 & w7584 ) | ( w7582 & w7584 ) ;
  assign w7586 = ( w839 & ~w7583 ) | ( w839 & w7585 ) | ( ~w7583 & w7585 ) ;
  assign w7587 = \pi017 ^ w7586 ;
  assign w7588 = ( w7325 & w7448 ) | ( w7325 & w7449 ) | ( w7448 & w7449 ) ;
  assign w7589 = ( w7326 & w7438 ) | ( w7326 & w7446 ) | ( w7438 & w7446 ) ;
  assign w7590 = ~\pi096 & w1944 ;
  assign w7591 = \pi095 & w2072 ;
  assign w7592 = ( w1944 & ~w7590 ) | ( w1944 & w7591 ) | ( ~w7590 & w7591 ) ;
  assign w7593 = ~\pi097 & w1946 ;
  assign w7594 = w2673 | w7592 ;
  assign w7595 = ( w1947 & w7592 ) | ( w1947 & w7594 ) | ( w7592 & w7594 ) ;
  assign w7596 = ( w1946 & ~w7593 ) | ( w1946 & w7595 ) | ( ~w7593 & w7595 ) ;
  assign w7597 = \pi029 ^ w7596 ;
  assign w7598 = ( w7188 & w7396 ) | ( w7188 & w7404 ) | ( w7396 & w7404 ) ;
  assign w7599 = ~\pi084 & w3635 ;
  assign w7600 = \pi083 & w3817 ;
  assign w7601 = ( w3635 & ~w7599 ) | ( w3635 & w7600 ) | ( ~w7599 & w7600 ) ;
  assign w7602 = ~\pi085 & w3637 ;
  assign w7603 = w1274 | w7601 ;
  assign w7604 = ( w3638 & w7601 ) | ( w3638 & w7603 ) | ( w7601 & w7603 ) ;
  assign w7605 = ( w3637 & ~w7602 ) | ( w3637 & w7604 ) | ( ~w7602 & w7604 ) ;
  assign w7606 = \pi041 ^ w7605 ;
  assign w7607 = ( w7329 & w7337 ) | ( w7329 & w7394 ) | ( w7337 & w7394 ) ;
  assign w7608 = ~\pi081 & w4141 ;
  assign w7609 = \pi080 & w4334 ;
  assign w7610 = ( w4141 & ~w7608 ) | ( w4141 & w7609 ) | ( ~w7608 & w7609 ) ;
  assign w7611 = ~\pi082 & w4143 ;
  assign w7612 = w1008 | w7610 ;
  assign w7613 = ( w4144 & w7610 ) | ( w4144 & w7612 ) | ( w7610 & w7612 ) ;
  assign w7614 = ( w4143 & ~w7611 ) | ( w4143 & w7613 ) | ( ~w7611 & w7613 ) ;
  assign w7615 = \pi044 ^ w7614 ;
  assign w7616 = ( w7166 & w7345 ) | ( w7166 & w7392 ) | ( w7345 & w7392 ) ;
  assign w7617 = ~\pi078 & w4654 ;
  assign w7618 = \pi077 & w4876 ;
  assign w7619 = ( w4654 & ~w7617 ) | ( w4654 & w7618 ) | ( ~w7617 & w7618 ) ;
  assign w7620 = ~\pi079 & w4656 ;
  assign w7621 = w730 | w7619 ;
  assign w7622 = ( w4657 & w7619 ) | ( w4657 & w7621 ) | ( w7619 & w7621 ) ;
  assign w7623 = ( w4656 & ~w7620 ) | ( w4656 & w7622 ) | ( ~w7620 & w7622 ) ;
  assign w7624 = \pi047 ^ w7623 ;
  assign w7625 = ( w7346 & w7354 ) | ( w7346 & w7390 ) | ( w7354 & w7390 ) ;
  assign w7626 = ~\pi075 & w5209 ;
  assign w7627 = \pi074 & w5433 ;
  assign w7628 = ( w5209 & ~w7626 ) | ( w5209 & w7627 ) | ( ~w7626 & w7627 ) ;
  assign w7629 = ~\pi076 & w5211 ;
  assign w7630 = w538 | w7628 ;
  assign w7631 = ( w5212 & w7628 ) | ( w5212 & w7630 ) | ( w7628 & w7630 ) ;
  assign w7632 = ( w5211 & ~w7629 ) | ( w5211 & w7631 ) | ( ~w7629 & w7631 ) ;
  assign w7633 = \pi050 ^ w7632 ;
  assign w7634 = ( w7355 & w7380 ) | ( w7355 & w7388 ) | ( w7380 & w7388 ) ;
  assign w7635 = ~\pi069 & w6466 ;
  assign w7636 = \pi068 & w6702 ;
  assign w7637 = ( w6466 & ~w7635 ) | ( w6466 & w7636 ) | ( ~w7635 & w7636 ) ;
  assign w7638 = ~\pi070 & w6468 ;
  assign w7639 = w271 | w7637 ;
  assign w7640 = ( w6469 & w7637 ) | ( w6469 & w7639 ) | ( w7637 & w7639 ) ;
  assign w7641 = ( w6468 & ~w7638 ) | ( w6468 & w7640 ) | ( ~w7638 & w7640 ) ;
  assign w7642 = \pi056 ^ w7641 ;
  assign w7643 = ~\pi066 & w7135 ;
  assign w7644 = \pi065 & w7359 ;
  assign w7645 = ( w7135 & ~w7643 ) | ( w7135 & w7644 ) | ( ~w7643 & w7644 ) ;
  assign w7646 = ~\pi067 & w7137 ;
  assign w7647 = w160 | w7645 ;
  assign w7648 = ( w7138 & w7645 ) | ( w7138 & w7647 ) | ( w7645 & w7647 ) ;
  assign w7649 = ( w7137 & ~w7646 ) | ( w7137 & w7648 ) | ( ~w7646 & w7648 ) ;
  assign w7650 = \pi059 ^ w7649 ;
  assign w7651 = w7368 ^ w7650 ;
  assign w7652 = \pi059 ^ \pi060 ;
  assign w7653 = \pi064 & w7652 ;
  assign w7654 = w7651 ^ w7653 ;
  assign w7655 = w7378 ^ w7654 ;
  assign w7656 = w7642 ^ w7655 ;
  assign w7657 = ~\pi072 & w5802 ;
  assign w7658 = \pi071 & w6052 ;
  assign w7659 = ( w5802 & ~w7657 ) | ( w5802 & w7658 ) | ( ~w7657 & w7658 ) ;
  assign w7660 = ~\pi073 & w5804 ;
  assign w7661 = w404 | w7659 ;
  assign w7662 = ( w5805 & w7659 ) | ( w5805 & w7661 ) | ( w7659 & w7661 ) ;
  assign w7663 = ( w5804 & ~w7660 ) | ( w5804 & w7662 ) | ( ~w7660 & w7662 ) ;
  assign w7664 = \pi053 ^ w7663 ;
  assign w7665 = w7634 ^ w7656 ;
  assign w7666 = w7664 ^ w7665 ;
  assign w7667 = w7625 ^ w7666 ;
  assign w7668 = w7633 ^ w7667 ;
  assign w7669 = w7616 ^ w7668 ;
  assign w7670 = w7624 ^ w7669 ;
  assign w7671 = w7607 ^ w7670 ;
  assign w7672 = w7615 ^ w7671 ;
  assign w7673 = w7598 ^ w7672 ;
  assign w7674 = w7606 ^ w7673 ;
  assign w7675 = ~\pi087 & w3178 ;
  assign w7676 = \pi086 & w3340 ;
  assign w7677 = ( w3178 & ~w7675 ) | ( w3178 & w7676 ) | ( ~w7675 & w7676 ) ;
  assign w7678 = ~\pi088 & w3180 ;
  assign w7679 = w1574 | w7677 ;
  assign w7680 = ( w3181 & w7677 ) | ( w3181 & w7679 ) | ( w7677 & w7679 ) ;
  assign w7681 = ( w3180 & ~w7678 ) | ( w3180 & w7680 ) | ( ~w7678 & w7680 ) ;
  assign w7682 = \pi038 ^ w7681 ;
  assign w7683 = ( w7328 & w7406 ) | ( w7328 & w7414 ) | ( w7406 & w7414 ) ;
  assign w7684 = w7674 ^ w7683 ;
  assign w7685 = w7682 ^ w7684 ;
  assign w7686 = ~\pi090 & w2712 ;
  assign w7687 = \pi089 & w2872 ;
  assign w7688 = ( w2712 & ~w7686 ) | ( w2712 & w7687 ) | ( ~w7686 & w7687 ) ;
  assign w7689 = ~\pi091 & w2714 ;
  assign w7690 = w1908 | w7688 ;
  assign w7691 = ( w2715 & w7688 ) | ( w2715 & w7690 ) | ( w7688 & w7690 ) ;
  assign w7692 = ( w2714 & ~w7689 ) | ( w2714 & w7691 ) | ( ~w7689 & w7691 ) ;
  assign w7693 = \pi035 ^ w7692 ;
  assign w7694 = ( w7416 & w7424 ) | ( w7416 & w7425 ) | ( w7424 & w7425 ) ;
  assign w7695 = w7685 ^ w7694 ;
  assign w7696 = w7693 ^ w7695 ;
  assign w7697 = ~\pi093 & w2310 ;
  assign w7698 = \pi092 & w2443 ;
  assign w7699 = ( w2310 & ~w7697 ) | ( w2310 & w7698 ) | ( ~w7697 & w7698 ) ;
  assign w7700 = ~\pi094 & w2312 ;
  assign w7701 = w2274 | w7699 ;
  assign w7702 = ( w2313 & w7699 ) | ( w2313 & w7701 ) | ( w7699 & w7701 ) ;
  assign w7703 = ( w2312 & ~w7700 ) | ( w2312 & w7702 ) | ( ~w7700 & w7702 ) ;
  assign w7704 = \pi032 ^ w7703 ;
  assign w7705 = w7436 ^ w7696 ;
  assign w7706 = w7704 ^ w7705 ;
  assign w7707 = w7589 ^ w7706 ;
  assign w7708 = w7597 ^ w7707 ;
  assign w7709 = ~\pi099 & w1629 ;
  assign w7710 = \pi098 & w1722 ;
  assign w7711 = ( w1629 & ~w7709 ) | ( w1629 & w7710 ) | ( ~w7709 & w7710 ) ;
  assign w7712 = ~\pi100 & w1631 ;
  assign w7713 = w3104 | w7711 ;
  assign w7714 = ( w1632 & w7711 ) | ( w1632 & w7713 ) | ( w7711 & w7713 ) ;
  assign w7715 = ( w1631 & ~w7712 ) | ( w1631 & w7714 ) | ( ~w7712 & w7714 ) ;
  assign w7716 = \pi026 ^ w7715 ;
  assign w7717 = w7588 ^ w7708 ;
  assign w7718 = w7716 ^ w7717 ;
  assign w7719 = ~\pi102 & w1313 ;
  assign w7720 = \pi101 & w1417 ;
  assign w7721 = ( w1313 & ~w7719 ) | ( w1313 & w7720 ) | ( ~w7719 & w7720 ) ;
  assign w7722 = ~\pi103 & w1315 ;
  assign w7723 = w3437 | w7721 ;
  assign w7724 = ( w1316 & w7721 ) | ( w1316 & w7723 ) | ( w7721 & w7723 ) ;
  assign w7725 = ( w1315 & ~w7722 ) | ( w1315 & w7724 ) | ( ~w7722 & w7724 ) ;
  assign w7726 = \pi023 ^ w7725 ;
  assign w7727 = ( w7451 & w7459 ) | ( w7451 & w7460 ) | ( w7459 & w7460 ) ;
  assign w7728 = w7718 ^ w7727 ;
  assign w7729 = w7726 ^ w7728 ;
  assign w7730 = ~\pi105 & w1044 ;
  assign w7731 = \pi104 & w1138 ;
  assign w7732 = ( w1044 & ~w7730 ) | ( w1044 & w7731 ) | ( ~w7730 & w7731 ) ;
  assign w7733 = ~\pi106 & w1046 ;
  assign w7734 = w4068 | w7732 ;
  assign w7735 = ( w1047 & w7732 ) | ( w1047 & w7734 ) | ( w7732 & w7734 ) ;
  assign w7736 = ( w1046 & ~w7733 ) | ( w1046 & w7735 ) | ( ~w7733 & w7735 ) ;
  assign w7737 = \pi020 ^ w7736 ;
  assign w7738 = w7471 ^ w7729 ;
  assign w7739 = w7737 ^ w7738 ;
  assign w7740 = w7579 ^ w7739 ;
  assign w7741 = w7587 ^ w7740 ;
  assign w7742 = w7570 ^ w7741 ;
  assign w7743 = w7578 ^ w7742 ;
  assign w7744 = w7561 ^ w7743 ;
  assign w7745 = w7569 ^ w7744 ;
  assign w7746 = w7552 ^ w7745 ;
  assign w7747 = w7560 ^ w7746 ;
  assign w7748 = w7543 ^ w7747 ;
  assign w7749 = w7551 ^ w7748 ;
  assign w7750 = w7526 ^ w7749 ;
  assign w7751 = w7527 ^ w7750 ;
  assign w7752 = ~\pi118 & w305 ;
  assign w7753 = \pi117 & w328 ;
  assign w7754 = ( w305 & ~w7752 ) | ( w305 & w7753 ) | ( ~w7752 & w7753 ) ;
  assign w7755 = ~\pi119 & w307 ;
  assign w7756 = w6616 | w7754 ;
  assign w7757 = ( w308 & w7754 ) | ( w308 & w7756 ) | ( w7754 & w7756 ) ;
  assign w7758 = ( w307 & ~w7755 ) | ( w307 & w7757 ) | ( ~w7755 & w7757 ) ;
  assign w7759 = \pi008 ^ w7758 ;
  assign w7760 = ( w7561 & w7569 ) | ( w7561 & w7743 ) | ( w7569 & w7743 ) ;
  assign w7761 = ~\pi115 & w432 ;
  assign w7762 = \pi114 & w486 ;
  assign w7763 = ( w432 & ~w7761 ) | ( w432 & w7762 ) | ( ~w7761 & w7762 ) ;
  assign w7764 = ~\pi116 & w434 ;
  assign w7765 = w5976 | w7763 ;
  assign w7766 = ( w435 & w7763 ) | ( w435 & w7765 ) | ( w7763 & w7765 ) ;
  assign w7767 = ( w434 & ~w7764 ) | ( w434 & w7766 ) | ( ~w7764 & w7766 ) ;
  assign w7768 = \pi011 ^ w7767 ;
  assign w7769 = ( w7570 & w7578 ) | ( w7570 & w7741 ) | ( w7578 & w7741 ) ;
  assign w7770 = ~\pi112 & w601 ;
  assign w7771 = \pi111 & w683 ;
  assign w7772 = ( w601 & ~w7770 ) | ( w601 & w7771 ) | ( ~w7770 & w7771 ) ;
  assign w7773 = ~\pi113 & w603 ;
  assign w7774 = w5366 | w7772 ;
  assign w7775 = ( w604 & w7772 ) | ( w604 & w7774 ) | ( w7772 & w7774 ) ;
  assign w7776 = ( w603 & ~w7773 ) | ( w603 & w7775 ) | ( ~w7773 & w7775 ) ;
  assign w7777 = \pi014 ^ w7776 ;
  assign w7778 = ( w7579 & w7587 ) | ( w7579 & w7739 ) | ( w7587 & w7739 ) ;
  assign w7779 = ( w7471 & w7729 ) | ( w7471 & w7737 ) | ( w7729 & w7737 ) ;
  assign w7780 = ( w7589 & w7597 ) | ( w7589 & w7706 ) | ( w7597 & w7706 ) ;
  assign w7781 = ( w7436 & w7696 ) | ( w7436 & w7704 ) | ( w7696 & w7704 ) ;
  assign w7782 = ( w7607 & w7615 ) | ( w7607 & w7670 ) | ( w7615 & w7670 ) ;
  assign w7783 = ( w7625 & w7633 ) | ( w7625 & w7666 ) | ( w7633 & w7666 ) ;
  assign w7784 = ~\pi073 & w5802 ;
  assign w7785 = \pi072 & w6052 ;
  assign w7786 = ( w5802 & ~w7784 ) | ( w5802 & w7785 ) | ( ~w7784 & w7785 ) ;
  assign w7787 = ~\pi074 & w5804 ;
  assign w7788 = w465 | w7786 ;
  assign w7789 = ( w5805 & w7786 ) | ( w5805 & w7788 ) | ( w7786 & w7788 ) ;
  assign w7790 = ( w5804 & ~w7787 ) | ( w5804 & w7789 ) | ( ~w7787 & w7789 ) ;
  assign w7791 = \pi053 ^ w7790 ;
  assign w7792 = ( w7378 & w7642 ) | ( w7378 & w7654 ) | ( w7642 & w7654 ) ;
  assign w7793 = ~\pi070 & w6466 ;
  assign w7794 = \pi069 & w6702 ;
  assign w7795 = ( w6466 & ~w7793 ) | ( w6466 & w7794 ) | ( ~w7793 & w7794 ) ;
  assign w7796 = ~\pi071 & w6468 ;
  assign w7797 = w290 | w7795 ;
  assign w7798 = ( w6469 & w7795 ) | ( w6469 & w7797 ) | ( w7795 & w7797 ) ;
  assign w7799 = ( w6468 & ~w7796 ) | ( w6468 & w7798 ) | ( ~w7796 & w7798 ) ;
  assign w7800 = \pi056 ^ w7799 ;
  assign w7801 = ( w7368 & w7650 ) | ( w7368 & w7653 ) | ( w7650 & w7653 ) ;
  assign w7802 = ~\pi067 & w7135 ;
  assign w7803 = \pi066 & w7359 ;
  assign w7804 = ( w7135 & ~w7802 ) | ( w7135 & w7803 ) | ( ~w7802 & w7803 ) ;
  assign w7805 = ~\pi068 & w7137 ;
  assign w7806 = w182 | w7804 ;
  assign w7807 = ( w7138 & w7804 ) | ( w7138 & w7806 ) | ( w7804 & w7806 ) ;
  assign w7808 = ( w7137 & ~w7805 ) | ( w7137 & w7807 ) | ( ~w7805 & w7807 ) ;
  assign w7809 = \pi059 ^ w7808 ;
  assign w7810 = ( \pi059 & \pi060 ) | ( \pi059 & \pi061 ) | ( \pi060 & \pi061 ) ;
  assign w7811 = \pi061 ^ w7810 ;
  assign w7812 = \pi061 ^ \pi062 ;
  assign w7813 = w7652 & ~w7812 ;
  assign w7814 = w7652 & w7812 ;
  assign w7815 = ( \pi059 & \pi060 ) | ( \pi059 & ~\pi062 ) | ( \pi060 & ~\pi062 ) ;
  assign w7816 = \pi062 & ~\pi064 ;
  assign w7817 = ~\pi065 & w7816 ;
  assign w7818 = ( \pi059 & \pi060 ) | ( \pi059 & ~w7817 ) | ( \pi060 & ~w7817 ) ;
  assign w7819 = ( \pi061 & \pi062 ) | ( \pi061 & ~w7818 ) | ( \pi062 & ~w7818 ) ;
  assign w7820 = ( \pi061 & ~w7816 ) | ( \pi061 & w7818 ) | ( ~w7816 & w7818 ) ;
  assign w7821 = ( w7815 & w7819 ) | ( w7815 & ~w7820 ) | ( w7819 & ~w7820 ) ;
  assign w7822 = ( \pi059 & \pi060 ) | ( \pi059 & \pi065 ) | ( \pi060 & \pi065 ) ;
  assign w7823 = \pi059 & \pi060 ;
  assign w7824 = \pi064 ^ w7823 ;
  assign w7825 = ( \pi061 & w7823 ) | ( \pi061 & w7824 ) | ( w7823 & w7824 ) ;
  assign w7826 = w7822 ^ w7825 ;
  assign w7827 = w7801 ^ w7809 ;
  assign w7828 = w7826 ^ w7827 ;
  assign w7829 = w7792 ^ w7828 ;
  assign w7830 = w7800 ^ w7829 ;
  assign w7831 = ( w7634 & w7656 ) | ( w7634 & w7664 ) | ( w7656 & w7664 ) ;
  assign w7832 = w7830 ^ w7831 ;
  assign w7833 = w7791 ^ w7832 ;
  assign w7834 = ~\pi076 & w5209 ;
  assign w7835 = \pi075 & w5433 ;
  assign w7836 = ( w5209 & ~w7834 ) | ( w5209 & w7835 ) | ( ~w7834 & w7835 ) ;
  assign w7837 = ~\pi077 & w5211 ;
  assign w7838 = w644 | w7836 ;
  assign w7839 = ( w5212 & w7836 ) | ( w5212 & w7838 ) | ( w7836 & w7838 ) ;
  assign w7840 = ( w5211 & ~w7837 ) | ( w5211 & w7839 ) | ( ~w7837 & w7839 ) ;
  assign w7841 = \pi050 ^ w7840 ;
  assign w7842 = ( w7783 & w7833 ) | ( w7783 & w7841 ) | ( w7833 & w7841 ) ;
  assign w7843 = w7783 ^ w7833 ;
  assign w7844 = w7841 ^ w7843 ;
  assign w7845 = ~\pi079 & w4654 ;
  assign w7846 = \pi078 & w4876 ;
  assign w7847 = ( w4654 & ~w7845 ) | ( w4654 & w7846 ) | ( ~w7845 & w7846 ) ;
  assign w7848 = ~\pi080 & w4656 ;
  assign w7849 = w794 | w7847 ;
  assign w7850 = ( w4657 & w7847 ) | ( w4657 & w7849 ) | ( w7847 & w7849 ) ;
  assign w7851 = ( w4656 & ~w7848 ) | ( w4656 & w7850 ) | ( ~w7848 & w7850 ) ;
  assign w7852 = \pi047 ^ w7851 ;
  assign w7853 = ( w7616 & w7624 ) | ( w7616 & w7668 ) | ( w7624 & w7668 ) ;
  assign w7854 = w7844 ^ w7853 ;
  assign w7855 = w7852 ^ w7854 ;
  assign w7856 = ~\pi082 & w4141 ;
  assign w7857 = \pi081 & w4334 ;
  assign w7858 = ( w4141 & ~w7856 ) | ( w4141 & w7857 ) | ( ~w7856 & w7857 ) ;
  assign w7859 = ~\pi083 & w4143 ;
  assign w7860 = w1099 | w7858 ;
  assign w7861 = ( w4144 & w7858 ) | ( w4144 & w7860 ) | ( w7858 & w7860 ) ;
  assign w7862 = ( w4143 & ~w7859 ) | ( w4143 & w7861 ) | ( ~w7859 & w7861 ) ;
  assign w7863 = \pi044 ^ w7862 ;
  assign w7864 = ( w7782 & w7855 ) | ( w7782 & w7863 ) | ( w7855 & w7863 ) ;
  assign w7865 = w7782 ^ w7855 ;
  assign w7866 = w7863 ^ w7865 ;
  assign w7867 = ~\pi085 & w3635 ;
  assign w7868 = \pi084 & w3817 ;
  assign w7869 = ( w3635 & ~w7867 ) | ( w3635 & w7868 ) | ( ~w7867 & w7868 ) ;
  assign w7870 = ~\pi086 & w3637 ;
  assign w7871 = w1379 | w7869 ;
  assign w7872 = ( w3638 & w7869 ) | ( w3638 & w7871 ) | ( w7869 & w7871 ) ;
  assign w7873 = ( w3637 & ~w7870 ) | ( w3637 & w7872 ) | ( ~w7870 & w7872 ) ;
  assign w7874 = \pi041 ^ w7873 ;
  assign w7875 = ( w7598 & w7606 ) | ( w7598 & w7672 ) | ( w7606 & w7672 ) ;
  assign w7876 = w7866 ^ w7875 ;
  assign w7877 = w7874 ^ w7876 ;
  assign w7878 = ~\pi088 & w3178 ;
  assign w7879 = \pi087 & w3340 ;
  assign w7880 = ( w3178 & ~w7878 ) | ( w3178 & w7879 ) | ( ~w7878 & w7879 ) ;
  assign w7881 = ~\pi089 & w3180 ;
  assign w7882 = w1595 | w7880 ;
  assign w7883 = ( w3181 & w7880 ) | ( w3181 & w7882 ) | ( w7880 & w7882 ) ;
  assign w7884 = ( w3180 & ~w7881 ) | ( w3180 & w7883 ) | ( ~w7881 & w7883 ) ;
  assign w7885 = \pi038 ^ w7884 ;
  assign w7886 = ( w7674 & w7682 ) | ( w7674 & w7683 ) | ( w7682 & w7683 ) ;
  assign w7887 = w7877 ^ w7886 ;
  assign w7888 = w7885 ^ w7887 ;
  assign w7889 = ~\pi091 & w2712 ;
  assign w7890 = \pi090 & w2872 ;
  assign w7891 = ( w2712 & ~w7889 ) | ( w2712 & w7890 ) | ( ~w7889 & w7890 ) ;
  assign w7892 = ~\pi092 & w2714 ;
  assign w7893 = w2033 | w7891 ;
  assign w7894 = ( w2715 & w7891 ) | ( w2715 & w7893 ) | ( w7891 & w7893 ) ;
  assign w7895 = ( w2714 & ~w7892 ) | ( w2714 & w7894 ) | ( ~w7892 & w7894 ) ;
  assign w7896 = \pi035 ^ w7895 ;
  assign w7897 = ( w7685 & w7693 ) | ( w7685 & w7694 ) | ( w7693 & w7694 ) ;
  assign w7898 = w7888 ^ w7897 ;
  assign w7899 = w7896 ^ w7898 ;
  assign w7900 = ~\pi094 & w2310 ;
  assign w7901 = \pi093 & w2443 ;
  assign w7902 = ( w2310 & ~w7900 ) | ( w2310 & w7901 ) | ( ~w7900 & w7901 ) ;
  assign w7903 = ~\pi095 & w2312 ;
  assign w7904 = w2409 | w7902 ;
  assign w7905 = ( w2313 & w7902 ) | ( w2313 & w7904 ) | ( w7902 & w7904 ) ;
  assign w7906 = ( w2312 & ~w7903 ) | ( w2312 & w7905 ) | ( ~w7903 & w7905 ) ;
  assign w7907 = \pi032 ^ w7906 ;
  assign w7908 = w7781 ^ w7899 ;
  assign w7909 = w7907 ^ w7908 ;
  assign w7910 = ~\pi097 & w1944 ;
  assign w7911 = \pi096 & w2072 ;
  assign w7912 = ( w1944 & ~w7910 ) | ( w1944 & w7911 ) | ( ~w7910 & w7911 ) ;
  assign w7913 = ~\pi098 & w1946 ;
  assign w7914 = w2824 | w7912 ;
  assign w7915 = ( w1947 & w7912 ) | ( w1947 & w7914 ) | ( w7912 & w7914 ) ;
  assign w7916 = ( w1946 & ~w7913 ) | ( w1946 & w7915 ) | ( ~w7913 & w7915 ) ;
  assign w7917 = \pi029 ^ w7916 ;
  assign w7918 = w7780 ^ w7909 ;
  assign w7919 = w7917 ^ w7918 ;
  assign w7920 = ~\pi100 & w1629 ;
  assign w7921 = \pi099 & w1722 ;
  assign w7922 = ( w1629 & ~w7920 ) | ( w1629 & w7921 ) | ( ~w7920 & w7921 ) ;
  assign w7923 = ~\pi101 & w1631 ;
  assign w7924 = w3264 | w7922 ;
  assign w7925 = ( w1632 & w7922 ) | ( w1632 & w7924 ) | ( w7922 & w7924 ) ;
  assign w7926 = ( w1631 & ~w7923 ) | ( w1631 & w7925 ) | ( ~w7923 & w7925 ) ;
  assign w7927 = \pi026 ^ w7926 ;
  assign w7928 = ( w7588 & w7708 ) | ( w7588 & w7716 ) | ( w7708 & w7716 ) ;
  assign w7929 = w7919 ^ w7928 ;
  assign w7930 = w7927 ^ w7929 ;
  assign w7931 = ~\pi103 & w1313 ;
  assign w7932 = \pi102 & w1417 ;
  assign w7933 = ( w1313 & ~w7931 ) | ( w1313 & w7932 ) | ( ~w7931 & w7932 ) ;
  assign w7934 = ~\pi104 & w1315 ;
  assign w7935 = w3740 | w7933 ;
  assign w7936 = ( w1316 & w7933 ) | ( w1316 & w7935 ) | ( w7933 & w7935 ) ;
  assign w7937 = ( w1315 & ~w7934 ) | ( w1315 & w7936 ) | ( ~w7934 & w7936 ) ;
  assign w7938 = \pi023 ^ w7937 ;
  assign w7939 = ( w7718 & w7726 ) | ( w7718 & w7727 ) | ( w7726 & w7727 ) ;
  assign w7940 = w7930 ^ w7939 ;
  assign w7941 = w7938 ^ w7940 ;
  assign w7942 = ~\pi106 & w1044 ;
  assign w7943 = \pi105 & w1138 ;
  assign w7944 = ( w1044 & ~w7942 ) | ( w1044 & w7943 ) | ( ~w7942 & w7943 ) ;
  assign w7945 = ~\pi107 & w1046 ;
  assign w7946 = w4087 | w7944 ;
  assign w7947 = ( w1047 & w7944 ) | ( w1047 & w7946 ) | ( w7944 & w7946 ) ;
  assign w7948 = ( w1046 & ~w7945 ) | ( w1046 & w7947 ) | ( ~w7945 & w7947 ) ;
  assign w7949 = \pi020 ^ w7948 ;
  assign w7950 = ( w7779 & w7941 ) | ( w7779 & w7949 ) | ( w7941 & w7949 ) ;
  assign w7951 = w7779 ^ w7941 ;
  assign w7952 = w7949 ^ w7951 ;
  assign w7953 = ~\pi109 & w837 ;
  assign w7954 = \pi108 & w902 ;
  assign w7955 = ( w837 & ~w7953 ) | ( w837 & w7954 ) | ( ~w7953 & w7954 ) ;
  assign w7956 = ~\pi110 & w839 ;
  assign w7957 = w4792 | w7955 ;
  assign w7958 = ( w840 & w7955 ) | ( w840 & w7957 ) | ( w7955 & w7957 ) ;
  assign w7959 = ( w839 & ~w7956 ) | ( w839 & w7958 ) | ( ~w7956 & w7958 ) ;
  assign w7960 = \pi017 ^ w7959 ;
  assign w7961 = w7778 ^ w7952 ;
  assign w7962 = w7960 ^ w7961 ;
  assign w7963 = w7769 ^ w7962 ;
  assign w7964 = w7777 ^ w7963 ;
  assign w7965 = w7760 ^ w7964 ;
  assign w7966 = w7768 ^ w7965 ;
  assign w7967 = ( w7552 & w7560 ) | ( w7552 & w7745 ) | ( w7560 & w7745 ) ;
  assign w7968 = w7966 ^ w7967 ;
  assign w7969 = w7759 ^ w7968 ;
  assign w7970 = ~\pi121 & w189 ;
  assign w7971 = \pi120 & w229 ;
  assign w7972 = ( w189 & ~w7970 ) | ( w189 & w7971 ) | ( ~w7970 & w7971 ) ;
  assign w7973 = ~\pi122 & w191 ;
  assign w7974 = w7069 | w7972 ;
  assign w7975 = ( w192 & w7972 ) | ( w192 & w7974 ) | ( w7972 & w7974 ) ;
  assign w7976 = ( w191 & ~w7973 ) | ( w191 & w7975 ) | ( ~w7973 & w7975 ) ;
  assign w7977 = \pi005 ^ w7976 ;
  assign w7978 = ( ~\pi002 & \pi124 ) | ( ~\pi002 & \pi125 ) | ( \pi124 & \pi125 ) ;
  assign w7979 = \pi000 ^ w7978 ;
  assign w7980 = ( \pi002 & \pi125 ) | ( \pi002 & ~w7979 ) | ( \pi125 & ~w7979 ) ;
  assign w7981 = ( \pi002 & \pi124 ) | ( \pi002 & w7979 ) | ( \pi124 & w7979 ) ;
  assign w7982 = \pi001 & w7981 ;
  assign w7983 = ( ~\pi000 & \pi123 ) | ( ~\pi000 & w7982 ) | ( \pi123 & w7982 ) ;
  assign w7984 = ( \pi001 & \pi002 ) | ( \pi001 & ~w7983 ) | ( \pi002 & ~w7983 ) ;
  assign w7985 = ( w7980 & w7982 ) | ( w7980 & ~w7984 ) | ( w7982 & ~w7984 ) ;
  assign w7986 = ( \pi123 & \pi124 ) | ( \pi123 & w7536 ) | ( \pi124 & w7536 ) ;
  assign w7987 = \pi124 ^ w7986 ;
  assign w7988 = \pi125 ^ w7987 ;
  assign w7989 = \pi002 ^ w7985 ;
  assign w7990 = \pi000 & ~w7985 ;
  assign w7991 = w7988 & w7990 ;
  assign w7992 = \pi001 ^ w7991 ;
  assign w7993 = ( \pi001 & w7989 ) | ( \pi001 & ~w7992 ) | ( w7989 & ~w7992 ) ;
  assign w7994 = w7969 ^ w7993 ;
  assign w7995 = w7977 ^ w7994 ;
  assign w7996 = ( w7543 & w7551 ) | ( w7543 & w7747 ) | ( w7551 & w7747 ) ;
  assign w7997 = ( w7526 & w7527 ) | ( w7526 & w7749 ) | ( w7527 & w7749 ) ;
  assign w7998 = w7995 ^ w7997 ;
  assign w7999 = w7996 ^ w7998 ;
  assign w8000 = ( w7995 & w7996 ) | ( w7995 & w7997 ) | ( w7996 & w7997 ) ;
  assign w8001 = ( w7969 & w7977 ) | ( w7969 & w7993 ) | ( w7977 & w7993 ) ;
  assign w8002 = ( w7760 & w7768 ) | ( w7760 & w7964 ) | ( w7768 & w7964 ) ;
  assign w8003 = ( w7769 & w7777 ) | ( w7769 & w7962 ) | ( w7777 & w7962 ) ;
  assign w8004 = ~\pi113 & w601 ;
  assign w8005 = \pi112 & w683 ;
  assign w8006 = ( w601 & ~w8004 ) | ( w601 & w8005 ) | ( ~w8004 & w8005 ) ;
  assign w8007 = ~\pi114 & w603 ;
  assign w8008 = w5565 | w8006 ;
  assign w8009 = ( w604 & w8006 ) | ( w604 & w8008 ) | ( w8006 & w8008 ) ;
  assign w8010 = ( w603 & ~w8007 ) | ( w603 & w8009 ) | ( ~w8007 & w8009 ) ;
  assign w8011 = \pi014 ^ w8010 ;
  assign w8012 = ( w7778 & w7952 ) | ( w7778 & w7960 ) | ( w7952 & w7960 ) ;
  assign w8013 = ( w7930 & w7938 ) | ( w7930 & w7939 ) | ( w7938 & w7939 ) ;
  assign w8014 = ( w7781 & w7899 ) | ( w7781 & w7907 ) | ( w7899 & w7907 ) ;
  assign w8015 = ( w7866 & w7874 ) | ( w7866 & w7875 ) | ( w7874 & w7875 ) ;
  assign w8016 = ( w7844 & w7852 ) | ( w7844 & w7853 ) | ( w7852 & w7853 ) ;
  assign w8017 = ~\pi080 & w4654 ;
  assign w8018 = \pi079 & w4876 ;
  assign w8019 = ( w4654 & ~w8017 ) | ( w4654 & w8018 ) | ( ~w8017 & w8018 ) ;
  assign w8020 = ~\pi081 & w4656 ;
  assign w8021 = w874 | w8019 ;
  assign w8022 = ( w4657 & w8019 ) | ( w4657 & w8021 ) | ( w8019 & w8021 ) ;
  assign w8023 = ( w4656 & ~w8020 ) | ( w4656 & w8022 ) | ( ~w8020 & w8022 ) ;
  assign w8024 = \pi047 ^ w8023 ;
  assign w8025 = ~\pi077 & w5209 ;
  assign w8026 = \pi076 & w5433 ;
  assign w8027 = ( w5209 & ~w8025 ) | ( w5209 & w8026 ) | ( ~w8025 & w8026 ) ;
  assign w8028 = ~\pi078 & w5211 ;
  assign w8029 = w665 | w8027 ;
  assign w8030 = ( w5212 & w8027 ) | ( w5212 & w8029 ) | ( w8027 & w8029 ) ;
  assign w8031 = ( w5211 & ~w8028 ) | ( w5211 & w8030 ) | ( ~w8028 & w8030 ) ;
  assign w8032 = \pi050 ^ w8031 ;
  assign w8033 = ( w7791 & w7830 ) | ( w7791 & w7831 ) | ( w7830 & w7831 ) ;
  assign w8034 = ~\pi074 & w5802 ;
  assign w8035 = \pi073 & w6052 ;
  assign w8036 = ( w5802 & ~w8034 ) | ( w5802 & w8035 ) | ( ~w8034 & w8035 ) ;
  assign w8037 = ~\pi075 & w5804 ;
  assign w8038 = w519 | w8036 ;
  assign w8039 = ( w5805 & w8036 ) | ( w5805 & w8038 ) | ( w8036 & w8038 ) ;
  assign w8040 = ( w5804 & ~w8037 ) | ( w5804 & w8039 ) | ( ~w8037 & w8039 ) ;
  assign w8041 = \pi053 ^ w8040 ;
  assign w8042 = ( w7792 & w7800 ) | ( w7792 & w7828 ) | ( w7800 & w7828 ) ;
  assign w8043 = ( w7801 & w7809 ) | ( w7801 & w7826 ) | ( w7809 & w7826 ) ;
  assign w8044 = ( \pi060 & ~\pi061 ) | ( \pi060 & \pi062 ) | ( ~\pi061 & \pi062 ) ;
  assign w8045 = ( \pi059 & \pi060 ) | ( \pi059 & w8044 ) | ( \pi060 & w8044 ) ;
  assign w8046 = w8044 ^ w8045 ;
  assign w8047 = \pi064 & w8046 ;
  assign w8048 = ( \pi066 & w7813 ) | ( \pi066 & w8047 ) | ( w7813 & w8047 ) ;
  assign w8049 = \pi065 | w8048 ;
  assign w8050 = ( w7811 & w8048 ) | ( w7811 & w8049 ) | ( w8048 & w8049 ) ;
  assign w8051 = w8047 | w8050 ;
  assign w8052 = ~w134 & w7814 ;
  assign w8053 = ( w7814 & w8051 ) | ( w7814 & ~w8052 ) | ( w8051 & ~w8052 ) ;
  assign w8054 = \pi062 ^ w8053 ;
  assign w8055 = w7821 & w8054 ;
  assign w8056 = w7821 ^ w8054 ;
  assign w8057 = ~\pi068 & w7135 ;
  assign w8058 = \pi067 & w7359 ;
  assign w8059 = ( w7135 & ~w8057 ) | ( w7135 & w8058 ) | ( ~w8057 & w8058 ) ;
  assign w8060 = ~\pi069 & w7137 ;
  assign w8061 = w221 | w8059 ;
  assign w8062 = ( w7138 & w8059 ) | ( w7138 & w8061 ) | ( w8059 & w8061 ) ;
  assign w8063 = ( w7137 & ~w8060 ) | ( w7137 & w8062 ) | ( ~w8060 & w8062 ) ;
  assign w8064 = \pi059 ^ w8063 ;
  assign w8065 = ( w8043 & w8056 ) | ( w8043 & w8064 ) | ( w8056 & w8064 ) ;
  assign w8066 = w8043 ^ w8056 ;
  assign w8067 = w8064 ^ w8066 ;
  assign w8068 = ~\pi071 & w6466 ;
  assign w8069 = \pi070 & w6702 ;
  assign w8070 = ( w6466 & ~w8068 ) | ( w6466 & w8069 ) | ( ~w8068 & w8069 ) ;
  assign w8071 = ~\pi072 & w6468 ;
  assign w8072 = w361 | w8070 ;
  assign w8073 = ( w6469 & w8070 ) | ( w6469 & w8072 ) | ( w8070 & w8072 ) ;
  assign w8074 = ( w6468 & ~w8071 ) | ( w6468 & w8073 ) | ( ~w8071 & w8073 ) ;
  assign w8075 = \pi056 ^ w8074 ;
  assign w8076 = w8042 ^ w8067 ;
  assign w8077 = w8075 ^ w8076 ;
  assign w8078 = w8033 ^ w8077 ;
  assign w8079 = w8041 ^ w8078 ;
  assign w8080 = w7842 ^ w8079 ;
  assign w8081 = w8032 ^ w8080 ;
  assign w8082 = w8016 ^ w8081 ;
  assign w8083 = w8024 ^ w8082 ;
  assign w8084 = ~\pi083 & w4141 ;
  assign w8085 = \pi082 & w4334 ;
  assign w8086 = ( w4141 & ~w8084 ) | ( w4141 & w8085 ) | ( ~w8084 & w8085 ) ;
  assign w8087 = ~\pi084 & w4143 ;
  assign w8088 = w1188 | w8086 ;
  assign w8089 = ( w4144 & w8086 ) | ( w4144 & w8088 ) | ( w8086 & w8088 ) ;
  assign w8090 = ( w4143 & ~w8087 ) | ( w4143 & w8089 ) | ( ~w8087 & w8089 ) ;
  assign w8091 = \pi044 ^ w8090 ;
  assign w8092 = w7864 ^ w8083 ;
  assign w8093 = w8091 ^ w8092 ;
  assign w8094 = ~\pi086 & w3635 ;
  assign w8095 = \pi085 & w3817 ;
  assign w8096 = ( w3635 & ~w8094 ) | ( w3635 & w8095 ) | ( ~w8094 & w8095 ) ;
  assign w8097 = ~\pi087 & w3637 ;
  assign w8098 = w1477 | w8096 ;
  assign w8099 = ( w3638 & w8096 ) | ( w3638 & w8098 ) | ( w8096 & w8098 ) ;
  assign w8100 = ( w3637 & ~w8097 ) | ( w3637 & w8099 ) | ( ~w8097 & w8099 ) ;
  assign w8101 = \pi041 ^ w8100 ;
  assign w8102 = w8015 ^ w8093 ;
  assign w8103 = w8101 ^ w8102 ;
  assign w8104 = ~\pi089 & w3178 ;
  assign w8105 = \pi088 & w3340 ;
  assign w8106 = ( w3178 & ~w8104 ) | ( w3178 & w8105 ) | ( ~w8104 & w8105 ) ;
  assign w8107 = ~\pi090 & w3180 ;
  assign w8108 = w1801 | w8106 ;
  assign w8109 = ( w3181 & w8106 ) | ( w3181 & w8108 ) | ( w8106 & w8108 ) ;
  assign w8110 = ( w3180 & ~w8107 ) | ( w3180 & w8109 ) | ( ~w8107 & w8109 ) ;
  assign w8111 = \pi038 ^ w8110 ;
  assign w8112 = ( w7877 & w7885 ) | ( w7877 & w7886 ) | ( w7885 & w7886 ) ;
  assign w8113 = w8103 ^ w8112 ;
  assign w8114 = w8111 ^ w8113 ;
  assign w8115 = ~\pi092 & w2712 ;
  assign w8116 = \pi091 & w2872 ;
  assign w8117 = ( w2712 & ~w8115 ) | ( w2712 & w8116 ) | ( ~w8115 & w8116 ) ;
  assign w8118 = ~\pi093 & w2714 ;
  assign w8119 = w2155 | w8117 ;
  assign w8120 = ( w2715 & w8117 ) | ( w2715 & w8119 ) | ( w8117 & w8119 ) ;
  assign w8121 = ( w2714 & ~w8118 ) | ( w2714 & w8120 ) | ( ~w8118 & w8120 ) ;
  assign w8122 = \pi035 ^ w8121 ;
  assign w8123 = ( w7888 & w7896 ) | ( w7888 & w7897 ) | ( w7896 & w7897 ) ;
  assign w8124 = w8114 ^ w8123 ;
  assign w8125 = w8122 ^ w8124 ;
  assign w8126 = ~\pi095 & w2310 ;
  assign w8127 = \pi094 & w2443 ;
  assign w8128 = ( w2310 & ~w8126 ) | ( w2310 & w8127 ) | ( ~w8126 & w8127 ) ;
  assign w8129 = ~\pi096 & w2312 ;
  assign w8130 = w2546 | w8128 ;
  assign w8131 = ( w2313 & w8128 ) | ( w2313 & w8130 ) | ( w8128 & w8130 ) ;
  assign w8132 = ( w2312 & ~w8129 ) | ( w2312 & w8131 ) | ( ~w8129 & w8131 ) ;
  assign w8133 = \pi032 ^ w8132 ;
  assign w8134 = ( w8014 & w8125 ) | ( w8014 & w8133 ) | ( w8125 & w8133 ) ;
  assign w8135 = w8014 ^ w8125 ;
  assign w8136 = w8133 ^ w8135 ;
  assign w8137 = ~\pi098 & w1944 ;
  assign w8138 = \pi097 & w2072 ;
  assign w8139 = ( w1944 & ~w8137 ) | ( w1944 & w8138 ) | ( ~w8137 & w8138 ) ;
  assign w8140 = ~\pi099 & w1946 ;
  assign w8141 = w2966 | w8139 ;
  assign w8142 = ( w1947 & w8139 ) | ( w1947 & w8141 ) | ( w8139 & w8141 ) ;
  assign w8143 = ( w1946 & ~w8140 ) | ( w1946 & w8142 ) | ( ~w8140 & w8142 ) ;
  assign w8144 = \pi029 ^ w8143 ;
  assign w8145 = ( w7780 & w7909 ) | ( w7780 & w7917 ) | ( w7909 & w7917 ) ;
  assign w8146 = w8136 ^ w8145 ;
  assign w8147 = w8144 ^ w8146 ;
  assign w8148 = ~\pi101 & w1629 ;
  assign w8149 = \pi100 & w1722 ;
  assign w8150 = ( w1629 & ~w8148 ) | ( w1629 & w8149 ) | ( ~w8148 & w8149 ) ;
  assign w8151 = ~\pi102 & w1631 ;
  assign w8152 = w3284 | w8150 ;
  assign w8153 = ( w1632 & w8150 ) | ( w1632 & w8152 ) | ( w8150 & w8152 ) ;
  assign w8154 = ( w1631 & ~w8151 ) | ( w1631 & w8153 ) | ( ~w8151 & w8153 ) ;
  assign w8155 = \pi026 ^ w8154 ;
  assign w8156 = ( w7919 & w7927 ) | ( w7919 & w7928 ) | ( w7927 & w7928 ) ;
  assign w8157 = w8147 ^ w8156 ;
  assign w8158 = w8155 ^ w8157 ;
  assign w8159 = ~\pi104 & w1313 ;
  assign w8160 = \pi103 & w1417 ;
  assign w8161 = ( w1313 & ~w8159 ) | ( w1313 & w8160 ) | ( ~w8159 & w8160 ) ;
  assign w8162 = ~\pi105 & w1315 ;
  assign w8163 = w3905 | w8161 ;
  assign w8164 = ( w1316 & w8161 ) | ( w1316 & w8163 ) | ( w8161 & w8163 ) ;
  assign w8165 = ( w1315 & ~w8162 ) | ( w1315 & w8164 ) | ( ~w8162 & w8164 ) ;
  assign w8166 = \pi023 ^ w8165 ;
  assign w8167 = ( w8013 & w8158 ) | ( w8013 & w8166 ) | ( w8158 & w8166 ) ;
  assign w8168 = w8013 ^ w8158 ;
  assign w8169 = w8166 ^ w8168 ;
  assign w8170 = ~\pi107 & w1044 ;
  assign w8171 = \pi106 & w1138 ;
  assign w8172 = ( w1044 & ~w8170 ) | ( w1044 & w8171 ) | ( ~w8170 & w8171 ) ;
  assign w8173 = ~\pi108 & w1046 ;
  assign w8174 = w4425 | w8172 ;
  assign w8175 = ( w1047 & w8172 ) | ( w1047 & w8174 ) | ( w8172 & w8174 ) ;
  assign w8176 = ( w1046 & ~w8173 ) | ( w1046 & w8175 ) | ( ~w8173 & w8175 ) ;
  assign w8177 = \pi020 ^ w8176 ;
  assign w8178 = w7950 ^ w8169 ;
  assign w8179 = w8177 ^ w8178 ;
  assign w8180 = ~\pi110 & w837 ;
  assign w8181 = \pi109 & w902 ;
  assign w8182 = ( w837 & ~w8180 ) | ( w837 & w8181 ) | ( ~w8180 & w8181 ) ;
  assign w8183 = ~\pi111 & w839 ;
  assign w8184 = w4811 | w8182 ;
  assign w8185 = ( w840 & w8182 ) | ( w840 & w8184 ) | ( w8182 & w8184 ) ;
  assign w8186 = ( w839 & ~w8183 ) | ( w839 & w8185 ) | ( ~w8183 & w8185 ) ;
  assign w8187 = \pi017 ^ w8186 ;
  assign w8188 = w8012 ^ w8179 ;
  assign w8189 = w8187 ^ w8188 ;
  assign w8190 = w8003 ^ w8189 ;
  assign w8191 = w8011 ^ w8190 ;
  assign w8192 = ~\pi116 & w432 ;
  assign w8193 = \pi115 & w486 ;
  assign w8194 = ( w432 & ~w8192 ) | ( w432 & w8193 ) | ( ~w8192 & w8193 ) ;
  assign w8195 = ~\pi117 & w434 ;
  assign w8196 = w6185 | w8194 ;
  assign w8197 = ( w435 & w8194 ) | ( w435 & w8196 ) | ( w8194 & w8196 ) ;
  assign w8198 = ( w434 & ~w8195 ) | ( w434 & w8197 ) | ( ~w8195 & w8197 ) ;
  assign w8199 = \pi011 ^ w8198 ;
  assign w8200 = w8002 ^ w8191 ;
  assign w8201 = w8199 ^ w8200 ;
  assign w8202 = ~\pi119 & w305 ;
  assign w8203 = \pi118 & w328 ;
  assign w8204 = ( w305 & ~w8202 ) | ( w305 & w8203 ) | ( ~w8202 & w8203 ) ;
  assign w8205 = ~\pi120 & w307 ;
  assign w8206 = w6634 | w8204 ;
  assign w8207 = ( w308 & w8204 ) | ( w308 & w8206 ) | ( w8204 & w8206 ) ;
  assign w8208 = ( w307 & ~w8205 ) | ( w307 & w8207 ) | ( ~w8205 & w8207 ) ;
  assign w8209 = \pi008 ^ w8208 ;
  assign w8210 = ~\pi122 & w189 ;
  assign w8211 = \pi121 & w229 ;
  assign w8212 = ( w189 & ~w8210 ) | ( w189 & w8211 ) | ( ~w8210 & w8211 ) ;
  assign w8213 = ~\pi123 & w191 ;
  assign w8214 = w7516 | w8212 ;
  assign w8215 = ( w192 & w8212 ) | ( w192 & w8214 ) | ( w8212 & w8214 ) ;
  assign w8216 = ( w191 & ~w8213 ) | ( w191 & w8215 ) | ( ~w8213 & w8215 ) ;
  assign w8217 = \pi005 ^ w8216 ;
  assign w8218 = w8201 ^ w8217 ;
  assign w8219 = w8209 ^ w8218 ;
  assign w8220 = ( w7759 & w7966 ) | ( w7759 & w7967 ) | ( w7966 & w7967 ) ;
  assign w8221 = ( ~\pi002 & \pi125 ) | ( ~\pi002 & \pi126 ) | ( \pi125 & \pi126 ) ;
  assign w8222 = \pi000 ^ w8221 ;
  assign w8223 = ( \pi002 & \pi126 ) | ( \pi002 & ~w8222 ) | ( \pi126 & ~w8222 ) ;
  assign w8224 = ( \pi002 & \pi125 ) | ( \pi002 & w8222 ) | ( \pi125 & w8222 ) ;
  assign w8225 = \pi001 & w8224 ;
  assign w8226 = ( ~\pi000 & \pi124 ) | ( ~\pi000 & w8225 ) | ( \pi124 & w8225 ) ;
  assign w8227 = ( \pi001 & \pi002 ) | ( \pi001 & ~w8226 ) | ( \pi002 & ~w8226 ) ;
  assign w8228 = ( w8223 & w8225 ) | ( w8223 & ~w8227 ) | ( w8225 & ~w8227 ) ;
  assign w8229 = ( \pi124 & \pi125 ) | ( \pi124 & w7986 ) | ( \pi125 & w7986 ) ;
  assign w8230 = \pi125 ^ w8229 ;
  assign w8231 = \pi126 ^ w8230 ;
  assign w8232 = \pi002 ^ w8228 ;
  assign w8233 = \pi000 & ~w8228 ;
  assign w8234 = w8231 & w8233 ;
  assign w8235 = \pi001 ^ w8234 ;
  assign w8236 = ( \pi001 & w8232 ) | ( \pi001 & ~w8235 ) | ( w8232 & ~w8235 ) ;
  assign w8237 = w8219 ^ w8220 ;
  assign w8238 = w8236 ^ w8237 ;
  assign w8239 = w8000 ^ w8001 ;
  assign w8240 = w8238 ^ w8239 ;
  assign w8241 = ( w8003 & w8011 ) | ( w8003 & w8189 ) | ( w8011 & w8189 ) ;
  assign w8242 = ~\pi114 & w601 ;
  assign w8243 = \pi113 & w683 ;
  assign w8244 = ( w601 & ~w8242 ) | ( w601 & w8243 ) | ( ~w8242 & w8243 ) ;
  assign w8245 = ~\pi115 & w603 ;
  assign w8246 = w5585 | w8244 ;
  assign w8247 = ( w604 & w8244 ) | ( w604 & w8246 ) | ( w8244 & w8246 ) ;
  assign w8248 = ( w603 & ~w8245 ) | ( w603 & w8247 ) | ( ~w8245 & w8247 ) ;
  assign w8249 = \pi014 ^ w8248 ;
  assign w8250 = ( w8012 & w8179 ) | ( w8012 & w8187 ) | ( w8179 & w8187 ) ;
  assign w8251 = ~\pi111 & w837 ;
  assign w8252 = \pi110 & w902 ;
  assign w8253 = ( w837 & ~w8251 ) | ( w837 & w8252 ) | ( ~w8251 & w8252 ) ;
  assign w8254 = ~\pi112 & w839 ;
  assign w8255 = w4999 | w8253 ;
  assign w8256 = ( w840 & w8253 ) | ( w840 & w8255 ) | ( w8253 & w8255 ) ;
  assign w8257 = ( w839 & ~w8254 ) | ( w839 & w8256 ) | ( ~w8254 & w8256 ) ;
  assign w8258 = \pi017 ^ w8257 ;
  assign w8259 = ( w7950 & w8169 ) | ( w7950 & w8177 ) | ( w8169 & w8177 ) ;
  assign w8260 = ~\pi108 & w1044 ;
  assign w8261 = \pi107 & w1138 ;
  assign w8262 = ( w1044 & ~w8260 ) | ( w1044 & w8261 ) | ( ~w8260 & w8261 ) ;
  assign w8263 = ~\pi109 & w1046 ;
  assign w8264 = w4599 | w8262 ;
  assign w8265 = ( w1047 & w8262 ) | ( w1047 & w8264 ) | ( w8262 & w8264 ) ;
  assign w8266 = ( w1046 & ~w8263 ) | ( w1046 & w8265 ) | ( ~w8263 & w8265 ) ;
  assign w8267 = \pi020 ^ w8266 ;
  assign w8268 = ~\pi105 & w1313 ;
  assign w8269 = \pi104 & w1417 ;
  assign w8270 = ( w1313 & ~w8268 ) | ( w1313 & w8269 ) | ( ~w8268 & w8269 ) ;
  assign w8271 = ~\pi106 & w1315 ;
  assign w8272 = w4068 | w8270 ;
  assign w8273 = ( w1316 & w8270 ) | ( w1316 & w8272 ) | ( w8270 & w8272 ) ;
  assign w8274 = ( w1315 & ~w8271 ) | ( w1315 & w8273 ) | ( ~w8271 & w8273 ) ;
  assign w8275 = \pi023 ^ w8274 ;
  assign w8276 = ( w8147 & w8155 ) | ( w8147 & w8156 ) | ( w8155 & w8156 ) ;
  assign w8277 = ( w8136 & w8144 ) | ( w8136 & w8145 ) | ( w8144 & w8145 ) ;
  assign w8278 = ~\pi096 & w2310 ;
  assign w8279 = \pi095 & w2443 ;
  assign w8280 = ( w2310 & ~w8278 ) | ( w2310 & w8279 ) | ( ~w8278 & w8279 ) ;
  assign w8281 = ~\pi097 & w2312 ;
  assign w8282 = w2673 | w8280 ;
  assign w8283 = ( w2313 & w8280 ) | ( w2313 & w8282 ) | ( w8280 & w8282 ) ;
  assign w8284 = ( w2312 & ~w8281 ) | ( w2312 & w8283 ) | ( ~w8281 & w8283 ) ;
  assign w8285 = \pi032 ^ w8284 ;
  assign w8286 = ( w7864 & w8083 ) | ( w7864 & w8091 ) | ( w8083 & w8091 ) ;
  assign w8287 = ~\pi084 & w4141 ;
  assign w8288 = \pi083 & w4334 ;
  assign w8289 = ( w4141 & ~w8287 ) | ( w4141 & w8288 ) | ( ~w8287 & w8288 ) ;
  assign w8290 = ~\pi085 & w4143 ;
  assign w8291 = w1274 | w8289 ;
  assign w8292 = ( w4144 & w8289 ) | ( w4144 & w8291 ) | ( w8289 & w8291 ) ;
  assign w8293 = ( w4143 & ~w8290 ) | ( w4143 & w8292 ) | ( ~w8290 & w8292 ) ;
  assign w8294 = \pi044 ^ w8293 ;
  assign w8295 = ( w8016 & w8024 ) | ( w8016 & w8081 ) | ( w8024 & w8081 ) ;
  assign w8296 = ~\pi078 & w5209 ;
  assign w8297 = \pi077 & w5433 ;
  assign w8298 = ( w5209 & ~w8296 ) | ( w5209 & w8297 ) | ( ~w8296 & w8297 ) ;
  assign w8299 = ~\pi079 & w5211 ;
  assign w8300 = w730 | w8298 ;
  assign w8301 = ( w5212 & w8298 ) | ( w5212 & w8300 ) | ( w8298 & w8300 ) ;
  assign w8302 = ( w5211 & ~w8299 ) | ( w5211 & w8301 ) | ( ~w8299 & w8301 ) ;
  assign w8303 = \pi050 ^ w8302 ;
  assign w8304 = ( w8033 & w8041 ) | ( w8033 & w8077 ) | ( w8041 & w8077 ) ;
  assign w8305 = ( w8042 & w8067 ) | ( w8042 & w8075 ) | ( w8067 & w8075 ) ;
  assign w8306 = ~\pi072 & w6466 ;
  assign w8307 = \pi071 & w6702 ;
  assign w8308 = ( w6466 & ~w8306 ) | ( w6466 & w8307 ) | ( ~w8306 & w8307 ) ;
  assign w8309 = ~\pi073 & w6468 ;
  assign w8310 = w404 | w8308 ;
  assign w8311 = ( w6469 & w8308 ) | ( w6469 & w8310 ) | ( w8308 & w8310 ) ;
  assign w8312 = ( w6468 & ~w8309 ) | ( w6468 & w8311 ) | ( ~w8309 & w8311 ) ;
  assign w8313 = \pi056 ^ w8312 ;
  assign w8314 = ~\pi066 & w7811 ;
  assign w8315 = \pi065 & w8046 ;
  assign w8316 = ( w7811 & ~w8314 ) | ( w7811 & w8315 ) | ( ~w8314 & w8315 ) ;
  assign w8317 = ~\pi067 & w7813 ;
  assign w8318 = w160 | w8316 ;
  assign w8319 = ( w7814 & w8316 ) | ( w7814 & w8318 ) | ( w8316 & w8318 ) ;
  assign w8320 = ( w7813 & ~w8317 ) | ( w7813 & w8319 ) | ( ~w8317 & w8319 ) ;
  assign w8321 = \pi062 ^ w8320 ;
  assign w8322 = w8055 ^ w8321 ;
  assign w8323 = \pi062 ^ \pi063 ;
  assign w8324 = \pi064 & w8323 ;
  assign w8325 = w8322 ^ w8324 ;
  assign w8326 = ~\pi069 & w7135 ;
  assign w8327 = \pi068 & w7359 ;
  assign w8328 = ( w7135 & ~w8326 ) | ( w7135 & w8327 ) | ( ~w8326 & w8327 ) ;
  assign w8329 = ~\pi070 & w7137 ;
  assign w8330 = w271 | w8328 ;
  assign w8331 = ( w7138 & w8328 ) | ( w7138 & w8330 ) | ( w8328 & w8330 ) ;
  assign w8332 = ( w7137 & ~w8329 ) | ( w7137 & w8331 ) | ( ~w8329 & w8331 ) ;
  assign w8333 = \pi059 ^ w8332 ;
  assign w8334 = w8065 ^ w8325 ;
  assign w8335 = w8333 ^ w8334 ;
  assign w8336 = w8305 ^ w8335 ;
  assign w8337 = w8313 ^ w8336 ;
  assign w8338 = ~\pi075 & w5802 ;
  assign w8339 = \pi074 & w6052 ;
  assign w8340 = ( w5802 & ~w8338 ) | ( w5802 & w8339 ) | ( ~w8338 & w8339 ) ;
  assign w8341 = ~\pi076 & w5804 ;
  assign w8342 = w538 | w8340 ;
  assign w8343 = ( w5805 & w8340 ) | ( w5805 & w8342 ) | ( w8340 & w8342 ) ;
  assign w8344 = ( w5804 & ~w8341 ) | ( w5804 & w8343 ) | ( ~w8341 & w8343 ) ;
  assign w8345 = \pi053 ^ w8344 ;
  assign w8346 = w8304 ^ w8337 ;
  assign w8347 = w8345 ^ w8346 ;
  assign w8348 = ( w7842 & w8032 ) | ( w7842 & w8079 ) | ( w8032 & w8079 ) ;
  assign w8349 = w8347 ^ w8348 ;
  assign w8350 = w8303 ^ w8349 ;
  assign w8351 = ~\pi081 & w4654 ;
  assign w8352 = \pi080 & w4876 ;
  assign w8353 = ( w4654 & ~w8351 ) | ( w4654 & w8352 ) | ( ~w8351 & w8352 ) ;
  assign w8354 = ~\pi082 & w4656 ;
  assign w8355 = w1008 | w8353 ;
  assign w8356 = ( w4657 & w8353 ) | ( w4657 & w8355 ) | ( w8353 & w8355 ) ;
  assign w8357 = ( w4656 & ~w8354 ) | ( w4656 & w8356 ) | ( ~w8354 & w8356 ) ;
  assign w8358 = \pi047 ^ w8357 ;
  assign w8359 = w8295 ^ w8350 ;
  assign w8360 = w8358 ^ w8359 ;
  assign w8361 = w8286 ^ w8360 ;
  assign w8362 = w8294 ^ w8361 ;
  assign w8363 = ~\pi087 & w3635 ;
  assign w8364 = \pi086 & w3817 ;
  assign w8365 = ( w3635 & ~w8363 ) | ( w3635 & w8364 ) | ( ~w8363 & w8364 ) ;
  assign w8366 = ~\pi088 & w3637 ;
  assign w8367 = w1574 | w8365 ;
  assign w8368 = ( w3638 & w8365 ) | ( w3638 & w8367 ) | ( w8365 & w8367 ) ;
  assign w8369 = ( w3637 & ~w8366 ) | ( w3637 & w8368 ) | ( ~w8366 & w8368 ) ;
  assign w8370 = \pi041 ^ w8369 ;
  assign w8371 = ( w8015 & w8093 ) | ( w8015 & w8101 ) | ( w8093 & w8101 ) ;
  assign w8372 = w8362 ^ w8371 ;
  assign w8373 = w8370 ^ w8372 ;
  assign w8374 = ~\pi090 & w3178 ;
  assign w8375 = \pi089 & w3340 ;
  assign w8376 = ( w3178 & ~w8374 ) | ( w3178 & w8375 ) | ( ~w8374 & w8375 ) ;
  assign w8377 = ~\pi091 & w3180 ;
  assign w8378 = w1908 | w8376 ;
  assign w8379 = ( w3181 & w8376 ) | ( w3181 & w8378 ) | ( w8376 & w8378 ) ;
  assign w8380 = ( w3180 & ~w8377 ) | ( w3180 & w8379 ) | ( ~w8377 & w8379 ) ;
  assign w8381 = \pi038 ^ w8380 ;
  assign w8382 = ( w8103 & w8111 ) | ( w8103 & w8112 ) | ( w8111 & w8112 ) ;
  assign w8383 = w8373 ^ w8382 ;
  assign w8384 = w8381 ^ w8383 ;
  assign w8385 = ~\pi093 & w2712 ;
  assign w8386 = \pi092 & w2872 ;
  assign w8387 = ( w2712 & ~w8385 ) | ( w2712 & w8386 ) | ( ~w8385 & w8386 ) ;
  assign w8388 = ~\pi094 & w2714 ;
  assign w8389 = w2274 | w8387 ;
  assign w8390 = ( w2715 & w8387 ) | ( w2715 & w8389 ) | ( w8387 & w8389 ) ;
  assign w8391 = ( w2714 & ~w8388 ) | ( w2714 & w8390 ) | ( ~w8388 & w8390 ) ;
  assign w8392 = \pi035 ^ w8391 ;
  assign w8393 = ( w8114 & w8122 ) | ( w8114 & w8123 ) | ( w8122 & w8123 ) ;
  assign w8394 = w8384 ^ w8393 ;
  assign w8395 = w8392 ^ w8394 ;
  assign w8396 = w8134 ^ w8395 ;
  assign w8397 = w8285 ^ w8396 ;
  assign w8398 = ~\pi099 & w1944 ;
  assign w8399 = \pi098 & w2072 ;
  assign w8400 = ( w1944 & ~w8398 ) | ( w1944 & w8399 ) | ( ~w8398 & w8399 ) ;
  assign w8401 = ~\pi100 & w1946 ;
  assign w8402 = w3104 | w8400 ;
  assign w8403 = ( w1947 & w8400 ) | ( w1947 & w8402 ) | ( w8400 & w8402 ) ;
  assign w8404 = ( w1946 & ~w8401 ) | ( w1946 & w8403 ) | ( ~w8401 & w8403 ) ;
  assign w8405 = \pi029 ^ w8404 ;
  assign w8406 = w8277 ^ w8397 ;
  assign w8407 = w8405 ^ w8406 ;
  assign w8408 = ~\pi102 & w1629 ;
  assign w8409 = \pi101 & w1722 ;
  assign w8410 = ( w1629 & ~w8408 ) | ( w1629 & w8409 ) | ( ~w8408 & w8409 ) ;
  assign w8411 = ~\pi103 & w1631 ;
  assign w8412 = w3437 | w8410 ;
  assign w8413 = ( w1632 & w8410 ) | ( w1632 & w8412 ) | ( w8410 & w8412 ) ;
  assign w8414 = ( w1631 & ~w8411 ) | ( w1631 & w8413 ) | ( ~w8411 & w8413 ) ;
  assign w8415 = \pi026 ^ w8414 ;
  assign w8416 = w8276 ^ w8407 ;
  assign w8417 = w8415 ^ w8416 ;
  assign w8418 = w8167 ^ w8417 ;
  assign w8419 = w8275 ^ w8418 ;
  assign w8420 = w8259 ^ w8419 ;
  assign w8421 = w8267 ^ w8420 ;
  assign w8422 = w8250 ^ w8421 ;
  assign w8423 = w8258 ^ w8422 ;
  assign w8424 = w8241 ^ w8423 ;
  assign w8425 = w8249 ^ w8424 ;
  assign w8426 = ~\pi117 & w432 ;
  assign w8427 = \pi116 & w486 ;
  assign w8428 = ( w432 & ~w8426 ) | ( w432 & w8427 ) | ( ~w8426 & w8427 ) ;
  assign w8429 = ~\pi118 & w434 ;
  assign w8430 = w6206 | w8428 ;
  assign w8431 = ( w435 & w8428 ) | ( w435 & w8430 ) | ( w8428 & w8430 ) ;
  assign w8432 = ( w434 & ~w8429 ) | ( w434 & w8431 ) | ( ~w8429 & w8431 ) ;
  assign w8433 = \pi011 ^ w8432 ;
  assign w8434 = ( w8002 & w8191 ) | ( w8002 & w8199 ) | ( w8191 & w8199 ) ;
  assign w8435 = w8425 ^ w8434 ;
  assign w8436 = w8433 ^ w8435 ;
  assign w8437 = ~\pi120 & w305 ;
  assign w8438 = \pi119 & w328 ;
  assign w8439 = ( w305 & ~w8437 ) | ( w305 & w8438 ) | ( ~w8437 & w8438 ) ;
  assign w8440 = ~\pi121 & w307 ;
  assign w8441 = w7050 | w8439 ;
  assign w8442 = ( w308 & w8439 ) | ( w308 & w8441 ) | ( w8439 & w8441 ) ;
  assign w8443 = ( w307 & ~w8440 ) | ( w307 & w8442 ) | ( ~w8440 & w8442 ) ;
  assign w8444 = \pi008 ^ w8443 ;
  assign w8445 = ~\pi123 & w189 ;
  assign w8446 = \pi122 & w229 ;
  assign w8447 = ( w189 & ~w8445 ) | ( w189 & w8446 ) | ( ~w8445 & w8446 ) ;
  assign w8448 = ~\pi124 & w191 ;
  assign w8449 = w7538 | w8447 ;
  assign w8450 = ( w192 & w8447 ) | ( w192 & w8449 ) | ( w8447 & w8449 ) ;
  assign w8451 = ( w191 & ~w8448 ) | ( w191 & w8450 ) | ( ~w8448 & w8450 ) ;
  assign w8452 = \pi005 ^ w8451 ;
  assign w8453 = w8436 ^ w8452 ;
  assign w8454 = w8444 ^ w8453 ;
  assign w8455 = ( w8201 & w8209 ) | ( w8201 & w8217 ) | ( w8209 & w8217 ) ;
  assign w8456 = ( ~\pi002 & \pi126 ) | ( ~\pi002 & \pi127 ) | ( \pi126 & \pi127 ) ;
  assign w8457 = \pi000 ^ w8456 ;
  assign w8458 = ( \pi002 & \pi127 ) | ( \pi002 & ~w8457 ) | ( \pi127 & ~w8457 ) ;
  assign w8459 = ( \pi002 & \pi126 ) | ( \pi002 & w8457 ) | ( \pi126 & w8457 ) ;
  assign w8460 = \pi001 & w8459 ;
  assign w8461 = ( ~\pi000 & \pi125 ) | ( ~\pi000 & w8460 ) | ( \pi125 & w8460 ) ;
  assign w8462 = ( \pi001 & \pi002 ) | ( \pi001 & ~w8461 ) | ( \pi002 & ~w8461 ) ;
  assign w8463 = ( w8458 & w8460 ) | ( w8458 & ~w8462 ) | ( w8460 & ~w8462 ) ;
  assign w8464 = ( \pi125 & \pi126 ) | ( \pi125 & w8229 ) | ( \pi126 & w8229 ) ;
  assign w8465 = \pi126 ^ w8464 ;
  assign w8466 = \pi127 ^ w8465 ;
  assign w8467 = \pi002 ^ w8463 ;
  assign w8468 = \pi000 & ~w8463 ;
  assign w8469 = w8466 & w8468 ;
  assign w8470 = \pi001 ^ w8469 ;
  assign w8471 = ( \pi001 & w8467 ) | ( \pi001 & ~w8470 ) | ( w8467 & ~w8470 ) ;
  assign w8472 = w8454 ^ w8455 ;
  assign w8473 = w8471 ^ w8472 ;
  assign w8474 = ( w8219 & w8220 ) | ( w8219 & w8236 ) | ( w8220 & w8236 ) ;
  assign w8475 = ( w8000 & w8001 ) | ( w8000 & w8238 ) | ( w8001 & w8238 ) ;
  assign w8476 = w8473 ^ w8475 ;
  assign w8477 = w8474 ^ w8476 ;
  assign w8478 = ( w8473 & w8474 ) | ( w8473 & w8475 ) | ( w8474 & w8475 ) ;
  assign w8479 = ( w8454 & w8455 ) | ( w8454 & w8471 ) | ( w8455 & w8471 ) ;
  assign w8480 = ( \pi126 & \pi127 ) | ( \pi126 & w8464 ) | ( \pi127 & w8464 ) ;
  assign w8481 = \pi127 & w8480 ;
  assign w8482 = \pi000 & \pi002 ;
  assign w8483 = \pi000 & w8480 ;
  assign w8484 = \pi127 ^ w8483 ;
  assign w8485 = \pi002 | w8484 ;
  assign w8486 = \pi001 & w8485 ;
  assign w8487 = ( \pi002 & \pi127 ) | ( \pi002 & w8482 ) | ( \pi127 & w8482 ) ;
  assign w8488 = ( w8482 & w8486 ) | ( w8482 & ~w8487 ) | ( w8486 & ~w8487 ) ;
  assign w8489 = ~\pi001 & \pi002 ;
  assign w8490 = ( \pi126 & \pi127 ) | ( \pi126 & ~w8464 ) | ( \pi127 & ~w8464 ) ;
  assign w8491 = \pi000 & w8490 ;
  assign w8492 = \pi126 ^ w8491 ;
  assign w8493 = w8489 & ~w8492 ;
  assign w8494 = w8488 | w8493 ;
  assign w8495 = ( w8436 & w8444 ) | ( w8436 & w8452 ) | ( w8444 & w8452 ) ;
  assign w8496 = ( w8425 & w8433 ) | ( w8425 & w8434 ) | ( w8433 & w8434 ) ;
  assign w8497 = ~\pi118 & w432 ;
  assign w8498 = \pi117 & w486 ;
  assign w8499 = ( w432 & ~w8497 ) | ( w432 & w8498 ) | ( ~w8497 & w8498 ) ;
  assign w8500 = ~\pi119 & w434 ;
  assign w8501 = w6616 | w8499 ;
  assign w8502 = ( w435 & w8499 ) | ( w435 & w8501 ) | ( w8499 & w8501 ) ;
  assign w8503 = ( w434 & ~w8500 ) | ( w434 & w8502 ) | ( ~w8500 & w8502 ) ;
  assign w8504 = \pi011 ^ w8503 ;
  assign w8505 = ( w8241 & w8249 ) | ( w8241 & w8423 ) | ( w8249 & w8423 ) ;
  assign w8506 = ~\pi115 & w601 ;
  assign w8507 = \pi114 & w683 ;
  assign w8508 = ( w601 & ~w8506 ) | ( w601 & w8507 ) | ( ~w8506 & w8507 ) ;
  assign w8509 = ~\pi116 & w603 ;
  assign w8510 = w5976 | w8508 ;
  assign w8511 = ( w604 & w8508 ) | ( w604 & w8510 ) | ( w8508 & w8510 ) ;
  assign w8512 = ( w603 & ~w8509 ) | ( w603 & w8511 ) | ( ~w8509 & w8511 ) ;
  assign w8513 = \pi014 ^ w8512 ;
  assign w8514 = ( w8250 & w8258 ) | ( w8250 & w8421 ) | ( w8258 & w8421 ) ;
  assign w8515 = ~\pi112 & w837 ;
  assign w8516 = \pi111 & w902 ;
  assign w8517 = ( w837 & ~w8515 ) | ( w837 & w8516 ) | ( ~w8515 & w8516 ) ;
  assign w8518 = ~\pi113 & w839 ;
  assign w8519 = w5366 | w8517 ;
  assign w8520 = ( w840 & w8517 ) | ( w840 & w8519 ) | ( w8517 & w8519 ) ;
  assign w8521 = ( w839 & ~w8518 ) | ( w839 & w8520 ) | ( ~w8518 & w8520 ) ;
  assign w8522 = \pi017 ^ w8521 ;
  assign w8523 = ( w8259 & w8267 ) | ( w8259 & w8419 ) | ( w8267 & w8419 ) ;
  assign w8524 = ~\pi109 & w1044 ;
  assign w8525 = \pi108 & w1138 ;
  assign w8526 = ( w1044 & ~w8524 ) | ( w1044 & w8525 ) | ( ~w8524 & w8525 ) ;
  assign w8527 = ~\pi110 & w1046 ;
  assign w8528 = w4792 | w8526 ;
  assign w8529 = ( w1047 & w8526 ) | ( w1047 & w8528 ) | ( w8526 & w8528 ) ;
  assign w8530 = ( w1046 & ~w8527 ) | ( w1046 & w8529 ) | ( ~w8527 & w8529 ) ;
  assign w8531 = \pi020 ^ w8530 ;
  assign w8532 = ( w8167 & w8275 ) | ( w8167 & w8417 ) | ( w8275 & w8417 ) ;
  assign w8533 = ~\pi097 & w2310 ;
  assign w8534 = \pi096 & w2443 ;
  assign w8535 = ( w2310 & ~w8533 ) | ( w2310 & w8534 ) | ( ~w8533 & w8534 ) ;
  assign w8536 = ~\pi098 & w2312 ;
  assign w8537 = w2824 | w8535 ;
  assign w8538 = ( w2313 & w8535 ) | ( w2313 & w8537 ) | ( w8535 & w8537 ) ;
  assign w8539 = ( w2312 & ~w8536 ) | ( w2312 & w8538 ) | ( ~w8536 & w8538 ) ;
  assign w8540 = \pi032 ^ w8539 ;
  assign w8541 = ~\pi085 & w4141 ;
  assign w8542 = \pi084 & w4334 ;
  assign w8543 = ( w4141 & ~w8541 ) | ( w4141 & w8542 ) | ( ~w8541 & w8542 ) ;
  assign w8544 = ~\pi086 & w4143 ;
  assign w8545 = w1379 | w8543 ;
  assign w8546 = ( w4144 & w8543 ) | ( w4144 & w8545 ) | ( w8543 & w8545 ) ;
  assign w8547 = ( w4143 & ~w8544 ) | ( w4143 & w8546 ) | ( ~w8544 & w8546 ) ;
  assign w8548 = \pi044 ^ w8547 ;
  assign w8549 = ~\pi079 & w5209 ;
  assign w8550 = \pi078 & w5433 ;
  assign w8551 = ( w5209 & ~w8549 ) | ( w5209 & w8550 ) | ( ~w8549 & w8550 ) ;
  assign w8552 = ~\pi080 & w5211 ;
  assign w8553 = w794 | w8551 ;
  assign w8554 = ( w5212 & w8551 ) | ( w5212 & w8553 ) | ( w8551 & w8553 ) ;
  assign w8555 = ( w5211 & ~w8552 ) | ( w5211 & w8554 ) | ( ~w8552 & w8554 ) ;
  assign w8556 = \pi050 ^ w8555 ;
  assign w8557 = ~\pi073 & w6466 ;
  assign w8558 = \pi072 & w6702 ;
  assign w8559 = ( w6466 & ~w8557 ) | ( w6466 & w8558 ) | ( ~w8557 & w8558 ) ;
  assign w8560 = ~\pi074 & w6468 ;
  assign w8561 = w465 | w8559 ;
  assign w8562 = ( w6469 & w8559 ) | ( w6469 & w8561 ) | ( w8559 & w8561 ) ;
  assign w8563 = ( w6468 & ~w8560 ) | ( w6468 & w8562 ) | ( ~w8560 & w8562 ) ;
  assign w8564 = \pi056 ^ w8563 ;
  assign w8565 = ( w8065 & w8325 ) | ( w8065 & w8333 ) | ( w8325 & w8333 ) ;
  assign w8566 = ~\pi067 & w7811 ;
  assign w8567 = \pi066 & w8046 ;
  assign w8568 = ( w7811 & ~w8566 ) | ( w7811 & w8567 ) | ( ~w8566 & w8567 ) ;
  assign w8569 = ~\pi068 & w7813 ;
  assign w8570 = w182 | w8568 ;
  assign w8571 = ( w7814 & w8568 ) | ( w7814 & w8570 ) | ( w8568 & w8570 ) ;
  assign w8572 = ( w7813 & ~w8569 ) | ( w7813 & w8571 ) | ( ~w8569 & w8571 ) ;
  assign w8573 = \pi062 ^ w8572 ;
  assign w8574 = ( w8055 & w8321 ) | ( w8055 & w8324 ) | ( w8321 & w8324 ) ;
  assign w8575 = w8573 ^ w8574 ;
  assign w8576 = ( \pi062 & \pi063 ) | ( \pi062 & \pi065 ) | ( \pi063 & \pi065 ) ;
  assign w8577 = \pi063 & ~\pi064 ;
  assign w8578 = \pi062 & w8577 ;
  assign w8579 = w8576 ^ w8578 ;
  assign w8580 = w8575 ^ w8579 ;
  assign w8581 = ~\pi070 & w7135 ;
  assign w8582 = \pi069 & w7359 ;
  assign w8583 = ( w7135 & ~w8581 ) | ( w7135 & w8582 ) | ( ~w8581 & w8582 ) ;
  assign w8584 = ~\pi071 & w7137 ;
  assign w8585 = w290 | w8583 ;
  assign w8586 = ( w7138 & w8583 ) | ( w7138 & w8585 ) | ( w8583 & w8585 ) ;
  assign w8587 = ( w7137 & ~w8584 ) | ( w7137 & w8586 ) | ( ~w8584 & w8586 ) ;
  assign w8588 = \pi059 ^ w8587 ;
  assign w8589 = w8565 ^ w8580 ;
  assign w8590 = w8588 ^ w8589 ;
  assign w8591 = ( w8305 & w8313 ) | ( w8305 & w8335 ) | ( w8313 & w8335 ) ;
  assign w8592 = w8590 ^ w8591 ;
  assign w8593 = w8564 ^ w8592 ;
  assign w8594 = ~\pi076 & w5802 ;
  assign w8595 = \pi075 & w6052 ;
  assign w8596 = ( w5802 & ~w8594 ) | ( w5802 & w8595 ) | ( ~w8594 & w8595 ) ;
  assign w8597 = ~\pi077 & w5804 ;
  assign w8598 = w644 | w8596 ;
  assign w8599 = ( w5805 & w8596 ) | ( w5805 & w8598 ) | ( w8596 & w8598 ) ;
  assign w8600 = ( w5804 & ~w8597 ) | ( w5804 & w8599 ) | ( ~w8597 & w8599 ) ;
  assign w8601 = \pi053 ^ w8600 ;
  assign w8602 = ( w8304 & w8337 ) | ( w8304 & w8345 ) | ( w8337 & w8345 ) ;
  assign w8603 = w8593 ^ w8602 ;
  assign w8604 = w8601 ^ w8603 ;
  assign w8605 = ( w8303 & w8347 ) | ( w8303 & w8348 ) | ( w8347 & w8348 ) ;
  assign w8606 = w8604 ^ w8605 ;
  assign w8607 = w8556 ^ w8606 ;
  assign w8608 = ~\pi082 & w4654 ;
  assign w8609 = \pi081 & w4876 ;
  assign w8610 = ( w4654 & ~w8608 ) | ( w4654 & w8609 ) | ( ~w8608 & w8609 ) ;
  assign w8611 = ~\pi083 & w4656 ;
  assign w8612 = w1099 | w8610 ;
  assign w8613 = ( w4657 & w8610 ) | ( w4657 & w8612 ) | ( w8610 & w8612 ) ;
  assign w8614 = ( w4656 & ~w8611 ) | ( w4656 & w8613 ) | ( ~w8611 & w8613 ) ;
  assign w8615 = \pi047 ^ w8614 ;
  assign w8616 = ( w8295 & w8350 ) | ( w8295 & w8358 ) | ( w8350 & w8358 ) ;
  assign w8617 = w8607 ^ w8616 ;
  assign w8618 = w8615 ^ w8617 ;
  assign w8619 = ( w8286 & w8294 ) | ( w8286 & w8360 ) | ( w8294 & w8360 ) ;
  assign w8620 = w8618 ^ w8619 ;
  assign w8621 = w8548 ^ w8620 ;
  assign w8622 = ~\pi088 & w3635 ;
  assign w8623 = \pi087 & w3817 ;
  assign w8624 = ( w3635 & ~w8622 ) | ( w3635 & w8623 ) | ( ~w8622 & w8623 ) ;
  assign w8625 = ~\pi089 & w3637 ;
  assign w8626 = w1595 | w8624 ;
  assign w8627 = ( w3638 & w8624 ) | ( w3638 & w8626 ) | ( w8624 & w8626 ) ;
  assign w8628 = ( w3637 & ~w8625 ) | ( w3637 & w8627 ) | ( ~w8625 & w8627 ) ;
  assign w8629 = \pi041 ^ w8628 ;
  assign w8630 = ( w8362 & w8370 ) | ( w8362 & w8371 ) | ( w8370 & w8371 ) ;
  assign w8631 = w8621 ^ w8630 ;
  assign w8632 = w8629 ^ w8631 ;
  assign w8633 = ~\pi091 & w3178 ;
  assign w8634 = \pi090 & w3340 ;
  assign w8635 = ( w3178 & ~w8633 ) | ( w3178 & w8634 ) | ( ~w8633 & w8634 ) ;
  assign w8636 = ~\pi092 & w3180 ;
  assign w8637 = w2033 | w8635 ;
  assign w8638 = ( w3181 & w8635 ) | ( w3181 & w8637 ) | ( w8635 & w8637 ) ;
  assign w8639 = ( w3180 & ~w8636 ) | ( w3180 & w8638 ) | ( ~w8636 & w8638 ) ;
  assign w8640 = \pi038 ^ w8639 ;
  assign w8641 = ( w8373 & w8381 ) | ( w8373 & w8382 ) | ( w8381 & w8382 ) ;
  assign w8642 = w8632 ^ w8641 ;
  assign w8643 = w8640 ^ w8642 ;
  assign w8644 = ~\pi094 & w2712 ;
  assign w8645 = \pi093 & w2872 ;
  assign w8646 = ( w2712 & ~w8644 ) | ( w2712 & w8645 ) | ( ~w8644 & w8645 ) ;
  assign w8647 = ~\pi095 & w2714 ;
  assign w8648 = w2409 | w8646 ;
  assign w8649 = ( w2715 & w8646 ) | ( w2715 & w8648 ) | ( w8646 & w8648 ) ;
  assign w8650 = ( w2714 & ~w8647 ) | ( w2714 & w8649 ) | ( ~w8647 & w8649 ) ;
  assign w8651 = \pi035 ^ w8650 ;
  assign w8652 = ( w8384 & w8392 ) | ( w8384 & w8393 ) | ( w8392 & w8393 ) ;
  assign w8653 = w8643 ^ w8652 ;
  assign w8654 = w8651 ^ w8653 ;
  assign w8655 = ( w8134 & w8285 ) | ( w8134 & w8395 ) | ( w8285 & w8395 ) ;
  assign w8656 = w8654 ^ w8655 ;
  assign w8657 = w8540 ^ w8656 ;
  assign w8658 = ~\pi100 & w1944 ;
  assign w8659 = \pi099 & w2072 ;
  assign w8660 = ( w1944 & ~w8658 ) | ( w1944 & w8659 ) | ( ~w8658 & w8659 ) ;
  assign w8661 = ~\pi101 & w1946 ;
  assign w8662 = w3264 | w8660 ;
  assign w8663 = ( w1947 & w8660 ) | ( w1947 & w8662 ) | ( w8660 & w8662 ) ;
  assign w8664 = ( w1946 & ~w8661 ) | ( w1946 & w8663 ) | ( ~w8661 & w8663 ) ;
  assign w8665 = \pi029 ^ w8664 ;
  assign w8666 = ( w8277 & w8397 ) | ( w8277 & w8405 ) | ( w8397 & w8405 ) ;
  assign w8667 = w8657 ^ w8666 ;
  assign w8668 = w8665 ^ w8667 ;
  assign w8669 = ~\pi103 & w1629 ;
  assign w8670 = \pi102 & w1722 ;
  assign w8671 = ( w1629 & ~w8669 ) | ( w1629 & w8670 ) | ( ~w8669 & w8670 ) ;
  assign w8672 = ~\pi104 & w1631 ;
  assign w8673 = w3740 | w8671 ;
  assign w8674 = ( w1632 & w8671 ) | ( w1632 & w8673 ) | ( w8671 & w8673 ) ;
  assign w8675 = ( w1631 & ~w8672 ) | ( w1631 & w8674 ) | ( ~w8672 & w8674 ) ;
  assign w8676 = \pi026 ^ w8675 ;
  assign w8677 = ( w8276 & w8407 ) | ( w8276 & w8415 ) | ( w8407 & w8415 ) ;
  assign w8678 = w8668 ^ w8677 ;
  assign w8679 = w8676 ^ w8678 ;
  assign w8680 = ~\pi106 & w1313 ;
  assign w8681 = \pi105 & w1417 ;
  assign w8682 = ( w1313 & ~w8680 ) | ( w1313 & w8681 ) | ( ~w8680 & w8681 ) ;
  assign w8683 = ~\pi107 & w1315 ;
  assign w8684 = w4087 | w8682 ;
  assign w8685 = ( w1316 & w8682 ) | ( w1316 & w8684 ) | ( w8682 & w8684 ) ;
  assign w8686 = ( w1315 & ~w8683 ) | ( w1315 & w8685 ) | ( ~w8683 & w8685 ) ;
  assign w8687 = \pi023 ^ w8686 ;
  assign w8688 = w8532 ^ w8679 ;
  assign w8689 = w8687 ^ w8688 ;
  assign w8690 = w8523 ^ w8689 ;
  assign w8691 = w8531 ^ w8690 ;
  assign w8692 = w8514 ^ w8691 ;
  assign w8693 = w8522 ^ w8692 ;
  assign w8694 = w8505 ^ w8693 ;
  assign w8695 = w8513 ^ w8694 ;
  assign w8696 = w8496 ^ w8695 ;
  assign w8697 = w8504 ^ w8696 ;
  assign w8698 = ~\pi121 & w305 ;
  assign w8699 = \pi120 & w328 ;
  assign w8700 = ( w305 & ~w8698 ) | ( w305 & w8699 ) | ( ~w8698 & w8699 ) ;
  assign w8701 = ~\pi122 & w307 ;
  assign w8702 = w7069 | w8700 ;
  assign w8703 = ( w308 & w8700 ) | ( w308 & w8702 ) | ( w8700 & w8702 ) ;
  assign w8704 = ( w307 & ~w8701 ) | ( w307 & w8703 ) | ( ~w8701 & w8703 ) ;
  assign w8705 = \pi008 ^ w8704 ;
  assign w8706 = ~\pi124 & w189 ;
  assign w8707 = \pi123 & w229 ;
  assign w8708 = ( w189 & ~w8706 ) | ( w189 & w8707 ) | ( ~w8706 & w8707 ) ;
  assign w8709 = ~\pi125 & w191 ;
  assign w8710 = w7988 | w8708 ;
  assign w8711 = ( w192 & w8708 ) | ( w192 & w8710 ) | ( w8708 & w8710 ) ;
  assign w8712 = ( w191 & ~w8709 ) | ( w191 & w8711 ) | ( ~w8709 & w8711 ) ;
  assign w8713 = \pi005 ^ w8712 ;
  assign w8714 = w8697 ^ w8713 ;
  assign w8715 = w8705 ^ w8714 ;
  assign w8716 = w8495 ^ w8715 ;
  assign w8717 = w8494 ^ w8716 ;
  assign w8718 = w8478 ^ w8717 ;
  assign w8719 = w8479 ^ w8718 ;
  assign w8720 = ~\pi116 & w601 ;
  assign w8721 = \pi115 & w683 ;
  assign w8722 = ( w601 & ~w8720 ) | ( w601 & w8721 ) | ( ~w8720 & w8721 ) ;
  assign w8723 = ~\pi117 & w603 ;
  assign w8724 = w6185 | w8722 ;
  assign w8725 = ( w604 & w8722 ) | ( w604 & w8724 ) | ( w8722 & w8724 ) ;
  assign w8726 = ( w603 & ~w8723 ) | ( w603 & w8725 ) | ( ~w8723 & w8725 ) ;
  assign w8727 = \pi014 ^ w8726 ;
  assign w8728 = ( w8514 & w8522 ) | ( w8514 & w8691 ) | ( w8522 & w8691 ) ;
  assign w8729 = ( w8523 & w8531 ) | ( w8523 & w8689 ) | ( w8531 & w8689 ) ;
  assign w8730 = ~\pi110 & w1044 ;
  assign w8731 = \pi109 & w1138 ;
  assign w8732 = ( w1044 & ~w8730 ) | ( w1044 & w8731 ) | ( ~w8730 & w8731 ) ;
  assign w8733 = ~\pi111 & w1046 ;
  assign w8734 = w4811 | w8732 ;
  assign w8735 = ( w1047 & w8732 ) | ( w1047 & w8734 ) | ( w8732 & w8734 ) ;
  assign w8736 = ( w1046 & ~w8733 ) | ( w1046 & w8735 ) | ( ~w8733 & w8735 ) ;
  assign w8737 = \pi020 ^ w8736 ;
  assign w8738 = ( w8668 & w8676 ) | ( w8668 & w8677 ) | ( w8676 & w8677 ) ;
  assign w8739 = ( w8643 & w8651 ) | ( w8643 & w8652 ) | ( w8651 & w8652 ) ;
  assign w8740 = ( w8548 & w8618 ) | ( w8548 & w8619 ) | ( w8618 & w8619 ) ;
  assign w8741 = ( w8607 & w8615 ) | ( w8607 & w8616 ) | ( w8615 & w8616 ) ;
  assign w8742 = ( w8556 & w8604 ) | ( w8556 & w8605 ) | ( w8604 & w8605 ) ;
  assign w8743 = ( w8593 & w8601 ) | ( w8593 & w8602 ) | ( w8601 & w8602 ) ;
  assign w8744 = ~\pi077 & w5802 ;
  assign w8745 = \pi076 & w6052 ;
  assign w8746 = ( w5802 & ~w8744 ) | ( w5802 & w8745 ) | ( ~w8744 & w8745 ) ;
  assign w8747 = ~\pi078 & w5804 ;
  assign w8748 = w665 | w8746 ;
  assign w8749 = ( w5805 & w8746 ) | ( w5805 & w8748 ) | ( w8746 & w8748 ) ;
  assign w8750 = ( w5804 & ~w8747 ) | ( w5804 & w8749 ) | ( ~w8747 & w8749 ) ;
  assign w8751 = \pi053 ^ w8750 ;
  assign w8752 = ( w8564 & w8590 ) | ( w8564 & w8591 ) | ( w8590 & w8591 ) ;
  assign w8753 = ( w8565 & w8580 ) | ( w8565 & w8588 ) | ( w8580 & w8588 ) ;
  assign w8754 = ~\pi068 & w7811 ;
  assign w8755 = \pi067 & w8046 ;
  assign w8756 = ( w7811 & ~w8754 ) | ( w7811 & w8755 ) | ( ~w8754 & w8755 ) ;
  assign w8757 = ~\pi069 & w7813 ;
  assign w8758 = w221 | w8756 ;
  assign w8759 = ( w7814 & w8756 ) | ( w7814 & w8758 ) | ( w8756 & w8758 ) ;
  assign w8760 = ( w7813 & ~w8757 ) | ( w7813 & w8759 ) | ( ~w8757 & w8759 ) ;
  assign w8761 = \pi062 ^ w8760 ;
  assign w8762 = \pi063 & \pi064 ;
  assign w8763 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w8762 ) | ( \pi063 & w8762 ) ;
  assign w8764 = ( \pi062 & ~\pi063 ) | ( \pi062 & w8762 ) | ( ~\pi063 & w8762 ) ;
  assign w8765 = ( \pi065 & w8763 ) | ( \pi065 & w8764 ) | ( w8763 & w8764 ) ;
  assign w8766 = ( w8573 & w8574 ) | ( w8573 & w8765 ) | ( w8574 & w8765 ) ;
  assign w8767 = w8761 ^ w8766 ;
  assign w8768 = ( \pi062 & \pi063 ) | ( \pi062 & \pi066 ) | ( \pi063 & \pi066 ) ;
  assign w8769 = \pi063 & ~\pi065 ;
  assign w8770 = \pi062 & w8769 ;
  assign w8771 = w8768 ^ w8770 ;
  assign w8772 = w8767 ^ w8771 ;
  assign w8773 = ~\pi071 & w7135 ;
  assign w8774 = \pi070 & w7359 ;
  assign w8775 = ( w7135 & ~w8773 ) | ( w7135 & w8774 ) | ( ~w8773 & w8774 ) ;
  assign w8776 = ~\pi072 & w7137 ;
  assign w8777 = w361 | w8775 ;
  assign w8778 = ( w7138 & w8775 ) | ( w7138 & w8777 ) | ( w8775 & w8777 ) ;
  assign w8779 = ( w7137 & ~w8776 ) | ( w7137 & w8778 ) | ( ~w8776 & w8778 ) ;
  assign w8780 = \pi059 ^ w8779 ;
  assign w8781 = ( w8753 & w8772 ) | ( w8753 & w8780 ) | ( w8772 & w8780 ) ;
  assign w8782 = w8753 ^ w8772 ;
  assign w8783 = w8780 ^ w8782 ;
  assign w8784 = ~\pi074 & w6466 ;
  assign w8785 = \pi073 & w6702 ;
  assign w8786 = ( w6466 & ~w8784 ) | ( w6466 & w8785 ) | ( ~w8784 & w8785 ) ;
  assign w8787 = ~\pi075 & w6468 ;
  assign w8788 = w519 | w8786 ;
  assign w8789 = ( w6469 & w8786 ) | ( w6469 & w8788 ) | ( w8786 & w8788 ) ;
  assign w8790 = ( w6468 & ~w8787 ) | ( w6468 & w8789 ) | ( ~w8787 & w8789 ) ;
  assign w8791 = \pi056 ^ w8790 ;
  assign w8792 = w8752 ^ w8783 ;
  assign w8793 = w8791 ^ w8792 ;
  assign w8794 = w8743 ^ w8793 ;
  assign w8795 = w8751 ^ w8794 ;
  assign w8796 = ~\pi080 & w5209 ;
  assign w8797 = \pi079 & w5433 ;
  assign w8798 = ( w5209 & ~w8796 ) | ( w5209 & w8797 ) | ( ~w8796 & w8797 ) ;
  assign w8799 = ~\pi081 & w5211 ;
  assign w8800 = w874 | w8798 ;
  assign w8801 = ( w5212 & w8798 ) | ( w5212 & w8800 ) | ( w8798 & w8800 ) ;
  assign w8802 = ( w5211 & ~w8799 ) | ( w5211 & w8801 ) | ( ~w8799 & w8801 ) ;
  assign w8803 = \pi050 ^ w8802 ;
  assign w8804 = w8742 ^ w8795 ;
  assign w8805 = w8803 ^ w8804 ;
  assign w8806 = ~\pi083 & w4654 ;
  assign w8807 = \pi082 & w4876 ;
  assign w8808 = ( w4654 & ~w8806 ) | ( w4654 & w8807 ) | ( ~w8806 & w8807 ) ;
  assign w8809 = ~\pi084 & w4656 ;
  assign w8810 = w1188 | w8808 ;
  assign w8811 = ( w4657 & w8808 ) | ( w4657 & w8810 ) | ( w8808 & w8810 ) ;
  assign w8812 = ( w4656 & ~w8809 ) | ( w4656 & w8811 ) | ( ~w8809 & w8811 ) ;
  assign w8813 = \pi047 ^ w8812 ;
  assign w8814 = w8741 ^ w8805 ;
  assign w8815 = w8813 ^ w8814 ;
  assign w8816 = ~\pi086 & w4141 ;
  assign w8817 = \pi085 & w4334 ;
  assign w8818 = ( w4141 & ~w8816 ) | ( w4141 & w8817 ) | ( ~w8816 & w8817 ) ;
  assign w8819 = ~\pi087 & w4143 ;
  assign w8820 = w1477 | w8818 ;
  assign w8821 = ( w4144 & w8818 ) | ( w4144 & w8820 ) | ( w8818 & w8820 ) ;
  assign w8822 = ( w4143 & ~w8819 ) | ( w4143 & w8821 ) | ( ~w8819 & w8821 ) ;
  assign w8823 = \pi044 ^ w8822 ;
  assign w8824 = w8740 ^ w8815 ;
  assign w8825 = w8823 ^ w8824 ;
  assign w8826 = ~\pi089 & w3635 ;
  assign w8827 = \pi088 & w3817 ;
  assign w8828 = ( w3635 & ~w8826 ) | ( w3635 & w8827 ) | ( ~w8826 & w8827 ) ;
  assign w8829 = ~\pi090 & w3637 ;
  assign w8830 = w1801 | w8828 ;
  assign w8831 = ( w3638 & w8828 ) | ( w3638 & w8830 ) | ( w8828 & w8830 ) ;
  assign w8832 = ( w3637 & ~w8829 ) | ( w3637 & w8831 ) | ( ~w8829 & w8831 ) ;
  assign w8833 = \pi041 ^ w8832 ;
  assign w8834 = ( w8621 & w8629 ) | ( w8621 & w8630 ) | ( w8629 & w8630 ) ;
  assign w8835 = w8825 ^ w8834 ;
  assign w8836 = w8833 ^ w8835 ;
  assign w8837 = ~\pi092 & w3178 ;
  assign w8838 = \pi091 & w3340 ;
  assign w8839 = ( w3178 & ~w8837 ) | ( w3178 & w8838 ) | ( ~w8837 & w8838 ) ;
  assign w8840 = ~\pi093 & w3180 ;
  assign w8841 = w2155 | w8839 ;
  assign w8842 = ( w3181 & w8839 ) | ( w3181 & w8841 ) | ( w8839 & w8841 ) ;
  assign w8843 = ( w3180 & ~w8840 ) | ( w3180 & w8842 ) | ( ~w8840 & w8842 ) ;
  assign w8844 = \pi038 ^ w8843 ;
  assign w8845 = ( w8632 & w8640 ) | ( w8632 & w8641 ) | ( w8640 & w8641 ) ;
  assign w8846 = w8836 ^ w8845 ;
  assign w8847 = w8844 ^ w8846 ;
  assign w8848 = ~\pi095 & w2712 ;
  assign w8849 = \pi094 & w2872 ;
  assign w8850 = ( w2712 & ~w8848 ) | ( w2712 & w8849 ) | ( ~w8848 & w8849 ) ;
  assign w8851 = ~\pi096 & w2714 ;
  assign w8852 = w2546 | w8850 ;
  assign w8853 = ( w2715 & w8850 ) | ( w2715 & w8852 ) | ( w8850 & w8852 ) ;
  assign w8854 = ( w2714 & ~w8851 ) | ( w2714 & w8853 ) | ( ~w8851 & w8853 ) ;
  assign w8855 = \pi035 ^ w8854 ;
  assign w8856 = ( w8739 & w8847 ) | ( w8739 & w8855 ) | ( w8847 & w8855 ) ;
  assign w8857 = w8739 ^ w8847 ;
  assign w8858 = w8855 ^ w8857 ;
  assign w8859 = ~\pi098 & w2310 ;
  assign w8860 = \pi097 & w2443 ;
  assign w8861 = ( w2310 & ~w8859 ) | ( w2310 & w8860 ) | ( ~w8859 & w8860 ) ;
  assign w8862 = ~\pi099 & w2312 ;
  assign w8863 = w2966 | w8861 ;
  assign w8864 = ( w2313 & w8861 ) | ( w2313 & w8863 ) | ( w8861 & w8863 ) ;
  assign w8865 = ( w2312 & ~w8862 ) | ( w2312 & w8864 ) | ( ~w8862 & w8864 ) ;
  assign w8866 = \pi032 ^ w8865 ;
  assign w8867 = ( w8540 & w8654 ) | ( w8540 & w8655 ) | ( w8654 & w8655 ) ;
  assign w8868 = w8858 ^ w8867 ;
  assign w8869 = w8866 ^ w8868 ;
  assign w8870 = ~\pi101 & w1944 ;
  assign w8871 = \pi100 & w2072 ;
  assign w8872 = ( w1944 & ~w8870 ) | ( w1944 & w8871 ) | ( ~w8870 & w8871 ) ;
  assign w8873 = ~\pi102 & w1946 ;
  assign w8874 = w3284 | w8872 ;
  assign w8875 = ( w1947 & w8872 ) | ( w1947 & w8874 ) | ( w8872 & w8874 ) ;
  assign w8876 = ( w1946 & ~w8873 ) | ( w1946 & w8875 ) | ( ~w8873 & w8875 ) ;
  assign w8877 = \pi029 ^ w8876 ;
  assign w8878 = ( w8657 & w8665 ) | ( w8657 & w8666 ) | ( w8665 & w8666 ) ;
  assign w8879 = w8869 ^ w8878 ;
  assign w8880 = w8877 ^ w8879 ;
  assign w8881 = ~\pi104 & w1629 ;
  assign w8882 = \pi103 & w1722 ;
  assign w8883 = ( w1629 & ~w8881 ) | ( w1629 & w8882 ) | ( ~w8881 & w8882 ) ;
  assign w8884 = ~\pi105 & w1631 ;
  assign w8885 = w3905 | w8883 ;
  assign w8886 = ( w1632 & w8883 ) | ( w1632 & w8885 ) | ( w8883 & w8885 ) ;
  assign w8887 = ( w1631 & ~w8884 ) | ( w1631 & w8886 ) | ( ~w8884 & w8886 ) ;
  assign w8888 = \pi026 ^ w8887 ;
  assign w8889 = ( w8738 & w8880 ) | ( w8738 & w8888 ) | ( w8880 & w8888 ) ;
  assign w8890 = w8738 ^ w8880 ;
  assign w8891 = w8888 ^ w8890 ;
  assign w8892 = ~\pi107 & w1313 ;
  assign w8893 = \pi106 & w1417 ;
  assign w8894 = ( w1313 & ~w8892 ) | ( w1313 & w8893 ) | ( ~w8892 & w8893 ) ;
  assign w8895 = ~\pi108 & w1315 ;
  assign w8896 = w4425 | w8894 ;
  assign w8897 = ( w1316 & w8894 ) | ( w1316 & w8896 ) | ( w8894 & w8896 ) ;
  assign w8898 = ( w1315 & ~w8895 ) | ( w1315 & w8897 ) | ( ~w8895 & w8897 ) ;
  assign w8899 = \pi023 ^ w8898 ;
  assign w8900 = ( w8532 & w8679 ) | ( w8532 & w8687 ) | ( w8679 & w8687 ) ;
  assign w8901 = w8891 ^ w8900 ;
  assign w8902 = w8899 ^ w8901 ;
  assign w8903 = w8729 ^ w8902 ;
  assign w8904 = w8737 ^ w8903 ;
  assign w8905 = ~\pi113 & w837 ;
  assign w8906 = \pi112 & w902 ;
  assign w8907 = ( w837 & ~w8905 ) | ( w837 & w8906 ) | ( ~w8905 & w8906 ) ;
  assign w8908 = ~\pi114 & w839 ;
  assign w8909 = w5565 | w8907 ;
  assign w8910 = ( w840 & w8907 ) | ( w840 & w8909 ) | ( w8907 & w8909 ) ;
  assign w8911 = ( w839 & ~w8908 ) | ( w839 & w8910 ) | ( ~w8908 & w8910 ) ;
  assign w8912 = \pi017 ^ w8911 ;
  assign w8913 = w8728 ^ w8904 ;
  assign w8914 = w8912 ^ w8913 ;
  assign w8915 = ( w8505 & w8513 ) | ( w8505 & w8693 ) | ( w8513 & w8693 ) ;
  assign w8916 = w8914 ^ w8915 ;
  assign w8917 = w8727 ^ w8916 ;
  assign w8918 = ~\pi119 & w432 ;
  assign w8919 = \pi118 & w486 ;
  assign w8920 = ( w432 & ~w8918 ) | ( w432 & w8919 ) | ( ~w8918 & w8919 ) ;
  assign w8921 = ~\pi120 & w434 ;
  assign w8922 = w6634 | w8920 ;
  assign w8923 = ( w435 & w8920 ) | ( w435 & w8922 ) | ( w8920 & w8922 ) ;
  assign w8924 = ( w434 & ~w8921 ) | ( w434 & w8923 ) | ( ~w8921 & w8923 ) ;
  assign w8925 = \pi011 ^ w8924 ;
  assign w8926 = ~\pi122 & w305 ;
  assign w8927 = \pi121 & w328 ;
  assign w8928 = ( w305 & ~w8926 ) | ( w305 & w8927 ) | ( ~w8926 & w8927 ) ;
  assign w8929 = ~\pi123 & w307 ;
  assign w8930 = w7516 | w8928 ;
  assign w8931 = ( w308 & w8928 ) | ( w308 & w8930 ) | ( w8928 & w8930 ) ;
  assign w8932 = ( w307 & ~w8929 ) | ( w307 & w8931 ) | ( ~w8929 & w8931 ) ;
  assign w8933 = \pi008 ^ w8932 ;
  assign w8934 = w8917 ^ w8933 ;
  assign w8935 = w8925 ^ w8934 ;
  assign w8936 = ( w8496 & w8504 ) | ( w8496 & w8695 ) | ( w8504 & w8695 ) ;
  assign w8937 = ~\pi125 & w189 ;
  assign w8938 = \pi124 & w229 ;
  assign w8939 = ( w189 & ~w8937 ) | ( w189 & w8938 ) | ( ~w8937 & w8938 ) ;
  assign w8940 = ~\pi126 & w191 ;
  assign w8941 = w8231 | w8939 ;
  assign w8942 = ( w192 & w8939 ) | ( w192 & w8941 ) | ( w8939 & w8941 ) ;
  assign w8943 = ( w191 & ~w8940 ) | ( w191 & w8942 ) | ( ~w8940 & w8942 ) ;
  assign w8944 = \pi005 ^ w8943 ;
  assign w8945 = w8935 ^ w8936 ;
  assign w8946 = w8944 ^ w8945 ;
  assign w8947 = ( w8697 & w8705 ) | ( w8697 & w8713 ) | ( w8705 & w8713 ) ;
  assign w8948 = \pi002 & ~w8481 ;
  assign w8949 = ( \pi000 & \pi002 ) | ( \pi000 & w8481 ) | ( \pi002 & w8481 ) ;
  assign w8950 = ~\pi000 & \pi127 ;
  assign w8951 = ( \pi000 & ~\pi001 ) | ( \pi000 & w8950 ) | ( ~\pi001 & w8950 ) ;
  assign w8952 = ( w8948 & w8949 ) | ( w8948 & ~w8951 ) | ( w8949 & ~w8951 ) ;
  assign w8953 = w8946 ^ w8947 ;
  assign w8954 = w8952 ^ w8953 ;
  assign w8955 = ( w8494 & w8495 ) | ( w8494 & w8715 ) | ( w8495 & w8715 ) ;
  assign w8956 = ( w8478 & w8479 ) | ( w8478 & w8717 ) | ( w8479 & w8717 ) ;
  assign w8957 = w8954 ^ w8956 ;
  assign w8958 = w8955 ^ w8957 ;
  assign w8959 = ( w8935 & w8936 ) | ( w8935 & w8944 ) | ( w8936 & w8944 ) ;
  assign w8960 = ~\pi126 & w189 ;
  assign w8961 = \pi125 & w229 ;
  assign w8962 = ( w189 & ~w8960 ) | ( w189 & w8961 ) | ( ~w8960 & w8961 ) ;
  assign w8963 = ~\pi127 & w191 ;
  assign w8964 = w8466 | w8962 ;
  assign w8965 = ( w192 & w8962 ) | ( w192 & w8964 ) | ( w8962 & w8964 ) ;
  assign w8966 = ( w191 & ~w8963 ) | ( w191 & w8965 ) | ( ~w8963 & w8965 ) ;
  assign w8967 = \pi005 ^ w8966 ;
  assign w8968 = ~\pi120 & w432 ;
  assign w8969 = \pi119 & w486 ;
  assign w8970 = ( w432 & ~w8968 ) | ( w432 & w8969 ) | ( ~w8968 & w8969 ) ;
  assign w8971 = ~\pi121 & w434 ;
  assign w8972 = w7050 | w8970 ;
  assign w8973 = ( w435 & w8970 ) | ( w435 & w8972 ) | ( w8970 & w8972 ) ;
  assign w8974 = ( w434 & ~w8971 ) | ( w434 & w8973 ) | ( ~w8971 & w8973 ) ;
  assign w8975 = \pi011 ^ w8974 ;
  assign w8976 = ( w8727 & w8914 ) | ( w8727 & w8915 ) | ( w8914 & w8915 ) ;
  assign w8977 = ~\pi114 & w837 ;
  assign w8978 = \pi113 & w902 ;
  assign w8979 = ( w837 & ~w8977 ) | ( w837 & w8978 ) | ( ~w8977 & w8978 ) ;
  assign w8980 = ~\pi115 & w839 ;
  assign w8981 = w5585 | w8979 ;
  assign w8982 = ( w840 & w8979 ) | ( w840 & w8981 ) | ( w8979 & w8981 ) ;
  assign w8983 = ( w839 & ~w8980 ) | ( w839 & w8982 ) | ( ~w8980 & w8982 ) ;
  assign w8984 = \pi017 ^ w8983 ;
  assign w8985 = ( w8729 & w8737 ) | ( w8729 & w8902 ) | ( w8737 & w8902 ) ;
  assign w8986 = ~\pi111 & w1044 ;
  assign w8987 = \pi110 & w1138 ;
  assign w8988 = ( w1044 & ~w8986 ) | ( w1044 & w8987 ) | ( ~w8986 & w8987 ) ;
  assign w8989 = ~\pi112 & w1046 ;
  assign w8990 = w4999 | w8988 ;
  assign w8991 = ( w1047 & w8988 ) | ( w1047 & w8990 ) | ( w8988 & w8990 ) ;
  assign w8992 = ( w1046 & ~w8989 ) | ( w1046 & w8991 ) | ( ~w8989 & w8991 ) ;
  assign w8993 = \pi020 ^ w8992 ;
  assign w8994 = ( w8891 & w8899 ) | ( w8891 & w8900 ) | ( w8899 & w8900 ) ;
  assign w8995 = w8993 ^ w8994 ;
  assign w8996 = ~\pi108 & w1313 ;
  assign w8997 = \pi107 & w1417 ;
  assign w8998 = ( w1313 & ~w8996 ) | ( w1313 & w8997 ) | ( ~w8996 & w8997 ) ;
  assign w8999 = ~\pi109 & w1315 ;
  assign w9000 = w4599 | w8998 ;
  assign w9001 = ( w1316 & w8998 ) | ( w1316 & w9000 ) | ( w8998 & w9000 ) ;
  assign w9002 = ( w1315 & ~w8999 ) | ( w1315 & w9001 ) | ( ~w8999 & w9001 ) ;
  assign w9003 = \pi023 ^ w9002 ;
  assign w9004 = ~\pi105 & w1629 ;
  assign w9005 = \pi104 & w1722 ;
  assign w9006 = ( w1629 & ~w9004 ) | ( w1629 & w9005 ) | ( ~w9004 & w9005 ) ;
  assign w9007 = ~\pi106 & w1631 ;
  assign w9008 = w4068 | w9006 ;
  assign w9009 = ( w1632 & w9006 ) | ( w1632 & w9008 ) | ( w9006 & w9008 ) ;
  assign w9010 = ( w1631 & ~w9007 ) | ( w1631 & w9009 ) | ( ~w9007 & w9009 ) ;
  assign w9011 = \pi026 ^ w9010 ;
  assign w9012 = ( w8869 & w8877 ) | ( w8869 & w8878 ) | ( w8877 & w8878 ) ;
  assign w9013 = w9011 ^ w9012 ;
  assign w9014 = ( w8858 & w8866 ) | ( w8858 & w8867 ) | ( w8866 & w8867 ) ;
  assign w9015 = \pi101 & w2072 ;
  assign w9016 = ( \pi103 & w1946 ) | ( \pi103 & w9015 ) | ( w1946 & w9015 ) ;
  assign w9017 = \pi102 | w9016 ;
  assign w9018 = ( w1944 & w9016 ) | ( w1944 & w9017 ) | ( w9016 & w9017 ) ;
  assign w9019 = w9015 | w9018 ;
  assign w9020 = ~\pi096 & w2712 ;
  assign w9021 = \pi095 & w2872 ;
  assign w9022 = ( w2712 & ~w9020 ) | ( w2712 & w9021 ) | ( ~w9020 & w9021 ) ;
  assign w9023 = ~\pi097 & w2714 ;
  assign w9024 = w2673 | w9022 ;
  assign w9025 = ( w2715 & w9022 ) | ( w2715 & w9024 ) | ( w9022 & w9024 ) ;
  assign w9026 = ( w2714 & ~w9023 ) | ( w2714 & w9025 ) | ( ~w9023 & w9025 ) ;
  assign w9027 = \pi035 ^ w9026 ;
  assign w9028 = ~\pi087 & w4141 ;
  assign w9029 = \pi086 & w4334 ;
  assign w9030 = ( w4141 & ~w9028 ) | ( w4141 & w9029 ) | ( ~w9028 & w9029 ) ;
  assign w9031 = ~\pi088 & w4143 ;
  assign w9032 = w1574 | w9030 ;
  assign w9033 = ( w4144 & w9030 ) | ( w4144 & w9032 ) | ( w9030 & w9032 ) ;
  assign w9034 = ( w4143 & ~w9031 ) | ( w4143 & w9033 ) | ( ~w9031 & w9033 ) ;
  assign w9035 = \pi044 ^ w9034 ;
  assign w9036 = ~\pi078 & w5802 ;
  assign w9037 = \pi077 & w6052 ;
  assign w9038 = ( w5802 & ~w9036 ) | ( w5802 & w9037 ) | ( ~w9036 & w9037 ) ;
  assign w9039 = ~\pi079 & w5804 ;
  assign w9040 = w730 | w9038 ;
  assign w9041 = ( w5805 & w9038 ) | ( w5805 & w9040 ) | ( w9038 & w9040 ) ;
  assign w9042 = ( w5804 & ~w9039 ) | ( w5804 & w9041 ) | ( ~w9039 & w9041 ) ;
  assign w9043 = \pi053 ^ w9042 ;
  assign w9044 = ( w8752 & w8783 ) | ( w8752 & w8791 ) | ( w8783 & w8791 ) ;
  assign w9045 = \pi063 & \pi065 ;
  assign w9046 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w9045 ) | ( \pi063 & w9045 ) ;
  assign w9047 = ( \pi062 & ~\pi063 ) | ( \pi062 & w9045 ) | ( ~\pi063 & w9045 ) ;
  assign w9048 = ( \pi066 & w9046 ) | ( \pi066 & w9047 ) | ( w9046 & w9047 ) ;
  assign w9049 = ( w8761 & w8766 ) | ( w8761 & w9048 ) | ( w8766 & w9048 ) ;
  assign w9050 = ~\pi069 & w7811 ;
  assign w9051 = \pi068 & w8046 ;
  assign w9052 = ( w7811 & ~w9050 ) | ( w7811 & w9051 ) | ( ~w9050 & w9051 ) ;
  assign w9053 = ~\pi070 & w7813 ;
  assign w9054 = ~w271 & w7814 ;
  assign w9055 = ( w7814 & w9052 ) | ( w7814 & ~w9054 ) | ( w9052 & ~w9054 ) ;
  assign w9056 = ( w7813 & ~w9053 ) | ( w7813 & w9055 ) | ( ~w9053 & w9055 ) ;
  assign w9057 = \pi002 ^ w9056 ;
  assign w9058 = \pi062 ^ \pi067 ;
  assign w9059 = \pi063 ^ \pi067 ;
  assign w9060 = \pi062 & ~\pi066 ;
  assign w9061 = ( w9058 & ~w9059 ) | ( w9058 & w9060 ) | ( ~w9059 & w9060 ) ;
  assign w9062 = w9057 ^ w9061 ;
  assign w9063 = ~\pi072 & w7135 ;
  assign w9064 = \pi071 & w7359 ;
  assign w9065 = ( w7135 & ~w9063 ) | ( w7135 & w9064 ) | ( ~w9063 & w9064 ) ;
  assign w9066 = ~\pi073 & w7137 ;
  assign w9067 = w404 | w9065 ;
  assign w9068 = ( w7138 & w9065 ) | ( w7138 & w9067 ) | ( w9065 & w9067 ) ;
  assign w9069 = ( w7137 & ~w9066 ) | ( w7137 & w9068 ) | ( ~w9066 & w9068 ) ;
  assign w9070 = \pi059 ^ w9069 ;
  assign w9071 = w9049 ^ w9062 ;
  assign w9072 = w9070 ^ w9071 ;
  assign w9073 = ~\pi075 & w6466 ;
  assign w9074 = \pi074 & w6702 ;
  assign w9075 = ( w6466 & ~w9073 ) | ( w6466 & w9074 ) | ( ~w9073 & w9074 ) ;
  assign w9076 = ~\pi076 & w6468 ;
  assign w9077 = w538 | w9075 ;
  assign w9078 = ( w6469 & w9075 ) | ( w6469 & w9077 ) | ( w9075 & w9077 ) ;
  assign w9079 = ( w6468 & ~w9076 ) | ( w6468 & w9078 ) | ( ~w9076 & w9078 ) ;
  assign w9080 = \pi056 ^ w9079 ;
  assign w9081 = w8781 ^ w9072 ;
  assign w9082 = w9080 ^ w9081 ;
  assign w9083 = w9044 ^ w9082 ;
  assign w9084 = w9043 ^ w9083 ;
  assign w9085 = ( w8743 & w8751 ) | ( w8743 & w8793 ) | ( w8751 & w8793 ) ;
  assign w9086 = ~\pi081 & w5209 ;
  assign w9087 = \pi080 & w5433 ;
  assign w9088 = ( w5209 & ~w9086 ) | ( w5209 & w9087 ) | ( ~w9086 & w9087 ) ;
  assign w9089 = ~\pi082 & w5211 ;
  assign w9090 = w1008 | w9088 ;
  assign w9091 = ( w5212 & w9088 ) | ( w5212 & w9090 ) | ( w9088 & w9090 ) ;
  assign w9092 = ( w5211 & ~w9089 ) | ( w5211 & w9091 ) | ( ~w9089 & w9091 ) ;
  assign w9093 = \pi050 ^ w9092 ;
  assign w9094 = w9084 ^ w9085 ;
  assign w9095 = w9093 ^ w9094 ;
  assign w9096 = ( w8742 & w8795 ) | ( w8742 & w8803 ) | ( w8795 & w8803 ) ;
  assign w9097 = ~\pi084 & w4654 ;
  assign w9098 = \pi083 & w4876 ;
  assign w9099 = ( w4654 & ~w9097 ) | ( w4654 & w9098 ) | ( ~w9097 & w9098 ) ;
  assign w9100 = ~\pi085 & w4656 ;
  assign w9101 = w1274 | w9099 ;
  assign w9102 = ( w4657 & w9099 ) | ( w4657 & w9101 ) | ( w9099 & w9101 ) ;
  assign w9103 = ( w4656 & ~w9100 ) | ( w4656 & w9102 ) | ( ~w9100 & w9102 ) ;
  assign w9104 = \pi047 ^ w9103 ;
  assign w9105 = w9095 ^ w9096 ;
  assign w9106 = w9104 ^ w9105 ;
  assign w9107 = ( w8741 & w8805 ) | ( w8741 & w8813 ) | ( w8805 & w8813 ) ;
  assign w9108 = w9106 ^ w9107 ;
  assign w9109 = w9035 ^ w9108 ;
  assign w9110 = ( w8740 & w8815 ) | ( w8740 & w8823 ) | ( w8815 & w8823 ) ;
  assign w9111 = ~\pi090 & w3635 ;
  assign w9112 = \pi089 & w3817 ;
  assign w9113 = ( w3635 & ~w9111 ) | ( w3635 & w9112 ) | ( ~w9111 & w9112 ) ;
  assign w9114 = ~\pi091 & w3637 ;
  assign w9115 = w1908 | w9113 ;
  assign w9116 = ( w3638 & w9113 ) | ( w3638 & w9115 ) | ( w9113 & w9115 ) ;
  assign w9117 = ( w3637 & ~w9114 ) | ( w3637 & w9116 ) | ( ~w9114 & w9116 ) ;
  assign w9118 = \pi041 ^ w9117 ;
  assign w9119 = w9109 ^ w9110 ;
  assign w9120 = w9118 ^ w9119 ;
  assign w9121 = ( w8825 & w8833 ) | ( w8825 & w8834 ) | ( w8833 & w8834 ) ;
  assign w9122 = ~\pi093 & w3178 ;
  assign w9123 = \pi092 & w3340 ;
  assign w9124 = ( w3178 & ~w9122 ) | ( w3178 & w9123 ) | ( ~w9122 & w9123 ) ;
  assign w9125 = ~\pi094 & w3180 ;
  assign w9126 = w2274 | w9124 ;
  assign w9127 = ( w3181 & w9124 ) | ( w3181 & w9126 ) | ( w9124 & w9126 ) ;
  assign w9128 = ( w3180 & ~w9125 ) | ( w3180 & w9127 ) | ( ~w9125 & w9127 ) ;
  assign w9129 = \pi038 ^ w9128 ;
  assign w9130 = w9120 ^ w9121 ;
  assign w9131 = w9129 ^ w9130 ;
  assign w9132 = ( w8836 & w8844 ) | ( w8836 & w8845 ) | ( w8844 & w8845 ) ;
  assign w9133 = w9131 ^ w9132 ;
  assign w9134 = w9027 ^ w9133 ;
  assign w9135 = \pi098 & w2443 ;
  assign w9136 = ( \pi100 & w2312 ) | ( \pi100 & w9135 ) | ( w2312 & w9135 ) ;
  assign w9137 = \pi099 | w9136 ;
  assign w9138 = ( w2310 & w9136 ) | ( w2310 & w9137 ) | ( w9136 & w9137 ) ;
  assign w9139 = w9135 | w9138 ;
  assign w9140 = w2313 & ~w3104 ;
  assign w9141 = ( w2313 & w9139 ) | ( w2313 & ~w9140 ) | ( w9139 & ~w9140 ) ;
  assign w9142 = w8856 ^ w9141 ;
  assign w9143 = \pi032 ^ w9134 ;
  assign w9144 = w9142 ^ w9143 ;
  assign w9145 = w1947 & ~w3437 ;
  assign w9146 = ( w1947 & w9019 ) | ( w1947 & ~w9145 ) | ( w9019 & ~w9145 ) ;
  assign w9147 = w9014 ^ w9146 ;
  assign w9148 = \pi029 ^ w9144 ;
  assign w9149 = w9147 ^ w9148 ;
  assign w9150 = w9003 ^ w9149 ;
  assign w9151 = w8889 ^ w9150 ;
  assign w9152 = w9013 ^ w9151 ;
  assign w9153 = w8984 ^ w9152 ;
  assign w9154 = w8985 ^ w9153 ;
  assign w9155 = w8995 ^ w9154 ;
  assign w9156 = ( w8728 & w8904 ) | ( w8728 & w8912 ) | ( w8904 & w8912 ) ;
  assign w9157 = \pi116 & w683 ;
  assign w9158 = ( \pi118 & w603 ) | ( \pi118 & w9157 ) | ( w603 & w9157 ) ;
  assign w9159 = \pi117 | w9158 ;
  assign w9160 = ( w601 & w9158 ) | ( w601 & w9159 ) | ( w9158 & w9159 ) ;
  assign w9161 = w9157 | w9160 ;
  assign w9162 = w604 & ~w6206 ;
  assign w9163 = ( w604 & w9161 ) | ( w604 & ~w9162 ) | ( w9161 & ~w9162 ) ;
  assign w9164 = w9156 ^ w9163 ;
  assign w9165 = \pi014 ^ w9155 ;
  assign w9166 = w9164 ^ w9165 ;
  assign w9167 = w8976 ^ w9166 ;
  assign w9168 = w8975 ^ w9167 ;
  assign w9169 = ~\pi123 & w305 ;
  assign w9170 = \pi122 & w328 ;
  assign w9171 = ( w305 & ~w9169 ) | ( w305 & w9170 ) | ( ~w9169 & w9170 ) ;
  assign w9172 = ~\pi124 & w307 ;
  assign w9173 = w7538 | w9171 ;
  assign w9174 = ( w308 & w9171 ) | ( w308 & w9173 ) | ( w9171 & w9173 ) ;
  assign w9175 = ( w307 & ~w9172 ) | ( w307 & w9174 ) | ( ~w9172 & w9174 ) ;
  assign w9176 = \pi008 ^ w9175 ;
  assign w9177 = ( w8917 & w8925 ) | ( w8917 & w8933 ) | ( w8925 & w8933 ) ;
  assign w9178 = w9168 ^ w9177 ;
  assign w9179 = w9176 ^ w9178 ;
  assign w9180 = w8959 ^ w9179 ;
  assign w9181 = w8967 ^ w9180 ;
  assign w9182 = ( w8946 & w8947 ) | ( w8946 & w8952 ) | ( w8947 & w8952 ) ;
  assign w9183 = ( w8954 & w8955 ) | ( w8954 & w8956 ) | ( w8955 & w8956 ) ;
  assign w9184 = w9181 ^ w9183 ;
  assign w9185 = w9182 ^ w9184 ;
  assign w9186 = ( w9181 & w9182 ) | ( w9181 & w9183 ) | ( w9182 & w9183 ) ;
  assign w9187 = ( w8959 & w8967 ) | ( w8959 & w9179 ) | ( w8967 & w9179 ) ;
  assign w9188 = ~\pi118 & w601 ;
  assign w9189 = \pi117 & w683 ;
  assign w9190 = ( w601 & ~w9188 ) | ( w601 & w9189 ) | ( ~w9188 & w9189 ) ;
  assign w9191 = ~\pi119 & w603 ;
  assign w9192 = w6616 | w9190 ;
  assign w9193 = ( w604 & w9190 ) | ( w604 & w9192 ) | ( w9190 & w9192 ) ;
  assign w9194 = ( w603 & ~w9191 ) | ( w603 & w9193 ) | ( ~w9191 & w9193 ) ;
  assign w9195 = \pi014 ^ w9194 ;
  assign w9196 = w8995 ^ w9152 ;
  assign w9197 = ( w8984 & w8985 ) | ( w8984 & w9196 ) | ( w8985 & w9196 ) ;
  assign w9198 = ~\pi112 & w1044 ;
  assign w9199 = \pi111 & w1138 ;
  assign w9200 = ( w1044 & ~w9198 ) | ( w1044 & w9199 ) | ( ~w9198 & w9199 ) ;
  assign w9201 = ~\pi113 & w1046 ;
  assign w9202 = w5366 | w9200 ;
  assign w9203 = ( w1047 & w9200 ) | ( w1047 & w9202 ) | ( w9200 & w9202 ) ;
  assign w9204 = ( w1046 & ~w9201 ) | ( w1046 & w9203 ) | ( ~w9201 & w9203 ) ;
  assign w9205 = \pi020 ^ w9204 ;
  assign w9206 = w9013 ^ w9149 ;
  assign w9207 = ( w8889 & w9003 ) | ( w8889 & w9206 ) | ( w9003 & w9206 ) ;
  assign w9208 = ~\pi106 & w1629 ;
  assign w9209 = \pi105 & w1722 ;
  assign w9210 = ( w1629 & ~w9208 ) | ( w1629 & w9209 ) | ( ~w9208 & w9209 ) ;
  assign w9211 = ~\pi107 & w1631 ;
  assign w9212 = w4087 | w9210 ;
  assign w9213 = ( w1632 & w9210 ) | ( w1632 & w9212 ) | ( w9210 & w9212 ) ;
  assign w9214 = ( w1631 & ~w9211 ) | ( w1631 & w9213 ) | ( ~w9211 & w9213 ) ;
  assign w9215 = \pi026 ^ w9214 ;
  assign w9216 = w3437 | w9019 ;
  assign w9217 = ( w1947 & w9019 ) | ( w1947 & w9216 ) | ( w9019 & w9216 ) ;
  assign w9218 = \pi029 ^ w9217 ;
  assign w9219 = ( w9014 & w9144 ) | ( w9014 & w9218 ) | ( w9144 & w9218 ) ;
  assign w9220 = ( w9027 & w9131 ) | ( w9027 & w9132 ) | ( w9131 & w9132 ) ;
  assign w9221 = \pi099 & w2443 ;
  assign w9222 = ( \pi101 & w2312 ) | ( \pi101 & w9221 ) | ( w2312 & w9221 ) ;
  assign w9223 = \pi100 | w9222 ;
  assign w9224 = ( w2310 & w9222 ) | ( w2310 & w9223 ) | ( w9222 & w9223 ) ;
  assign w9225 = w9221 | w9224 ;
  assign w9226 = ~\pi097 & w2712 ;
  assign w9227 = \pi096 & w2872 ;
  assign w9228 = ( w2712 & ~w9226 ) | ( w2712 & w9227 ) | ( ~w9226 & w9227 ) ;
  assign w9229 = ~\pi098 & w2714 ;
  assign w9230 = w2824 | w9228 ;
  assign w9231 = ( w2715 & w9228 ) | ( w2715 & w9230 ) | ( w9228 & w9230 ) ;
  assign w9232 = ( w2714 & ~w9229 ) | ( w2714 & w9231 ) | ( ~w9229 & w9231 ) ;
  assign w9233 = \pi035 ^ w9232 ;
  assign w9234 = ( w9120 & w9121 ) | ( w9120 & w9129 ) | ( w9121 & w9129 ) ;
  assign w9235 = ~\pi079 & w5802 ;
  assign w9236 = \pi078 & w6052 ;
  assign w9237 = ( w5802 & ~w9235 ) | ( w5802 & w9236 ) | ( ~w9235 & w9236 ) ;
  assign w9238 = ~\pi080 & w5804 ;
  assign w9239 = w794 | w9237 ;
  assign w9240 = ( w5805 & w9237 ) | ( w5805 & w9239 ) | ( w9237 & w9239 ) ;
  assign w9241 = ( w5804 & ~w9238 ) | ( w5804 & w9240 ) | ( ~w9238 & w9240 ) ;
  assign w9242 = \pi053 ^ w9241 ;
  assign w9243 = ~\pi070 & w7811 ;
  assign w9244 = \pi069 & w8046 ;
  assign w9245 = ( w7811 & ~w9243 ) | ( w7811 & w9244 ) | ( ~w9243 & w9244 ) ;
  assign w9246 = ~\pi071 & w7813 ;
  assign w9247 = w290 | w9245 ;
  assign w9248 = ( w7814 & w9245 ) | ( w7814 & w9247 ) | ( w9245 & w9247 ) ;
  assign w9249 = ( w7813 & ~w9246 ) | ( w7813 & w9248 ) | ( ~w9246 & w9248 ) ;
  assign w9250 = \pi062 ^ w9249 ;
  assign w9251 = \pi002 ^ w9250 ;
  assign w9252 = ( \pi062 & \pi063 ) | ( \pi062 & \pi068 ) | ( \pi063 & \pi068 ) ;
  assign w9253 = \pi063 & ~\pi067 ;
  assign w9254 = \pi062 & w9253 ;
  assign w9255 = w9252 ^ w9254 ;
  assign w9256 = w9251 ^ w9255 ;
  assign w9257 = \pi062 ^ w9056 ;
  assign w9258 = ~\pi066 & w8768 ;
  assign w9259 = ( \pi062 & \pi063 ) | ( \pi062 & \pi067 ) | ( \pi063 & \pi067 ) ;
  assign w9260 = w9258 ^ w9259 ;
  assign w9261 = ( \pi002 & w9257 ) | ( \pi002 & w9260 ) | ( w9257 & w9260 ) ;
  assign w9262 = ~\pi073 & w7135 ;
  assign w9263 = \pi072 & w7359 ;
  assign w9264 = ( w7135 & ~w9262 ) | ( w7135 & w9263 ) | ( ~w9262 & w9263 ) ;
  assign w9265 = ~\pi074 & w7137 ;
  assign w9266 = w465 | w9264 ;
  assign w9267 = ( w7138 & w9264 ) | ( w7138 & w9266 ) | ( w9264 & w9266 ) ;
  assign w9268 = ( w7137 & ~w9265 ) | ( w7137 & w9267 ) | ( ~w9265 & w9267 ) ;
  assign w9269 = \pi059 ^ w9268 ;
  assign w9270 = w9256 ^ w9261 ;
  assign w9271 = w9269 ^ w9270 ;
  assign w9272 = ( w9049 & w9062 ) | ( w9049 & w9070 ) | ( w9062 & w9070 ) ;
  assign w9273 = ~\pi076 & w6466 ;
  assign w9274 = \pi075 & w6702 ;
  assign w9275 = ( w6466 & ~w9273 ) | ( w6466 & w9274 ) | ( ~w9273 & w9274 ) ;
  assign w9276 = ~\pi077 & w6468 ;
  assign w9277 = w644 | w9275 ;
  assign w9278 = ( w6469 & w9275 ) | ( w6469 & w9277 ) | ( w9275 & w9277 ) ;
  assign w9279 = ( w6468 & ~w9276 ) | ( w6468 & w9278 ) | ( ~w9276 & w9278 ) ;
  assign w9280 = \pi056 ^ w9279 ;
  assign w9281 = w9271 ^ w9272 ;
  assign w9282 = w9280 ^ w9281 ;
  assign w9283 = ( w8781 & w9072 ) | ( w8781 & w9080 ) | ( w9072 & w9080 ) ;
  assign w9284 = w9282 ^ w9283 ;
  assign w9285 = w9242 ^ w9284 ;
  assign w9286 = ( w9043 & w9044 ) | ( w9043 & w9082 ) | ( w9044 & w9082 ) ;
  assign w9287 = ~\pi082 & w5209 ;
  assign w9288 = \pi081 & w5433 ;
  assign w9289 = ( w5209 & ~w9287 ) | ( w5209 & w9288 ) | ( ~w9287 & w9288 ) ;
  assign w9290 = ~\pi083 & w5211 ;
  assign w9291 = w1099 | w9289 ;
  assign w9292 = ( w5212 & w9289 ) | ( w5212 & w9291 ) | ( w9289 & w9291 ) ;
  assign w9293 = ( w5211 & ~w9290 ) | ( w5211 & w9292 ) | ( ~w9290 & w9292 ) ;
  assign w9294 = \pi050 ^ w9293 ;
  assign w9295 = w9285 ^ w9286 ;
  assign w9296 = w9294 ^ w9295 ;
  assign w9297 = ( w9084 & w9085 ) | ( w9084 & w9093 ) | ( w9085 & w9093 ) ;
  assign w9298 = ~\pi085 & w4654 ;
  assign w9299 = \pi084 & w4876 ;
  assign w9300 = ( w4654 & ~w9298 ) | ( w4654 & w9299 ) | ( ~w9298 & w9299 ) ;
  assign w9301 = ~\pi086 & w4656 ;
  assign w9302 = w1379 | w9300 ;
  assign w9303 = ( w4657 & w9300 ) | ( w4657 & w9302 ) | ( w9300 & w9302 ) ;
  assign w9304 = ( w4656 & ~w9301 ) | ( w4656 & w9303 ) | ( ~w9301 & w9303 ) ;
  assign w9305 = \pi047 ^ w9304 ;
  assign w9306 = w9296 ^ w9297 ;
  assign w9307 = w9305 ^ w9306 ;
  assign w9308 = ( w9095 & w9096 ) | ( w9095 & w9104 ) | ( w9096 & w9104 ) ;
  assign w9309 = ~\pi088 & w4141 ;
  assign w9310 = \pi087 & w4334 ;
  assign w9311 = ( w4141 & ~w9309 ) | ( w4141 & w9310 ) | ( ~w9309 & w9310 ) ;
  assign w9312 = ~\pi089 & w4143 ;
  assign w9313 = w1595 | w9311 ;
  assign w9314 = ( w4144 & w9311 ) | ( w4144 & w9313 ) | ( w9311 & w9313 ) ;
  assign w9315 = ( w4143 & ~w9312 ) | ( w4143 & w9314 ) | ( ~w9312 & w9314 ) ;
  assign w9316 = \pi044 ^ w9315 ;
  assign w9317 = w9307 ^ w9308 ;
  assign w9318 = w9316 ^ w9317 ;
  assign w9319 = ( w9035 & w9106 ) | ( w9035 & w9107 ) | ( w9106 & w9107 ) ;
  assign w9320 = ~\pi091 & w3635 ;
  assign w9321 = \pi090 & w3817 ;
  assign w9322 = ( w3635 & ~w9320 ) | ( w3635 & w9321 ) | ( ~w9320 & w9321 ) ;
  assign w9323 = ~\pi092 & w3637 ;
  assign w9324 = w2033 | w9322 ;
  assign w9325 = ( w3638 & w9322 ) | ( w3638 & w9324 ) | ( w9322 & w9324 ) ;
  assign w9326 = ( w3637 & ~w9323 ) | ( w3637 & w9325 ) | ( ~w9323 & w9325 ) ;
  assign w9327 = \pi041 ^ w9326 ;
  assign w9328 = w9318 ^ w9319 ;
  assign w9329 = w9327 ^ w9328 ;
  assign w9330 = ( w9109 & w9110 ) | ( w9109 & w9118 ) | ( w9110 & w9118 ) ;
  assign w9331 = ~\pi094 & w3178 ;
  assign w9332 = \pi093 & w3340 ;
  assign w9333 = ( w3178 & ~w9331 ) | ( w3178 & w9332 ) | ( ~w9331 & w9332 ) ;
  assign w9334 = ~\pi095 & w3180 ;
  assign w9335 = w2409 | w9333 ;
  assign w9336 = ( w3181 & w9333 ) | ( w3181 & w9335 ) | ( w9333 & w9335 ) ;
  assign w9337 = ( w3180 & ~w9334 ) | ( w3180 & w9336 ) | ( ~w9334 & w9336 ) ;
  assign w9338 = \pi038 ^ w9337 ;
  assign w9339 = w9329 ^ w9330 ;
  assign w9340 = w9338 ^ w9339 ;
  assign w9341 = w9234 ^ w9340 ;
  assign w9342 = w9233 ^ w9341 ;
  assign w9343 = w2313 & ~w3264 ;
  assign w9344 = ( w2313 & w9225 ) | ( w2313 & ~w9343 ) | ( w9225 & ~w9343 ) ;
  assign w9345 = w9220 ^ w9344 ;
  assign w9346 = \pi032 ^ w9342 ;
  assign w9347 = w9345 ^ w9346 ;
  assign w9348 = w3104 | w9139 ;
  assign w9349 = ( w2313 & w9139 ) | ( w2313 & w9348 ) | ( w9139 & w9348 ) ;
  assign w9350 = \pi032 ^ w9349 ;
  assign w9351 = ( w8856 & w9134 ) | ( w8856 & w9350 ) | ( w9134 & w9350 ) ;
  assign w9352 = \pi102 & w2072 ;
  assign w9353 = ( \pi104 & w1946 ) | ( \pi104 & w9352 ) | ( w1946 & w9352 ) ;
  assign w9354 = \pi103 | w9353 ;
  assign w9355 = ( w1944 & w9353 ) | ( w1944 & w9354 ) | ( w9353 & w9354 ) ;
  assign w9356 = w9352 | w9355 ;
  assign w9357 = w1947 & ~w3740 ;
  assign w9358 = ( w1947 & w9356 ) | ( w1947 & ~w9357 ) | ( w9356 & ~w9357 ) ;
  assign w9359 = w9351 ^ w9358 ;
  assign w9360 = \pi029 ^ w9347 ;
  assign w9361 = w9359 ^ w9360 ;
  assign w9362 = w9219 ^ w9361 ;
  assign w9363 = w9215 ^ w9362 ;
  assign w9364 = ~\pi109 & w1313 ;
  assign w9365 = \pi108 & w1417 ;
  assign w9366 = ( w1313 & ~w9364 ) | ( w1313 & w9365 ) | ( ~w9364 & w9365 ) ;
  assign w9367 = ~\pi110 & w1315 ;
  assign w9368 = w4792 | w9366 ;
  assign w9369 = ( w1316 & w9366 ) | ( w1316 & w9368 ) | ( w9366 & w9368 ) ;
  assign w9370 = ( w1315 & ~w9367 ) | ( w1315 & w9369 ) | ( ~w9367 & w9369 ) ;
  assign w9371 = \pi023 ^ w9370 ;
  assign w9372 = ( w9011 & w9012 ) | ( w9011 & w9149 ) | ( w9012 & w9149 ) ;
  assign w9373 = w9363 ^ w9372 ;
  assign w9374 = w9371 ^ w9373 ;
  assign w9375 = w9207 ^ w9374 ;
  assign w9376 = w9205 ^ w9375 ;
  assign w9377 = ~\pi115 & w837 ;
  assign w9378 = \pi114 & w902 ;
  assign w9379 = ( w837 & ~w9377 ) | ( w837 & w9378 ) | ( ~w9377 & w9378 ) ;
  assign w9380 = ~\pi116 & w839 ;
  assign w9381 = w5976 | w9379 ;
  assign w9382 = ( w840 & w9379 ) | ( w840 & w9381 ) | ( w9379 & w9381 ) ;
  assign w9383 = ( w839 & ~w9380 ) | ( w839 & w9382 ) | ( ~w9380 & w9382 ) ;
  assign w9384 = \pi017 ^ w9383 ;
  assign w9385 = ( w8993 & w8994 ) | ( w8993 & w9152 ) | ( w8994 & w9152 ) ;
  assign w9386 = w9376 ^ w9385 ;
  assign w9387 = w9384 ^ w9386 ;
  assign w9388 = w9197 ^ w9387 ;
  assign w9389 = w9195 ^ w9388 ;
  assign w9390 = w6206 | w9161 ;
  assign w9391 = ( w604 & w9161 ) | ( w604 & w9390 ) | ( w9161 & w9390 ) ;
  assign w9392 = \pi014 ^ w9391 ;
  assign w9393 = ( w9155 & w9156 ) | ( w9155 & w9392 ) | ( w9156 & w9392 ) ;
  assign w9394 = \pi120 & w486 ;
  assign w9395 = ( \pi122 & w434 ) | ( \pi122 & w9394 ) | ( w434 & w9394 ) ;
  assign w9396 = \pi121 | w9395 ;
  assign w9397 = ( w432 & w9395 ) | ( w432 & w9396 ) | ( w9395 & w9396 ) ;
  assign w9398 = w9394 | w9397 ;
  assign w9399 = w435 & ~w7069 ;
  assign w9400 = ( w435 & w9398 ) | ( w435 & ~w9399 ) | ( w9398 & ~w9399 ) ;
  assign w9401 = w9393 ^ w9400 ;
  assign w9402 = \pi011 ^ w9389 ;
  assign w9403 = w9401 ^ w9402 ;
  assign w9404 = ( w8975 & w8976 ) | ( w8975 & w9166 ) | ( w8976 & w9166 ) ;
  assign w9405 = \pi123 & w328 ;
  assign w9406 = ( \pi125 & w307 ) | ( \pi125 & w9405 ) | ( w307 & w9405 ) ;
  assign w9407 = \pi124 | w9406 ;
  assign w9408 = ( w305 & w9406 ) | ( w305 & w9407 ) | ( w9406 & w9407 ) ;
  assign w9409 = w9405 | w9408 ;
  assign w9410 = w308 & ~w7988 ;
  assign w9411 = ( w308 & w9409 ) | ( w308 & ~w9410 ) | ( w9409 & ~w9410 ) ;
  assign w9412 = w9404 ^ w9411 ;
  assign w9413 = \pi008 ^ w9403 ;
  assign w9414 = w9412 ^ w9413 ;
  assign w9415 = ( w9168 & w9176 ) | ( w9168 & w9177 ) | ( w9176 & w9177 ) ;
  assign w9416 = \pi127 & w189 ;
  assign w9417 = ( \pi126 & ~w192 ) | ( \pi126 & w8490 ) | ( ~w192 & w8490 ) ;
  assign w9418 = \pi126 & ~w229 ;
  assign w9419 = ( ~\pi126 & w9417 ) | ( ~\pi126 & w9418 ) | ( w9417 & w9418 ) ;
  assign w9420 = \pi126 | w8490 ;
  assign w9421 = ( w9416 & ~w9419 ) | ( w9416 & w9420 ) | ( ~w9419 & w9420 ) ;
  assign w9422 = \pi005 ^ w9421 ;
  assign w9423 = w9414 ^ w9422 ;
  assign w9424 = w9415 ^ w9423 ;
  assign w9425 = w9186 ^ w9187 ;
  assign w9426 = w9424 ^ w9425 ;
  assign w9427 = ( w9186 & w9187 ) | ( w9186 & w9424 ) | ( w9187 & w9424 ) ;
  assign w9428 = ( w9414 & w9415 ) | ( w9414 & w9422 ) | ( w9415 & w9422 ) ;
  assign w9429 = w7988 | w9409 ;
  assign w9430 = ( w308 & w9409 ) | ( w308 & w9429 ) | ( w9409 & w9429 ) ;
  assign w9431 = \pi008 ^ w9430 ;
  assign w9432 = ( w9403 & w9404 ) | ( w9403 & w9431 ) | ( w9404 & w9431 ) ;
  assign w9433 = w192 & w8481 ;
  assign w9434 = w229 | w9433 ;
  assign w9435 = ( \pi127 & w9433 ) | ( \pi127 & w9434 ) | ( w9433 & w9434 ) ;
  assign w9436 = \pi005 ^ w9435 ;
  assign w9437 = ~\pi122 & w432 ;
  assign w9438 = \pi121 & w486 ;
  assign w9439 = ( w432 & ~w9437 ) | ( w432 & w9438 ) | ( ~w9437 & w9438 ) ;
  assign w9440 = ~\pi123 & w434 ;
  assign w9441 = w7516 | w9439 ;
  assign w9442 = ( w435 & w9439 ) | ( w435 & w9441 ) | ( w9439 & w9441 ) ;
  assign w9443 = ( w434 & ~w9440 ) | ( w434 & w9442 ) | ( ~w9440 & w9442 ) ;
  assign w9444 = \pi011 ^ w9443 ;
  assign w9445 = ( w9195 & w9197 ) | ( w9195 & w9387 ) | ( w9197 & w9387 ) ;
  assign w9446 = ~\pi119 & w601 ;
  assign w9447 = \pi118 & w683 ;
  assign w9448 = ( w601 & ~w9446 ) | ( w601 & w9447 ) | ( ~w9446 & w9447 ) ;
  assign w9449 = ~\pi120 & w603 ;
  assign w9450 = w6634 | w9448 ;
  assign w9451 = ( w604 & w9448 ) | ( w604 & w9450 ) | ( w9448 & w9450 ) ;
  assign w9452 = ( w603 & ~w9449 ) | ( w603 & w9451 ) | ( ~w9449 & w9451 ) ;
  assign w9453 = \pi014 ^ w9452 ;
  assign w9454 = ( w9376 & w9384 ) | ( w9376 & w9385 ) | ( w9384 & w9385 ) ;
  assign w9455 = ( w9205 & w9207 ) | ( w9205 & w9374 ) | ( w9207 & w9374 ) ;
  assign w9456 = \pi115 & w902 ;
  assign w9457 = ( \pi117 & w839 ) | ( \pi117 & w9456 ) | ( w839 & w9456 ) ;
  assign w9458 = \pi116 | w9457 ;
  assign w9459 = ( w837 & w9457 ) | ( w837 & w9458 ) | ( w9457 & w9458 ) ;
  assign w9460 = w9456 | w9459 ;
  assign w9461 = ~\pi113 & w1044 ;
  assign w9462 = \pi112 & w1138 ;
  assign w9463 = ( w1044 & ~w9461 ) | ( w1044 & w9462 ) | ( ~w9461 & w9462 ) ;
  assign w9464 = ~\pi114 & w1046 ;
  assign w9465 = w5565 | w9463 ;
  assign w9466 = ( w1047 & w9463 ) | ( w1047 & w9465 ) | ( w9463 & w9465 ) ;
  assign w9467 = ( w1046 & ~w9464 ) | ( w1046 & w9466 ) | ( ~w9464 & w9466 ) ;
  assign w9468 = \pi020 ^ w9467 ;
  assign w9469 = ( w9363 & w9371 ) | ( w9363 & w9372 ) | ( w9371 & w9372 ) ;
  assign w9470 = ~\pi110 & w1313 ;
  assign w9471 = \pi109 & w1417 ;
  assign w9472 = ( w1313 & ~w9470 ) | ( w1313 & w9471 ) | ( ~w9470 & w9471 ) ;
  assign w9473 = ~\pi111 & w1315 ;
  assign w9474 = w4811 | w9472 ;
  assign w9475 = ( w1316 & w9472 ) | ( w1316 & w9474 ) | ( w9472 & w9474 ) ;
  assign w9476 = ( w1315 & ~w9473 ) | ( w1315 & w9475 ) | ( ~w9473 & w9475 ) ;
  assign w9477 = \pi023 ^ w9476 ;
  assign w9478 = ( w9215 & w9219 ) | ( w9215 & w9361 ) | ( w9219 & w9361 ) ;
  assign w9479 = ~\pi104 & w1944 ;
  assign w9480 = \pi103 & w2072 ;
  assign w9481 = ( w1944 & ~w9479 ) | ( w1944 & w9480 ) | ( ~w9479 & w9480 ) ;
  assign w9482 = ~\pi105 & w1946 ;
  assign w9483 = w3905 | w9481 ;
  assign w9484 = ( w1947 & w9481 ) | ( w1947 & w9483 ) | ( w9481 & w9483 ) ;
  assign w9485 = ( w1946 & ~w9482 ) | ( w1946 & w9484 ) | ( ~w9482 & w9484 ) ;
  assign w9486 = \pi029 ^ w9485 ;
  assign w9487 = w3264 | w9225 ;
  assign w9488 = ( w2313 & w9225 ) | ( w2313 & w9487 ) | ( w9225 & w9487 ) ;
  assign w9489 = \pi032 ^ w9488 ;
  assign w9490 = ( w9220 & w9342 ) | ( w9220 & w9489 ) | ( w9342 & w9489 ) ;
  assign w9491 = ~\pi098 & w2712 ;
  assign w9492 = \pi097 & w2872 ;
  assign w9493 = ( w2712 & ~w9491 ) | ( w2712 & w9492 ) | ( ~w9491 & w9492 ) ;
  assign w9494 = ~\pi099 & w2714 ;
  assign w9495 = w2966 | w9493 ;
  assign w9496 = ( w2715 & w9493 ) | ( w2715 & w9495 ) | ( w9493 & w9495 ) ;
  assign w9497 = ( w2714 & ~w9494 ) | ( w2714 & w9496 ) | ( ~w9494 & w9496 ) ;
  assign w9498 = \pi035 ^ w9497 ;
  assign w9499 = ~\pi086 & w4654 ;
  assign w9500 = \pi085 & w4876 ;
  assign w9501 = ( w4654 & ~w9499 ) | ( w4654 & w9500 ) | ( ~w9499 & w9500 ) ;
  assign w9502 = ~\pi087 & w4656 ;
  assign w9503 = w1477 | w9501 ;
  assign w9504 = ( w4657 & w9501 ) | ( w4657 & w9503 ) | ( w9501 & w9503 ) ;
  assign w9505 = ( w4656 & ~w9502 ) | ( w4656 & w9504 ) | ( ~w9502 & w9504 ) ;
  assign w9506 = \pi047 ^ w9505 ;
  assign w9507 = ~\pi077 & w6466 ;
  assign w9508 = \pi076 & w6702 ;
  assign w9509 = ( w6466 & ~w9507 ) | ( w6466 & w9508 ) | ( ~w9507 & w9508 ) ;
  assign w9510 = ~\pi078 & w6468 ;
  assign w9511 = w665 | w9509 ;
  assign w9512 = ( w6469 & w9509 ) | ( w6469 & w9511 ) | ( w9509 & w9511 ) ;
  assign w9513 = ( w6468 & ~w9510 ) | ( w6468 & w9512 ) | ( ~w9510 & w9512 ) ;
  assign w9514 = \pi056 ^ w9513 ;
  assign w9515 = ~\pi071 & w7811 ;
  assign w9516 = \pi070 & w8046 ;
  assign w9517 = ( w7811 & ~w9515 ) | ( w7811 & w9516 ) | ( ~w9515 & w9516 ) ;
  assign w9518 = ~\pi072 & w7813 ;
  assign w9519 = w361 | w9517 ;
  assign w9520 = ( w7814 & w9517 ) | ( w7814 & w9519 ) | ( w9517 & w9519 ) ;
  assign w9521 = ( w7813 & ~w9518 ) | ( w7813 & w9520 ) | ( ~w9518 & w9520 ) ;
  assign w9522 = \pi062 ^ w9521 ;
  assign w9523 = \pi002 ^ w9522 ;
  assign w9524 = ( \pi062 & \pi063 ) | ( \pi062 & \pi069 ) | ( \pi063 & \pi069 ) ;
  assign w9525 = \pi063 & ~\pi068 ;
  assign w9526 = \pi062 & w9525 ;
  assign w9527 = w9524 ^ w9526 ;
  assign w9528 = w9523 ^ w9527 ;
  assign w9529 = \pi063 & \pi067 ;
  assign w9530 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w9529 ) | ( \pi063 & w9529 ) ;
  assign w9531 = ( \pi062 & ~\pi063 ) | ( \pi062 & w9529 ) | ( ~\pi063 & w9529 ) ;
  assign w9532 = ( \pi068 & w9530 ) | ( \pi068 & w9531 ) | ( w9530 & w9531 ) ;
  assign w9533 = ( \pi002 & w9250 ) | ( \pi002 & w9532 ) | ( w9250 & w9532 ) ;
  assign w9534 = ~\pi074 & w7135 ;
  assign w9535 = \pi073 & w7359 ;
  assign w9536 = ( w7135 & ~w9534 ) | ( w7135 & w9535 ) | ( ~w9534 & w9535 ) ;
  assign w9537 = ~\pi075 & w7137 ;
  assign w9538 = w519 | w9536 ;
  assign w9539 = ( w7138 & w9536 ) | ( w7138 & w9538 ) | ( w9536 & w9538 ) ;
  assign w9540 = ( w7137 & ~w9537 ) | ( w7137 & w9539 ) | ( ~w9537 & w9539 ) ;
  assign w9541 = \pi059 ^ w9540 ;
  assign w9542 = w9528 ^ w9533 ;
  assign w9543 = w9541 ^ w9542 ;
  assign w9544 = ( w9256 & w9261 ) | ( w9256 & w9269 ) | ( w9261 & w9269 ) ;
  assign w9545 = w9514 ^ w9543 ;
  assign w9546 = w9544 ^ w9545 ;
  assign w9547 = ( w9271 & w9272 ) | ( w9271 & w9280 ) | ( w9272 & w9280 ) ;
  assign w9548 = ~\pi080 & w5802 ;
  assign w9549 = \pi079 & w6052 ;
  assign w9550 = ( w5802 & ~w9548 ) | ( w5802 & w9549 ) | ( ~w9548 & w9549 ) ;
  assign w9551 = ~\pi081 & w5804 ;
  assign w9552 = w874 | w9550 ;
  assign w9553 = ( w5805 & w9550 ) | ( w5805 & w9552 ) | ( w9550 & w9552 ) ;
  assign w9554 = ( w5804 & ~w9551 ) | ( w5804 & w9553 ) | ( ~w9551 & w9553 ) ;
  assign w9555 = \pi053 ^ w9554 ;
  assign w9556 = w9546 ^ w9547 ;
  assign w9557 = w9555 ^ w9556 ;
  assign w9558 = ( w9242 & w9282 ) | ( w9242 & w9283 ) | ( w9282 & w9283 ) ;
  assign w9559 = ~\pi083 & w5209 ;
  assign w9560 = \pi082 & w5433 ;
  assign w9561 = ( w5209 & ~w9559 ) | ( w5209 & w9560 ) | ( ~w9559 & w9560 ) ;
  assign w9562 = ~\pi084 & w5211 ;
  assign w9563 = w1188 | w9561 ;
  assign w9564 = ( w5212 & w9561 ) | ( w5212 & w9563 ) | ( w9561 & w9563 ) ;
  assign w9565 = ( w5211 & ~w9562 ) | ( w5211 & w9564 ) | ( ~w9562 & w9564 ) ;
  assign w9566 = \pi050 ^ w9565 ;
  assign w9567 = w9557 ^ w9558 ;
  assign w9568 = w9566 ^ w9567 ;
  assign w9569 = ( w9285 & w9286 ) | ( w9285 & w9294 ) | ( w9286 & w9294 ) ;
  assign w9570 = w9568 ^ w9569 ;
  assign w9571 = w9506 ^ w9570 ;
  assign w9572 = ( w9296 & w9297 ) | ( w9296 & w9305 ) | ( w9297 & w9305 ) ;
  assign w9573 = ~\pi089 & w4141 ;
  assign w9574 = \pi088 & w4334 ;
  assign w9575 = ( w4141 & ~w9573 ) | ( w4141 & w9574 ) | ( ~w9573 & w9574 ) ;
  assign w9576 = ~\pi090 & w4143 ;
  assign w9577 = w1801 | w9575 ;
  assign w9578 = ( w4144 & w9575 ) | ( w4144 & w9577 ) | ( w9575 & w9577 ) ;
  assign w9579 = ( w4143 & ~w9576 ) | ( w4143 & w9578 ) | ( ~w9576 & w9578 ) ;
  assign w9580 = \pi044 ^ w9579 ;
  assign w9581 = w9571 ^ w9572 ;
  assign w9582 = w9580 ^ w9581 ;
  assign w9583 = ( w9307 & w9308 ) | ( w9307 & w9316 ) | ( w9308 & w9316 ) ;
  assign w9584 = ~\pi092 & w3635 ;
  assign w9585 = \pi091 & w3817 ;
  assign w9586 = ( w3635 & ~w9584 ) | ( w3635 & w9585 ) | ( ~w9584 & w9585 ) ;
  assign w9587 = ~\pi093 & w3637 ;
  assign w9588 = w2155 | w9586 ;
  assign w9589 = ( w3638 & w9586 ) | ( w3638 & w9588 ) | ( w9586 & w9588 ) ;
  assign w9590 = ( w3637 & ~w9587 ) | ( w3637 & w9589 ) | ( ~w9587 & w9589 ) ;
  assign w9591 = \pi041 ^ w9590 ;
  assign w9592 = w9582 ^ w9583 ;
  assign w9593 = w9591 ^ w9592 ;
  assign w9594 = ( w9318 & w9319 ) | ( w9318 & w9327 ) | ( w9319 & w9327 ) ;
  assign w9595 = ~\pi095 & w3178 ;
  assign w9596 = \pi094 & w3340 ;
  assign w9597 = ( w3178 & ~w9595 ) | ( w3178 & w9596 ) | ( ~w9595 & w9596 ) ;
  assign w9598 = ~\pi096 & w3180 ;
  assign w9599 = w2546 | w9597 ;
  assign w9600 = ( w3181 & w9597 ) | ( w3181 & w9599 ) | ( w9597 & w9599 ) ;
  assign w9601 = ( w3180 & ~w9598 ) | ( w3180 & w9600 ) | ( ~w9598 & w9600 ) ;
  assign w9602 = \pi038 ^ w9601 ;
  assign w9603 = w9593 ^ w9594 ;
  assign w9604 = w9602 ^ w9603 ;
  assign w9605 = ( w9329 & w9330 ) | ( w9329 & w9338 ) | ( w9330 & w9338 ) ;
  assign w9606 = w9604 ^ w9605 ;
  assign w9607 = w9498 ^ w9606 ;
  assign w9608 = ( w9233 & w9234 ) | ( w9233 & w9340 ) | ( w9234 & w9340 ) ;
  assign w9609 = \pi100 & w2443 ;
  assign w9610 = ( \pi102 & w2312 ) | ( \pi102 & w9609 ) | ( w2312 & w9609 ) ;
  assign w9611 = \pi101 | w9610 ;
  assign w9612 = ( w2310 & w9610 ) | ( w2310 & w9611 ) | ( w9610 & w9611 ) ;
  assign w9613 = w9609 | w9612 ;
  assign w9614 = w2313 & ~w3284 ;
  assign w9615 = ( w2313 & w9613 ) | ( w2313 & ~w9614 ) | ( w9613 & ~w9614 ) ;
  assign w9616 = w9608 ^ w9615 ;
  assign w9617 = \pi032 ^ w9607 ;
  assign w9618 = w9616 ^ w9617 ;
  assign w9619 = w9490 ^ w9618 ;
  assign w9620 = w9486 ^ w9619 ;
  assign w9621 = w3740 | w9356 ;
  assign w9622 = ( w1947 & w9356 ) | ( w1947 & w9621 ) | ( w9356 & w9621 ) ;
  assign w9623 = \pi029 ^ w9622 ;
  assign w9624 = ( w9347 & w9351 ) | ( w9347 & w9623 ) | ( w9351 & w9623 ) ;
  assign w9625 = \pi106 & w1722 ;
  assign w9626 = ( \pi108 & w1631 ) | ( \pi108 & w9625 ) | ( w1631 & w9625 ) ;
  assign w9627 = \pi107 | w9626 ;
  assign w9628 = ( w1629 & w9626 ) | ( w1629 & w9627 ) | ( w9626 & w9627 ) ;
  assign w9629 = w9625 | w9628 ;
  assign w9630 = w1632 & ~w4425 ;
  assign w9631 = ( w1632 & w9629 ) | ( w1632 & ~w9630 ) | ( w9629 & ~w9630 ) ;
  assign w9632 = w9624 ^ w9631 ;
  assign w9633 = \pi026 ^ w9620 ;
  assign w9634 = w9632 ^ w9633 ;
  assign w9635 = w9478 ^ w9634 ;
  assign w9636 = w9477 ^ w9635 ;
  assign w9637 = w9469 ^ w9636 ;
  assign w9638 = w9468 ^ w9637 ;
  assign w9639 = w840 & ~w6185 ;
  assign w9640 = ( w840 & w9460 ) | ( w840 & ~w9639 ) | ( w9460 & ~w9639 ) ;
  assign w9641 = w9455 ^ w9640 ;
  assign w9642 = \pi017 ^ w9638 ;
  assign w9643 = w9641 ^ w9642 ;
  assign w9644 = w9454 ^ w9643 ;
  assign w9645 = w9453 ^ w9644 ;
  assign w9646 = w9445 ^ w9645 ;
  assign w9647 = w9444 ^ w9646 ;
  assign w9648 = w7069 | w9398 ;
  assign w9649 = ( w435 & w9398 ) | ( w435 & w9648 ) | ( w9398 & w9648 ) ;
  assign w9650 = \pi011 ^ w9649 ;
  assign w9651 = ( w9389 & w9393 ) | ( w9389 & w9650 ) | ( w9393 & w9650 ) ;
  assign w9652 = \pi124 & w328 ;
  assign w9653 = ( \pi126 & w307 ) | ( \pi126 & w9652 ) | ( w307 & w9652 ) ;
  assign w9654 = \pi125 | w9653 ;
  assign w9655 = ( w305 & w9653 ) | ( w305 & w9654 ) | ( w9653 & w9654 ) ;
  assign w9656 = w9652 | w9655 ;
  assign w9657 = w308 & ~w8231 ;
  assign w9658 = ( w308 & w9656 ) | ( w308 & ~w9657 ) | ( w9656 & ~w9657 ) ;
  assign w9659 = w9651 ^ w9658 ;
  assign w9660 = \pi008 ^ w9647 ;
  assign w9661 = w9659 ^ w9660 ;
  assign w9662 = w9432 ^ w9661 ;
  assign w9663 = w9436 ^ w9662 ;
  assign w9664 = w9427 ^ w9428 ;
  assign w9665 = w9663 ^ w9664 ;
  assign w9666 = ( w9427 & w9428 ) | ( w9427 & w9663 ) | ( w9428 & w9663 ) ;
  assign w9667 = ( w9432 & w9436 ) | ( w9432 & w9661 ) | ( w9436 & w9661 ) ;
  assign w9668 = w8231 | w9656 ;
  assign w9669 = ( w308 & w9656 ) | ( w308 & w9668 ) | ( w9656 & w9668 ) ;
  assign w9670 = \pi008 ^ w9669 ;
  assign w9671 = ( w9647 & w9651 ) | ( w9647 & w9670 ) | ( w9651 & w9670 ) ;
  assign w9672 = ~\pi126 & w305 ;
  assign w9673 = \pi125 & w328 ;
  assign w9674 = ( w305 & ~w9672 ) | ( w305 & w9673 ) | ( ~w9672 & w9673 ) ;
  assign w9675 = ~\pi127 & w307 ;
  assign w9676 = w8466 | w9674 ;
  assign w9677 = ( w308 & w9674 ) | ( w308 & w9676 ) | ( w9674 & w9676 ) ;
  assign w9678 = ( w307 & ~w9675 ) | ( w307 & w9677 ) | ( ~w9675 & w9677 ) ;
  assign w9679 = \pi008 ^ w9678 ;
  assign w9680 = ~\pi123 & w432 ;
  assign w9681 = \pi122 & w486 ;
  assign w9682 = ( w432 & ~w9680 ) | ( w432 & w9681 ) | ( ~w9680 & w9681 ) ;
  assign w9683 = ~\pi124 & w434 ;
  assign w9684 = w7538 | w9682 ;
  assign w9685 = ( w435 & w9682 ) | ( w435 & w9684 ) | ( w9682 & w9684 ) ;
  assign w9686 = ( w434 & ~w9683 ) | ( w434 & w9685 ) | ( ~w9683 & w9685 ) ;
  assign w9687 = \pi011 ^ w9686 ;
  assign w9688 = ( w9444 & w9445 ) | ( w9444 & w9645 ) | ( w9445 & w9645 ) ;
  assign w9689 = w6185 | w9460 ;
  assign w9690 = ( w840 & w9460 ) | ( w840 & w9689 ) | ( w9460 & w9689 ) ;
  assign w9691 = \pi017 ^ w9690 ;
  assign w9692 = ( w9455 & w9638 ) | ( w9455 & w9691 ) | ( w9638 & w9691 ) ;
  assign w9693 = ~\pi117 & w837 ;
  assign w9694 = \pi116 & w902 ;
  assign w9695 = ( w837 & ~w9693 ) | ( w837 & w9694 ) | ( ~w9693 & w9694 ) ;
  assign w9696 = ~\pi118 & w839 ;
  assign w9697 = w6206 | w9695 ;
  assign w9698 = ( w840 & w9695 ) | ( w840 & w9697 ) | ( w9695 & w9697 ) ;
  assign w9699 = ( w839 & ~w9696 ) | ( w839 & w9698 ) | ( ~w9696 & w9698 ) ;
  assign w9700 = \pi017 ^ w9699 ;
  assign w9701 = ~\pi111 & w1313 ;
  assign w9702 = \pi110 & w1417 ;
  assign w9703 = ( w1313 & ~w9701 ) | ( w1313 & w9702 ) | ( ~w9701 & w9702 ) ;
  assign w9704 = ~\pi112 & w1315 ;
  assign w9705 = w4999 | w9703 ;
  assign w9706 = ( w1316 & w9703 ) | ( w1316 & w9705 ) | ( w9703 & w9705 ) ;
  assign w9707 = ( w1315 & ~w9704 ) | ( w1315 & w9706 ) | ( ~w9704 & w9706 ) ;
  assign w9708 = \pi023 ^ w9707 ;
  assign w9709 = ( w9477 & w9478 ) | ( w9477 & w9634 ) | ( w9478 & w9634 ) ;
  assign w9710 = w4425 | w9629 ;
  assign w9711 = ( w1632 & w9629 ) | ( w1632 & w9710 ) | ( w9629 & w9710 ) ;
  assign w9712 = \pi026 ^ w9711 ;
  assign w9713 = ( w9620 & w9624 ) | ( w9620 & w9712 ) | ( w9624 & w9712 ) ;
  assign w9714 = ~\pi108 & w1629 ;
  assign w9715 = \pi107 & w1722 ;
  assign w9716 = ( w1629 & ~w9714 ) | ( w1629 & w9715 ) | ( ~w9714 & w9715 ) ;
  assign w9717 = ~\pi109 & w1631 ;
  assign w9718 = w4599 | w9716 ;
  assign w9719 = ( w1632 & w9716 ) | ( w1632 & w9718 ) | ( w9716 & w9718 ) ;
  assign w9720 = ( w1631 & ~w9717 ) | ( w1631 & w9719 ) | ( ~w9717 & w9719 ) ;
  assign w9721 = \pi026 ^ w9720 ;
  assign w9722 = ~\pi105 & w1944 ;
  assign w9723 = \pi104 & w2072 ;
  assign w9724 = ( w1944 & ~w9722 ) | ( w1944 & w9723 ) | ( ~w9722 & w9723 ) ;
  assign w9725 = ~\pi106 & w1946 ;
  assign w9726 = w4068 | w9724 ;
  assign w9727 = ( w1947 & w9724 ) | ( w1947 & w9726 ) | ( w9724 & w9726 ) ;
  assign w9728 = ( w1946 & ~w9725 ) | ( w1946 & w9727 ) | ( ~w9725 & w9727 ) ;
  assign w9729 = \pi029 ^ w9728 ;
  assign w9730 = ( w9486 & w9490 ) | ( w9486 & w9618 ) | ( w9490 & w9618 ) ;
  assign w9731 = ( w9498 & w9604 ) | ( w9498 & w9605 ) | ( w9604 & w9605 ) ;
  assign w9732 = ( w9593 & w9594 ) | ( w9593 & w9602 ) | ( w9594 & w9602 ) ;
  assign w9733 = ( w9582 & w9583 ) | ( w9582 & w9591 ) | ( w9583 & w9591 ) ;
  assign w9734 = ( w9506 & w9568 ) | ( w9506 & w9569 ) | ( w9568 & w9569 ) ;
  assign w9735 = ( w9557 & w9558 ) | ( w9557 & w9566 ) | ( w9558 & w9566 ) ;
  assign w9736 = ( w9528 & w9533 ) | ( w9528 & w9541 ) | ( w9533 & w9541 ) ;
  assign w9737 = ~\pi075 & w7135 ;
  assign w9738 = \pi074 & w7359 ;
  assign w9739 = ( w7135 & ~w9737 ) | ( w7135 & w9738 ) | ( ~w9737 & w9738 ) ;
  assign w9740 = ~\pi076 & w7137 ;
  assign w9741 = w538 | w9739 ;
  assign w9742 = ( w7138 & w9739 ) | ( w7138 & w9741 ) | ( w9739 & w9741 ) ;
  assign w9743 = ( w7137 & ~w9740 ) | ( w7137 & w9742 ) | ( ~w9740 & w9742 ) ;
  assign w9744 = \pi059 ^ w9743 ;
  assign w9745 = \pi063 & \pi068 ;
  assign w9746 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w9745 ) | ( \pi063 & w9745 ) ;
  assign w9747 = ( \pi062 & ~\pi063 ) | ( \pi062 & w9745 ) | ( ~\pi063 & w9745 ) ;
  assign w9748 = ( \pi069 & w9746 ) | ( \pi069 & w9747 ) | ( w9746 & w9747 ) ;
  assign w9749 = ( \pi002 & w9522 ) | ( \pi002 & w9748 ) | ( w9522 & w9748 ) ;
  assign w9750 = \pi002 ^ \pi005 ;
  assign w9751 = ( \pi062 & \pi063 ) | ( \pi062 & \pi070 ) | ( \pi063 & \pi070 ) ;
  assign w9752 = \pi063 & ~\pi069 ;
  assign w9753 = \pi062 & w9752 ;
  assign w9754 = w9751 ^ w9753 ;
  assign w9755 = w9750 ^ w9754 ;
  assign w9756 = ~\pi072 & w7811 ;
  assign w9757 = \pi071 & w8046 ;
  assign w9758 = ( w7811 & ~w9756 ) | ( w7811 & w9757 ) | ( ~w9756 & w9757 ) ;
  assign w9759 = ~\pi073 & w7813 ;
  assign w9760 = w404 | w9758 ;
  assign w9761 = ( w7814 & w9758 ) | ( w7814 & w9760 ) | ( w9758 & w9760 ) ;
  assign w9762 = ( w7813 & ~w9759 ) | ( w7813 & w9761 ) | ( ~w9759 & w9761 ) ;
  assign w9763 = \pi062 ^ w9762 ;
  assign w9764 = w9749 ^ w9763 ;
  assign w9765 = w9755 ^ w9764 ;
  assign w9766 = w9736 ^ w9765 ;
  assign w9767 = w9744 ^ w9766 ;
  assign w9768 = ~\pi078 & w6466 ;
  assign w9769 = \pi077 & w6702 ;
  assign w9770 = ( w6466 & ~w9768 ) | ( w6466 & w9769 ) | ( ~w9768 & w9769 ) ;
  assign w9771 = ~\pi079 & w6468 ;
  assign w9772 = w730 | w9770 ;
  assign w9773 = ( w6469 & w9770 ) | ( w6469 & w9772 ) | ( w9770 & w9772 ) ;
  assign w9774 = ( w6468 & ~w9771 ) | ( w6468 & w9773 ) | ( ~w9771 & w9773 ) ;
  assign w9775 = \pi056 ^ w9774 ;
  assign w9776 = ( w9514 & w9543 ) | ( w9514 & w9544 ) | ( w9543 & w9544 ) ;
  assign w9777 = w9767 ^ w9776 ;
  assign w9778 = w9775 ^ w9777 ;
  assign w9779 = ~\pi081 & w5802 ;
  assign w9780 = \pi080 & w6052 ;
  assign w9781 = ( w5802 & ~w9779 ) | ( w5802 & w9780 ) | ( ~w9779 & w9780 ) ;
  assign w9782 = ~\pi082 & w5804 ;
  assign w9783 = w1008 | w9781 ;
  assign w9784 = ( w5805 & w9781 ) | ( w5805 & w9783 ) | ( w9781 & w9783 ) ;
  assign w9785 = ( w5804 & ~w9782 ) | ( w5804 & w9784 ) | ( ~w9782 & w9784 ) ;
  assign w9786 = \pi053 ^ w9785 ;
  assign w9787 = ( w9546 & w9547 ) | ( w9546 & w9555 ) | ( w9547 & w9555 ) ;
  assign w9788 = w9778 ^ w9787 ;
  assign w9789 = w9786 ^ w9788 ;
  assign w9790 = ~\pi084 & w5209 ;
  assign w9791 = \pi083 & w5433 ;
  assign w9792 = ( w5209 & ~w9790 ) | ( w5209 & w9791 ) | ( ~w9790 & w9791 ) ;
  assign w9793 = ~\pi085 & w5211 ;
  assign w9794 = w1274 | w9792 ;
  assign w9795 = ( w5212 & w9792 ) | ( w5212 & w9794 ) | ( w9792 & w9794 ) ;
  assign w9796 = ( w5211 & ~w9793 ) | ( w5211 & w9795 ) | ( ~w9793 & w9795 ) ;
  assign w9797 = \pi050 ^ w9796 ;
  assign w9798 = w9735 ^ w9789 ;
  assign w9799 = w9797 ^ w9798 ;
  assign w9800 = ~\pi087 & w4654 ;
  assign w9801 = \pi086 & w4876 ;
  assign w9802 = ( w4654 & ~w9800 ) | ( w4654 & w9801 ) | ( ~w9800 & w9801 ) ;
  assign w9803 = ~\pi088 & w4656 ;
  assign w9804 = w1574 | w9802 ;
  assign w9805 = ( w4657 & w9802 ) | ( w4657 & w9804 ) | ( w9802 & w9804 ) ;
  assign w9806 = ( w4656 & ~w9803 ) | ( w4656 & w9805 ) | ( ~w9803 & w9805 ) ;
  assign w9807 = \pi047 ^ w9806 ;
  assign w9808 = w9734 ^ w9799 ;
  assign w9809 = w9807 ^ w9808 ;
  assign w9810 = ~\pi090 & w4141 ;
  assign w9811 = \pi089 & w4334 ;
  assign w9812 = ( w4141 & ~w9810 ) | ( w4141 & w9811 ) | ( ~w9810 & w9811 ) ;
  assign w9813 = ~\pi091 & w4143 ;
  assign w9814 = w1908 | w9812 ;
  assign w9815 = ( w4144 & w9812 ) | ( w4144 & w9814 ) | ( w9812 & w9814 ) ;
  assign w9816 = ( w4143 & ~w9813 ) | ( w4143 & w9815 ) | ( ~w9813 & w9815 ) ;
  assign w9817 = \pi044 ^ w9816 ;
  assign w9818 = ( w9571 & w9572 ) | ( w9571 & w9580 ) | ( w9572 & w9580 ) ;
  assign w9819 = w9809 ^ w9818 ;
  assign w9820 = w9817 ^ w9819 ;
  assign w9821 = ~\pi093 & w3635 ;
  assign w9822 = \pi092 & w3817 ;
  assign w9823 = ( w3635 & ~w9821 ) | ( w3635 & w9822 ) | ( ~w9821 & w9822 ) ;
  assign w9824 = ~\pi094 & w3637 ;
  assign w9825 = w2274 | w9823 ;
  assign w9826 = ( w3638 & w9823 ) | ( w3638 & w9825 ) | ( w9823 & w9825 ) ;
  assign w9827 = ( w3637 & ~w9824 ) | ( w3637 & w9826 ) | ( ~w9824 & w9826 ) ;
  assign w9828 = \pi041 ^ w9827 ;
  assign w9829 = ( w9733 & w9820 ) | ( w9733 & w9828 ) | ( w9820 & w9828 ) ;
  assign w9830 = w9733 ^ w9820 ;
  assign w9831 = w9828 ^ w9830 ;
  assign w9832 = ~\pi096 & w3178 ;
  assign w9833 = \pi095 & w3340 ;
  assign w9834 = ( w3178 & ~w9832 ) | ( w3178 & w9833 ) | ( ~w9832 & w9833 ) ;
  assign w9835 = ~\pi097 & w3180 ;
  assign w9836 = w2673 | w9834 ;
  assign w9837 = ( w3181 & w9834 ) | ( w3181 & w9836 ) | ( w9834 & w9836 ) ;
  assign w9838 = ( w3180 & ~w9835 ) | ( w3180 & w9837 ) | ( ~w9835 & w9837 ) ;
  assign w9839 = \pi038 ^ w9838 ;
  assign w9840 = w9732 ^ w9831 ;
  assign w9841 = w9839 ^ w9840 ;
  assign w9842 = ~\pi099 & w2712 ;
  assign w9843 = \pi098 & w2872 ;
  assign w9844 = ( w2712 & ~w9842 ) | ( w2712 & w9843 ) | ( ~w9842 & w9843 ) ;
  assign w9845 = ~\pi100 & w2714 ;
  assign w9846 = w3104 | w9844 ;
  assign w9847 = ( w2715 & w9844 ) | ( w2715 & w9846 ) | ( w9844 & w9846 ) ;
  assign w9848 = ( w2714 & ~w9845 ) | ( w2714 & w9847 ) | ( ~w9845 & w9847 ) ;
  assign w9849 = \pi035 ^ w9848 ;
  assign w9850 = w9731 ^ w9841 ;
  assign w9851 = w9849 ^ w9850 ;
  assign w9852 = ~\pi102 & w2310 ;
  assign w9853 = \pi101 & w2443 ;
  assign w9854 = ( w2310 & ~w9852 ) | ( w2310 & w9853 ) | ( ~w9852 & w9853 ) ;
  assign w9855 = ~\pi103 & w2312 ;
  assign w9856 = w3437 | w9854 ;
  assign w9857 = ( w2313 & w9854 ) | ( w2313 & w9856 ) | ( w9854 & w9856 ) ;
  assign w9858 = ( w2312 & ~w9855 ) | ( w2312 & w9857 ) | ( ~w9855 & w9857 ) ;
  assign w9859 = \pi032 ^ w9858 ;
  assign w9860 = w3284 | w9613 ;
  assign w9861 = ( w2313 & w9613 ) | ( w2313 & w9860 ) | ( w9613 & w9860 ) ;
  assign w9862 = \pi032 ^ w9861 ;
  assign w9863 = ( w9607 & w9608 ) | ( w9607 & w9862 ) | ( w9608 & w9862 ) ;
  assign w9864 = w9851 ^ w9863 ;
  assign w9865 = w9859 ^ w9864 ;
  assign w9866 = w9730 ^ w9865 ;
  assign w9867 = w9729 ^ w9866 ;
  assign w9868 = w9713 ^ w9867 ;
  assign w9869 = w9721 ^ w9868 ;
  assign w9870 = w9709 ^ w9869 ;
  assign w9871 = w9708 ^ w9870 ;
  assign w9872 = ~\pi114 & w1044 ;
  assign w9873 = \pi113 & w1138 ;
  assign w9874 = ( w1044 & ~w9872 ) | ( w1044 & w9873 ) | ( ~w9872 & w9873 ) ;
  assign w9875 = ~\pi115 & w1046 ;
  assign w9876 = w5585 | w9874 ;
  assign w9877 = ( w1047 & w9874 ) | ( w1047 & w9876 ) | ( w9874 & w9876 ) ;
  assign w9878 = ( w1046 & ~w9875 ) | ( w1046 & w9877 ) | ( ~w9875 & w9877 ) ;
  assign w9879 = \pi020 ^ w9878 ;
  assign w9880 = ( w9468 & w9469 ) | ( w9468 & w9636 ) | ( w9469 & w9636 ) ;
  assign w9881 = w9871 ^ w9880 ;
  assign w9882 = w9879 ^ w9881 ;
  assign w9883 = w9692 ^ w9882 ;
  assign w9884 = w9700 ^ w9883 ;
  assign w9885 = ~\pi120 & w601 ;
  assign w9886 = \pi119 & w683 ;
  assign w9887 = ( w601 & ~w9885 ) | ( w601 & w9886 ) | ( ~w9885 & w9886 ) ;
  assign w9888 = ~\pi121 & w603 ;
  assign w9889 = w7050 | w9887 ;
  assign w9890 = ( w604 & w9887 ) | ( w604 & w9889 ) | ( w9887 & w9889 ) ;
  assign w9891 = ( w603 & ~w9888 ) | ( w603 & w9890 ) | ( ~w9888 & w9890 ) ;
  assign w9892 = \pi014 ^ w9891 ;
  assign w9893 = ( w9453 & w9454 ) | ( w9453 & w9643 ) | ( w9454 & w9643 ) ;
  assign w9894 = w9884 ^ w9893 ;
  assign w9895 = w9892 ^ w9894 ;
  assign w9896 = w9688 ^ w9895 ;
  assign w9897 = w9687 ^ w9896 ;
  assign w9898 = w9671 ^ w9897 ;
  assign w9899 = w9679 ^ w9898 ;
  assign w9900 = w9666 ^ w9667 ;
  assign w9901 = w9899 ^ w9900 ;
  assign w9902 = ( w9687 & w9688 ) | ( w9687 & w9895 ) | ( w9688 & w9895 ) ;
  assign w9903 = \pi127 & w305 ;
  assign w9904 = ( \pi126 & ~w308 ) | ( \pi126 & w8490 ) | ( ~w308 & w8490 ) ;
  assign w9905 = \pi126 & ~w328 ;
  assign w9906 = ( ~\pi126 & w9904 ) | ( ~\pi126 & w9905 ) | ( w9904 & w9905 ) ;
  assign w9907 = ( w9420 & w9903 ) | ( w9420 & ~w9906 ) | ( w9903 & ~w9906 ) ;
  assign w9908 = ~\pi124 & w432 ;
  assign w9909 = \pi123 & w486 ;
  assign w9910 = ( w432 & ~w9908 ) | ( w432 & w9909 ) | ( ~w9908 & w9909 ) ;
  assign w9911 = ~\pi125 & w434 ;
  assign w9912 = w7988 | w9910 ;
  assign w9913 = ( w435 & w9910 ) | ( w435 & w9912 ) | ( w9910 & w9912 ) ;
  assign w9914 = ( w434 & ~w9911 ) | ( w434 & w9913 ) | ( ~w9911 & w9913 ) ;
  assign w9915 = \pi011 ^ w9914 ;
  assign w9916 = ( w9884 & w9892 ) | ( w9884 & w9893 ) | ( w9892 & w9893 ) ;
  assign w9917 = w9915 ^ w9916 ;
  assign w9918 = ( w9692 & w9700 ) | ( w9692 & w9882 ) | ( w9700 & w9882 ) ;
  assign w9919 = \pi120 & w683 ;
  assign w9920 = ( \pi122 & w603 ) | ( \pi122 & w9919 ) | ( w603 & w9919 ) ;
  assign w9921 = \pi121 | w9920 ;
  assign w9922 = ( w601 & w9920 ) | ( w601 & w9921 ) | ( w9920 & w9921 ) ;
  assign w9923 = w9919 | w9922 ;
  assign w9924 = ~w604 & w7069 ;
  assign w9925 = ( w7069 & w9923 ) | ( w7069 & ~w9924 ) | ( w9923 & ~w9924 ) ;
  assign w9926 = \pi014 ^ w9925 ;
  assign w9927 = ~\pi118 & w837 ;
  assign w9928 = \pi117 & w902 ;
  assign w9929 = ( w837 & ~w9927 ) | ( w837 & w9928 ) | ( ~w9927 & w9928 ) ;
  assign w9930 = ~\pi119 & w839 ;
  assign w9931 = w6616 | w9929 ;
  assign w9932 = ( w840 & w9929 ) | ( w840 & w9931 ) | ( w9929 & w9931 ) ;
  assign w9933 = ( w839 & ~w9930 ) | ( w839 & w9932 ) | ( ~w9930 & w9932 ) ;
  assign w9934 = \pi017 ^ w9933 ;
  assign w9935 = ( w9871 & w9879 ) | ( w9871 & w9880 ) | ( w9879 & w9880 ) ;
  assign w9936 = w9934 ^ w9935 ;
  assign w9937 = ~\pi115 & w1044 ;
  assign w9938 = \pi114 & w1138 ;
  assign w9939 = ( w1044 & ~w9937 ) | ( w1044 & w9938 ) | ( ~w9937 & w9938 ) ;
  assign w9940 = ~\pi116 & w1046 ;
  assign w9941 = w5976 | w9939 ;
  assign w9942 = ( w1047 & w9939 ) | ( w1047 & w9941 ) | ( w9939 & w9941 ) ;
  assign w9943 = ( w1046 & ~w9940 ) | ( w1046 & w9942 ) | ( ~w9940 & w9942 ) ;
  assign w9944 = \pi020 ^ w9943 ;
  assign w9945 = ( w9708 & w9709 ) | ( w9708 & w9869 ) | ( w9709 & w9869 ) ;
  assign w9946 = ~\pi112 & w1313 ;
  assign w9947 = \pi111 & w1417 ;
  assign w9948 = ( w1313 & ~w9946 ) | ( w1313 & w9947 ) | ( ~w9946 & w9947 ) ;
  assign w9949 = ~\pi113 & w1315 ;
  assign w9950 = w5366 | w9948 ;
  assign w9951 = ( w1316 & w9948 ) | ( w1316 & w9950 ) | ( w9948 & w9950 ) ;
  assign w9952 = ( w1315 & ~w9949 ) | ( w1315 & w9951 ) | ( ~w9949 & w9951 ) ;
  assign w9953 = \pi023 ^ w9952 ;
  assign w9954 = ( w9713 & w9721 ) | ( w9713 & w9867 ) | ( w9721 & w9867 ) ;
  assign w9955 = ( w9729 & w9730 ) | ( w9729 & w9865 ) | ( w9730 & w9865 ) ;
  assign w9956 = \pi108 & w1722 ;
  assign w9957 = ( \pi110 & w1631 ) | ( \pi110 & w9956 ) | ( w1631 & w9956 ) ;
  assign w9958 = \pi109 | w9957 ;
  assign w9959 = ( w1629 & w9957 ) | ( w1629 & w9958 ) | ( w9957 & w9958 ) ;
  assign w9960 = w9956 | w9959 ;
  assign w9961 = ~\pi106 & w1944 ;
  assign w9962 = \pi105 & w2072 ;
  assign w9963 = ( w1944 & ~w9961 ) | ( w1944 & w9962 ) | ( ~w9961 & w9962 ) ;
  assign w9964 = ~\pi107 & w1946 ;
  assign w9965 = w4087 | w9963 ;
  assign w9966 = ( w1947 & w9963 ) | ( w1947 & w9965 ) | ( w9963 & w9965 ) ;
  assign w9967 = ( w1946 & ~w9964 ) | ( w1946 & w9966 ) | ( ~w9964 & w9966 ) ;
  assign w9968 = \pi029 ^ w9967 ;
  assign w9969 = ( w9851 & w9859 ) | ( w9851 & w9863 ) | ( w9859 & w9863 ) ;
  assign w9970 = ~\pi103 & w2310 ;
  assign w9971 = \pi102 & w2443 ;
  assign w9972 = ( w2310 & ~w9970 ) | ( w2310 & w9971 ) | ( ~w9970 & w9971 ) ;
  assign w9973 = ~\pi104 & w2312 ;
  assign w9974 = w3740 | w9972 ;
  assign w9975 = ( w2313 & w9972 ) | ( w2313 & w9974 ) | ( w9972 & w9974 ) ;
  assign w9976 = ( w2312 & ~w9973 ) | ( w2312 & w9975 ) | ( ~w9973 & w9975 ) ;
  assign w9977 = \pi032 ^ w9976 ;
  assign w9978 = ( w9731 & w9841 ) | ( w9731 & w9849 ) | ( w9841 & w9849 ) ;
  assign w9979 = ~\pi100 & w2712 ;
  assign w9980 = \pi099 & w2872 ;
  assign w9981 = ( w2712 & ~w9979 ) | ( w2712 & w9980 ) | ( ~w9979 & w9980 ) ;
  assign w9982 = ~\pi101 & w2714 ;
  assign w9983 = w3264 | w9981 ;
  assign w9984 = ( w2715 & w9981 ) | ( w2715 & w9983 ) | ( w9981 & w9983 ) ;
  assign w9985 = ( w2714 & ~w9982 ) | ( w2714 & w9984 ) | ( ~w9982 & w9984 ) ;
  assign w9986 = \pi035 ^ w9985 ;
  assign w9987 = ( w9732 & w9831 ) | ( w9732 & w9839 ) | ( w9831 & w9839 ) ;
  assign w9988 = ~\pi097 & w3178 ;
  assign w9989 = \pi096 & w3340 ;
  assign w9990 = ( w3178 & ~w9988 ) | ( w3178 & w9989 ) | ( ~w9988 & w9989 ) ;
  assign w9991 = ~\pi098 & w3180 ;
  assign w9992 = w2824 | w9990 ;
  assign w9993 = ( w3181 & w9990 ) | ( w3181 & w9992 ) | ( w9990 & w9992 ) ;
  assign w9994 = ( w3180 & ~w9991 ) | ( w3180 & w9993 ) | ( ~w9991 & w9993 ) ;
  assign w9995 = \pi038 ^ w9994 ;
  assign w9996 = ( w9749 & w9755 ) | ( w9749 & w9763 ) | ( w9755 & w9763 ) ;
  assign w9997 = \pi063 & \pi069 ;
  assign w9998 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w9997 ) | ( \pi063 & w9997 ) ;
  assign w9999 = ( \pi062 & ~\pi063 ) | ( \pi062 & w9997 ) | ( ~\pi063 & w9997 ) ;
  assign w10000 = ( \pi070 & w9998 ) | ( \pi070 & w9999 ) | ( w9998 & w9999 ) ;
  assign w10001 = ( \pi002 & \pi005 ) | ( \pi002 & ~w10000 ) | ( \pi005 & ~w10000 ) ;
  assign w10002 = ~\pi073 & w7811 ;
  assign w10003 = \pi072 & w8046 ;
  assign w10004 = ( w7811 & ~w10002 ) | ( w7811 & w10003 ) | ( ~w10002 & w10003 ) ;
  assign w10005 = ~\pi074 & w7813 ;
  assign w10006 = ~w465 & w7814 ;
  assign w10007 = ( w7814 & w10004 ) | ( w7814 & ~w10006 ) | ( w10004 & ~w10006 ) ;
  assign w10008 = ( w7813 & ~w10005 ) | ( w7813 & w10007 ) | ( ~w10005 & w10007 ) ;
  assign w10009 = w10001 ^ w10008 ;
  assign w10010 = \pi062 ^ \pi071 ;
  assign w10011 = \pi063 ^ \pi071 ;
  assign w10012 = \pi062 & ~\pi070 ;
  assign w10013 = ( w10010 & ~w10011 ) | ( w10010 & w10012 ) | ( ~w10011 & w10012 ) ;
  assign w10014 = w10009 ^ w10013 ;
  assign w10015 = ~\pi076 & w7135 ;
  assign w10016 = \pi075 & w7359 ;
  assign w10017 = ( w7135 & ~w10015 ) | ( w7135 & w10016 ) | ( ~w10015 & w10016 ) ;
  assign w10018 = ~\pi077 & w7137 ;
  assign w10019 = w644 | w10017 ;
  assign w10020 = ( w7138 & w10017 ) | ( w7138 & w10019 ) | ( w10017 & w10019 ) ;
  assign w10021 = ( w7137 & ~w10018 ) | ( w7137 & w10020 ) | ( ~w10018 & w10020 ) ;
  assign w10022 = \pi059 ^ w10021 ;
  assign w10023 = w9996 ^ w10014 ;
  assign w10024 = w10022 ^ w10023 ;
  assign w10025 = ( w9736 & w9744 ) | ( w9736 & w9765 ) | ( w9744 & w9765 ) ;
  assign w10026 = ~\pi079 & w6466 ;
  assign w10027 = \pi078 & w6702 ;
  assign w10028 = ( w6466 & ~w10026 ) | ( w6466 & w10027 ) | ( ~w10026 & w10027 ) ;
  assign w10029 = ~\pi080 & w6468 ;
  assign w10030 = w794 | w10028 ;
  assign w10031 = ( w6469 & w10028 ) | ( w6469 & w10030 ) | ( w10028 & w10030 ) ;
  assign w10032 = ( w6468 & ~w10029 ) | ( w6468 & w10031 ) | ( ~w10029 & w10031 ) ;
  assign w10033 = \pi056 ^ w10032 ;
  assign w10034 = w10024 ^ w10025 ;
  assign w10035 = w10033 ^ w10034 ;
  assign w10036 = ( w9767 & w9775 ) | ( w9767 & w9776 ) | ( w9775 & w9776 ) ;
  assign w10037 = ~\pi082 & w5802 ;
  assign w10038 = \pi081 & w6052 ;
  assign w10039 = ( w5802 & ~w10037 ) | ( w5802 & w10038 ) | ( ~w10037 & w10038 ) ;
  assign w10040 = ~\pi083 & w5804 ;
  assign w10041 = w1099 | w10039 ;
  assign w10042 = ( w5805 & w10039 ) | ( w5805 & w10041 ) | ( w10039 & w10041 ) ;
  assign w10043 = ( w5804 & ~w10040 ) | ( w5804 & w10042 ) | ( ~w10040 & w10042 ) ;
  assign w10044 = \pi053 ^ w10043 ;
  assign w10045 = w10035 ^ w10036 ;
  assign w10046 = w10044 ^ w10045 ;
  assign w10047 = ( w9778 & w9786 ) | ( w9778 & w9787 ) | ( w9786 & w9787 ) ;
  assign w10048 = ~\pi085 & w5209 ;
  assign w10049 = \pi084 & w5433 ;
  assign w10050 = ( w5209 & ~w10048 ) | ( w5209 & w10049 ) | ( ~w10048 & w10049 ) ;
  assign w10051 = ~\pi086 & w5211 ;
  assign w10052 = w1379 | w10050 ;
  assign w10053 = ( w5212 & w10050 ) | ( w5212 & w10052 ) | ( w10050 & w10052 ) ;
  assign w10054 = ( w5211 & ~w10051 ) | ( w5211 & w10053 ) | ( ~w10051 & w10053 ) ;
  assign w10055 = \pi050 ^ w10054 ;
  assign w10056 = w10046 ^ w10047 ;
  assign w10057 = w10055 ^ w10056 ;
  assign w10058 = ( w9735 & w9789 ) | ( w9735 & w9797 ) | ( w9789 & w9797 ) ;
  assign w10059 = ~\pi088 & w4654 ;
  assign w10060 = \pi087 & w4876 ;
  assign w10061 = ( w4654 & ~w10059 ) | ( w4654 & w10060 ) | ( ~w10059 & w10060 ) ;
  assign w10062 = ~\pi089 & w4656 ;
  assign w10063 = w1595 | w10061 ;
  assign w10064 = ( w4657 & w10061 ) | ( w4657 & w10063 ) | ( w10061 & w10063 ) ;
  assign w10065 = ( w4656 & ~w10062 ) | ( w4656 & w10064 ) | ( ~w10062 & w10064 ) ;
  assign w10066 = \pi047 ^ w10065 ;
  assign w10067 = w10057 ^ w10058 ;
  assign w10068 = w10066 ^ w10067 ;
  assign w10069 = ( w9734 & w9799 ) | ( w9734 & w9807 ) | ( w9799 & w9807 ) ;
  assign w10070 = ~\pi091 & w4141 ;
  assign w10071 = \pi090 & w4334 ;
  assign w10072 = ( w4141 & ~w10070 ) | ( w4141 & w10071 ) | ( ~w10070 & w10071 ) ;
  assign w10073 = ~\pi092 & w4143 ;
  assign w10074 = w2033 | w10072 ;
  assign w10075 = ( w4144 & w10072 ) | ( w4144 & w10074 ) | ( w10072 & w10074 ) ;
  assign w10076 = ( w4143 & ~w10073 ) | ( w4143 & w10075 ) | ( ~w10073 & w10075 ) ;
  assign w10077 = \pi044 ^ w10076 ;
  assign w10078 = w10068 ^ w10069 ;
  assign w10079 = w10077 ^ w10078 ;
  assign w10080 = ( w9809 & w9817 ) | ( w9809 & w9818 ) | ( w9817 & w9818 ) ;
  assign w10081 = ~\pi094 & w3635 ;
  assign w10082 = \pi093 & w3817 ;
  assign w10083 = ( w3635 & ~w10081 ) | ( w3635 & w10082 ) | ( ~w10081 & w10082 ) ;
  assign w10084 = ~\pi095 & w3637 ;
  assign w10085 = w2409 | w10083 ;
  assign w10086 = ( w3638 & w10083 ) | ( w3638 & w10085 ) | ( w10083 & w10085 ) ;
  assign w10087 = ( w3637 & ~w10084 ) | ( w3637 & w10086 ) | ( ~w10084 & w10086 ) ;
  assign w10088 = \pi041 ^ w10087 ;
  assign w10089 = w10079 ^ w10080 ;
  assign w10090 = w10088 ^ w10089 ;
  assign w10091 = w9829 ^ w10090 ;
  assign w10092 = w9995 ^ w10091 ;
  assign w10093 = w9987 ^ w10092 ;
  assign w10094 = w9986 ^ w10093 ;
  assign w10095 = w9978 ^ w10094 ;
  assign w10096 = w9977 ^ w10095 ;
  assign w10097 = w9969 ^ w10096 ;
  assign w10098 = w9968 ^ w10097 ;
  assign w10099 = w1632 & ~w4792 ;
  assign w10100 = ( w1632 & w9960 ) | ( w1632 & ~w10099 ) | ( w9960 & ~w10099 ) ;
  assign w10101 = w9955 ^ w10100 ;
  assign w10102 = \pi026 ^ w10098 ;
  assign w10103 = w10101 ^ w10102 ;
  assign w10104 = w9954 ^ w10103 ;
  assign w10105 = w9953 ^ w10104 ;
  assign w10106 = w9945 ^ w10105 ;
  assign w10107 = w9944 ^ w10106 ;
  assign w10108 = w9926 ^ w10107 ;
  assign w10109 = w9918 ^ w10108 ;
  assign w10110 = w9936 ^ w10109 ;
  assign w10111 = w9917 ^ w10110 ;
  assign w10112 = w9902 ^ w9907 ;
  assign w10113 = \pi008 ^ w10112 ;
  assign w10114 = w10111 ^ w10113 ;
  assign w10115 = ( w9671 & w9679 ) | ( w9671 & w9897 ) | ( w9679 & w9897 ) ;
  assign w10116 = ( w9666 & w9667 ) | ( w9666 & w9899 ) | ( w9667 & w9899 ) ;
  assign w10117 = w10115 ^ w10116 ;
  assign w10118 = w10114 ^ w10117 ;
  assign w10119 = ( w10114 & w10115 ) | ( w10114 & w10116 ) | ( w10115 & w10116 ) ;
  assign w10120 = \pi008 ^ w9907 ;
  assign w10121 = ( w9902 & w10111 ) | ( w9902 & w10120 ) | ( w10111 & w10120 ) ;
  assign w10122 = ( w9915 & w9916 ) | ( w9915 & w10110 ) | ( w9916 & w10110 ) ;
  assign w10123 = w308 & w8481 ;
  assign w10124 = w328 | w10123 ;
  assign w10125 = ( \pi127 & w10123 ) | ( \pi127 & w10124 ) | ( w10123 & w10124 ) ;
  assign w10126 = \pi008 ^ w10125 ;
  assign w10127 = ~\pi119 & w837 ;
  assign w10128 = \pi118 & w902 ;
  assign w10129 = ( w837 & ~w10127 ) | ( w837 & w10128 ) | ( ~w10127 & w10128 ) ;
  assign w10130 = ~\pi120 & w839 ;
  assign w10131 = w6634 | w10129 ;
  assign w10132 = ( w840 & w10129 ) | ( w840 & w10131 ) | ( w10129 & w10131 ) ;
  assign w10133 = ( w839 & ~w10130 ) | ( w839 & w10132 ) | ( ~w10130 & w10132 ) ;
  assign w10134 = \pi017 ^ w10133 ;
  assign w10135 = ( w9944 & w9945 ) | ( w9944 & w10105 ) | ( w9945 & w10105 ) ;
  assign w10136 = ~\pi113 & w1313 ;
  assign w10137 = \pi112 & w1417 ;
  assign w10138 = ( w1313 & ~w10136 ) | ( w1313 & w10137 ) | ( ~w10136 & w10137 ) ;
  assign w10139 = ~\pi114 & w1315 ;
  assign w10140 = w5565 | w10138 ;
  assign w10141 = ( w1316 & w10138 ) | ( w1316 & w10140 ) | ( w10138 & w10140 ) ;
  assign w10142 = ( w1315 & ~w10139 ) | ( w1315 & w10141 ) | ( ~w10139 & w10141 ) ;
  assign w10143 = \pi023 ^ w10142 ;
  assign w10144 = w4792 | w9960 ;
  assign w10145 = ( w1632 & w9960 ) | ( w1632 & w10144 ) | ( w9960 & w10144 ) ;
  assign w10146 = \pi026 ^ w10145 ;
  assign w10147 = ( w9955 & w10098 ) | ( w9955 & w10146 ) | ( w10098 & w10146 ) ;
  assign w10148 = ~\pi110 & w1629 ;
  assign w10149 = \pi109 & w1722 ;
  assign w10150 = ( w1629 & ~w10148 ) | ( w1629 & w10149 ) | ( ~w10148 & w10149 ) ;
  assign w10151 = ~\pi111 & w1631 ;
  assign w10152 = w4811 | w10150 ;
  assign w10153 = ( w1632 & w10150 ) | ( w1632 & w10152 ) | ( w10150 & w10152 ) ;
  assign w10154 = ( w1631 & ~w10151 ) | ( w1631 & w10153 ) | ( ~w10151 & w10153 ) ;
  assign w10155 = \pi026 ^ w10154 ;
  assign w10156 = ( w9968 & w9969 ) | ( w9968 & w10096 ) | ( w9969 & w10096 ) ;
  assign w10157 = ~\pi104 & w2310 ;
  assign w10158 = \pi103 & w2443 ;
  assign w10159 = ( w2310 & ~w10157 ) | ( w2310 & w10158 ) | ( ~w10157 & w10158 ) ;
  assign w10160 = ~\pi105 & w2312 ;
  assign w10161 = w3905 | w10159 ;
  assign w10162 = ( w2313 & w10159 ) | ( w2313 & w10161 ) | ( w10159 & w10161 ) ;
  assign w10163 = ( w2312 & ~w10160 ) | ( w2312 & w10162 ) | ( ~w10160 & w10162 ) ;
  assign w10164 = \pi032 ^ w10163 ;
  assign w10165 = ( w9986 & w9987 ) | ( w9986 & w10092 ) | ( w9987 & w10092 ) ;
  assign w10166 = ~\pi098 & w3178 ;
  assign w10167 = \pi097 & w3340 ;
  assign w10168 = ( w3178 & ~w10166 ) | ( w3178 & w10167 ) | ( ~w10166 & w10167 ) ;
  assign w10169 = ~\pi099 & w3180 ;
  assign w10170 = w2966 | w10168 ;
  assign w10171 = ( w3181 & w10168 ) | ( w3181 & w10170 ) | ( w10168 & w10170 ) ;
  assign w10172 = ( w3180 & ~w10169 ) | ( w3180 & w10171 ) | ( ~w10169 & w10171 ) ;
  assign w10173 = \pi038 ^ w10172 ;
  assign w10174 = ~\pi089 & w4654 ;
  assign w10175 = \pi088 & w4876 ;
  assign w10176 = ( w4654 & ~w10174 ) | ( w4654 & w10175 ) | ( ~w10174 & w10175 ) ;
  assign w10177 = ~\pi090 & w4656 ;
  assign w10178 = w1801 | w10176 ;
  assign w10179 = ( w4657 & w10176 ) | ( w4657 & w10178 ) | ( w10176 & w10178 ) ;
  assign w10180 = ( w4656 & ~w10177 ) | ( w4656 & w10179 ) | ( ~w10177 & w10179 ) ;
  assign w10181 = \pi047 ^ w10180 ;
  assign w10182 = ( w10046 & w10047 ) | ( w10046 & w10055 ) | ( w10047 & w10055 ) ;
  assign w10183 = ~\pi086 & w5209 ;
  assign w10184 = \pi085 & w5433 ;
  assign w10185 = ( w5209 & ~w10183 ) | ( w5209 & w10184 ) | ( ~w10183 & w10184 ) ;
  assign w10186 = ~\pi087 & w5211 ;
  assign w10187 = w1477 | w10185 ;
  assign w10188 = ( w5212 & w10185 ) | ( w5212 & w10187 ) | ( w10185 & w10187 ) ;
  assign w10189 = ( w5211 & ~w10186 ) | ( w5211 & w10188 ) | ( ~w10186 & w10188 ) ;
  assign w10190 = \pi050 ^ w10189 ;
  assign w10191 = ( w10035 & w10036 ) | ( w10035 & w10044 ) | ( w10036 & w10044 ) ;
  assign w10192 = ( w9996 & w10014 ) | ( w9996 & w10022 ) | ( w10014 & w10022 ) ;
  assign w10193 = \pi062 ^ w10008 ;
  assign w10194 = ( \pi062 & \pi063 ) | ( \pi062 & \pi071 ) | ( \pi063 & \pi071 ) ;
  assign w10195 = \pi062 & \pi070 ;
  assign w10196 = ( ~\pi062 & w10194 ) | ( ~\pi062 & w10195 ) | ( w10194 & w10195 ) ;
  assign w10197 = ( ~\pi063 & w10194 ) | ( ~\pi063 & w10196 ) | ( w10194 & w10196 ) ;
  assign w10198 = ( w10001 & ~w10193 ) | ( w10001 & w10197 ) | ( ~w10193 & w10197 ) ;
  assign w10199 = \pi071 & w10198 ;
  assign w10200 = ( \pi063 & ~\pi070 ) | ( \pi063 & w10199 ) | ( ~\pi070 & w10199 ) ;
  assign w10201 = ( \pi062 & ~\pi063 ) | ( \pi062 & w10200 ) | ( ~\pi063 & w10200 ) ;
  assign w10202 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi072 ) | ( \pi063 & ~\pi072 ) ;
  assign w10203 = ( \pi071 & ~w10198 ) | ( \pi071 & w10202 ) | ( ~w10198 & w10202 ) ;
  assign w10204 = ( \pi063 & w10198 ) | ( \pi063 & ~w10199 ) | ( w10198 & ~w10199 ) ;
  assign w10205 = ( ~\pi062 & \pi071 ) | ( ~\pi062 & w10204 ) | ( \pi071 & w10204 ) ;
  assign w10206 = ( w10201 & ~w10203 ) | ( w10201 & w10205 ) | ( ~w10203 & w10205 ) ;
  assign w10207 = \pi070 ^ \pi072 ;
  assign w10208 = ( \pi062 & \pi063 ) | ( \pi062 & ~w10207 ) | ( \pi063 & ~w10207 ) ;
  assign w10209 = \pi070 ^ \pi071 ;
  assign w10210 = \pi062 & ~w10209 ;
  assign w10211 = ( \pi063 & ~w10209 ) | ( \pi063 & w10210 ) | ( ~w10209 & w10210 ) ;
  assign w10212 = w10198 ^ w10211 ;
  assign w10213 = w10208 ^ w10212 ;
  assign w10214 = ~\pi074 & w7811 ;
  assign w10215 = \pi073 & w8046 ;
  assign w10216 = ( w7811 & ~w10214 ) | ( w7811 & w10215 ) | ( ~w10214 & w10215 ) ;
  assign w10217 = ~\pi075 & w7813 ;
  assign w10218 = w519 | w10216 ;
  assign w10219 = ( w7814 & w10216 ) | ( w7814 & w10218 ) | ( w10216 & w10218 ) ;
  assign w10220 = ( w7813 & ~w10217 ) | ( w7813 & w10219 ) | ( ~w10217 & w10219 ) ;
  assign w10221 = \pi062 ^ w10220 ;
  assign w10222 = ~\pi077 & w7135 ;
  assign w10223 = \pi076 & w7359 ;
  assign w10224 = ( w7135 & ~w10222 ) | ( w7135 & w10223 ) | ( ~w10222 & w10223 ) ;
  assign w10225 = ~\pi078 & w7137 ;
  assign w10226 = w665 | w10224 ;
  assign w10227 = ( w7138 & w10224 ) | ( w7138 & w10226 ) | ( w10224 & w10226 ) ;
  assign w10228 = ( w7137 & ~w10225 ) | ( w7137 & w10227 ) | ( ~w10225 & w10227 ) ;
  assign w10229 = \pi059 ^ w10228 ;
  assign w10230 = w10213 ^ w10229 ;
  assign w10231 = w10221 ^ w10230 ;
  assign w10232 = ~\pi080 & w6466 ;
  assign w10233 = \pi079 & w6702 ;
  assign w10234 = ( w6466 & ~w10232 ) | ( w6466 & w10233 ) | ( ~w10232 & w10233 ) ;
  assign w10235 = ~\pi081 & w6468 ;
  assign w10236 = w874 | w10234 ;
  assign w10237 = ( w6469 & w10234 ) | ( w6469 & w10236 ) | ( w10234 & w10236 ) ;
  assign w10238 = ( w6468 & ~w10235 ) | ( w6468 & w10237 ) | ( ~w10235 & w10237 ) ;
  assign w10239 = \pi056 ^ w10238 ;
  assign w10240 = w10192 ^ w10231 ;
  assign w10241 = w10239 ^ w10240 ;
  assign w10242 = ( w10024 & w10025 ) | ( w10024 & w10033 ) | ( w10025 & w10033 ) ;
  assign w10243 = ~\pi083 & w5802 ;
  assign w10244 = \pi082 & w6052 ;
  assign w10245 = ( w5802 & ~w10243 ) | ( w5802 & w10244 ) | ( ~w10243 & w10244 ) ;
  assign w10246 = ~\pi084 & w5804 ;
  assign w10247 = w1188 | w10245 ;
  assign w10248 = ( w5805 & w10245 ) | ( w5805 & w10247 ) | ( w10245 & w10247 ) ;
  assign w10249 = ( w5804 & ~w10246 ) | ( w5804 & w10248 ) | ( ~w10246 & w10248 ) ;
  assign w10250 = \pi053 ^ w10249 ;
  assign w10251 = w10241 ^ w10242 ;
  assign w10252 = w10250 ^ w10251 ;
  assign w10253 = w10191 ^ w10252 ;
  assign w10254 = w10190 ^ w10253 ;
  assign w10255 = w10182 ^ w10254 ;
  assign w10256 = w10181 ^ w10255 ;
  assign w10257 = ( w10057 & w10058 ) | ( w10057 & w10066 ) | ( w10058 & w10066 ) ;
  assign w10258 = ~\pi092 & w4141 ;
  assign w10259 = \pi091 & w4334 ;
  assign w10260 = ( w4141 & ~w10258 ) | ( w4141 & w10259 ) | ( ~w10258 & w10259 ) ;
  assign w10261 = ~\pi093 & w4143 ;
  assign w10262 = w2155 | w10260 ;
  assign w10263 = ( w4144 & w10260 ) | ( w4144 & w10262 ) | ( w10260 & w10262 ) ;
  assign w10264 = ( w4143 & ~w10261 ) | ( w4143 & w10263 ) | ( ~w10261 & w10263 ) ;
  assign w10265 = \pi044 ^ w10264 ;
  assign w10266 = w10256 ^ w10257 ;
  assign w10267 = w10265 ^ w10266 ;
  assign w10268 = ( w10068 & w10069 ) | ( w10068 & w10077 ) | ( w10069 & w10077 ) ;
  assign w10269 = ~\pi095 & w3635 ;
  assign w10270 = \pi094 & w3817 ;
  assign w10271 = ( w3635 & ~w10269 ) | ( w3635 & w10270 ) | ( ~w10269 & w10270 ) ;
  assign w10272 = ~\pi096 & w3637 ;
  assign w10273 = w2546 | w10271 ;
  assign w10274 = ( w3638 & w10271 ) | ( w3638 & w10273 ) | ( w10271 & w10273 ) ;
  assign w10275 = ( w3637 & ~w10272 ) | ( w3637 & w10274 ) | ( ~w10272 & w10274 ) ;
  assign w10276 = \pi041 ^ w10275 ;
  assign w10277 = w10267 ^ w10268 ;
  assign w10278 = w10276 ^ w10277 ;
  assign w10279 = ( w10079 & w10080 ) | ( w10079 & w10088 ) | ( w10080 & w10088 ) ;
  assign w10280 = w10278 ^ w10279 ;
  assign w10281 = w10173 ^ w10280 ;
  assign w10282 = ( w9829 & w9995 ) | ( w9829 & w10090 ) | ( w9995 & w10090 ) ;
  assign w10283 = w10281 ^ w10282 ;
  assign w10284 = ~\pi101 & w2712 ;
  assign w10285 = \pi100 & w2872 ;
  assign w10286 = ( w2712 & ~w10284 ) | ( w2712 & w10285 ) | ( ~w10284 & w10285 ) ;
  assign w10287 = ~\pi102 & w2714 ;
  assign w10288 = w3284 | w10286 ;
  assign w10289 = ( w2715 & w10286 ) | ( w2715 & w10288 ) | ( w10286 & w10288 ) ;
  assign w10290 = ( w2714 & ~w10287 ) | ( w2714 & w10289 ) | ( ~w10287 & w10289 ) ;
  assign w10291 = \pi035 ^ w10290 ;
  assign w10292 = w10164 ^ w10291 ;
  assign w10293 = w10165 ^ w10292 ;
  assign w10294 = w10283 ^ w10293 ;
  assign w10295 = ( w9977 & w9978 ) | ( w9977 & w10094 ) | ( w9978 & w10094 ) ;
  assign w10296 = \pi106 & w2072 ;
  assign w10297 = ( \pi108 & w1946 ) | ( \pi108 & w10296 ) | ( w1946 & w10296 ) ;
  assign w10298 = \pi107 | w10297 ;
  assign w10299 = ( w1944 & w10297 ) | ( w1944 & w10298 ) | ( w10297 & w10298 ) ;
  assign w10300 = w10296 | w10299 ;
  assign w10301 = w1947 & ~w4425 ;
  assign w10302 = ( w1947 & w10300 ) | ( w1947 & ~w10301 ) | ( w10300 & ~w10301 ) ;
  assign w10303 = w10295 ^ w10302 ;
  assign w10304 = \pi029 ^ w10294 ;
  assign w10305 = w10303 ^ w10304 ;
  assign w10306 = w10156 ^ w10305 ;
  assign w10307 = w10155 ^ w10306 ;
  assign w10308 = w10147 ^ w10307 ;
  assign w10309 = w10143 ^ w10308 ;
  assign w10310 = ( w9953 & w9954 ) | ( w9953 & w10103 ) | ( w9954 & w10103 ) ;
  assign w10311 = \pi115 & w1138 ;
  assign w10312 = ( \pi117 & w1046 ) | ( \pi117 & w10311 ) | ( w1046 & w10311 ) ;
  assign w10313 = \pi116 | w10312 ;
  assign w10314 = ( w1044 & w10312 ) | ( w1044 & w10313 ) | ( w10312 & w10313 ) ;
  assign w10315 = w10311 | w10314 ;
  assign w10316 = w1047 & ~w6185 ;
  assign w10317 = ( w1047 & w10315 ) | ( w1047 & ~w10316 ) | ( w10315 & ~w10316 ) ;
  assign w10318 = w10310 ^ w10317 ;
  assign w10319 = \pi020 ^ w10309 ;
  assign w10320 = w10318 ^ w10319 ;
  assign w10321 = w10135 ^ w10320 ;
  assign w10322 = w10134 ^ w10321 ;
  assign w10323 = ~\pi122 & w601 ;
  assign w10324 = \pi121 & w683 ;
  assign w10325 = ( w601 & ~w10323 ) | ( w601 & w10324 ) | ( ~w10323 & w10324 ) ;
  assign w10326 = ~\pi123 & w603 ;
  assign w10327 = w7516 | w10325 ;
  assign w10328 = ( w604 & w10325 ) | ( w604 & w10327 ) | ( w10325 & w10327 ) ;
  assign w10329 = ( w603 & ~w10326 ) | ( w603 & w10328 ) | ( ~w10326 & w10328 ) ;
  assign w10330 = \pi014 ^ w10329 ;
  assign w10331 = ( w9934 & w9935 ) | ( w9934 & w10107 ) | ( w9935 & w10107 ) ;
  assign w10332 = w10322 ^ w10331 ;
  assign w10333 = w10330 ^ w10332 ;
  assign w10334 = w9936 ^ w10107 ;
  assign w10335 = ( w9918 & w9926 ) | ( w9918 & w10334 ) | ( w9926 & w10334 ) ;
  assign w10336 = \pi124 & w486 ;
  assign w10337 = ( \pi126 & w434 ) | ( \pi126 & w10336 ) | ( w434 & w10336 ) ;
  assign w10338 = \pi125 | w10337 ;
  assign w10339 = ( w432 & w10337 ) | ( w432 & w10338 ) | ( w10337 & w10338 ) ;
  assign w10340 = w10336 | w10339 ;
  assign w10341 = w435 & ~w8231 ;
  assign w10342 = ( w435 & w10340 ) | ( w435 & ~w10341 ) | ( w10340 & ~w10341 ) ;
  assign w10343 = w10335 ^ w10342 ;
  assign w10344 = \pi011 ^ w10333 ;
  assign w10345 = w10343 ^ w10344 ;
  assign w10346 = w10122 ^ w10345 ;
  assign w10347 = w10126 ^ w10346 ;
  assign w10348 = w10119 ^ w10121 ;
  assign w10349 = w10347 ^ w10348 ;
  assign w10350 = ( w10119 & w10121 ) | ( w10119 & w10347 ) | ( w10121 & w10347 ) ;
  assign w10351 = ( w10122 & w10126 ) | ( w10122 & w10345 ) | ( w10126 & w10345 ) ;
  assign w10352 = w8231 | w10340 ;
  assign w10353 = ( w435 & w10340 ) | ( w435 & w10352 ) | ( w10340 & w10352 ) ;
  assign w10354 = \pi011 ^ w10353 ;
  assign w10355 = ( w10333 & w10335 ) | ( w10333 & w10354 ) | ( w10335 & w10354 ) ;
  assign w10356 = ~\pi126 & w432 ;
  assign w10357 = \pi125 & w486 ;
  assign w10358 = ( w432 & ~w10356 ) | ( w432 & w10357 ) | ( ~w10356 & w10357 ) ;
  assign w10359 = ~\pi127 & w434 ;
  assign w10360 = w8466 | w10358 ;
  assign w10361 = ( w435 & w10358 ) | ( w435 & w10360 ) | ( w10358 & w10360 ) ;
  assign w10362 = ( w434 & ~w10359 ) | ( w434 & w10361 ) | ( ~w10359 & w10361 ) ;
  assign w10363 = \pi011 ^ w10362 ;
  assign w10364 = ( w10322 & w10330 ) | ( w10322 & w10331 ) | ( w10330 & w10331 ) ;
  assign w10365 = ~\pi123 & w601 ;
  assign w10366 = \pi122 & w683 ;
  assign w10367 = ( w601 & ~w10365 ) | ( w601 & w10366 ) | ( ~w10365 & w10366 ) ;
  assign w10368 = ~\pi124 & w603 ;
  assign w10369 = w7538 | w10367 ;
  assign w10370 = ( w604 & w10367 ) | ( w604 & w10369 ) | ( w10367 & w10369 ) ;
  assign w10371 = ( w603 & ~w10368 ) | ( w603 & w10370 ) | ( ~w10368 & w10370 ) ;
  assign w10372 = \pi014 ^ w10371 ;
  assign w10373 = ~\pi120 & w837 ;
  assign w10374 = \pi119 & w902 ;
  assign w10375 = ( w837 & ~w10373 ) | ( w837 & w10374 ) | ( ~w10373 & w10374 ) ;
  assign w10376 = ~\pi121 & w839 ;
  assign w10377 = w7050 | w10375 ;
  assign w10378 = ( w840 & w10375 ) | ( w840 & w10377 ) | ( w10375 & w10377 ) ;
  assign w10379 = ( w839 & ~w10376 ) | ( w839 & w10378 ) | ( ~w10376 & w10378 ) ;
  assign w10380 = \pi017 ^ w10379 ;
  assign w10381 = ( w10134 & w10135 ) | ( w10134 & w10320 ) | ( w10135 & w10320 ) ;
  assign w10382 = w10380 ^ w10381 ;
  assign w10383 = w6185 | w10315 ;
  assign w10384 = ( w1047 & w10315 ) | ( w1047 & w10383 ) | ( w10315 & w10383 ) ;
  assign w10385 = \pi020 ^ w10384 ;
  assign w10386 = ( w10309 & w10310 ) | ( w10309 & w10385 ) | ( w10310 & w10385 ) ;
  assign w10387 = ~\pi117 & w1044 ;
  assign w10388 = \pi116 & w1138 ;
  assign w10389 = ( w1044 & ~w10387 ) | ( w1044 & w10388 ) | ( ~w10387 & w10388 ) ;
  assign w10390 = ~\pi118 & w1046 ;
  assign w10391 = w6206 | w10389 ;
  assign w10392 = ( w1047 & w10389 ) | ( w1047 & w10391 ) | ( w10389 & w10391 ) ;
  assign w10393 = ( w1046 & ~w10390 ) | ( w1046 & w10392 ) | ( ~w10390 & w10392 ) ;
  assign w10394 = \pi020 ^ w10393 ;
  assign w10395 = ~\pi111 & w1629 ;
  assign w10396 = \pi110 & w1722 ;
  assign w10397 = ( w1629 & ~w10395 ) | ( w1629 & w10396 ) | ( ~w10395 & w10396 ) ;
  assign w10398 = ~\pi112 & w1631 ;
  assign w10399 = w4999 | w10397 ;
  assign w10400 = ( w1632 & w10397 ) | ( w1632 & w10399 ) | ( w10397 & w10399 ) ;
  assign w10401 = ( w1631 & ~w10398 ) | ( w1631 & w10400 ) | ( ~w10398 & w10400 ) ;
  assign w10402 = \pi026 ^ w10401 ;
  assign w10403 = ( w10155 & w10156 ) | ( w10155 & w10305 ) | ( w10156 & w10305 ) ;
  assign w10404 = w4425 | w10300 ;
  assign w10405 = ( w1947 & w10300 ) | ( w1947 & w10404 ) | ( w10300 & w10404 ) ;
  assign w10406 = \pi029 ^ w10405 ;
  assign w10407 = ( w10294 & w10295 ) | ( w10294 & w10406 ) | ( w10295 & w10406 ) ;
  assign w10408 = ~\pi108 & w1944 ;
  assign w10409 = \pi107 & w2072 ;
  assign w10410 = ( w1944 & ~w10408 ) | ( w1944 & w10409 ) | ( ~w10408 & w10409 ) ;
  assign w10411 = ~\pi109 & w1946 ;
  assign w10412 = w4599 | w10410 ;
  assign w10413 = ( w1947 & w10410 ) | ( w1947 & w10412 ) | ( w10410 & w10412 ) ;
  assign w10414 = ( w1946 & ~w10411 ) | ( w1946 & w10413 ) | ( ~w10411 & w10413 ) ;
  assign w10415 = \pi029 ^ w10414 ;
  assign w10416 = w10283 ^ w10291 ;
  assign w10417 = ( w10164 & w10165 ) | ( w10164 & w10416 ) | ( w10165 & w10416 ) ;
  assign w10418 = ~\pi105 & w2310 ;
  assign w10419 = \pi104 & w2443 ;
  assign w10420 = ( w2310 & ~w10418 ) | ( w2310 & w10419 ) | ( ~w10418 & w10419 ) ;
  assign w10421 = ~\pi106 & w2312 ;
  assign w10422 = w4068 | w10420 ;
  assign w10423 = ( w2313 & w10420 ) | ( w2313 & w10422 ) | ( w10420 & w10422 ) ;
  assign w10424 = ( w2312 & ~w10421 ) | ( w2312 & w10423 ) | ( ~w10421 & w10423 ) ;
  assign w10425 = \pi032 ^ w10424 ;
  assign w10426 = ( w10173 & w10278 ) | ( w10173 & w10279 ) | ( w10278 & w10279 ) ;
  assign w10427 = ( w10267 & w10268 ) | ( w10267 & w10276 ) | ( w10268 & w10276 ) ;
  assign w10428 = ( w10256 & w10257 ) | ( w10256 & w10265 ) | ( w10257 & w10265 ) ;
  assign w10429 = ( w10190 & w10191 ) | ( w10190 & w10252 ) | ( w10191 & w10252 ) ;
  assign w10430 = ~\pi087 & w5209 ;
  assign w10431 = \pi086 & w5433 ;
  assign w10432 = ( w5209 & ~w10430 ) | ( w5209 & w10431 ) | ( ~w10430 & w10431 ) ;
  assign w10433 = ~\pi088 & w5211 ;
  assign w10434 = w1574 | w10432 ;
  assign w10435 = ( w5212 & w10432 ) | ( w5212 & w10434 ) | ( w10432 & w10434 ) ;
  assign w10436 = ( w5211 & ~w10433 ) | ( w5211 & w10435 ) | ( ~w10433 & w10435 ) ;
  assign w10437 = \pi050 ^ w10436 ;
  assign w10438 = ~\pi081 & w6466 ;
  assign w10439 = \pi080 & w6702 ;
  assign w10440 = ( w6466 & ~w10438 ) | ( w6466 & w10439 ) | ( ~w10438 & w10439 ) ;
  assign w10441 = ~\pi082 & w6468 ;
  assign w10442 = w1008 | w10440 ;
  assign w10443 = ( w6469 & w10440 ) | ( w6469 & w10442 ) | ( w10440 & w10442 ) ;
  assign w10444 = ( w6468 & ~w10441 ) | ( w6468 & w10443 ) | ( ~w10441 & w10443 ) ;
  assign w10445 = \pi056 ^ w10444 ;
  assign w10446 = ( w10213 & w10221 ) | ( w10213 & w10229 ) | ( w10221 & w10229 ) ;
  assign w10447 = ~\pi075 & w7811 ;
  assign w10448 = \pi074 & w8046 ;
  assign w10449 = ( w7811 & ~w10447 ) | ( w7811 & w10448 ) | ( ~w10447 & w10448 ) ;
  assign w10450 = ~\pi076 & w7813 ;
  assign w10451 = w538 | w10449 ;
  assign w10452 = ( w7814 & w10449 ) | ( w7814 & w10451 ) | ( w10449 & w10451 ) ;
  assign w10453 = ( w7813 & ~w10450 ) | ( w7813 & w10452 ) | ( ~w10450 & w10452 ) ;
  assign w10454 = \pi062 ^ w10453 ;
  assign w10455 = \pi071 ^ \pi073 ;
  assign w10456 = ( \pi062 & \pi063 ) | ( \pi062 & ~w10455 ) | ( \pi063 & ~w10455 ) ;
  assign w10457 = \pi071 ^ \pi072 ;
  assign w10458 = \pi062 & ~w10457 ;
  assign w10459 = ( \pi063 & ~w10457 ) | ( \pi063 & w10458 ) | ( ~w10457 & w10458 ) ;
  assign w10460 = \pi008 ^ w10459 ;
  assign w10461 = w10456 ^ w10460 ;
  assign w10462 = w10206 ^ w10454 ;
  assign w10463 = w10461 ^ w10462 ;
  assign w10464 = ~\pi078 & w7135 ;
  assign w10465 = \pi077 & w7359 ;
  assign w10466 = ( w7135 & ~w10464 ) | ( w7135 & w10465 ) | ( ~w10464 & w10465 ) ;
  assign w10467 = ~\pi079 & w7137 ;
  assign w10468 = w730 | w10466 ;
  assign w10469 = ( w7138 & w10466 ) | ( w7138 & w10468 ) | ( w10466 & w10468 ) ;
  assign w10470 = ( w7137 & ~w10467 ) | ( w7137 & w10469 ) | ( ~w10467 & w10469 ) ;
  assign w10471 = \pi059 ^ w10470 ;
  assign w10472 = w10446 ^ w10463 ;
  assign w10473 = w10471 ^ w10472 ;
  assign w10474 = ( w10192 & w10231 ) | ( w10192 & w10239 ) | ( w10231 & w10239 ) ;
  assign w10475 = w10473 ^ w10474 ;
  assign w10476 = w10445 ^ w10475 ;
  assign w10477 = ~\pi084 & w5802 ;
  assign w10478 = \pi083 & w6052 ;
  assign w10479 = ( w5802 & ~w10477 ) | ( w5802 & w10478 ) | ( ~w10477 & w10478 ) ;
  assign w10480 = ~\pi085 & w5804 ;
  assign w10481 = w1274 | w10479 ;
  assign w10482 = ( w5805 & w10479 ) | ( w5805 & w10481 ) | ( w10479 & w10481 ) ;
  assign w10483 = ( w5804 & ~w10480 ) | ( w5804 & w10482 ) | ( ~w10480 & w10482 ) ;
  assign w10484 = \pi053 ^ w10483 ;
  assign w10485 = ( w10241 & w10242 ) | ( w10241 & w10250 ) | ( w10242 & w10250 ) ;
  assign w10486 = w10476 ^ w10485 ;
  assign w10487 = w10484 ^ w10486 ;
  assign w10488 = w10429 ^ w10487 ;
  assign w10489 = w10437 ^ w10488 ;
  assign w10490 = ~\pi090 & w4654 ;
  assign w10491 = \pi089 & w4876 ;
  assign w10492 = ( w4654 & ~w10490 ) | ( w4654 & w10491 ) | ( ~w10490 & w10491 ) ;
  assign w10493 = ~\pi091 & w4656 ;
  assign w10494 = w1908 | w10492 ;
  assign w10495 = ( w4657 & w10492 ) | ( w4657 & w10494 ) | ( w10492 & w10494 ) ;
  assign w10496 = ( w4656 & ~w10493 ) | ( w4656 & w10495 ) | ( ~w10493 & w10495 ) ;
  assign w10497 = \pi047 ^ w10496 ;
  assign w10498 = ( w10181 & w10182 ) | ( w10181 & w10254 ) | ( w10182 & w10254 ) ;
  assign w10499 = w10489 ^ w10498 ;
  assign w10500 = w10497 ^ w10499 ;
  assign w10501 = ~\pi093 & w4141 ;
  assign w10502 = \pi092 & w4334 ;
  assign w10503 = ( w4141 & ~w10501 ) | ( w4141 & w10502 ) | ( ~w10501 & w10502 ) ;
  assign w10504 = ~\pi094 & w4143 ;
  assign w10505 = w2274 | w10503 ;
  assign w10506 = ( w4144 & w10503 ) | ( w4144 & w10505 ) | ( w10503 & w10505 ) ;
  assign w10507 = ( w4143 & ~w10504 ) | ( w4143 & w10506 ) | ( ~w10504 & w10506 ) ;
  assign w10508 = \pi044 ^ w10507 ;
  assign w10509 = ( w10428 & w10500 ) | ( w10428 & w10508 ) | ( w10500 & w10508 ) ;
  assign w10510 = w10428 ^ w10500 ;
  assign w10511 = w10508 ^ w10510 ;
  assign w10512 = ~\pi096 & w3635 ;
  assign w10513 = \pi095 & w3817 ;
  assign w10514 = ( w3635 & ~w10512 ) | ( w3635 & w10513 ) | ( ~w10512 & w10513 ) ;
  assign w10515 = ~\pi097 & w3637 ;
  assign w10516 = w2673 | w10514 ;
  assign w10517 = ( w3638 & w10514 ) | ( w3638 & w10516 ) | ( w10514 & w10516 ) ;
  assign w10518 = ( w3637 & ~w10515 ) | ( w3637 & w10517 ) | ( ~w10515 & w10517 ) ;
  assign w10519 = \pi041 ^ w10518 ;
  assign w10520 = w10427 ^ w10511 ;
  assign w10521 = w10519 ^ w10520 ;
  assign w10522 = ~\pi099 & w3178 ;
  assign w10523 = \pi098 & w3340 ;
  assign w10524 = ( w3178 & ~w10522 ) | ( w3178 & w10523 ) | ( ~w10522 & w10523 ) ;
  assign w10525 = ~\pi100 & w3180 ;
  assign w10526 = w3104 | w10524 ;
  assign w10527 = ( w3181 & w10524 ) | ( w3181 & w10526 ) | ( w10524 & w10526 ) ;
  assign w10528 = ( w3180 & ~w10525 ) | ( w3180 & w10527 ) | ( ~w10525 & w10527 ) ;
  assign w10529 = \pi038 ^ w10528 ;
  assign w10530 = w10426 ^ w10521 ;
  assign w10531 = w10529 ^ w10530 ;
  assign w10532 = ~\pi102 & w2712 ;
  assign w10533 = \pi101 & w2872 ;
  assign w10534 = ( w2712 & ~w10532 ) | ( w2712 & w10533 ) | ( ~w10532 & w10533 ) ;
  assign w10535 = ~\pi103 & w2714 ;
  assign w10536 = w3437 | w10534 ;
  assign w10537 = ( w2715 & w10534 ) | ( w2715 & w10536 ) | ( w10534 & w10536 ) ;
  assign w10538 = ( w2714 & ~w10535 ) | ( w2714 & w10537 ) | ( ~w10535 & w10537 ) ;
  assign w10539 = \pi035 ^ w10538 ;
  assign w10540 = ( w10281 & w10282 ) | ( w10281 & w10291 ) | ( w10282 & w10291 ) ;
  assign w10541 = w10531 ^ w10540 ;
  assign w10542 = w10539 ^ w10541 ;
  assign w10543 = w10417 ^ w10542 ;
  assign w10544 = w10425 ^ w10543 ;
  assign w10545 = w10407 ^ w10544 ;
  assign w10546 = w10415 ^ w10545 ;
  assign w10547 = w10403 ^ w10546 ;
  assign w10548 = w10402 ^ w10547 ;
  assign w10549 = ~\pi114 & w1313 ;
  assign w10550 = \pi113 & w1417 ;
  assign w10551 = ( w1313 & ~w10549 ) | ( w1313 & w10550 ) | ( ~w10549 & w10550 ) ;
  assign w10552 = ~\pi115 & w1315 ;
  assign w10553 = w5585 | w10551 ;
  assign w10554 = ( w1316 & w10551 ) | ( w1316 & w10553 ) | ( w10551 & w10553 ) ;
  assign w10555 = ( w1315 & ~w10552 ) | ( w1315 & w10554 ) | ( ~w10552 & w10554 ) ;
  assign w10556 = \pi023 ^ w10555 ;
  assign w10557 = ( w10143 & w10147 ) | ( w10143 & w10307 ) | ( w10147 & w10307 ) ;
  assign w10558 = w10548 ^ w10557 ;
  assign w10559 = w10556 ^ w10558 ;
  assign w10560 = w10386 ^ w10559 ;
  assign w10561 = w10394 ^ w10560 ;
  assign w10562 = w10372 ^ w10561 ;
  assign w10563 = w10364 ^ w10562 ;
  assign w10564 = w10382 ^ w10563 ;
  assign w10565 = w10355 ^ w10564 ;
  assign w10566 = w10363 ^ w10565 ;
  assign w10567 = w10350 ^ w10351 ;
  assign w10568 = w10566 ^ w10567 ;
  assign w10569 = ( w10350 & w10351 ) | ( w10350 & w10566 ) | ( w10351 & w10566 ) ;
  assign w10570 = ( w10355 & w10363 ) | ( w10355 & w10564 ) | ( w10363 & w10564 ) ;
  assign w10571 = ~\pi124 & w601 ;
  assign w10572 = \pi123 & w683 ;
  assign w10573 = ( w601 & ~w10571 ) | ( w601 & w10572 ) | ( ~w10571 & w10572 ) ;
  assign w10574 = ~\pi125 & w603 ;
  assign w10575 = w7988 | w10573 ;
  assign w10576 = ( w604 & w10573 ) | ( w604 & w10575 ) | ( w10573 & w10575 ) ;
  assign w10577 = ( w603 & ~w10574 ) | ( w603 & w10576 ) | ( ~w10574 & w10576 ) ;
  assign w10578 = \pi014 ^ w10577 ;
  assign w10579 = ( w10380 & w10381 ) | ( w10380 & w10561 ) | ( w10381 & w10561 ) ;
  assign w10580 = ~\pi118 & w1044 ;
  assign w10581 = \pi117 & w1138 ;
  assign w10582 = ( w1044 & ~w10580 ) | ( w1044 & w10581 ) | ( ~w10580 & w10581 ) ;
  assign w10583 = ~\pi119 & w1046 ;
  assign w10584 = w6616 | w10582 ;
  assign w10585 = ( w1047 & w10582 ) | ( w1047 & w10584 ) | ( w10582 & w10584 ) ;
  assign w10586 = ( w1046 & ~w10583 ) | ( w1046 & w10585 ) | ( ~w10583 & w10585 ) ;
  assign w10587 = \pi020 ^ w10586 ;
  assign w10588 = ( w10548 & w10556 ) | ( w10548 & w10557 ) | ( w10556 & w10557 ) ;
  assign w10589 = ~\pi115 & w1313 ;
  assign w10590 = \pi114 & w1417 ;
  assign w10591 = ( w1313 & ~w10589 ) | ( w1313 & w10590 ) | ( ~w10589 & w10590 ) ;
  assign w10592 = ~\pi116 & w1315 ;
  assign w10593 = w5976 | w10591 ;
  assign w10594 = ( w1316 & w10591 ) | ( w1316 & w10593 ) | ( w10591 & w10593 ) ;
  assign w10595 = ( w1315 & ~w10592 ) | ( w1315 & w10594 ) | ( ~w10592 & w10594 ) ;
  assign w10596 = \pi023 ^ w10595 ;
  assign w10597 = ( w10402 & w10403 ) | ( w10402 & w10546 ) | ( w10403 & w10546 ) ;
  assign w10598 = w10596 ^ w10597 ;
  assign w10599 = ~\pi112 & w1629 ;
  assign w10600 = \pi111 & w1722 ;
  assign w10601 = ( w1629 & ~w10599 ) | ( w1629 & w10600 ) | ( ~w10599 & w10600 ) ;
  assign w10602 = ~\pi113 & w1631 ;
  assign w10603 = w5366 | w10601 ;
  assign w10604 = ( w1632 & w10601 ) | ( w1632 & w10603 ) | ( w10601 & w10603 ) ;
  assign w10605 = ( w1631 & ~w10602 ) | ( w1631 & w10604 ) | ( ~w10602 & w10604 ) ;
  assign w10606 = \pi026 ^ w10605 ;
  assign w10607 = ( w10407 & w10415 ) | ( w10407 & w10544 ) | ( w10415 & w10544 ) ;
  assign w10608 = ~\pi106 & w2310 ;
  assign w10609 = \pi105 & w2443 ;
  assign w10610 = ( w2310 & ~w10608 ) | ( w2310 & w10609 ) | ( ~w10608 & w10609 ) ;
  assign w10611 = ~\pi107 & w2312 ;
  assign w10612 = w4087 | w10610 ;
  assign w10613 = ( w2313 & w10610 ) | ( w2313 & w10612 ) | ( w10610 & w10612 ) ;
  assign w10614 = ( w2312 & ~w10611 ) | ( w2312 & w10613 ) | ( ~w10611 & w10613 ) ;
  assign w10615 = \pi032 ^ w10614 ;
  assign w10616 = ( w10531 & w10539 ) | ( w10531 & w10540 ) | ( w10539 & w10540 ) ;
  assign w10617 = ~\pi103 & w2712 ;
  assign w10618 = \pi102 & w2872 ;
  assign w10619 = ( w2712 & ~w10617 ) | ( w2712 & w10618 ) | ( ~w10617 & w10618 ) ;
  assign w10620 = ~\pi104 & w2714 ;
  assign w10621 = w3740 | w10619 ;
  assign w10622 = ( w2715 & w10619 ) | ( w2715 & w10621 ) | ( w10619 & w10621 ) ;
  assign w10623 = ( w2714 & ~w10620 ) | ( w2714 & w10622 ) | ( ~w10620 & w10622 ) ;
  assign w10624 = \pi035 ^ w10623 ;
  assign w10625 = ( w10426 & w10521 ) | ( w10426 & w10529 ) | ( w10521 & w10529 ) ;
  assign w10626 = ~\pi100 & w3178 ;
  assign w10627 = \pi099 & w3340 ;
  assign w10628 = ( w3178 & ~w10626 ) | ( w3178 & w10627 ) | ( ~w10626 & w10627 ) ;
  assign w10629 = ~\pi101 & w3180 ;
  assign w10630 = w3264 | w10628 ;
  assign w10631 = ( w3181 & w10628 ) | ( w3181 & w10630 ) | ( w10628 & w10630 ) ;
  assign w10632 = ( w3180 & ~w10629 ) | ( w3180 & w10631 ) | ( ~w10629 & w10631 ) ;
  assign w10633 = \pi038 ^ w10632 ;
  assign w10634 = ( w10427 & w10511 ) | ( w10427 & w10519 ) | ( w10511 & w10519 ) ;
  assign w10635 = ~\pi097 & w3635 ;
  assign w10636 = \pi096 & w3817 ;
  assign w10637 = ( w3635 & ~w10635 ) | ( w3635 & w10636 ) | ( ~w10635 & w10636 ) ;
  assign w10638 = ~\pi098 & w3637 ;
  assign w10639 = w2824 | w10637 ;
  assign w10640 = ( w3638 & w10637 ) | ( w3638 & w10639 ) | ( w10637 & w10639 ) ;
  assign w10641 = ( w3637 & ~w10638 ) | ( w3637 & w10640 ) | ( ~w10638 & w10640 ) ;
  assign w10642 = \pi041 ^ w10641 ;
  assign w10643 = ~\pi076 & w7811 ;
  assign w10644 = \pi075 & w8046 ;
  assign w10645 = ( w7811 & ~w10643 ) | ( w7811 & w10644 ) | ( ~w10643 & w10644 ) ;
  assign w10646 = ~\pi077 & w7813 ;
  assign w10647 = w644 | w10645 ;
  assign w10648 = ( w7814 & w10645 ) | ( w7814 & w10647 ) | ( w10645 & w10647 ) ;
  assign w10649 = ( w7813 & ~w10646 ) | ( w7813 & w10648 ) | ( ~w10646 & w10648 ) ;
  assign w10650 = \pi062 ^ w10649 ;
  assign w10651 = ( \pi062 & \pi063 ) | ( \pi062 & \pi074 ) | ( \pi063 & \pi074 ) ;
  assign w10652 = \pi063 & ~\pi073 ;
  assign w10653 = w10651 & ~w10652 ;
  assign w10654 = ( ~\pi062 & w10651 ) | ( ~\pi062 & w10653 ) | ( w10651 & w10653 ) ;
  assign w10655 = \pi062 | \pi063 ;
  assign w10656 = \pi062 ^ w10011 ;
  assign w10657 = ( \pi071 & \pi073 ) | ( \pi071 & w10656 ) | ( \pi073 & w10656 ) ;
  assign w10658 = ( ~\pi008 & \pi072 ) | ( ~\pi008 & w10657 ) | ( \pi072 & w10657 ) ;
  assign w10659 = w10655 & w10658 ;
  assign w10660 = w10650 ^ w10654 ;
  assign w10661 = w10659 ^ w10660 ;
  assign w10662 = ( w10206 & ~w10454 ) | ( w10206 & w10461 ) | ( ~w10454 & w10461 ) ;
  assign w10663 = ~\pi079 & w7135 ;
  assign w10664 = \pi078 & w7359 ;
  assign w10665 = ( w7135 & ~w10663 ) | ( w7135 & w10664 ) | ( ~w10663 & w10664 ) ;
  assign w10666 = ~\pi080 & w7137 ;
  assign w10667 = w794 | w10665 ;
  assign w10668 = ( w7138 & w10665 ) | ( w7138 & w10667 ) | ( w10665 & w10667 ) ;
  assign w10669 = ( w7137 & ~w10666 ) | ( w7137 & w10668 ) | ( ~w10666 & w10668 ) ;
  assign w10670 = \pi059 ^ w10669 ;
  assign w10671 = w10661 ^ w10662 ;
  assign w10672 = w10670 ^ w10671 ;
  assign w10673 = ( w10446 & w10463 ) | ( w10446 & w10471 ) | ( w10463 & w10471 ) ;
  assign w10674 = ~\pi082 & w6466 ;
  assign w10675 = \pi081 & w6702 ;
  assign w10676 = ( w6466 & ~w10674 ) | ( w6466 & w10675 ) | ( ~w10674 & w10675 ) ;
  assign w10677 = ~\pi083 & w6468 ;
  assign w10678 = w1099 | w10676 ;
  assign w10679 = ( w6469 & w10676 ) | ( w6469 & w10678 ) | ( w10676 & w10678 ) ;
  assign w10680 = ( w6468 & ~w10677 ) | ( w6468 & w10679 ) | ( ~w10677 & w10679 ) ;
  assign w10681 = \pi056 ^ w10680 ;
  assign w10682 = w10672 ^ w10673 ;
  assign w10683 = w10681 ^ w10682 ;
  assign w10684 = ( w10445 & w10473 ) | ( w10445 & w10474 ) | ( w10473 & w10474 ) ;
  assign w10685 = ~\pi085 & w5802 ;
  assign w10686 = \pi084 & w6052 ;
  assign w10687 = ( w5802 & ~w10685 ) | ( w5802 & w10686 ) | ( ~w10685 & w10686 ) ;
  assign w10688 = ~\pi086 & w5804 ;
  assign w10689 = w1379 | w10687 ;
  assign w10690 = ( w5805 & w10687 ) | ( w5805 & w10689 ) | ( w10687 & w10689 ) ;
  assign w10691 = ( w5804 & ~w10688 ) | ( w5804 & w10690 ) | ( ~w10688 & w10690 ) ;
  assign w10692 = \pi053 ^ w10691 ;
  assign w10693 = w10683 ^ w10684 ;
  assign w10694 = w10692 ^ w10693 ;
  assign w10695 = ( w10476 & w10484 ) | ( w10476 & w10485 ) | ( w10484 & w10485 ) ;
  assign w10696 = ~\pi088 & w5209 ;
  assign w10697 = \pi087 & w5433 ;
  assign w10698 = ( w5209 & ~w10696 ) | ( w5209 & w10697 ) | ( ~w10696 & w10697 ) ;
  assign w10699 = ~\pi089 & w5211 ;
  assign w10700 = w1595 | w10698 ;
  assign w10701 = ( w5212 & w10698 ) | ( w5212 & w10700 ) | ( w10698 & w10700 ) ;
  assign w10702 = ( w5211 & ~w10699 ) | ( w5211 & w10701 ) | ( ~w10699 & w10701 ) ;
  assign w10703 = \pi050 ^ w10702 ;
  assign w10704 = w10694 ^ w10695 ;
  assign w10705 = w10703 ^ w10704 ;
  assign w10706 = ( w10429 & w10437 ) | ( w10429 & w10487 ) | ( w10437 & w10487 ) ;
  assign w10707 = ~\pi091 & w4654 ;
  assign w10708 = \pi090 & w4876 ;
  assign w10709 = ( w4654 & ~w10707 ) | ( w4654 & w10708 ) | ( ~w10707 & w10708 ) ;
  assign w10710 = ~\pi092 & w4656 ;
  assign w10711 = w2033 | w10709 ;
  assign w10712 = ( w4657 & w10709 ) | ( w4657 & w10711 ) | ( w10709 & w10711 ) ;
  assign w10713 = ( w4656 & ~w10710 ) | ( w4656 & w10712 ) | ( ~w10710 & w10712 ) ;
  assign w10714 = \pi047 ^ w10713 ;
  assign w10715 = w10705 ^ w10706 ;
  assign w10716 = w10714 ^ w10715 ;
  assign w10717 = ( w10489 & w10497 ) | ( w10489 & w10498 ) | ( w10497 & w10498 ) ;
  assign w10718 = ~\pi094 & w4141 ;
  assign w10719 = \pi093 & w4334 ;
  assign w10720 = ( w4141 & ~w10718 ) | ( w4141 & w10719 ) | ( ~w10718 & w10719 ) ;
  assign w10721 = ~\pi095 & w4143 ;
  assign w10722 = w2409 | w10720 ;
  assign w10723 = ( w4144 & w10720 ) | ( w4144 & w10722 ) | ( w10720 & w10722 ) ;
  assign w10724 = ( w4143 & ~w10721 ) | ( w4143 & w10723 ) | ( ~w10721 & w10723 ) ;
  assign w10725 = \pi044 ^ w10724 ;
  assign w10726 = w10716 ^ w10717 ;
  assign w10727 = w10725 ^ w10726 ;
  assign w10728 = w10509 ^ w10727 ;
  assign w10729 = w10642 ^ w10728 ;
  assign w10730 = w10634 ^ w10729 ;
  assign w10731 = w10633 ^ w10730 ;
  assign w10732 = w10625 ^ w10731 ;
  assign w10733 = w10624 ^ w10732 ;
  assign w10734 = w10616 ^ w10733 ;
  assign w10735 = w10615 ^ w10734 ;
  assign w10736 = ( w10417 & w10425 ) | ( w10417 & w10542 ) | ( w10425 & w10542 ) ;
  assign w10737 = \pi108 & w2072 ;
  assign w10738 = ( \pi110 & w1946 ) | ( \pi110 & w10737 ) | ( w1946 & w10737 ) ;
  assign w10739 = \pi109 | w10738 ;
  assign w10740 = ( w1944 & w10738 ) | ( w1944 & w10739 ) | ( w10738 & w10739 ) ;
  assign w10741 = w10737 | w10740 ;
  assign w10742 = w1947 & ~w4792 ;
  assign w10743 = ( w1947 & w10741 ) | ( w1947 & ~w10742 ) | ( w10741 & ~w10742 ) ;
  assign w10744 = w10736 ^ w10743 ;
  assign w10745 = \pi029 ^ w10735 ;
  assign w10746 = w10744 ^ w10745 ;
  assign w10747 = w10607 ^ w10746 ;
  assign w10748 = w10606 ^ w10747 ;
  assign w10749 = w10587 ^ w10748 ;
  assign w10750 = w10588 ^ w10749 ;
  assign w10751 = w10598 ^ w10750 ;
  assign w10752 = ( w10386 & w10394 ) | ( w10386 & w10559 ) | ( w10394 & w10559 ) ;
  assign w10753 = \pi120 & w902 ;
  assign w10754 = ( \pi122 & w839 ) | ( \pi122 & w10753 ) | ( w839 & w10753 ) ;
  assign w10755 = \pi121 | w10754 ;
  assign w10756 = ( w837 & w10754 ) | ( w837 & w10755 ) | ( w10754 & w10755 ) ;
  assign w10757 = w10753 | w10756 ;
  assign w10758 = w840 & ~w7069 ;
  assign w10759 = ( w840 & w10757 ) | ( w840 & ~w10758 ) | ( w10757 & ~w10758 ) ;
  assign w10760 = w10752 ^ w10759 ;
  assign w10761 = \pi017 ^ w10751 ;
  assign w10762 = w10760 ^ w10761 ;
  assign w10763 = w10579 ^ w10762 ;
  assign w10764 = w10578 ^ w10763 ;
  assign w10765 = w10382 ^ w10561 ;
  assign w10766 = ( w10364 & w10372 ) | ( w10364 & w10765 ) | ( w10372 & w10765 ) ;
  assign w10767 = \pi127 & w432 ;
  assign w10768 = ( \pi126 & ~w435 ) | ( \pi126 & w8490 ) | ( ~w435 & w8490 ) ;
  assign w10769 = \pi126 & ~w486 ;
  assign w10770 = ( ~\pi126 & w10768 ) | ( ~\pi126 & w10769 ) | ( w10768 & w10769 ) ;
  assign w10771 = ( w9420 & w10767 ) | ( w9420 & ~w10770 ) | ( w10767 & ~w10770 ) ;
  assign w10772 = \pi011 ^ w10771 ;
  assign w10773 = w10766 ^ w10772 ;
  assign w10774 = w10764 ^ w10773 ;
  assign w10775 = w10569 ^ w10570 ;
  assign w10776 = w10774 ^ w10775 ;
  assign w10777 = ( w10569 & w10570 ) | ( w10569 & w10774 ) | ( w10570 & w10774 ) ;
  assign w10778 = ( w10764 & w10766 ) | ( w10764 & w10772 ) | ( w10766 & w10772 ) ;
  assign w10779 = ( w10578 & w10579 ) | ( w10578 & w10762 ) | ( w10579 & w10762 ) ;
  assign w10780 = w435 & w8481 ;
  assign w10781 = w486 | w10780 ;
  assign w10782 = ( \pi127 & w10780 ) | ( \pi127 & w10781 ) | ( w10780 & w10781 ) ;
  assign w10783 = \pi011 ^ w10782 ;
  assign w10784 = w7069 | w10757 ;
  assign w10785 = ( w840 & w10757 ) | ( w840 & w10784 ) | ( w10757 & w10784 ) ;
  assign w10786 = \pi017 ^ w10785 ;
  assign w10787 = ( w10751 & w10752 ) | ( w10751 & w10786 ) | ( w10752 & w10786 ) ;
  assign w10788 = \pi124 & w683 ;
  assign w10789 = ( \pi126 & w603 ) | ( \pi126 & w10788 ) | ( w603 & w10788 ) ;
  assign w10790 = \pi125 | w10789 ;
  assign w10791 = ( w601 & w10789 ) | ( w601 & w10790 ) | ( w10789 & w10790 ) ;
  assign w10792 = w10788 | w10791 ;
  assign w10793 = ~w604 & w8231 ;
  assign w10794 = ( w8231 & w10792 ) | ( w8231 & ~w10793 ) | ( w10792 & ~w10793 ) ;
  assign w10795 = \pi014 ^ w10794 ;
  assign w10796 = ~\pi122 & w837 ;
  assign w10797 = \pi121 & w902 ;
  assign w10798 = ( w837 & ~w10796 ) | ( w837 & w10797 ) | ( ~w10796 & w10797 ) ;
  assign w10799 = ~\pi123 & w839 ;
  assign w10800 = w7516 | w10798 ;
  assign w10801 = ( w840 & w10798 ) | ( w840 & w10800 ) | ( w10798 & w10800 ) ;
  assign w10802 = ( w839 & ~w10799 ) | ( w839 & w10801 ) | ( ~w10799 & w10801 ) ;
  assign w10803 = \pi017 ^ w10802 ;
  assign w10804 = w10598 ^ w10748 ;
  assign w10805 = ( w10587 & w10588 ) | ( w10587 & w10804 ) | ( w10588 & w10804 ) ;
  assign w10806 = w10803 ^ w10805 ;
  assign w10807 = ~\pi119 & w1044 ;
  assign w10808 = \pi118 & w1138 ;
  assign w10809 = ( w1044 & ~w10807 ) | ( w1044 & w10808 ) | ( ~w10807 & w10808 ) ;
  assign w10810 = ~\pi120 & w1046 ;
  assign w10811 = w6634 | w10809 ;
  assign w10812 = ( w1047 & w10809 ) | ( w1047 & w10811 ) | ( w10809 & w10811 ) ;
  assign w10813 = ( w1046 & ~w10810 ) | ( w1046 & w10812 ) | ( ~w10810 & w10812 ) ;
  assign w10814 = \pi020 ^ w10813 ;
  assign w10815 = ( w10596 & w10597 ) | ( w10596 & w10748 ) | ( w10597 & w10748 ) ;
  assign w10816 = w4792 | w10741 ;
  assign w10817 = ( w1947 & w10741 ) | ( w1947 & w10816 ) | ( w10741 & w10816 ) ;
  assign w10818 = \pi029 ^ w10817 ;
  assign w10819 = ( w10735 & w10736 ) | ( w10735 & w10818 ) | ( w10736 & w10818 ) ;
  assign w10820 = \pi112 & w1722 ;
  assign w10821 = ( \pi114 & w1631 ) | ( \pi114 & w10820 ) | ( w1631 & w10820 ) ;
  assign w10822 = \pi113 | w10821 ;
  assign w10823 = ( w1629 & w10821 ) | ( w1629 & w10822 ) | ( w10821 & w10822 ) ;
  assign w10824 = w10820 | w10823 ;
  assign w10825 = ~w1632 & w5565 ;
  assign w10826 = ( w5565 & w10824 ) | ( w5565 & ~w10825 ) | ( w10824 & ~w10825 ) ;
  assign w10827 = \pi026 ^ w10826 ;
  assign w10828 = ~\pi110 & w1944 ;
  assign w10829 = \pi109 & w2072 ;
  assign w10830 = ( w1944 & ~w10828 ) | ( w1944 & w10829 ) | ( ~w10828 & w10829 ) ;
  assign w10831 = ~\pi111 & w1946 ;
  assign w10832 = w4811 | w10830 ;
  assign w10833 = ( w1947 & w10830 ) | ( w1947 & w10832 ) | ( w10830 & w10832 ) ;
  assign w10834 = ( w1946 & ~w10831 ) | ( w1946 & w10833 ) | ( ~w10831 & w10833 ) ;
  assign w10835 = \pi029 ^ w10834 ;
  assign w10836 = ( w10615 & w10616 ) | ( w10615 & w10733 ) | ( w10616 & w10733 ) ;
  assign w10837 = w10835 ^ w10836 ;
  assign w10838 = ( w10624 & w10625 ) | ( w10624 & w10731 ) | ( w10625 & w10731 ) ;
  assign w10839 = \pi106 & w2443 ;
  assign w10840 = ( \pi108 & w2312 ) | ( \pi108 & w10839 ) | ( w2312 & w10839 ) ;
  assign w10841 = \pi107 | w10840 ;
  assign w10842 = ( w2310 & w10840 ) | ( w2310 & w10841 ) | ( w10840 & w10841 ) ;
  assign w10843 = w10839 | w10842 ;
  assign w10844 = ~\pi104 & w2712 ;
  assign w10845 = \pi103 & w2872 ;
  assign w10846 = ( w2712 & ~w10844 ) | ( w2712 & w10845 ) | ( ~w10844 & w10845 ) ;
  assign w10847 = ~\pi105 & w2714 ;
  assign w10848 = w3905 | w10846 ;
  assign w10849 = ( w2715 & w10846 ) | ( w2715 & w10848 ) | ( w10846 & w10848 ) ;
  assign w10850 = ( w2714 & ~w10847 ) | ( w2714 & w10849 ) | ( ~w10847 & w10849 ) ;
  assign w10851 = \pi035 ^ w10850 ;
  assign w10852 = ( w10633 & w10634 ) | ( w10633 & w10729 ) | ( w10634 & w10729 ) ;
  assign w10853 = ~\pi098 & w3635 ;
  assign w10854 = \pi097 & w3817 ;
  assign w10855 = ( w3635 & ~w10853 ) | ( w3635 & w10854 ) | ( ~w10853 & w10854 ) ;
  assign w10856 = ~\pi099 & w3637 ;
  assign w10857 = w2966 | w10855 ;
  assign w10858 = ( w3638 & w10855 ) | ( w3638 & w10857 ) | ( w10855 & w10857 ) ;
  assign w10859 = ( w3637 & ~w10856 ) | ( w3637 & w10858 ) | ( ~w10856 & w10858 ) ;
  assign w10860 = \pi041 ^ w10859 ;
  assign w10861 = ( w10694 & w10695 ) | ( w10694 & w10703 ) | ( w10695 & w10703 ) ;
  assign w10862 = ~\pi089 & w5209 ;
  assign w10863 = \pi088 & w5433 ;
  assign w10864 = ( w5209 & ~w10862 ) | ( w5209 & w10863 ) | ( ~w10862 & w10863 ) ;
  assign w10865 = ~\pi090 & w5211 ;
  assign w10866 = w1801 | w10864 ;
  assign w10867 = ( w5212 & w10864 ) | ( w5212 & w10866 ) | ( w10864 & w10866 ) ;
  assign w10868 = ( w5211 & ~w10865 ) | ( w5211 & w10867 ) | ( ~w10865 & w10867 ) ;
  assign w10869 = \pi050 ^ w10868 ;
  assign w10870 = ( w10683 & w10684 ) | ( w10683 & w10692 ) | ( w10684 & w10692 ) ;
  assign w10871 = ~\pi086 & w5802 ;
  assign w10872 = \pi085 & w6052 ;
  assign w10873 = ( w5802 & ~w10871 ) | ( w5802 & w10872 ) | ( ~w10871 & w10872 ) ;
  assign w10874 = ~\pi087 & w5804 ;
  assign w10875 = w1477 | w10873 ;
  assign w10876 = ( w5805 & w10873 ) | ( w5805 & w10875 ) | ( w10873 & w10875 ) ;
  assign w10877 = ( w5804 & ~w10874 ) | ( w5804 & w10876 ) | ( ~w10874 & w10876 ) ;
  assign w10878 = \pi053 ^ w10877 ;
  assign w10879 = ( w10672 & w10673 ) | ( w10672 & w10681 ) | ( w10673 & w10681 ) ;
  assign w10880 = ( w10650 & ~w10654 ) | ( w10650 & w10659 ) | ( ~w10654 & w10659 ) ;
  assign w10881 = \pi073 ^ \pi075 ;
  assign w10882 = ( \pi062 & \pi063 ) | ( \pi062 & ~w10881 ) | ( \pi063 & ~w10881 ) ;
  assign w10883 = \pi073 ^ \pi074 ;
  assign w10884 = \pi062 & ~w10883 ;
  assign w10885 = ( \pi063 & ~w10883 ) | ( \pi063 & w10884 ) | ( ~w10883 & w10884 ) ;
  assign w10886 = w10880 ^ w10885 ;
  assign w10887 = w10882 ^ w10886 ;
  assign w10888 = ~\pi077 & w7811 ;
  assign w10889 = \pi076 & w8046 ;
  assign w10890 = ( w7811 & ~w10888 ) | ( w7811 & w10889 ) | ( ~w10888 & w10889 ) ;
  assign w10891 = ~\pi078 & w7813 ;
  assign w10892 = w665 | w10890 ;
  assign w10893 = ( w7814 & w10890 ) | ( w7814 & w10892 ) | ( w10890 & w10892 ) ;
  assign w10894 = ( w7813 & ~w10891 ) | ( w7813 & w10893 ) | ( ~w10891 & w10893 ) ;
  assign w10895 = \pi062 ^ w10894 ;
  assign w10896 = ~\pi080 & w7135 ;
  assign w10897 = \pi079 & w7359 ;
  assign w10898 = ( w7135 & ~w10896 ) | ( w7135 & w10897 ) | ( ~w10896 & w10897 ) ;
  assign w10899 = ~\pi081 & w7137 ;
  assign w10900 = w874 | w10898 ;
  assign w10901 = ( w7138 & w10898 ) | ( w7138 & w10900 ) | ( w10898 & w10900 ) ;
  assign w10902 = ( w7137 & ~w10899 ) | ( w7137 & w10901 ) | ( ~w10899 & w10901 ) ;
  assign w10903 = \pi059 ^ w10902 ;
  assign w10904 = w10887 ^ w10895 ;
  assign w10905 = w10903 ^ w10904 ;
  assign w10906 = ( w10661 & w10662 ) | ( w10661 & ~w10670 ) | ( w10662 & ~w10670 ) ;
  assign w10907 = ~\pi083 & w6466 ;
  assign w10908 = \pi082 & w6702 ;
  assign w10909 = ( w6466 & ~w10907 ) | ( w6466 & w10908 ) | ( ~w10907 & w10908 ) ;
  assign w10910 = ~\pi084 & w6468 ;
  assign w10911 = w1188 | w10909 ;
  assign w10912 = ( w6469 & w10909 ) | ( w6469 & w10911 ) | ( w10909 & w10911 ) ;
  assign w10913 = ( w6468 & ~w10910 ) | ( w6468 & w10912 ) | ( ~w10910 & w10912 ) ;
  assign w10914 = \pi056 ^ w10913 ;
  assign w10915 = w10905 ^ w10906 ;
  assign w10916 = w10914 ^ w10915 ;
  assign w10917 = w10879 ^ w10916 ;
  assign w10918 = w10878 ^ w10917 ;
  assign w10919 = w10870 ^ w10918 ;
  assign w10920 = w10869 ^ w10919 ;
  assign w10921 = ~\pi092 & w4654 ;
  assign w10922 = \pi091 & w4876 ;
  assign w10923 = ( w4654 & ~w10921 ) | ( w4654 & w10922 ) | ( ~w10921 & w10922 ) ;
  assign w10924 = ~\pi093 & w4656 ;
  assign w10925 = w2155 | w10923 ;
  assign w10926 = ( w4657 & w10923 ) | ( w4657 & w10925 ) | ( w10923 & w10925 ) ;
  assign w10927 = ( w4656 & ~w10924 ) | ( w4656 & w10926 ) | ( ~w10924 & w10926 ) ;
  assign w10928 = \pi047 ^ w10927 ;
  assign w10929 = w10861 ^ w10920 ;
  assign w10930 = w10928 ^ w10929 ;
  assign w10931 = ( w10705 & w10706 ) | ( w10705 & w10714 ) | ( w10706 & w10714 ) ;
  assign w10932 = ~\pi095 & w4141 ;
  assign w10933 = \pi094 & w4334 ;
  assign w10934 = ( w4141 & ~w10932 ) | ( w4141 & w10933 ) | ( ~w10932 & w10933 ) ;
  assign w10935 = ~\pi096 & w4143 ;
  assign w10936 = w2546 | w10934 ;
  assign w10937 = ( w4144 & w10934 ) | ( w4144 & w10936 ) | ( w10934 & w10936 ) ;
  assign w10938 = ( w4143 & ~w10935 ) | ( w4143 & w10937 ) | ( ~w10935 & w10937 ) ;
  assign w10939 = \pi044 ^ w10938 ;
  assign w10940 = w10930 ^ w10931 ;
  assign w10941 = w10939 ^ w10940 ;
  assign w10942 = ( w10716 & w10717 ) | ( w10716 & w10725 ) | ( w10717 & w10725 ) ;
  assign w10943 = w10941 ^ w10942 ;
  assign w10944 = w10860 ^ w10943 ;
  assign w10945 = ( w10509 & w10642 ) | ( w10509 & w10727 ) | ( w10642 & w10727 ) ;
  assign w10946 = ~\pi101 & w3178 ;
  assign w10947 = \pi100 & w3340 ;
  assign w10948 = ( w3178 & ~w10946 ) | ( w3178 & w10947 ) | ( ~w10946 & w10947 ) ;
  assign w10949 = ~\pi102 & w3180 ;
  assign w10950 = w3284 | w10948 ;
  assign w10951 = ( w3181 & w10948 ) | ( w3181 & w10950 ) | ( w10948 & w10950 ) ;
  assign w10952 = ( w3180 & ~w10949 ) | ( w3180 & w10951 ) | ( ~w10949 & w10951 ) ;
  assign w10953 = \pi038 ^ w10952 ;
  assign w10954 = w10944 ^ w10945 ;
  assign w10955 = w10953 ^ w10954 ;
  assign w10956 = w10852 ^ w10955 ;
  assign w10957 = w10851 ^ w10956 ;
  assign w10958 = w2313 & ~w4425 ;
  assign w10959 = ( w2313 & w10843 ) | ( w2313 & ~w10958 ) | ( w10843 & ~w10958 ) ;
  assign w10960 = w10838 ^ w10959 ;
  assign w10961 = \pi032 ^ w10957 ;
  assign w10962 = w10960 ^ w10961 ;
  assign w10963 = w10827 ^ w10962 ;
  assign w10964 = w10819 ^ w10963 ;
  assign w10965 = w10837 ^ w10964 ;
  assign w10966 = ( w10606 & w10607 ) | ( w10606 & w10746 ) | ( w10607 & w10746 ) ;
  assign w10967 = \pi115 & w1417 ;
  assign w10968 = ( \pi117 & w1315 ) | ( \pi117 & w10967 ) | ( w1315 & w10967 ) ;
  assign w10969 = \pi116 | w10968 ;
  assign w10970 = ( w1313 & w10968 ) | ( w1313 & w10969 ) | ( w10968 & w10969 ) ;
  assign w10971 = w10967 | w10970 ;
  assign w10972 = w1316 & ~w6185 ;
  assign w10973 = ( w1316 & w10971 ) | ( w1316 & ~w10972 ) | ( w10971 & ~w10972 ) ;
  assign w10974 = w10966 ^ w10973 ;
  assign w10975 = \pi023 ^ w10965 ;
  assign w10976 = w10974 ^ w10975 ;
  assign w10977 = w10815 ^ w10976 ;
  assign w10978 = w10814 ^ w10977 ;
  assign w10979 = w10795 ^ w10978 ;
  assign w10980 = w10787 ^ w10979 ;
  assign w10981 = w10806 ^ w10980 ;
  assign w10982 = w10779 ^ w10981 ;
  assign w10983 = w10783 ^ w10982 ;
  assign w10984 = w10777 ^ w10778 ;
  assign w10985 = w10983 ^ w10984 ;
  assign w10986 = ( w10777 & w10778 ) | ( w10777 & w10983 ) | ( w10778 & w10983 ) ;
  assign w10987 = ( w10779 & w10783 ) | ( w10779 & w10981 ) | ( w10783 & w10981 ) ;
  assign w10988 = w10806 ^ w10978 ;
  assign w10989 = ( w10787 & w10795 ) | ( w10787 & w10988 ) | ( w10795 & w10988 ) ;
  assign w10990 = ~\pi126 & w601 ;
  assign w10991 = \pi125 & w683 ;
  assign w10992 = ( w601 & ~w10990 ) | ( w601 & w10991 ) | ( ~w10990 & w10991 ) ;
  assign w10993 = ~\pi127 & w603 ;
  assign w10994 = w8466 | w10992 ;
  assign w10995 = ( w604 & w10992 ) | ( w604 & w10994 ) | ( w10992 & w10994 ) ;
  assign w10996 = ( w603 & ~w10993 ) | ( w603 & w10995 ) | ( ~w10993 & w10995 ) ;
  assign w10997 = \pi014 ^ w10996 ;
  assign w10998 = ( w10803 & w10805 ) | ( w10803 & w10978 ) | ( w10805 & w10978 ) ;
  assign w10999 = ~\pi123 & w837 ;
  assign w11000 = \pi122 & w902 ;
  assign w11001 = ( w837 & ~w10999 ) | ( w837 & w11000 ) | ( ~w10999 & w11000 ) ;
  assign w11002 = ~\pi124 & w839 ;
  assign w11003 = w7538 | w11001 ;
  assign w11004 = ( w840 & w11001 ) | ( w840 & w11003 ) | ( w11001 & w11003 ) ;
  assign w11005 = ( w839 & ~w11002 ) | ( w839 & w11004 ) | ( ~w11002 & w11004 ) ;
  assign w11006 = \pi017 ^ w11005 ;
  assign w11007 = ~\pi120 & w1044 ;
  assign w11008 = \pi119 & w1138 ;
  assign w11009 = ( w1044 & ~w11007 ) | ( w1044 & w11008 ) | ( ~w11007 & w11008 ) ;
  assign w11010 = ~\pi121 & w1046 ;
  assign w11011 = w7050 | w11009 ;
  assign w11012 = ( w1047 & w11009 ) | ( w1047 & w11011 ) | ( w11009 & w11011 ) ;
  assign w11013 = ( w1046 & ~w11010 ) | ( w1046 & w11012 ) | ( ~w11010 & w11012 ) ;
  assign w11014 = \pi020 ^ w11013 ;
  assign w11015 = ( w10814 & w10815 ) | ( w10814 & w10976 ) | ( w10815 & w10976 ) ;
  assign w11016 = w11014 ^ w11015 ;
  assign w11017 = w6185 | w10971 ;
  assign w11018 = ( w1316 & w10971 ) | ( w1316 & w11017 ) | ( w10971 & w11017 ) ;
  assign w11019 = \pi023 ^ w11018 ;
  assign w11020 = ( w10965 & w10966 ) | ( w10965 & w11019 ) | ( w10966 & w11019 ) ;
  assign w11021 = ~\pi117 & w1313 ;
  assign w11022 = \pi116 & w1417 ;
  assign w11023 = ( w1313 & ~w11021 ) | ( w1313 & w11022 ) | ( ~w11021 & w11022 ) ;
  assign w11024 = ~\pi118 & w1315 ;
  assign w11025 = w6206 | w11023 ;
  assign w11026 = ( w1316 & w11023 ) | ( w1316 & w11025 ) | ( w11023 & w11025 ) ;
  assign w11027 = ( w1315 & ~w11024 ) | ( w1315 & w11026 ) | ( ~w11024 & w11026 ) ;
  assign w11028 = \pi023 ^ w11027 ;
  assign w11029 = ~\pi114 & w1629 ;
  assign w11030 = \pi113 & w1722 ;
  assign w11031 = ( w1629 & ~w11029 ) | ( w1629 & w11030 ) | ( ~w11029 & w11030 ) ;
  assign w11032 = ~\pi115 & w1631 ;
  assign w11033 = w5585 | w11031 ;
  assign w11034 = ( w1632 & w11031 ) | ( w1632 & w11033 ) | ( w11031 & w11033 ) ;
  assign w11035 = ( w1631 & ~w11032 ) | ( w1631 & w11034 ) | ( ~w11032 & w11034 ) ;
  assign w11036 = \pi026 ^ w11035 ;
  assign w11037 = w10837 ^ w10962 ;
  assign w11038 = ( w10819 & w10827 ) | ( w10819 & w11037 ) | ( w10827 & w11037 ) ;
  assign w11039 = w11036 ^ w11038 ;
  assign w11040 = ( w10835 & w10836 ) | ( w10835 & w10962 ) | ( w10836 & w10962 ) ;
  assign w11041 = ~\pi111 & w1944 ;
  assign w11042 = \pi110 & w2072 ;
  assign w11043 = ( w1944 & ~w11041 ) | ( w1944 & w11042 ) | ( ~w11041 & w11042 ) ;
  assign w11044 = ~\pi112 & w1946 ;
  assign w11045 = w4999 | w11043 ;
  assign w11046 = ( w1947 & w11043 ) | ( w1947 & w11045 ) | ( w11043 & w11045 ) ;
  assign w11047 = ( w1946 & ~w11044 ) | ( w1946 & w11046 ) | ( ~w11044 & w11046 ) ;
  assign w11048 = \pi029 ^ w11047 ;
  assign w11049 = ( w10851 & w10852 ) | ( w10851 & w10955 ) | ( w10852 & w10955 ) ;
  assign w11050 = ( w10944 & w10945 ) | ( w10944 & w10953 ) | ( w10945 & w10953 ) ;
  assign w11051 = ( w10860 & w10941 ) | ( w10860 & w10942 ) | ( w10941 & w10942 ) ;
  assign w11052 = ( w10930 & w10931 ) | ( w10930 & w10939 ) | ( w10931 & w10939 ) ;
  assign w11053 = ( w10861 & w10920 ) | ( w10861 & w10928 ) | ( w10920 & w10928 ) ;
  assign w11054 = ( w10878 & w10879 ) | ( w10878 & w10916 ) | ( w10879 & w10916 ) ;
  assign w11055 = ~\pi087 & w5802 ;
  assign w11056 = \pi086 & w6052 ;
  assign w11057 = ( w5802 & ~w11055 ) | ( w5802 & w11056 ) | ( ~w11055 & w11056 ) ;
  assign w11058 = ~\pi088 & w5804 ;
  assign w11059 = w1574 | w11057 ;
  assign w11060 = ( w5805 & w11057 ) | ( w5805 & w11059 ) | ( w11057 & w11059 ) ;
  assign w11061 = ( w5804 & ~w11058 ) | ( w5804 & w11060 ) | ( ~w11058 & w11060 ) ;
  assign w11062 = \pi053 ^ w11061 ;
  assign w11063 = \pi074 | w10880 ;
  assign w11064 = ( \pi063 & \pi073 ) | ( \pi063 & ~w11063 ) | ( \pi073 & ~w11063 ) ;
  assign w11065 = ( \pi062 & ~\pi063 ) | ( \pi062 & w11064 ) | ( ~\pi063 & w11064 ) ;
  assign w11066 = ( \pi062 & \pi063 ) | ( \pi062 & \pi075 ) | ( \pi063 & \pi075 ) ;
  assign w11067 = ( ~\pi074 & w10880 ) | ( ~\pi074 & w11066 ) | ( w10880 & w11066 ) ;
  assign w11068 = ( \pi063 & ~w10880 ) | ( \pi063 & w11063 ) | ( ~w10880 & w11063 ) ;
  assign w11069 = ( \pi062 & \pi074 ) | ( \pi062 & ~w11068 ) | ( \pi074 & ~w11068 ) ;
  assign w11070 = ( ~w11065 & w11067 ) | ( ~w11065 & w11069 ) | ( w11067 & w11069 ) ;
  assign w11071 = ~\pi078 & w7811 ;
  assign w11072 = \pi077 & w8046 ;
  assign w11073 = ( w7811 & ~w11071 ) | ( w7811 & w11072 ) | ( ~w11071 & w11072 ) ;
  assign w11074 = ~\pi079 & w7813 ;
  assign w11075 = w730 | w11073 ;
  assign w11076 = ( w7814 & w11073 ) | ( w7814 & w11075 ) | ( w11073 & w11075 ) ;
  assign w11077 = ( w7813 & ~w11074 ) | ( w7813 & w11076 ) | ( ~w11074 & w11076 ) ;
  assign w11078 = \pi062 ^ w11077 ;
  assign w11079 = \pi011 ^ w10654 ;
  assign w11080 = ( \pi062 & \pi063 ) | ( \pi062 & \pi076 ) | ( \pi063 & \pi076 ) ;
  assign w11081 = \pi063 & ~\pi075 ;
  assign w11082 = \pi062 & w11081 ;
  assign w11083 = w11080 ^ w11082 ;
  assign w11084 = w11079 ^ w11083 ;
  assign w11085 = w11070 ^ w11078 ;
  assign w11086 = w11084 ^ w11085 ;
  assign w11087 = ~\pi081 & w7135 ;
  assign w11088 = \pi080 & w7359 ;
  assign w11089 = ( w7135 & ~w11087 ) | ( w7135 & w11088 ) | ( ~w11087 & w11088 ) ;
  assign w11090 = ~\pi082 & w7137 ;
  assign w11091 = w1008 | w11089 ;
  assign w11092 = ( w7138 & w11089 ) | ( w7138 & w11091 ) | ( w11089 & w11091 ) ;
  assign w11093 = ( w7137 & ~w11090 ) | ( w7137 & w11092 ) | ( ~w11090 & w11092 ) ;
  assign w11094 = \pi059 ^ w11093 ;
  assign w11095 = ( ~w10887 & w10895 ) | ( ~w10887 & w10903 ) | ( w10895 & w10903 ) ;
  assign w11096 = w11086 ^ w11095 ;
  assign w11097 = w11094 ^ w11096 ;
  assign w11098 = ~\pi084 & w6466 ;
  assign w11099 = \pi083 & w6702 ;
  assign w11100 = ( w6466 & ~w11098 ) | ( w6466 & w11099 ) | ( ~w11098 & w11099 ) ;
  assign w11101 = ~\pi085 & w6468 ;
  assign w11102 = w1274 | w11100 ;
  assign w11103 = ( w6469 & w11100 ) | ( w6469 & w11102 ) | ( w11100 & w11102 ) ;
  assign w11104 = ( w6468 & ~w11101 ) | ( w6468 & w11103 ) | ( ~w11101 & w11103 ) ;
  assign w11105 = \pi056 ^ w11104 ;
  assign w11106 = ( w10905 & w10906 ) | ( w10905 & ~w10914 ) | ( w10906 & ~w10914 ) ;
  assign w11107 = w11097 ^ w11106 ;
  assign w11108 = w11105 ^ w11107 ;
  assign w11109 = w11054 ^ w11108 ;
  assign w11110 = w11062 ^ w11109 ;
  assign w11111 = ~\pi090 & w5209 ;
  assign w11112 = \pi089 & w5433 ;
  assign w11113 = ( w5209 & ~w11111 ) | ( w5209 & w11112 ) | ( ~w11111 & w11112 ) ;
  assign w11114 = ~\pi091 & w5211 ;
  assign w11115 = w1908 | w11113 ;
  assign w11116 = ( w5212 & w11113 ) | ( w5212 & w11115 ) | ( w11113 & w11115 ) ;
  assign w11117 = ( w5211 & ~w11114 ) | ( w5211 & w11116 ) | ( ~w11114 & w11116 ) ;
  assign w11118 = \pi050 ^ w11117 ;
  assign w11119 = ( w10869 & w10870 ) | ( w10869 & w10918 ) | ( w10870 & w10918 ) ;
  assign w11120 = w11110 ^ w11119 ;
  assign w11121 = w11118 ^ w11120 ;
  assign w11122 = ~\pi093 & w4654 ;
  assign w11123 = \pi092 & w4876 ;
  assign w11124 = ( w4654 & ~w11122 ) | ( w4654 & w11123 ) | ( ~w11122 & w11123 ) ;
  assign w11125 = ~\pi094 & w4656 ;
  assign w11126 = w2274 | w11124 ;
  assign w11127 = ( w4657 & w11124 ) | ( w4657 & w11126 ) | ( w11124 & w11126 ) ;
  assign w11128 = ( w4656 & ~w11125 ) | ( w4656 & w11127 ) | ( ~w11125 & w11127 ) ;
  assign w11129 = \pi047 ^ w11128 ;
  assign w11130 = ( w11053 & w11121 ) | ( w11053 & w11129 ) | ( w11121 & w11129 ) ;
  assign w11131 = w11053 ^ w11121 ;
  assign w11132 = w11129 ^ w11131 ;
  assign w11133 = ~\pi096 & w4141 ;
  assign w11134 = \pi095 & w4334 ;
  assign w11135 = ( w4141 & ~w11133 ) | ( w4141 & w11134 ) | ( ~w11133 & w11134 ) ;
  assign w11136 = ~\pi097 & w4143 ;
  assign w11137 = w2673 | w11135 ;
  assign w11138 = ( w4144 & w11135 ) | ( w4144 & w11137 ) | ( w11135 & w11137 ) ;
  assign w11139 = ( w4143 & ~w11136 ) | ( w4143 & w11138 ) | ( ~w11136 & w11138 ) ;
  assign w11140 = \pi044 ^ w11139 ;
  assign w11141 = w11052 ^ w11132 ;
  assign w11142 = w11140 ^ w11141 ;
  assign w11143 = ~\pi099 & w3635 ;
  assign w11144 = \pi098 & w3817 ;
  assign w11145 = ( w3635 & ~w11143 ) | ( w3635 & w11144 ) | ( ~w11143 & w11144 ) ;
  assign w11146 = ~\pi100 & w3637 ;
  assign w11147 = w3104 | w11145 ;
  assign w11148 = ( w3638 & w11145 ) | ( w3638 & w11147 ) | ( w11145 & w11147 ) ;
  assign w11149 = ( w3637 & ~w11146 ) | ( w3637 & w11148 ) | ( ~w11146 & w11148 ) ;
  assign w11150 = \pi041 ^ w11149 ;
  assign w11151 = w11051 ^ w11142 ;
  assign w11152 = w11150 ^ w11151 ;
  assign w11153 = ~\pi102 & w3178 ;
  assign w11154 = \pi101 & w3340 ;
  assign w11155 = ( w3178 & ~w11153 ) | ( w3178 & w11154 ) | ( ~w11153 & w11154 ) ;
  assign w11156 = ~\pi103 & w3180 ;
  assign w11157 = w3437 | w11155 ;
  assign w11158 = ( w3181 & w11155 ) | ( w3181 & w11157 ) | ( w11155 & w11157 ) ;
  assign w11159 = ( w3180 & ~w11156 ) | ( w3180 & w11158 ) | ( ~w11156 & w11158 ) ;
  assign w11160 = \pi038 ^ w11159 ;
  assign w11161 = w11050 ^ w11152 ;
  assign w11162 = w11160 ^ w11161 ;
  assign w11163 = ~\pi105 & w2712 ;
  assign w11164 = \pi104 & w2872 ;
  assign w11165 = ( w2712 & ~w11163 ) | ( w2712 & w11164 ) | ( ~w11163 & w11164 ) ;
  assign w11166 = ~\pi106 & w2714 ;
  assign w11167 = w4068 | w11165 ;
  assign w11168 = ( w2715 & w11165 ) | ( w2715 & w11167 ) | ( w11165 & w11167 ) ;
  assign w11169 = ( w2714 & ~w11166 ) | ( w2714 & w11168 ) | ( ~w11166 & w11168 ) ;
  assign w11170 = \pi035 ^ w11169 ;
  assign w11171 = w11049 ^ w11162 ;
  assign w11172 = w11170 ^ w11171 ;
  assign w11173 = w4425 | w10843 ;
  assign w11174 = ( w2313 & w10843 ) | ( w2313 & w11173 ) | ( w10843 & w11173 ) ;
  assign w11175 = \pi032 ^ w11174 ;
  assign w11176 = ( w10838 & w10957 ) | ( w10838 & w11175 ) | ( w10957 & w11175 ) ;
  assign w11177 = ~\pi108 & w2310 ;
  assign w11178 = \pi107 & w2443 ;
  assign w11179 = ( w2310 & ~w11177 ) | ( w2310 & w11178 ) | ( ~w11177 & w11178 ) ;
  assign w11180 = ~\pi109 & w2312 ;
  assign w11181 = w4599 | w11179 ;
  assign w11182 = ( w2313 & w11179 ) | ( w2313 & w11181 ) | ( w11179 & w11181 ) ;
  assign w11183 = ( w2312 & ~w11180 ) | ( w2312 & w11182 ) | ( ~w11180 & w11182 ) ;
  assign w11184 = \pi032 ^ w11183 ;
  assign w11185 = w11176 ^ w11184 ;
  assign w11186 = w11048 ^ w11172 ;
  assign w11187 = w11040 ^ w11186 ;
  assign w11188 = w11185 ^ w11187 ;
  assign w11189 = w11028 ^ w11188 ;
  assign w11190 = w11020 ^ w11189 ;
  assign w11191 = w11039 ^ w11190 ;
  assign w11192 = w11006 ^ w11191 ;
  assign w11193 = w10998 ^ w11192 ;
  assign w11194 = w11016 ^ w11193 ;
  assign w11195 = w10989 ^ w11194 ;
  assign w11196 = w10997 ^ w11195 ;
  assign w11197 = w10986 ^ w10987 ;
  assign w11198 = w11196 ^ w11197 ;
  assign w11199 = ( w10986 & w10987 ) | ( w10986 & w11196 ) | ( w10987 & w11196 ) ;
  assign w11200 = ( w10989 & w10997 ) | ( w10989 & w11194 ) | ( w10997 & w11194 ) ;
  assign w11201 = ~\pi124 & w837 ;
  assign w11202 = \pi123 & w902 ;
  assign w11203 = ( w837 & ~w11201 ) | ( w837 & w11202 ) | ( ~w11201 & w11202 ) ;
  assign w11204 = ~\pi125 & w839 ;
  assign w11205 = w7988 | w11203 ;
  assign w11206 = ( w840 & w11203 ) | ( w840 & w11205 ) | ( w11203 & w11205 ) ;
  assign w11207 = ( w839 & ~w11204 ) | ( w839 & w11206 ) | ( ~w11204 & w11206 ) ;
  assign w11208 = \pi017 ^ w11207 ;
  assign w11209 = ( w11014 & w11015 ) | ( w11014 & w11191 ) | ( w11015 & w11191 ) ;
  assign w11210 = ~\pi118 & w1313 ;
  assign w11211 = \pi117 & w1417 ;
  assign w11212 = ( w1313 & ~w11210 ) | ( w1313 & w11211 ) | ( ~w11210 & w11211 ) ;
  assign w11213 = ~\pi119 & w1315 ;
  assign w11214 = w6616 | w11212 ;
  assign w11215 = ( w1316 & w11212 ) | ( w1316 & w11214 ) | ( w11212 & w11214 ) ;
  assign w11216 = ( w1315 & ~w11213 ) | ( w1315 & w11215 ) | ( ~w11213 & w11215 ) ;
  assign w11217 = \pi023 ^ w11216 ;
  assign w11218 = ( w11036 & w11038 ) | ( w11036 & w11188 ) | ( w11038 & w11188 ) ;
  assign w11219 = ~\pi112 & w1944 ;
  assign w11220 = \pi111 & w2072 ;
  assign w11221 = ( w1944 & ~w11219 ) | ( w1944 & w11220 ) | ( ~w11219 & w11220 ) ;
  assign w11222 = ~\pi113 & w1946 ;
  assign w11223 = w5366 | w11221 ;
  assign w11224 = ( w1947 & w11221 ) | ( w1947 & w11223 ) | ( w11221 & w11223 ) ;
  assign w11225 = ( w1946 & ~w11222 ) | ( w1946 & w11224 ) | ( ~w11222 & w11224 ) ;
  assign w11226 = \pi029 ^ w11225 ;
  assign w11227 = ( w11172 & w11176 ) | ( w11172 & w11184 ) | ( w11176 & w11184 ) ;
  assign w11228 = ~\pi106 & w2712 ;
  assign w11229 = \pi105 & w2872 ;
  assign w11230 = ( w2712 & ~w11228 ) | ( w2712 & w11229 ) | ( ~w11228 & w11229 ) ;
  assign w11231 = ~\pi107 & w2714 ;
  assign w11232 = w4087 | w11230 ;
  assign w11233 = ( w2715 & w11230 ) | ( w2715 & w11232 ) | ( w11230 & w11232 ) ;
  assign w11234 = ( w2714 & ~w11231 ) | ( w2714 & w11233 ) | ( ~w11231 & w11233 ) ;
  assign w11235 = \pi035 ^ w11234 ;
  assign w11236 = ( w11050 & w11152 ) | ( w11050 & w11160 ) | ( w11152 & w11160 ) ;
  assign w11237 = ~\pi103 & w3178 ;
  assign w11238 = \pi102 & w3340 ;
  assign w11239 = ( w3178 & ~w11237 ) | ( w3178 & w11238 ) | ( ~w11237 & w11238 ) ;
  assign w11240 = ~\pi104 & w3180 ;
  assign w11241 = w3740 | w11239 ;
  assign w11242 = ( w3181 & w11239 ) | ( w3181 & w11241 ) | ( w11239 & w11241 ) ;
  assign w11243 = ( w3180 & ~w11240 ) | ( w3180 & w11242 ) | ( ~w11240 & w11242 ) ;
  assign w11244 = \pi038 ^ w11243 ;
  assign w11245 = ( w11051 & w11142 ) | ( w11051 & w11150 ) | ( w11142 & w11150 ) ;
  assign w11246 = ~\pi100 & w3635 ;
  assign w11247 = \pi099 & w3817 ;
  assign w11248 = ( w3635 & ~w11246 ) | ( w3635 & w11247 ) | ( ~w11246 & w11247 ) ;
  assign w11249 = ~\pi101 & w3637 ;
  assign w11250 = w3264 | w11248 ;
  assign w11251 = ( w3638 & w11248 ) | ( w3638 & w11250 ) | ( w11248 & w11250 ) ;
  assign w11252 = ( w3637 & ~w11249 ) | ( w3637 & w11251 ) | ( ~w11249 & w11251 ) ;
  assign w11253 = \pi041 ^ w11252 ;
  assign w11254 = ( w11052 & w11132 ) | ( w11052 & w11140 ) | ( w11132 & w11140 ) ;
  assign w11255 = ~\pi097 & w4141 ;
  assign w11256 = \pi096 & w4334 ;
  assign w11257 = ( w4141 & ~w11255 ) | ( w4141 & w11256 ) | ( ~w11255 & w11256 ) ;
  assign w11258 = ~\pi098 & w4143 ;
  assign w11259 = w2824 | w11257 ;
  assign w11260 = ( w4144 & w11257 ) | ( w4144 & w11259 ) | ( w11257 & w11259 ) ;
  assign w11261 = ( w4143 & ~w11258 ) | ( w4143 & w11260 ) | ( ~w11258 & w11260 ) ;
  assign w11262 = \pi044 ^ w11261 ;
  assign w11263 = ~\pi094 & w4654 ;
  assign w11264 = \pi093 & w4876 ;
  assign w11265 = ( w4654 & ~w11263 ) | ( w4654 & w11264 ) | ( ~w11263 & w11264 ) ;
  assign w11266 = ~\pi095 & w4656 ;
  assign w11267 = w2409 | w11265 ;
  assign w11268 = ( w4657 & w11265 ) | ( w4657 & w11267 ) | ( w11265 & w11267 ) ;
  assign w11269 = ( w4656 & ~w11266 ) | ( w4656 & w11268 ) | ( ~w11266 & w11268 ) ;
  assign w11270 = \pi047 ^ w11269 ;
  assign w11271 = ( w11110 & w11118 ) | ( w11110 & w11119 ) | ( w11118 & w11119 ) ;
  assign w11272 = ( \pi062 & \pi063 ) | ( \pi062 & \pi077 ) | ( \pi063 & \pi077 ) ;
  assign w11273 = \pi063 & ~\pi076 ;
  assign w11274 = w11272 & ~w11273 ;
  assign w11275 = ( ~\pi062 & w11272 ) | ( ~\pi062 & w11274 ) | ( w11272 & w11274 ) ;
  assign w11276 = \pi063 & \pi075 ;
  assign w11277 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w11276 ) | ( \pi063 & w11276 ) ;
  assign w11278 = ( \pi062 & ~\pi063 ) | ( \pi062 & w11276 ) | ( ~\pi063 & w11276 ) ;
  assign w11279 = ( \pi076 & w11277 ) | ( \pi076 & w11278 ) | ( w11277 & w11278 ) ;
  assign w11280 = ( ~\pi011 & w10654 ) | ( ~\pi011 & w11279 ) | ( w10654 & w11279 ) ;
  assign w11281 = ~\pi079 & w7811 ;
  assign w11282 = \pi078 & w8046 ;
  assign w11283 = ( w7811 & ~w11281 ) | ( w7811 & w11282 ) | ( ~w11281 & w11282 ) ;
  assign w11284 = ~\pi080 & w7813 ;
  assign w11285 = w794 | w11283 ;
  assign w11286 = ( w7814 & w11283 ) | ( w7814 & w11285 ) | ( w11283 & w11285 ) ;
  assign w11287 = ( w7813 & ~w11284 ) | ( w7813 & w11286 ) | ( ~w11284 & w11286 ) ;
  assign w11288 = \pi062 ^ w11287 ;
  assign w11289 = w11280 ^ w11288 ;
  assign w11290 = w11275 ^ w11289 ;
  assign w11291 = ( w11070 & w11078 ) | ( w11070 & ~w11084 ) | ( w11078 & ~w11084 ) ;
  assign w11292 = ~\pi082 & w7135 ;
  assign w11293 = \pi081 & w7359 ;
  assign w11294 = ( w7135 & ~w11292 ) | ( w7135 & w11293 ) | ( ~w11292 & w11293 ) ;
  assign w11295 = ~\pi083 & w7137 ;
  assign w11296 = w1099 | w11294 ;
  assign w11297 = ( w7138 & w11294 ) | ( w7138 & w11296 ) | ( w11294 & w11296 ) ;
  assign w11298 = ( w7137 & ~w11295 ) | ( w7137 & w11297 ) | ( ~w11295 & w11297 ) ;
  assign w11299 = \pi059 ^ w11298 ;
  assign w11300 = w11290 ^ w11291 ;
  assign w11301 = w11299 ^ w11300 ;
  assign w11302 = ( ~w11086 & w11094 ) | ( ~w11086 & w11095 ) | ( w11094 & w11095 ) ;
  assign w11303 = ~\pi085 & w6466 ;
  assign w11304 = \pi084 & w6702 ;
  assign w11305 = ( w6466 & ~w11303 ) | ( w6466 & w11304 ) | ( ~w11303 & w11304 ) ;
  assign w11306 = ~\pi086 & w6468 ;
  assign w11307 = w1379 | w11305 ;
  assign w11308 = ( w6469 & w11305 ) | ( w6469 & w11307 ) | ( w11305 & w11307 ) ;
  assign w11309 = ( w6468 & ~w11306 ) | ( w6468 & w11308 ) | ( ~w11306 & w11308 ) ;
  assign w11310 = \pi056 ^ w11309 ;
  assign w11311 = w11301 ^ w11302 ;
  assign w11312 = w11310 ^ w11311 ;
  assign w11313 = ( w11097 & ~w11105 ) | ( w11097 & w11106 ) | ( ~w11105 & w11106 ) ;
  assign w11314 = ~\pi088 & w5802 ;
  assign w11315 = \pi087 & w6052 ;
  assign w11316 = ( w5802 & ~w11314 ) | ( w5802 & w11315 ) | ( ~w11314 & w11315 ) ;
  assign w11317 = ~\pi089 & w5804 ;
  assign w11318 = w1595 | w11316 ;
  assign w11319 = ( w5805 & w11316 ) | ( w5805 & w11318 ) | ( w11316 & w11318 ) ;
  assign w11320 = ( w5804 & ~w11317 ) | ( w5804 & w11319 ) | ( ~w11317 & w11319 ) ;
  assign w11321 = \pi053 ^ w11320 ;
  assign w11322 = w11312 ^ w11313 ;
  assign w11323 = w11321 ^ w11322 ;
  assign w11324 = ( w11054 & w11062 ) | ( w11054 & w11108 ) | ( w11062 & w11108 ) ;
  assign w11325 = ~\pi091 & w5209 ;
  assign w11326 = \pi090 & w5433 ;
  assign w11327 = ( w5209 & ~w11325 ) | ( w5209 & w11326 ) | ( ~w11325 & w11326 ) ;
  assign w11328 = ~\pi092 & w5211 ;
  assign w11329 = w2033 | w11327 ;
  assign w11330 = ( w5212 & w11327 ) | ( w5212 & w11329 ) | ( w11327 & w11329 ) ;
  assign w11331 = ( w5211 & ~w11328 ) | ( w5211 & w11330 ) | ( ~w11328 & w11330 ) ;
  assign w11332 = \pi050 ^ w11331 ;
  assign w11333 = w11323 ^ w11324 ;
  assign w11334 = w11332 ^ w11333 ;
  assign w11335 = w11271 ^ w11334 ;
  assign w11336 = w11270 ^ w11335 ;
  assign w11337 = w11130 ^ w11336 ;
  assign w11338 = w11262 ^ w11337 ;
  assign w11339 = w11254 ^ w11338 ;
  assign w11340 = w11253 ^ w11339 ;
  assign w11341 = w11245 ^ w11340 ;
  assign w11342 = w11244 ^ w11341 ;
  assign w11343 = w11236 ^ w11342 ;
  assign w11344 = w11235 ^ w11343 ;
  assign w11345 = ( w11049 & w11162 ) | ( w11049 & w11170 ) | ( w11162 & w11170 ) ;
  assign w11346 = \pi108 & w2443 ;
  assign w11347 = ( \pi110 & w2312 ) | ( \pi110 & w11346 ) | ( w2312 & w11346 ) ;
  assign w11348 = \pi109 | w11347 ;
  assign w11349 = ( w2310 & w11347 ) | ( w2310 & w11348 ) | ( w11347 & w11348 ) ;
  assign w11350 = w11346 | w11349 ;
  assign w11351 = w2313 & ~w4792 ;
  assign w11352 = ( w2313 & w11350 ) | ( w2313 & ~w11351 ) | ( w11350 & ~w11351 ) ;
  assign w11353 = w11345 ^ w11352 ;
  assign w11354 = \pi032 ^ w11344 ;
  assign w11355 = w11353 ^ w11354 ;
  assign w11356 = w11227 ^ w11355 ;
  assign w11357 = w11226 ^ w11356 ;
  assign w11358 = w11172 ^ w11185 ;
  assign w11359 = ( w11040 & w11048 ) | ( w11040 & w11358 ) | ( w11048 & w11358 ) ;
  assign w11360 = \pi114 & w1722 ;
  assign w11361 = ( \pi116 & w1631 ) | ( \pi116 & w11360 ) | ( w1631 & w11360 ) ;
  assign w11362 = \pi115 | w11361 ;
  assign w11363 = ( w1629 & w11361 ) | ( w1629 & w11362 ) | ( w11361 & w11362 ) ;
  assign w11364 = w11360 | w11363 ;
  assign w11365 = w1632 & ~w5976 ;
  assign w11366 = ( w1632 & w11364 ) | ( w1632 & ~w11365 ) | ( w11364 & ~w11365 ) ;
  assign w11367 = w11359 ^ w11366 ;
  assign w11368 = \pi026 ^ w11357 ;
  assign w11369 = w11367 ^ w11368 ;
  assign w11370 = w11218 ^ w11369 ;
  assign w11371 = w11217 ^ w11370 ;
  assign w11372 = w11039 ^ w11188 ;
  assign w11373 = ( w11020 & w11028 ) | ( w11020 & w11372 ) | ( w11028 & w11372 ) ;
  assign w11374 = \pi120 & w1138 ;
  assign w11375 = ( \pi122 & w1046 ) | ( \pi122 & w11374 ) | ( w1046 & w11374 ) ;
  assign w11376 = \pi121 | w11375 ;
  assign w11377 = ( w1044 & w11375 ) | ( w1044 & w11376 ) | ( w11375 & w11376 ) ;
  assign w11378 = w11374 | w11377 ;
  assign w11379 = w1047 & ~w7069 ;
  assign w11380 = ( w1047 & w11378 ) | ( w1047 & ~w11379 ) | ( w11378 & ~w11379 ) ;
  assign w11381 = w11373 ^ w11380 ;
  assign w11382 = \pi020 ^ w11371 ;
  assign w11383 = w11381 ^ w11382 ;
  assign w11384 = w11209 ^ w11383 ;
  assign w11385 = w11208 ^ w11384 ;
  assign w11386 = w11016 ^ w11191 ;
  assign w11387 = ( w10998 & w11006 ) | ( w10998 & w11386 ) | ( w11006 & w11386 ) ;
  assign w11388 = \pi127 & w601 ;
  assign w11389 = ( \pi126 & ~w604 ) | ( \pi126 & w8490 ) | ( ~w604 & w8490 ) ;
  assign w11390 = \pi126 & ~w683 ;
  assign w11391 = ( ~\pi126 & w11389 ) | ( ~\pi126 & w11390 ) | ( w11389 & w11390 ) ;
  assign w11392 = ( w9420 & w11388 ) | ( w9420 & ~w11391 ) | ( w11388 & ~w11391 ) ;
  assign w11393 = \pi014 ^ w11392 ;
  assign w11394 = w11387 ^ w11393 ;
  assign w11395 = w11385 ^ w11394 ;
  assign w11396 = w11199 ^ w11200 ;
  assign w11397 = w11395 ^ w11396 ;
  assign w11398 = ( w11199 & w11200 ) | ( w11199 & w11395 ) | ( w11200 & w11395 ) ;
  assign w11399 = ( w11385 & w11387 ) | ( w11385 & w11393 ) | ( w11387 & w11393 ) ;
  assign w11400 = ( w11208 & w11209 ) | ( w11208 & w11383 ) | ( w11209 & w11383 ) ;
  assign w11401 = w604 & w8481 ;
  assign w11402 = w683 | w11401 ;
  assign w11403 = ( \pi127 & w11401 ) | ( \pi127 & w11402 ) | ( w11401 & w11402 ) ;
  assign w11404 = \pi014 ^ w11403 ;
  assign w11405 = ~\pi122 & w1044 ;
  assign w11406 = \pi121 & w1138 ;
  assign w11407 = ( w1044 & ~w11405 ) | ( w1044 & w11406 ) | ( ~w11405 & w11406 ) ;
  assign w11408 = ~\pi123 & w1046 ;
  assign w11409 = w7516 | w11407 ;
  assign w11410 = ( w1047 & w11407 ) | ( w1047 & w11409 ) | ( w11407 & w11409 ) ;
  assign w11411 = ( w1046 & ~w11408 ) | ( w1046 & w11410 ) | ( ~w11408 & w11410 ) ;
  assign w11412 = \pi020 ^ w11411 ;
  assign w11413 = ( w11217 & w11218 ) | ( w11217 & w11369 ) | ( w11218 & w11369 ) ;
  assign w11414 = ~\pi119 & w1313 ;
  assign w11415 = \pi118 & w1417 ;
  assign w11416 = ( w1313 & ~w11414 ) | ( w1313 & w11415 ) | ( ~w11414 & w11415 ) ;
  assign w11417 = ~\pi120 & w1315 ;
  assign w11418 = w6634 | w11416 ;
  assign w11419 = ( w1316 & w11416 ) | ( w1316 & w11418 ) | ( w11416 & w11418 ) ;
  assign w11420 = ( w1315 & ~w11417 ) | ( w1315 & w11419 ) | ( ~w11417 & w11419 ) ;
  assign w11421 = \pi023 ^ w11420 ;
  assign w11422 = w5976 | w11364 ;
  assign w11423 = ( w1632 & w11364 ) | ( w1632 & w11422 ) | ( w11364 & w11422 ) ;
  assign w11424 = \pi026 ^ w11423 ;
  assign w11425 = ( w11357 & w11359 ) | ( w11357 & w11424 ) | ( w11359 & w11424 ) ;
  assign w11426 = w11421 ^ w11425 ;
  assign w11427 = ~\pi116 & w1629 ;
  assign w11428 = \pi115 & w1722 ;
  assign w11429 = ( w1629 & ~w11427 ) | ( w1629 & w11428 ) | ( ~w11427 & w11428 ) ;
  assign w11430 = ~\pi117 & w1631 ;
  assign w11431 = w6185 | w11429 ;
  assign w11432 = ( w1632 & w11429 ) | ( w1632 & w11431 ) | ( w11429 & w11431 ) ;
  assign w11433 = ( w1631 & ~w11430 ) | ( w1631 & w11432 ) | ( ~w11430 & w11432 ) ;
  assign w11434 = \pi026 ^ w11433 ;
  assign w11435 = ( w11226 & w11227 ) | ( w11226 & w11355 ) | ( w11227 & w11355 ) ;
  assign w11436 = ( w11235 & w11236 ) | ( w11235 & w11342 ) | ( w11236 & w11342 ) ;
  assign w11437 = \pi109 & w2443 ;
  assign w11438 = ( \pi111 & w2312 ) | ( \pi111 & w11437 ) | ( w2312 & w11437 ) ;
  assign w11439 = \pi110 | w11438 ;
  assign w11440 = ( w2310 & w11438 ) | ( w2310 & w11439 ) | ( w11438 & w11439 ) ;
  assign w11441 = w11437 | w11440 ;
  assign w11442 = ~\pi107 & w2712 ;
  assign w11443 = \pi106 & w2872 ;
  assign w11444 = ( w2712 & ~w11442 ) | ( w2712 & w11443 ) | ( ~w11442 & w11443 ) ;
  assign w11445 = ~\pi108 & w2714 ;
  assign w11446 = w4425 | w11444 ;
  assign w11447 = ( w2715 & w11444 ) | ( w2715 & w11446 ) | ( w11444 & w11446 ) ;
  assign w11448 = ( w2714 & ~w11445 ) | ( w2714 & w11447 ) | ( ~w11445 & w11447 ) ;
  assign w11449 = \pi035 ^ w11448 ;
  assign w11450 = ( w11244 & w11245 ) | ( w11244 & w11340 ) | ( w11245 & w11340 ) ;
  assign w11451 = ~\pi104 & w3178 ;
  assign w11452 = \pi103 & w3340 ;
  assign w11453 = ( w3178 & ~w11451 ) | ( w3178 & w11452 ) | ( ~w11451 & w11452 ) ;
  assign w11454 = ~\pi105 & w3180 ;
  assign w11455 = w3905 | w11453 ;
  assign w11456 = ( w3181 & w11453 ) | ( w3181 & w11455 ) | ( w11453 & w11455 ) ;
  assign w11457 = ( w3180 & ~w11454 ) | ( w3180 & w11456 ) | ( ~w11454 & w11456 ) ;
  assign w11458 = \pi038 ^ w11457 ;
  assign w11459 = ( w11253 & w11254 ) | ( w11253 & w11338 ) | ( w11254 & w11338 ) ;
  assign w11460 = ( w11270 & w11271 ) | ( w11270 & w11334 ) | ( w11271 & w11334 ) ;
  assign w11461 = ( w11312 & w11313 ) | ( w11312 & ~w11321 ) | ( w11313 & ~w11321 ) ;
  assign w11462 = ~\pi089 & w5802 ;
  assign w11463 = \pi088 & w6052 ;
  assign w11464 = ( w5802 & ~w11462 ) | ( w5802 & w11463 ) | ( ~w11462 & w11463 ) ;
  assign w11465 = ~\pi090 & w5804 ;
  assign w11466 = w1801 | w11464 ;
  assign w11467 = ( w5805 & w11464 ) | ( w5805 & w11466 ) | ( w11464 & w11466 ) ;
  assign w11468 = ( w5804 & ~w11465 ) | ( w5804 & w11467 ) | ( ~w11465 & w11467 ) ;
  assign w11469 = \pi053 ^ w11468 ;
  assign w11470 = ( ~w11301 & w11302 ) | ( ~w11301 & w11310 ) | ( w11302 & w11310 ) ;
  assign w11471 = ( ~w11275 & w11280 ) | ( ~w11275 & w11288 ) | ( w11280 & w11288 ) ;
  assign w11472 = ~\pi080 & w7811 ;
  assign w11473 = \pi079 & w8046 ;
  assign w11474 = ( w7811 & ~w11472 ) | ( w7811 & w11473 ) | ( ~w11472 & w11473 ) ;
  assign w11475 = ~\pi081 & w7813 ;
  assign w11476 = ~w874 & w7814 ;
  assign w11477 = ( w7814 & w11474 ) | ( w7814 & ~w11476 ) | ( w11474 & ~w11476 ) ;
  assign w11478 = ( w7813 & ~w11475 ) | ( w7813 & w11477 ) | ( ~w11475 & w11477 ) ;
  assign w11479 = ~\pi063 & \pi077 ;
  assign w11480 = ( \pi062 & ~w11273 ) | ( \pi062 & w11479 ) | ( ~w11273 & w11479 ) ;
  assign w11481 = w11478 ^ w11480 ;
  assign w11482 = \pi077 ^ w11481 ;
  assign w11483 = ( \pi063 & w11478 ) | ( \pi063 & ~w11479 ) | ( w11478 & ~w11479 ) ;
  assign w11484 = ( \pi062 & ~\pi063 ) | ( \pi062 & w11483 ) | ( ~\pi063 & w11483 ) ;
  assign w11485 = ( \pi062 & ~w11482 ) | ( \pi062 & w11484 ) | ( ~w11482 & w11484 ) ;
  assign w11486 = ( \pi063 & \pi078 ) | ( \pi063 & w11485 ) | ( \pi078 & w11485 ) ;
  assign w11487 = w11482 ^ w11486 ;
  assign w11488 = ~\pi083 & w7135 ;
  assign w11489 = \pi082 & w7359 ;
  assign w11490 = ( w7135 & ~w11488 ) | ( w7135 & w11489 ) | ( ~w11488 & w11489 ) ;
  assign w11491 = ~\pi084 & w7137 ;
  assign w11492 = w1188 | w11490 ;
  assign w11493 = ( w7138 & w11490 ) | ( w7138 & w11492 ) | ( w11490 & w11492 ) ;
  assign w11494 = ( w7137 & ~w11491 ) | ( w7137 & w11493 ) | ( ~w11491 & w11493 ) ;
  assign w11495 = \pi059 ^ w11494 ;
  assign w11496 = w11471 ^ w11487 ;
  assign w11497 = w11495 ^ w11496 ;
  assign w11498 = ( ~w11290 & w11291 ) | ( ~w11290 & w11299 ) | ( w11291 & w11299 ) ;
  assign w11499 = ~\pi086 & w6466 ;
  assign w11500 = \pi085 & w6702 ;
  assign w11501 = ( w6466 & ~w11499 ) | ( w6466 & w11500 ) | ( ~w11499 & w11500 ) ;
  assign w11502 = ~\pi087 & w6468 ;
  assign w11503 = w1477 | w11501 ;
  assign w11504 = ( w6469 & w11501 ) | ( w6469 & w11503 ) | ( w11501 & w11503 ) ;
  assign w11505 = ( w6468 & ~w11502 ) | ( w6468 & w11504 ) | ( ~w11502 & w11504 ) ;
  assign w11506 = \pi056 ^ w11505 ;
  assign w11507 = w11497 ^ w11498 ;
  assign w11508 = w11506 ^ w11507 ;
  assign w11509 = w11470 ^ w11508 ;
  assign w11510 = w11469 ^ w11509 ;
  assign w11511 = ~\pi092 & w5209 ;
  assign w11512 = \pi091 & w5433 ;
  assign w11513 = ( w5209 & ~w11511 ) | ( w5209 & w11512 ) | ( ~w11511 & w11512 ) ;
  assign w11514 = ~\pi093 & w5211 ;
  assign w11515 = w2155 | w11513 ;
  assign w11516 = ( w5212 & w11513 ) | ( w5212 & w11515 ) | ( w11513 & w11515 ) ;
  assign w11517 = ( w5211 & ~w11514 ) | ( w5211 & w11516 ) | ( ~w11514 & w11516 ) ;
  assign w11518 = \pi050 ^ w11517 ;
  assign w11519 = w11461 ^ w11510 ;
  assign w11520 = w11518 ^ w11519 ;
  assign w11521 = ( w11323 & w11324 ) | ( w11323 & w11332 ) | ( w11324 & w11332 ) ;
  assign w11522 = ~\pi095 & w4654 ;
  assign w11523 = \pi094 & w4876 ;
  assign w11524 = ( w4654 & ~w11522 ) | ( w4654 & w11523 ) | ( ~w11522 & w11523 ) ;
  assign w11525 = ~\pi096 & w4656 ;
  assign w11526 = w2546 | w11524 ;
  assign w11527 = ( w4657 & w11524 ) | ( w4657 & w11526 ) | ( w11524 & w11526 ) ;
  assign w11528 = ( w4656 & ~w11525 ) | ( w4656 & w11527 ) | ( ~w11525 & w11527 ) ;
  assign w11529 = \pi047 ^ w11528 ;
  assign w11530 = w11520 ^ w11521 ;
  assign w11531 = w11529 ^ w11530 ;
  assign w11532 = ~\pi098 & w4141 ;
  assign w11533 = \pi097 & w4334 ;
  assign w11534 = ( w4141 & ~w11532 ) | ( w4141 & w11533 ) | ( ~w11532 & w11533 ) ;
  assign w11535 = ~\pi099 & w4143 ;
  assign w11536 = w2966 | w11534 ;
  assign w11537 = ( w4144 & w11534 ) | ( w4144 & w11536 ) | ( w11534 & w11536 ) ;
  assign w11538 = ( w4143 & ~w11535 ) | ( w4143 & w11537 ) | ( ~w11535 & w11537 ) ;
  assign w11539 = \pi044 ^ w11538 ;
  assign w11540 = w11460 ^ w11531 ;
  assign w11541 = w11539 ^ w11540 ;
  assign w11542 = ( w11130 & w11262 ) | ( w11130 & w11336 ) | ( w11262 & w11336 ) ;
  assign w11543 = ~\pi101 & w3635 ;
  assign w11544 = \pi100 & w3817 ;
  assign w11545 = ( w3635 & ~w11543 ) | ( w3635 & w11544 ) | ( ~w11543 & w11544 ) ;
  assign w11546 = ~\pi102 & w3637 ;
  assign w11547 = w3284 | w11545 ;
  assign w11548 = ( w3638 & w11545 ) | ( w3638 & w11547 ) | ( w11545 & w11547 ) ;
  assign w11549 = ( w3637 & ~w11546 ) | ( w3637 & w11548 ) | ( ~w11546 & w11548 ) ;
  assign w11550 = \pi041 ^ w11549 ;
  assign w11551 = w11541 ^ w11542 ;
  assign w11552 = w11550 ^ w11551 ;
  assign w11553 = w11459 ^ w11552 ;
  assign w11554 = w11458 ^ w11553 ;
  assign w11555 = w11450 ^ w11554 ;
  assign w11556 = w11449 ^ w11555 ;
  assign w11557 = w2313 & ~w4811 ;
  assign w11558 = ( w2313 & w11441 ) | ( w2313 & ~w11557 ) | ( w11441 & ~w11557 ) ;
  assign w11559 = w11436 ^ w11558 ;
  assign w11560 = \pi032 ^ w11556 ;
  assign w11561 = w11559 ^ w11560 ;
  assign w11562 = w4792 | w11350 ;
  assign w11563 = ( w2313 & w11350 ) | ( w2313 & w11562 ) | ( w11350 & w11562 ) ;
  assign w11564 = \pi032 ^ w11563 ;
  assign w11565 = ( w11344 & w11345 ) | ( w11344 & w11564 ) | ( w11345 & w11564 ) ;
  assign w11566 = \pi112 & w2072 ;
  assign w11567 = ( \pi114 & w1946 ) | ( \pi114 & w11566 ) | ( w1946 & w11566 ) ;
  assign w11568 = \pi113 | w11567 ;
  assign w11569 = ( w1944 & w11567 ) | ( w1944 & w11568 ) | ( w11567 & w11568 ) ;
  assign w11570 = w11566 | w11569 ;
  assign w11571 = w1947 & ~w5565 ;
  assign w11572 = ( w1947 & w11570 ) | ( w1947 & ~w11571 ) | ( w11570 & ~w11571 ) ;
  assign w11573 = w11565 ^ w11572 ;
  assign w11574 = \pi029 ^ w11561 ;
  assign w11575 = w11573 ^ w11574 ;
  assign w11576 = w11435 ^ w11575 ;
  assign w11577 = w11434 ^ w11576 ;
  assign w11578 = w11412 ^ w11577 ;
  assign w11579 = w11413 ^ w11578 ;
  assign w11580 = w11426 ^ w11579 ;
  assign w11581 = w7069 | w11378 ;
  assign w11582 = ( w1047 & w11378 ) | ( w1047 & w11581 ) | ( w11378 & w11581 ) ;
  assign w11583 = \pi020 ^ w11582 ;
  assign w11584 = ( w11371 & w11373 ) | ( w11371 & w11583 ) | ( w11373 & w11583 ) ;
  assign w11585 = \pi124 & w902 ;
  assign w11586 = ( \pi126 & w839 ) | ( \pi126 & w11585 ) | ( w839 & w11585 ) ;
  assign w11587 = \pi125 | w11586 ;
  assign w11588 = ( w837 & w11586 ) | ( w837 & w11587 ) | ( w11586 & w11587 ) ;
  assign w11589 = w11585 | w11588 ;
  assign w11590 = w840 & ~w8231 ;
  assign w11591 = ( w840 & w11589 ) | ( w840 & ~w11590 ) | ( w11589 & ~w11590 ) ;
  assign w11592 = w11584 ^ w11591 ;
  assign w11593 = \pi017 ^ w11580 ;
  assign w11594 = w11592 ^ w11593 ;
  assign w11595 = w11400 ^ w11594 ;
  assign w11596 = w11404 ^ w11595 ;
  assign w11597 = w11398 ^ w11399 ;
  assign w11598 = w11596 ^ w11597 ;
  assign w11599 = w8231 | w11589 ;
  assign w11600 = ( w840 & w11589 ) | ( w840 & w11599 ) | ( w11589 & w11599 ) ;
  assign w11601 = \pi017 ^ w11600 ;
  assign w11602 = ( w11580 & w11584 ) | ( w11580 & w11601 ) | ( w11584 & w11601 ) ;
  assign w11603 = ~\pi126 & w837 ;
  assign w11604 = \pi125 & w902 ;
  assign w11605 = ( w837 & ~w11603 ) | ( w837 & w11604 ) | ( ~w11603 & w11604 ) ;
  assign w11606 = ~\pi127 & w839 ;
  assign w11607 = w8466 | w11605 ;
  assign w11608 = ( w840 & w11605 ) | ( w840 & w11607 ) | ( w11605 & w11607 ) ;
  assign w11609 = ( w839 & ~w11606 ) | ( w839 & w11608 ) | ( ~w11606 & w11608 ) ;
  assign w11610 = \pi017 ^ w11609 ;
  assign w11611 = ~\pi123 & w1044 ;
  assign w11612 = \pi122 & w1138 ;
  assign w11613 = ( w1044 & ~w11611 ) | ( w1044 & w11612 ) | ( ~w11611 & w11612 ) ;
  assign w11614 = ~\pi124 & w1046 ;
  assign w11615 = w7538 | w11613 ;
  assign w11616 = ( w1047 & w11613 ) | ( w1047 & w11615 ) | ( w11613 & w11615 ) ;
  assign w11617 = ( w1046 & ~w11614 ) | ( w1046 & w11616 ) | ( ~w11614 & w11616 ) ;
  assign w11618 = \pi020 ^ w11617 ;
  assign w11619 = w11426 ^ w11577 ;
  assign w11620 = ( w11412 & w11413 ) | ( w11412 & w11619 ) | ( w11413 & w11619 ) ;
  assign w11621 = w11618 ^ w11620 ;
  assign w11622 = ( w11421 & w11425 ) | ( w11421 & w11577 ) | ( w11425 & w11577 ) ;
  assign w11623 = ~\pi120 & w1313 ;
  assign w11624 = \pi119 & w1417 ;
  assign w11625 = ( w1313 & ~w11623 ) | ( w1313 & w11624 ) | ( ~w11623 & w11624 ) ;
  assign w11626 = ~\pi121 & w1315 ;
  assign w11627 = w7050 | w11625 ;
  assign w11628 = ( w1316 & w11625 ) | ( w1316 & w11627 ) | ( w11625 & w11627 ) ;
  assign w11629 = ( w1315 & ~w11626 ) | ( w1315 & w11628 ) | ( ~w11626 & w11628 ) ;
  assign w11630 = \pi023 ^ w11629 ;
  assign w11631 = ~\pi117 & w1629 ;
  assign w11632 = \pi116 & w1722 ;
  assign w11633 = ( w1629 & ~w11631 ) | ( w1629 & w11632 ) | ( ~w11631 & w11632 ) ;
  assign w11634 = ~\pi118 & w1631 ;
  assign w11635 = w6206 | w11633 ;
  assign w11636 = ( w1632 & w11633 ) | ( w1632 & w11635 ) | ( w11633 & w11635 ) ;
  assign w11637 = ( w1631 & ~w11634 ) | ( w1631 & w11636 ) | ( ~w11634 & w11636 ) ;
  assign w11638 = \pi026 ^ w11637 ;
  assign w11639 = ( w11434 & w11435 ) | ( w11434 & w11575 ) | ( w11435 & w11575 ) ;
  assign w11640 = w11638 ^ w11639 ;
  assign w11641 = ~\pi114 & w1944 ;
  assign w11642 = \pi113 & w2072 ;
  assign w11643 = ( w1944 & ~w11641 ) | ( w1944 & w11642 ) | ( ~w11641 & w11642 ) ;
  assign w11644 = ~\pi115 & w1946 ;
  assign w11645 = w5585 | w11643 ;
  assign w11646 = ( w1947 & w11643 ) | ( w1947 & w11645 ) | ( w11643 & w11645 ) ;
  assign w11647 = ( w1946 & ~w11644 ) | ( w1946 & w11646 ) | ( ~w11644 & w11646 ) ;
  assign w11648 = \pi029 ^ w11647 ;
  assign w11649 = w5565 | w11570 ;
  assign w11650 = ( w1947 & w11570 ) | ( w1947 & w11649 ) | ( w11570 & w11649 ) ;
  assign w11651 = \pi029 ^ w11650 ;
  assign w11652 = ( w11561 & w11565 ) | ( w11561 & w11651 ) | ( w11565 & w11651 ) ;
  assign w11653 = ( w11458 & w11459 ) | ( w11458 & w11552 ) | ( w11459 & w11552 ) ;
  assign w11654 = ( w11541 & w11542 ) | ( w11541 & w11550 ) | ( w11542 & w11550 ) ;
  assign w11655 = ( w11460 & w11531 ) | ( w11460 & w11539 ) | ( w11531 & w11539 ) ;
  assign w11656 = ( w11520 & w11521 ) | ( w11520 & w11529 ) | ( w11521 & w11529 ) ;
  assign w11657 = ( ~w11497 & w11498 ) | ( ~w11497 & w11506 ) | ( w11498 & w11506 ) ;
  assign w11658 = ( \pi062 & \pi063 ) | ( \pi062 & \pi079 ) | ( \pi063 & \pi079 ) ;
  assign w11659 = \pi078 | w8323 ;
  assign w11660 = w11658 & w11659 ;
  assign w11661 = \pi014 ^ w11660 ;
  assign w11662 = ~\pi081 & w7811 ;
  assign w11663 = \pi080 & w8046 ;
  assign w11664 = ( w7811 & ~w11662 ) | ( w7811 & w11663 ) | ( ~w11662 & w11663 ) ;
  assign w11665 = ~\pi082 & w7813 ;
  assign w11666 = w1008 | w11664 ;
  assign w11667 = ( w7814 & w11664 ) | ( w7814 & w11666 ) | ( w11664 & w11666 ) ;
  assign w11668 = ( w7813 & ~w11665 ) | ( w7813 & w11667 ) | ( ~w11665 & w11667 ) ;
  assign w11669 = \pi062 ^ w11668 ;
  assign w11670 = \pi063 ^ w11478 ;
  assign w11671 = ( \pi077 & ~\pi078 ) | ( \pi077 & w11670 ) | ( ~\pi078 & w11670 ) ;
  assign w11672 = w8323 ^ w11671 ;
  assign w11673 = ( \pi076 & \pi077 ) | ( \pi076 & ~w11478 ) | ( \pi077 & ~w11478 ) ;
  assign w11674 = ( \pi077 & w11670 ) | ( \pi077 & ~w11673 ) | ( w11670 & ~w11673 ) ;
  assign w11675 = ( ~w11671 & w11672 ) | ( ~w11671 & w11674 ) | ( w11672 & w11674 ) ;
  assign w11676 = w11275 ^ w11661 ;
  assign w11677 = w11669 ^ w11676 ;
  assign w11678 = w11675 ^ w11677 ;
  assign w11679 = ~\pi084 & w7135 ;
  assign w11680 = \pi083 & w7359 ;
  assign w11681 = ( w7135 & ~w11679 ) | ( w7135 & w11680 ) | ( ~w11679 & w11680 ) ;
  assign w11682 = ~\pi085 & w7137 ;
  assign w11683 = w1274 | w11681 ;
  assign w11684 = ( w7138 & w11681 ) | ( w7138 & w11683 ) | ( w11681 & w11683 ) ;
  assign w11685 = ( w7137 & ~w11682 ) | ( w7137 & w11684 ) | ( ~w11682 & w11684 ) ;
  assign w11686 = \pi059 ^ w11685 ;
  assign w11687 = ( w11471 & ~w11487 ) | ( w11471 & w11495 ) | ( ~w11487 & w11495 ) ;
  assign w11688 = w11678 ^ w11687 ;
  assign w11689 = w11686 ^ w11688 ;
  assign w11690 = ~\pi087 & w6466 ;
  assign w11691 = \pi086 & w6702 ;
  assign w11692 = ( w6466 & ~w11690 ) | ( w6466 & w11691 ) | ( ~w11690 & w11691 ) ;
  assign w11693 = ~\pi088 & w6468 ;
  assign w11694 = w1574 | w11692 ;
  assign w11695 = ( w6469 & w11692 ) | ( w6469 & w11694 ) | ( w11692 & w11694 ) ;
  assign w11696 = ( w6468 & ~w11693 ) | ( w6468 & w11695 ) | ( ~w11693 & w11695 ) ;
  assign w11697 = \pi056 ^ w11696 ;
  assign w11698 = ( w11657 & ~w11689 ) | ( w11657 & w11697 ) | ( ~w11689 & w11697 ) ;
  assign w11699 = w11657 ^ w11689 ;
  assign w11700 = w11697 ^ w11699 ;
  assign w11701 = ~\pi090 & w5802 ;
  assign w11702 = \pi089 & w6052 ;
  assign w11703 = ( w5802 & ~w11701 ) | ( w5802 & w11702 ) | ( ~w11701 & w11702 ) ;
  assign w11704 = ~\pi091 & w5804 ;
  assign w11705 = w1908 | w11703 ;
  assign w11706 = ( w5805 & w11703 ) | ( w5805 & w11705 ) | ( w11703 & w11705 ) ;
  assign w11707 = ( w5804 & ~w11704 ) | ( w5804 & w11706 ) | ( ~w11704 & w11706 ) ;
  assign w11708 = \pi053 ^ w11707 ;
  assign w11709 = ( w11469 & w11470 ) | ( w11469 & ~w11508 ) | ( w11470 & ~w11508 ) ;
  assign w11710 = w11700 ^ w11709 ;
  assign w11711 = w11708 ^ w11710 ;
  assign w11712 = ~\pi093 & w5209 ;
  assign w11713 = \pi092 & w5433 ;
  assign w11714 = ( w5209 & ~w11712 ) | ( w5209 & w11713 ) | ( ~w11712 & w11713 ) ;
  assign w11715 = ~\pi094 & w5211 ;
  assign w11716 = w2274 | w11714 ;
  assign w11717 = ( w5212 & w11714 ) | ( w5212 & w11716 ) | ( w11714 & w11716 ) ;
  assign w11718 = ( w5211 & ~w11715 ) | ( w5211 & w11717 ) | ( ~w11715 & w11717 ) ;
  assign w11719 = \pi050 ^ w11718 ;
  assign w11720 = ( w11461 & w11510 ) | ( w11461 & ~w11518 ) | ( w11510 & ~w11518 ) ;
  assign w11721 = w11711 ^ w11720 ;
  assign w11722 = w11719 ^ w11721 ;
  assign w11723 = ~\pi096 & w4654 ;
  assign w11724 = \pi095 & w4876 ;
  assign w11725 = ( w4654 & ~w11723 ) | ( w4654 & w11724 ) | ( ~w11723 & w11724 ) ;
  assign w11726 = ~\pi097 & w4656 ;
  assign w11727 = w2673 | w11725 ;
  assign w11728 = ( w4657 & w11725 ) | ( w4657 & w11727 ) | ( w11725 & w11727 ) ;
  assign w11729 = ( w4656 & ~w11726 ) | ( w4656 & w11728 ) | ( ~w11726 & w11728 ) ;
  assign w11730 = \pi047 ^ w11729 ;
  assign w11731 = w11656 ^ w11722 ;
  assign w11732 = w11730 ^ w11731 ;
  assign w11733 = ~\pi099 & w4141 ;
  assign w11734 = \pi098 & w4334 ;
  assign w11735 = ( w4141 & ~w11733 ) | ( w4141 & w11734 ) | ( ~w11733 & w11734 ) ;
  assign w11736 = ~\pi100 & w4143 ;
  assign w11737 = w3104 | w11735 ;
  assign w11738 = ( w4144 & w11735 ) | ( w4144 & w11737 ) | ( w11735 & w11737 ) ;
  assign w11739 = ( w4143 & ~w11736 ) | ( w4143 & w11738 ) | ( ~w11736 & w11738 ) ;
  assign w11740 = \pi044 ^ w11739 ;
  assign w11741 = w11655 ^ w11732 ;
  assign w11742 = w11740 ^ w11741 ;
  assign w11743 = ~\pi102 & w3635 ;
  assign w11744 = \pi101 & w3817 ;
  assign w11745 = ( w3635 & ~w11743 ) | ( w3635 & w11744 ) | ( ~w11743 & w11744 ) ;
  assign w11746 = ~\pi103 & w3637 ;
  assign w11747 = w3437 | w11745 ;
  assign w11748 = ( w3638 & w11745 ) | ( w3638 & w11747 ) | ( w11745 & w11747 ) ;
  assign w11749 = ( w3637 & ~w11746 ) | ( w3637 & w11748 ) | ( ~w11746 & w11748 ) ;
  assign w11750 = \pi041 ^ w11749 ;
  assign w11751 = w11654 ^ w11742 ;
  assign w11752 = w11750 ^ w11751 ;
  assign w11753 = ~\pi105 & w3178 ;
  assign w11754 = \pi104 & w3340 ;
  assign w11755 = ( w3178 & ~w11753 ) | ( w3178 & w11754 ) | ( ~w11753 & w11754 ) ;
  assign w11756 = ~\pi106 & w3180 ;
  assign w11757 = w4068 | w11755 ;
  assign w11758 = ( w3181 & w11755 ) | ( w3181 & w11757 ) | ( w11755 & w11757 ) ;
  assign w11759 = ( w3180 & ~w11756 ) | ( w3180 & w11758 ) | ( ~w11756 & w11758 ) ;
  assign w11760 = \pi038 ^ w11759 ;
  assign w11761 = w11653 ^ w11752 ;
  assign w11762 = w11760 ^ w11761 ;
  assign w11763 = ~\pi108 & w2712 ;
  assign w11764 = \pi107 & w2872 ;
  assign w11765 = ( w2712 & ~w11763 ) | ( w2712 & w11764 ) | ( ~w11763 & w11764 ) ;
  assign w11766 = ~\pi109 & w2714 ;
  assign w11767 = w4599 | w11765 ;
  assign w11768 = ( w2715 & w11765 ) | ( w2715 & w11767 ) | ( w11765 & w11767 ) ;
  assign w11769 = ( w2714 & ~w11766 ) | ( w2714 & w11768 ) | ( ~w11766 & w11768 ) ;
  assign w11770 = \pi035 ^ w11769 ;
  assign w11771 = ( w11449 & w11450 ) | ( w11449 & w11554 ) | ( w11450 & w11554 ) ;
  assign w11772 = w11762 ^ w11771 ;
  assign w11773 = w11770 ^ w11772 ;
  assign w11774 = w4811 | w11441 ;
  assign w11775 = ( w2313 & w11441 ) | ( w2313 & w11774 ) | ( w11441 & w11774 ) ;
  assign w11776 = \pi032 ^ w11775 ;
  assign w11777 = ( w11436 & w11556 ) | ( w11436 & w11776 ) | ( w11556 & w11776 ) ;
  assign w11778 = ~\pi111 & w2310 ;
  assign w11779 = \pi110 & w2443 ;
  assign w11780 = ( w2310 & ~w11778 ) | ( w2310 & w11779 ) | ( ~w11778 & w11779 ) ;
  assign w11781 = ~\pi112 & w2312 ;
  assign w11782 = w4999 | w11780 ;
  assign w11783 = ( w2313 & w11780 ) | ( w2313 & w11782 ) | ( w11780 & w11782 ) ;
  assign w11784 = ( w2312 & ~w11781 ) | ( w2312 & w11783 ) | ( ~w11781 & w11783 ) ;
  assign w11785 = \pi032 ^ w11784 ;
  assign w11786 = w11777 ^ w11785 ;
  assign w11787 = w11648 ^ w11773 ;
  assign w11788 = w11652 ^ w11787 ;
  assign w11789 = w11786 ^ w11788 ;
  assign w11790 = w11630 ^ w11789 ;
  assign w11791 = w11622 ^ w11790 ;
  assign w11792 = w11640 ^ w11791 ;
  assign w11793 = w11610 ^ w11792 ;
  assign w11794 = w11602 ^ w11793 ;
  assign w11795 = w11621 ^ w11794 ;
  assign w11796 = ( w11400 & w11404 ) | ( w11400 & w11594 ) | ( w11404 & w11594 ) ;
  assign w11797 = ( w11398 & w11399 ) | ( w11398 & w11596 ) | ( w11399 & w11596 ) ;
  assign w11798 = w11796 ^ w11797 ;
  assign w11799 = w11795 ^ w11798 ;
  assign w11800 = ( w11618 & w11620 ) | ( w11618 & w11792 ) | ( w11620 & w11792 ) ;
  assign w11801 = \pi127 & w837 ;
  assign w11802 = ( \pi126 & ~w840 ) | ( \pi126 & w8490 ) | ( ~w840 & w8490 ) ;
  assign w11803 = \pi126 & ~w902 ;
  assign w11804 = ( ~\pi126 & w11802 ) | ( ~\pi126 & w11803 ) | ( w11802 & w11803 ) ;
  assign w11805 = ( w9420 & w11801 ) | ( w9420 & ~w11804 ) | ( w11801 & ~w11804 ) ;
  assign w11806 = ~\pi124 & w1044 ;
  assign w11807 = \pi123 & w1138 ;
  assign w11808 = ( w1044 & ~w11806 ) | ( w1044 & w11807 ) | ( ~w11806 & w11807 ) ;
  assign w11809 = ~\pi125 & w1046 ;
  assign w11810 = w7988 | w11808 ;
  assign w11811 = ( w1047 & w11808 ) | ( w1047 & w11810 ) | ( w11808 & w11810 ) ;
  assign w11812 = ( w1046 & ~w11809 ) | ( w1046 & w11811 ) | ( ~w11809 & w11811 ) ;
  assign w11813 = \pi020 ^ w11812 ;
  assign w11814 = w11640 ^ w11789 ;
  assign w11815 = ( w11622 & w11630 ) | ( w11622 & w11814 ) | ( w11630 & w11814 ) ;
  assign w11816 = w11813 ^ w11815 ;
  assign w11817 = ( w11638 & w11639 ) | ( w11638 & w11789 ) | ( w11639 & w11789 ) ;
  assign w11818 = \pi120 & w1417 ;
  assign w11819 = ( \pi122 & w1315 ) | ( \pi122 & w11818 ) | ( w1315 & w11818 ) ;
  assign w11820 = \pi121 | w11819 ;
  assign w11821 = ( w1313 & w11819 ) | ( w1313 & w11820 ) | ( w11819 & w11820 ) ;
  assign w11822 = w11818 | w11821 ;
  assign w11823 = ~w1316 & w7069 ;
  assign w11824 = ( w7069 & w11822 ) | ( w7069 & ~w11823 ) | ( w11822 & ~w11823 ) ;
  assign w11825 = \pi023 ^ w11824 ;
  assign w11826 = ~\pi118 & w1629 ;
  assign w11827 = \pi117 & w1722 ;
  assign w11828 = ( w1629 & ~w11826 ) | ( w1629 & w11827 ) | ( ~w11826 & w11827 ) ;
  assign w11829 = ~\pi119 & w1631 ;
  assign w11830 = w6616 | w11828 ;
  assign w11831 = ( w1632 & w11828 ) | ( w1632 & w11830 ) | ( w11828 & w11830 ) ;
  assign w11832 = ( w1631 & ~w11829 ) | ( w1631 & w11831 ) | ( ~w11829 & w11831 ) ;
  assign w11833 = \pi026 ^ w11832 ;
  assign w11834 = w11773 ^ w11786 ;
  assign w11835 = ( w11648 & w11652 ) | ( w11648 & w11834 ) | ( w11652 & w11834 ) ;
  assign w11836 = w11833 ^ w11835 ;
  assign w11837 = ~\pi115 & w1944 ;
  assign w11838 = \pi114 & w2072 ;
  assign w11839 = ( w1944 & ~w11837 ) | ( w1944 & w11838 ) | ( ~w11837 & w11838 ) ;
  assign w11840 = ~\pi116 & w1946 ;
  assign w11841 = w5976 | w11839 ;
  assign w11842 = ( w1947 & w11839 ) | ( w1947 & w11841 ) | ( w11839 & w11841 ) ;
  assign w11843 = ( w1946 & ~w11840 ) | ( w1946 & w11842 ) | ( ~w11840 & w11842 ) ;
  assign w11844 = \pi029 ^ w11843 ;
  assign w11845 = ( w11773 & w11777 ) | ( w11773 & w11785 ) | ( w11777 & w11785 ) ;
  assign w11846 = ~\pi112 & w2310 ;
  assign w11847 = \pi111 & w2443 ;
  assign w11848 = ( w2310 & ~w11846 ) | ( w2310 & w11847 ) | ( ~w11846 & w11847 ) ;
  assign w11849 = ~\pi113 & w2312 ;
  assign w11850 = w5366 | w11848 ;
  assign w11851 = ( w2313 & w11848 ) | ( w2313 & w11850 ) | ( w11848 & w11850 ) ;
  assign w11852 = ( w2312 & ~w11849 ) | ( w2312 & w11851 ) | ( ~w11849 & w11851 ) ;
  assign w11853 = \pi032 ^ w11852 ;
  assign w11854 = ( w11762 & w11770 ) | ( w11762 & w11771 ) | ( w11770 & w11771 ) ;
  assign w11855 = w11853 ^ w11854 ;
  assign w11856 = ~\pi106 & w3178 ;
  assign w11857 = \pi105 & w3340 ;
  assign w11858 = ( w3178 & ~w11856 ) | ( w3178 & w11857 ) | ( ~w11856 & w11857 ) ;
  assign w11859 = ~\pi107 & w3180 ;
  assign w11860 = w4087 | w11858 ;
  assign w11861 = ( w3181 & w11858 ) | ( w3181 & w11860 ) | ( w11858 & w11860 ) ;
  assign w11862 = ( w3180 & ~w11859 ) | ( w3180 & w11861 ) | ( ~w11859 & w11861 ) ;
  assign w11863 = \pi038 ^ w11862 ;
  assign w11864 = ( w11654 & w11742 ) | ( w11654 & w11750 ) | ( w11742 & w11750 ) ;
  assign w11865 = ~\pi103 & w3635 ;
  assign w11866 = \pi102 & w3817 ;
  assign w11867 = ( w3635 & ~w11865 ) | ( w3635 & w11866 ) | ( ~w11865 & w11866 ) ;
  assign w11868 = ~\pi104 & w3637 ;
  assign w11869 = w3740 | w11867 ;
  assign w11870 = ( w3638 & w11867 ) | ( w3638 & w11869 ) | ( w11867 & w11869 ) ;
  assign w11871 = ( w3637 & ~w11868 ) | ( w3637 & w11870 ) | ( ~w11868 & w11870 ) ;
  assign w11872 = \pi041 ^ w11871 ;
  assign w11873 = ( w11655 & w11732 ) | ( w11655 & w11740 ) | ( w11732 & w11740 ) ;
  assign w11874 = ~\pi100 & w4141 ;
  assign w11875 = \pi099 & w4334 ;
  assign w11876 = ( w4141 & ~w11874 ) | ( w4141 & w11875 ) | ( ~w11874 & w11875 ) ;
  assign w11877 = ~\pi101 & w4143 ;
  assign w11878 = w3264 | w11876 ;
  assign w11879 = ( w4144 & w11876 ) | ( w4144 & w11878 ) | ( w11876 & w11878 ) ;
  assign w11880 = ( w4143 & ~w11877 ) | ( w4143 & w11879 ) | ( ~w11877 & w11879 ) ;
  assign w11881 = \pi044 ^ w11880 ;
  assign w11882 = ( w11656 & w11722 ) | ( w11656 & w11730 ) | ( w11722 & w11730 ) ;
  assign w11883 = ~\pi094 & w5209 ;
  assign w11884 = \pi093 & w5433 ;
  assign w11885 = ( w5209 & ~w11883 ) | ( w5209 & w11884 ) | ( ~w11883 & w11884 ) ;
  assign w11886 = ~\pi095 & w5211 ;
  assign w11887 = w2409 | w11885 ;
  assign w11888 = ( w5212 & w11885 ) | ( w5212 & w11887 ) | ( w11885 & w11887 ) ;
  assign w11889 = ( w5211 & ~w11886 ) | ( w5211 & w11888 ) | ( ~w11886 & w11888 ) ;
  assign w11890 = \pi050 ^ w11889 ;
  assign w11891 = ( w11669 & w11675 ) | ( w11669 & ~w11676 ) | ( w11675 & ~w11676 ) ;
  assign w11892 = \pi063 & \pi078 ;
  assign w11893 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w11892 ) | ( \pi063 & w11892 ) ;
  assign w11894 = ( \pi062 & ~\pi063 ) | ( \pi062 & w11892 ) | ( ~\pi063 & w11892 ) ;
  assign w11895 = ( \pi079 & w11893 ) | ( \pi079 & w11894 ) | ( w11893 & w11894 ) ;
  assign w11896 = ( ~\pi014 & w11275 ) | ( ~\pi014 & w11895 ) | ( w11275 & w11895 ) ;
  assign w11897 = ~\pi082 & w7811 ;
  assign w11898 = \pi081 & w8046 ;
  assign w11899 = ( w7811 & ~w11897 ) | ( w7811 & w11898 ) | ( ~w11897 & w11898 ) ;
  assign w11900 = ~\pi083 & w7813 ;
  assign w11901 = ~w1099 & w7814 ;
  assign w11902 = ( w7814 & w11899 ) | ( w7814 & ~w11901 ) | ( w11899 & ~w11901 ) ;
  assign w11903 = ( w7813 & ~w11900 ) | ( w7813 & w11902 ) | ( ~w11900 & w11902 ) ;
  assign w11904 = w11896 ^ w11903 ;
  assign w11905 = \pi062 ^ \pi080 ;
  assign w11906 = \pi063 ^ \pi080 ;
  assign w11907 = \pi062 & ~\pi079 ;
  assign w11908 = ( w11905 & ~w11906 ) | ( w11905 & w11907 ) | ( ~w11906 & w11907 ) ;
  assign w11909 = w11904 ^ w11908 ;
  assign w11910 = ~\pi085 & w7135 ;
  assign w11911 = \pi084 & w7359 ;
  assign w11912 = ( w7135 & ~w11910 ) | ( w7135 & w11911 ) | ( ~w11910 & w11911 ) ;
  assign w11913 = ~\pi086 & w7137 ;
  assign w11914 = w1379 | w11912 ;
  assign w11915 = ( w7138 & w11912 ) | ( w7138 & w11914 ) | ( w11912 & w11914 ) ;
  assign w11916 = ( w7137 & ~w11913 ) | ( w7137 & w11915 ) | ( ~w11913 & w11915 ) ;
  assign w11917 = \pi059 ^ w11916 ;
  assign w11918 = w11891 ^ w11909 ;
  assign w11919 = w11917 ^ w11918 ;
  assign w11920 = ( ~w11678 & w11686 ) | ( ~w11678 & w11687 ) | ( w11686 & w11687 ) ;
  assign w11921 = ~\pi088 & w6466 ;
  assign w11922 = \pi087 & w6702 ;
  assign w11923 = ( w6466 & ~w11921 ) | ( w6466 & w11922 ) | ( ~w11921 & w11922 ) ;
  assign w11924 = ~\pi089 & w6468 ;
  assign w11925 = w1595 | w11923 ;
  assign w11926 = ( w6469 & w11923 ) | ( w6469 & w11925 ) | ( w11923 & w11925 ) ;
  assign w11927 = ( w6468 & ~w11924 ) | ( w6468 & w11926 ) | ( ~w11924 & w11926 ) ;
  assign w11928 = \pi056 ^ w11927 ;
  assign w11929 = w11919 ^ w11920 ;
  assign w11930 = w11928 ^ w11929 ;
  assign w11931 = ~\pi091 & w5802 ;
  assign w11932 = \pi090 & w6052 ;
  assign w11933 = ( w5802 & ~w11931 ) | ( w5802 & w11932 ) | ( ~w11931 & w11932 ) ;
  assign w11934 = ~\pi092 & w5804 ;
  assign w11935 = w2033 | w11933 ;
  assign w11936 = ( w5805 & w11933 ) | ( w5805 & w11935 ) | ( w11933 & w11935 ) ;
  assign w11937 = ( w5804 & ~w11934 ) | ( w5804 & w11936 ) | ( ~w11934 & w11936 ) ;
  assign w11938 = \pi053 ^ w11937 ;
  assign w11939 = w11698 ^ w11930 ;
  assign w11940 = w11938 ^ w11939 ;
  assign w11941 = ( ~w11700 & w11708 ) | ( ~w11700 & w11709 ) | ( w11708 & w11709 ) ;
  assign w11942 = w11940 ^ w11941 ;
  assign w11943 = w11890 ^ w11942 ;
  assign w11944 = ( w11711 & ~w11719 ) | ( w11711 & w11720 ) | ( ~w11719 & w11720 ) ;
  assign w11945 = ~\pi097 & w4654 ;
  assign w11946 = \pi096 & w4876 ;
  assign w11947 = ( w4654 & ~w11945 ) | ( w4654 & w11946 ) | ( ~w11945 & w11946 ) ;
  assign w11948 = ~\pi098 & w4656 ;
  assign w11949 = w2824 | w11947 ;
  assign w11950 = ( w4657 & w11947 ) | ( w4657 & w11949 ) | ( w11947 & w11949 ) ;
  assign w11951 = ( w4656 & ~w11948 ) | ( w4656 & w11950 ) | ( ~w11948 & w11950 ) ;
  assign w11952 = \pi047 ^ w11951 ;
  assign w11953 = w11943 ^ w11944 ;
  assign w11954 = w11952 ^ w11953 ;
  assign w11955 = w11882 ^ w11954 ;
  assign w11956 = w11881 ^ w11955 ;
  assign w11957 = w11873 ^ w11956 ;
  assign w11958 = w11872 ^ w11957 ;
  assign w11959 = w11864 ^ w11958 ;
  assign w11960 = w11863 ^ w11959 ;
  assign w11961 = ( w11653 & w11752 ) | ( w11653 & w11760 ) | ( w11752 & w11760 ) ;
  assign w11962 = ~\pi109 & w2712 ;
  assign w11963 = \pi108 & w2872 ;
  assign w11964 = ( w2712 & ~w11962 ) | ( w2712 & w11963 ) | ( ~w11962 & w11963 ) ;
  assign w11965 = ~\pi110 & w2714 ;
  assign w11966 = w4792 | w11964 ;
  assign w11967 = ( w2715 & w11964 ) | ( w2715 & w11966 ) | ( w11964 & w11966 ) ;
  assign w11968 = ( w2714 & ~w11965 ) | ( w2714 & w11967 ) | ( ~w11965 & w11967 ) ;
  assign w11969 = \pi035 ^ w11968 ;
  assign w11970 = w11960 ^ w11961 ;
  assign w11971 = w11969 ^ w11970 ;
  assign w11972 = w11844 ^ w11971 ;
  assign w11973 = w11845 ^ w11972 ;
  assign w11974 = w11855 ^ w11973 ;
  assign w11975 = w11825 ^ w11974 ;
  assign w11976 = w11817 ^ w11975 ;
  assign w11977 = w11836 ^ w11976 ;
  assign w11978 = w11816 ^ w11977 ;
  assign w11979 = w11800 ^ w11805 ;
  assign w11980 = \pi017 ^ w11979 ;
  assign w11981 = w11978 ^ w11980 ;
  assign w11982 = w11621 ^ w11792 ;
  assign w11983 = ( w11602 & w11610 ) | ( w11602 & w11982 ) | ( w11610 & w11982 ) ;
  assign w11984 = ( w11795 & w11796 ) | ( w11795 & w11797 ) | ( w11796 & w11797 ) ;
  assign w11985 = w11983 ^ w11984 ;
  assign w11986 = w11981 ^ w11985 ;
  assign w11987 = ( w11981 & w11983 ) | ( w11981 & w11984 ) | ( w11983 & w11984 ) ;
  assign w11988 = \pi017 ^ w11805 ;
  assign w11989 = ( w11800 & w11978 ) | ( w11800 & w11988 ) | ( w11978 & w11988 ) ;
  assign w11990 = ( w11813 & w11815 ) | ( w11813 & w11977 ) | ( w11815 & w11977 ) ;
  assign w11991 = w840 & w8481 ;
  assign w11992 = w902 | w11991 ;
  assign w11993 = ( \pi127 & w11991 ) | ( \pi127 & w11992 ) | ( w11991 & w11992 ) ;
  assign w11994 = \pi017 ^ w11993 ;
  assign w11995 = ~\pi125 & w1044 ;
  assign w11996 = \pi124 & w1138 ;
  assign w11997 = ( w1044 & ~w11995 ) | ( w1044 & w11996 ) | ( ~w11995 & w11996 ) ;
  assign w11998 = ~\pi126 & w1046 ;
  assign w11999 = w8231 | w11997 ;
  assign w12000 = ( w1047 & w11997 ) | ( w1047 & w11999 ) | ( w11997 & w11999 ) ;
  assign w12001 = ( w1046 & ~w11998 ) | ( w1046 & w12000 ) | ( ~w11998 & w12000 ) ;
  assign w12002 = \pi020 ^ w12001 ;
  assign w12003 = w11836 ^ w11974 ;
  assign w12004 = ( w11817 & w11825 ) | ( w11817 & w12003 ) | ( w11825 & w12003 ) ;
  assign w12005 = ~\pi122 & w1313 ;
  assign w12006 = \pi121 & w1417 ;
  assign w12007 = ( w1313 & ~w12005 ) | ( w1313 & w12006 ) | ( ~w12005 & w12006 ) ;
  assign w12008 = ~\pi123 & w1315 ;
  assign w12009 = w7516 | w12007 ;
  assign w12010 = ( w1316 & w12007 ) | ( w1316 & w12009 ) | ( w12007 & w12009 ) ;
  assign w12011 = ( w1315 & ~w12008 ) | ( w1315 & w12010 ) | ( ~w12008 & w12010 ) ;
  assign w12012 = \pi023 ^ w12011 ;
  assign w12013 = ( w11833 & w11835 ) | ( w11833 & w11974 ) | ( w11835 & w11974 ) ;
  assign w12014 = ~\pi119 & w1629 ;
  assign w12015 = \pi118 & w1722 ;
  assign w12016 = ( w1629 & ~w12014 ) | ( w1629 & w12015 ) | ( ~w12014 & w12015 ) ;
  assign w12017 = ~\pi120 & w1631 ;
  assign w12018 = w6634 | w12016 ;
  assign w12019 = ( w1632 & w12016 ) | ( w1632 & w12018 ) | ( w12016 & w12018 ) ;
  assign w12020 = ( w1631 & ~w12017 ) | ( w1631 & w12019 ) | ( ~w12017 & w12019 ) ;
  assign w12021 = \pi026 ^ w12020 ;
  assign w12022 = w11855 ^ w11971 ;
  assign w12023 = ( w11844 & w11845 ) | ( w11844 & w12022 ) | ( w11845 & w12022 ) ;
  assign w12024 = w12021 ^ w12023 ;
  assign w12025 = ~\pi116 & w1944 ;
  assign w12026 = \pi115 & w2072 ;
  assign w12027 = ( w1944 & ~w12025 ) | ( w1944 & w12026 ) | ( ~w12025 & w12026 ) ;
  assign w12028 = ~\pi117 & w1946 ;
  assign w12029 = w6185 | w12027 ;
  assign w12030 = ( w1947 & w12027 ) | ( w1947 & w12029 ) | ( w12027 & w12029 ) ;
  assign w12031 = ( w1946 & ~w12028 ) | ( w1946 & w12030 ) | ( ~w12028 & w12030 ) ;
  assign w12032 = \pi029 ^ w12031 ;
  assign w12033 = ( w11853 & w11854 ) | ( w11853 & w11971 ) | ( w11854 & w11971 ) ;
  assign w12034 = ~\pi113 & w2310 ;
  assign w12035 = \pi112 & w2443 ;
  assign w12036 = ( w2310 & ~w12034 ) | ( w2310 & w12035 ) | ( ~w12034 & w12035 ) ;
  assign w12037 = ~\pi114 & w2312 ;
  assign w12038 = w5565 | w12036 ;
  assign w12039 = ( w2313 & w12036 ) | ( w2313 & w12038 ) | ( w12036 & w12038 ) ;
  assign w12040 = ( w2312 & ~w12037 ) | ( w2312 & w12039 ) | ( ~w12037 & w12039 ) ;
  assign w12041 = \pi032 ^ w12040 ;
  assign w12042 = ( w11960 & w11961 ) | ( w11960 & w11969 ) | ( w11961 & w11969 ) ;
  assign w12043 = w12041 ^ w12042 ;
  assign w12044 = ( w11863 & w11864 ) | ( w11863 & w11958 ) | ( w11864 & w11958 ) ;
  assign w12045 = ~\pi107 & w3178 ;
  assign w12046 = \pi106 & w3340 ;
  assign w12047 = ( w3178 & ~w12045 ) | ( w3178 & w12046 ) | ( ~w12045 & w12046 ) ;
  assign w12048 = ~\pi108 & w3180 ;
  assign w12049 = w4425 | w12047 ;
  assign w12050 = ( w3181 & w12047 ) | ( w3181 & w12049 ) | ( w12047 & w12049 ) ;
  assign w12051 = ( w3180 & ~w12048 ) | ( w3180 & w12050 ) | ( ~w12048 & w12050 ) ;
  assign w12052 = \pi038 ^ w12051 ;
  assign w12053 = ( w11872 & w11873 ) | ( w11872 & w11956 ) | ( w11873 & w11956 ) ;
  assign w12054 = ~\pi104 & w3635 ;
  assign w12055 = \pi103 & w3817 ;
  assign w12056 = ( w3635 & ~w12054 ) | ( w3635 & w12055 ) | ( ~w12054 & w12055 ) ;
  assign w12057 = ~\pi105 & w3637 ;
  assign w12058 = w3905 | w12056 ;
  assign w12059 = ( w3638 & w12056 ) | ( w3638 & w12058 ) | ( w12056 & w12058 ) ;
  assign w12060 = ( w3637 & ~w12057 ) | ( w3637 & w12059 ) | ( ~w12057 & w12059 ) ;
  assign w12061 = \pi041 ^ w12060 ;
  assign w12062 = ( w11881 & w11882 ) | ( w11881 & w11954 ) | ( w11882 & w11954 ) ;
  assign w12063 = ( ~w11919 & w11920 ) | ( ~w11919 & w11928 ) | ( w11920 & w11928 ) ;
  assign w12064 = ~\pi089 & w6466 ;
  assign w12065 = \pi088 & w6702 ;
  assign w12066 = ( w6466 & ~w12064 ) | ( w6466 & w12065 ) | ( ~w12064 & w12065 ) ;
  assign w12067 = ~\pi090 & w6468 ;
  assign w12068 = w1801 | w12066 ;
  assign w12069 = ( w6469 & w12066 ) | ( w6469 & w12068 ) | ( w12066 & w12068 ) ;
  assign w12070 = ( w6468 & ~w12067 ) | ( w6468 & w12069 ) | ( ~w12067 & w12069 ) ;
  assign w12071 = \pi056 ^ w12070 ;
  assign w12072 = ( w11891 & ~w11909 ) | ( w11891 & w11917 ) | ( ~w11909 & w11917 ) ;
  assign w12073 = ~\pi083 & w7811 ;
  assign w12074 = \pi082 & w8046 ;
  assign w12075 = ( w7811 & ~w12073 ) | ( w7811 & w12074 ) | ( ~w12073 & w12074 ) ;
  assign w12076 = ~\pi084 & w7813 ;
  assign w12077 = w1188 | w12075 ;
  assign w12078 = ( w7814 & w12075 ) | ( w7814 & w12077 ) | ( w12075 & w12077 ) ;
  assign w12079 = ( w7813 & ~w12076 ) | ( w7813 & w12078 ) | ( ~w12076 & w12078 ) ;
  assign w12080 = \pi062 ^ w12079 ;
  assign w12081 = \pi080 & ~w12080 ;
  assign w12082 = ( \pi063 & ~\pi079 ) | ( \pi063 & w12081 ) | ( ~\pi079 & w12081 ) ;
  assign w12083 = ( \pi062 & ~\pi063 ) | ( \pi062 & w12082 ) | ( ~\pi063 & w12082 ) ;
  assign w12084 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi081 ) | ( \pi063 & ~\pi081 ) ;
  assign w12085 = ( \pi080 & w12080 ) | ( \pi080 & w12084 ) | ( w12080 & w12084 ) ;
  assign w12086 = ( ~\pi063 & w12080 ) | ( ~\pi063 & w12081 ) | ( w12080 & w12081 ) ;
  assign w12087 = ( \pi062 & ~\pi080 ) | ( \pi062 & w12086 ) | ( ~\pi080 & w12086 ) ;
  assign w12088 = ( ~w12083 & w12085 ) | ( ~w12083 & w12087 ) | ( w12085 & w12087 ) ;
  assign w12089 = \pi079 ^ \pi081 ;
  assign w12090 = ( \pi062 & \pi063 ) | ( \pi062 & ~w12089 ) | ( \pi063 & ~w12089 ) ;
  assign w12091 = \pi079 ^ \pi080 ;
  assign w12092 = \pi062 & ~w12091 ;
  assign w12093 = ( \pi063 & ~w12091 ) | ( \pi063 & w12092 ) | ( ~w12091 & w12092 ) ;
  assign w12094 = w12080 ^ w12093 ;
  assign w12095 = w12090 ^ w12094 ;
  assign w12096 = \pi062 ^ w11903 ;
  assign w12097 = ( \pi062 & \pi063 ) | ( \pi062 & \pi080 ) | ( \pi063 & \pi080 ) ;
  assign w12098 = \pi062 & \pi079 ;
  assign w12099 = ( ~\pi062 & w12097 ) | ( ~\pi062 & w12098 ) | ( w12097 & w12098 ) ;
  assign w12100 = ( ~\pi063 & w12097 ) | ( ~\pi063 & w12099 ) | ( w12097 & w12099 ) ;
  assign w12101 = ( w11896 & w12096 ) | ( w11896 & ~w12100 ) | ( w12096 & ~w12100 ) ;
  assign w12102 = ~\pi086 & w7135 ;
  assign w12103 = \pi085 & w7359 ;
  assign w12104 = ( w7135 & ~w12102 ) | ( w7135 & w12103 ) | ( ~w12102 & w12103 ) ;
  assign w12105 = ~\pi087 & w7137 ;
  assign w12106 = w1477 | w12104 ;
  assign w12107 = ( w7138 & w12104 ) | ( w7138 & w12106 ) | ( w12104 & w12106 ) ;
  assign w12108 = ( w7137 & ~w12105 ) | ( w7137 & w12107 ) | ( ~w12105 & w12107 ) ;
  assign w12109 = \pi059 ^ w12108 ;
  assign w12110 = w12095 ^ w12101 ;
  assign w12111 = w12109 ^ w12110 ;
  assign w12112 = w12071 ^ w12072 ;
  assign w12113 = w12111 ^ w12112 ;
  assign w12114 = ~\pi092 & w5802 ;
  assign w12115 = \pi091 & w6052 ;
  assign w12116 = ( w5802 & ~w12114 ) | ( w5802 & w12115 ) | ( ~w12114 & w12115 ) ;
  assign w12117 = ~\pi093 & w5804 ;
  assign w12118 = w2155 | w12116 ;
  assign w12119 = ( w5805 & w12116 ) | ( w5805 & w12118 ) | ( w12116 & w12118 ) ;
  assign w12120 = ( w5804 & ~w12117 ) | ( w5804 & w12119 ) | ( ~w12117 & w12119 ) ;
  assign w12121 = \pi053 ^ w12120 ;
  assign w12122 = w12063 ^ w12113 ;
  assign w12123 = w12121 ^ w12122 ;
  assign w12124 = ( w11698 & ~w11930 ) | ( w11698 & w11938 ) | ( ~w11930 & w11938 ) ;
  assign w12125 = ~\pi095 & w5209 ;
  assign w12126 = \pi094 & w5433 ;
  assign w12127 = ( w5209 & ~w12125 ) | ( w5209 & w12126 ) | ( ~w12125 & w12126 ) ;
  assign w12128 = ~\pi096 & w5211 ;
  assign w12129 = w2546 | w12127 ;
  assign w12130 = ( w5212 & w12127 ) | ( w5212 & w12129 ) | ( w12127 & w12129 ) ;
  assign w12131 = ( w5211 & ~w12128 ) | ( w5211 & w12130 ) | ( ~w12128 & w12130 ) ;
  assign w12132 = \pi050 ^ w12131 ;
  assign w12133 = w12123 ^ w12124 ;
  assign w12134 = w12132 ^ w12133 ;
  assign w12135 = ( w11890 & ~w11940 ) | ( w11890 & w11941 ) | ( ~w11940 & w11941 ) ;
  assign w12136 = ~\pi098 & w4654 ;
  assign w12137 = \pi097 & w4876 ;
  assign w12138 = ( w4654 & ~w12136 ) | ( w4654 & w12137 ) | ( ~w12136 & w12137 ) ;
  assign w12139 = ~\pi099 & w4656 ;
  assign w12140 = w2966 | w12138 ;
  assign w12141 = ( w4657 & w12138 ) | ( w4657 & w12140 ) | ( w12138 & w12140 ) ;
  assign w12142 = ( w4656 & ~w12139 ) | ( w4656 & w12141 ) | ( ~w12139 & w12141 ) ;
  assign w12143 = \pi047 ^ w12142 ;
  assign w12144 = w12134 ^ w12135 ;
  assign w12145 = w12143 ^ w12144 ;
  assign w12146 = ( w11943 & w11944 ) | ( w11943 & ~w11952 ) | ( w11944 & ~w11952 ) ;
  assign w12147 = ~\pi101 & w4141 ;
  assign w12148 = \pi100 & w4334 ;
  assign w12149 = ( w4141 & ~w12147 ) | ( w4141 & w12148 ) | ( ~w12147 & w12148 ) ;
  assign w12150 = ~\pi102 & w4143 ;
  assign w12151 = w3284 | w12149 ;
  assign w12152 = ( w4144 & w12149 ) | ( w4144 & w12151 ) | ( w12149 & w12151 ) ;
  assign w12153 = ( w4143 & ~w12150 ) | ( w4143 & w12152 ) | ( ~w12150 & w12152 ) ;
  assign w12154 = \pi044 ^ w12153 ;
  assign w12155 = w12145 ^ w12146 ;
  assign w12156 = w12154 ^ w12155 ;
  assign w12157 = w12062 ^ w12156 ;
  assign w12158 = w12061 ^ w12157 ;
  assign w12159 = w12053 ^ w12158 ;
  assign w12160 = w12052 ^ w12159 ;
  assign w12161 = ~\pi110 & w2712 ;
  assign w12162 = \pi109 & w2872 ;
  assign w12163 = ( w2712 & ~w12161 ) | ( w2712 & w12162 ) | ( ~w12161 & w12162 ) ;
  assign w12164 = ~\pi111 & w2714 ;
  assign w12165 = w4811 | w12163 ;
  assign w12166 = ( w2715 & w12163 ) | ( w2715 & w12165 ) | ( w12163 & w12165 ) ;
  assign w12167 = ( w2714 & ~w12164 ) | ( w2714 & w12166 ) | ( ~w12164 & w12166 ) ;
  assign w12168 = \pi035 ^ w12167 ;
  assign w12169 = w12044 ^ w12160 ;
  assign w12170 = w12168 ^ w12169 ;
  assign w12171 = w12032 ^ w12170 ;
  assign w12172 = w12033 ^ w12171 ;
  assign w12173 = w12043 ^ w12172 ;
  assign w12174 = w12012 ^ w12173 ;
  assign w12175 = w12013 ^ w12174 ;
  assign w12176 = w12024 ^ w12175 ;
  assign w12177 = w12004 ^ w12176 ;
  assign w12178 = w12002 ^ w12177 ;
  assign w12179 = w11990 ^ w12178 ;
  assign w12180 = w11994 ^ w12179 ;
  assign w12181 = w11987 ^ w11989 ;
  assign w12182 = w12180 ^ w12181 ;
  assign w12183 = ( w11987 & w11989 ) | ( w11987 & w12180 ) | ( w11989 & w12180 ) ;
  assign w12184 = ( w11990 & w11994 ) | ( w11990 & w12178 ) | ( w11994 & w12178 ) ;
  assign w12185 = ( w12002 & w12004 ) | ( w12002 & w12176 ) | ( w12004 & w12176 ) ;
  assign w12186 = ~\pi126 & w1044 ;
  assign w12187 = \pi125 & w1138 ;
  assign w12188 = ( w1044 & ~w12186 ) | ( w1044 & w12187 ) | ( ~w12186 & w12187 ) ;
  assign w12189 = ~\pi127 & w1046 ;
  assign w12190 = w8466 | w12188 ;
  assign w12191 = ( w1047 & w12188 ) | ( w1047 & w12190 ) | ( w12188 & w12190 ) ;
  assign w12192 = ( w1046 & ~w12189 ) | ( w1046 & w12191 ) | ( ~w12189 & w12191 ) ;
  assign w12193 = \pi020 ^ w12192 ;
  assign w12194 = ~\pi123 & w1313 ;
  assign w12195 = \pi122 & w1417 ;
  assign w12196 = ( w1313 & ~w12194 ) | ( w1313 & w12195 ) | ( ~w12194 & w12195 ) ;
  assign w12197 = ~\pi124 & w1315 ;
  assign w12198 = w7538 | w12196 ;
  assign w12199 = ( w1316 & w12196 ) | ( w1316 & w12198 ) | ( w12196 & w12198 ) ;
  assign w12200 = ( w1315 & ~w12197 ) | ( w1315 & w12199 ) | ( ~w12197 & w12199 ) ;
  assign w12201 = \pi023 ^ w12200 ;
  assign w12202 = w12024 ^ w12173 ;
  assign w12203 = ( w12012 & w12013 ) | ( w12012 & w12202 ) | ( w12013 & w12202 ) ;
  assign w12204 = ~\pi117 & w1944 ;
  assign w12205 = \pi116 & w2072 ;
  assign w12206 = ( w1944 & ~w12204 ) | ( w1944 & w12205 ) | ( ~w12204 & w12205 ) ;
  assign w12207 = ~\pi118 & w1946 ;
  assign w12208 = w6206 | w12206 ;
  assign w12209 = ( w1947 & w12206 ) | ( w1947 & w12208 ) | ( w12206 & w12208 ) ;
  assign w12210 = ( w1946 & ~w12207 ) | ( w1946 & w12209 ) | ( ~w12207 & w12209 ) ;
  assign w12211 = \pi029 ^ w12210 ;
  assign w12212 = w12043 ^ w12170 ;
  assign w12213 = ( w12032 & w12033 ) | ( w12032 & w12212 ) | ( w12033 & w12212 ) ;
  assign w12214 = ( w12061 & w12062 ) | ( w12061 & w12156 ) | ( w12062 & w12156 ) ;
  assign w12215 = ( w12145 & w12146 ) | ( w12145 & ~w12154 ) | ( w12146 & ~w12154 ) ;
  assign w12216 = ( ~w12134 & w12135 ) | ( ~w12134 & w12143 ) | ( w12135 & w12143 ) ;
  assign w12217 = ~\pi090 & w6466 ;
  assign w12218 = \pi089 & w6702 ;
  assign w12219 = ( w6466 & ~w12217 ) | ( w6466 & w12218 ) | ( ~w12217 & w12218 ) ;
  assign w12220 = ~\pi091 & w6468 ;
  assign w12221 = w1908 | w12219 ;
  assign w12222 = ( w6469 & w12219 ) | ( w6469 & w12221 ) | ( w12219 & w12221 ) ;
  assign w12223 = ( w6468 & ~w12220 ) | ( w6468 & w12222 ) | ( ~w12220 & w12222 ) ;
  assign w12224 = \pi056 ^ w12223 ;
  assign w12225 = ( ~w12095 & w12101 ) | ( ~w12095 & w12109 ) | ( w12101 & w12109 ) ;
  assign w12226 = ~\pi084 & w7811 ;
  assign w12227 = \pi083 & w8046 ;
  assign w12228 = ( w7811 & ~w12226 ) | ( w7811 & w12227 ) | ( ~w12226 & w12227 ) ;
  assign w12229 = ~\pi085 & w7813 ;
  assign w12230 = w1274 | w12228 ;
  assign w12231 = ( w7814 & w12228 ) | ( w7814 & w12230 ) | ( w12228 & w12230 ) ;
  assign w12232 = ( w7813 & ~w12229 ) | ( w7813 & w12231 ) | ( ~w12229 & w12231 ) ;
  assign w12233 = \pi062 ^ w12232 ;
  assign w12234 = \pi080 ^ \pi082 ;
  assign w12235 = ( \pi062 & \pi063 ) | ( \pi062 & ~w12234 ) | ( \pi063 & ~w12234 ) ;
  assign w12236 = \pi062 & ~w873 ;
  assign w12237 = ( \pi063 & ~w873 ) | ( \pi063 & w12236 ) | ( ~w873 & w12236 ) ;
  assign w12238 = \pi017 ^ w12237 ;
  assign w12239 = w12235 ^ w12238 ;
  assign w12240 = w12088 ^ w12233 ;
  assign w12241 = w12239 ^ w12240 ;
  assign w12242 = ~\pi087 & w7135 ;
  assign w12243 = \pi086 & w7359 ;
  assign w12244 = ( w7135 & ~w12242 ) | ( w7135 & w12243 ) | ( ~w12242 & w12243 ) ;
  assign w12245 = ~\pi088 & w7137 ;
  assign w12246 = w1574 | w12244 ;
  assign w12247 = ( w7138 & w12244 ) | ( w7138 & w12246 ) | ( w12244 & w12246 ) ;
  assign w12248 = ( w7137 & ~w12245 ) | ( w7137 & w12247 ) | ( ~w12245 & w12247 ) ;
  assign w12249 = \pi059 ^ w12248 ;
  assign w12250 = w12225 ^ w12241 ;
  assign w12251 = w12249 ^ w12250 ;
  assign w12252 = ( w12071 & w12072 ) | ( w12071 & ~w12111 ) | ( w12072 & ~w12111 ) ;
  assign w12253 = w12251 ^ w12252 ;
  assign w12254 = w12224 ^ w12253 ;
  assign w12255 = ~\pi093 & w5802 ;
  assign w12256 = \pi092 & w6052 ;
  assign w12257 = ( w5802 & ~w12255 ) | ( w5802 & w12256 ) | ( ~w12255 & w12256 ) ;
  assign w12258 = ~\pi094 & w5804 ;
  assign w12259 = w2274 | w12257 ;
  assign w12260 = ( w5805 & w12257 ) | ( w5805 & w12259 ) | ( w12257 & w12259 ) ;
  assign w12261 = ( w5804 & ~w12258 ) | ( w5804 & w12260 ) | ( ~w12258 & w12260 ) ;
  assign w12262 = \pi053 ^ w12261 ;
  assign w12263 = ( w12063 & ~w12113 ) | ( w12063 & w12121 ) | ( ~w12113 & w12121 ) ;
  assign w12264 = w12254 ^ w12263 ;
  assign w12265 = w12262 ^ w12264 ;
  assign w12266 = ~\pi096 & w5209 ;
  assign w12267 = \pi095 & w5433 ;
  assign w12268 = ( w5209 & ~w12266 ) | ( w5209 & w12267 ) | ( ~w12266 & w12267 ) ;
  assign w12269 = ~\pi097 & w5211 ;
  assign w12270 = w2673 | w12268 ;
  assign w12271 = ( w5212 & w12268 ) | ( w5212 & w12270 ) | ( w12268 & w12270 ) ;
  assign w12272 = ( w5211 & ~w12269 ) | ( w5211 & w12271 ) | ( ~w12269 & w12271 ) ;
  assign w12273 = \pi050 ^ w12272 ;
  assign w12274 = ( ~w12123 & w12124 ) | ( ~w12123 & w12132 ) | ( w12124 & w12132 ) ;
  assign w12275 = w12265 ^ w12274 ;
  assign w12276 = w12273 ^ w12275 ;
  assign w12277 = ~\pi099 & w4654 ;
  assign w12278 = \pi098 & w4876 ;
  assign w12279 = ( w4654 & ~w12277 ) | ( w4654 & w12278 ) | ( ~w12277 & w12278 ) ;
  assign w12280 = ~\pi100 & w4656 ;
  assign w12281 = w3104 | w12279 ;
  assign w12282 = ( w4657 & w12279 ) | ( w4657 & w12281 ) | ( w12279 & w12281 ) ;
  assign w12283 = ( w4656 & ~w12280 ) | ( w4656 & w12282 ) | ( ~w12280 & w12282 ) ;
  assign w12284 = \pi047 ^ w12283 ;
  assign w12285 = w12216 ^ w12276 ;
  assign w12286 = w12284 ^ w12285 ;
  assign w12287 = ~\pi102 & w4141 ;
  assign w12288 = \pi101 & w4334 ;
  assign w12289 = ( w4141 & ~w12287 ) | ( w4141 & w12288 ) | ( ~w12287 & w12288 ) ;
  assign w12290 = ~\pi103 & w4143 ;
  assign w12291 = w3437 | w12289 ;
  assign w12292 = ( w4144 & w12289 ) | ( w4144 & w12291 ) | ( w12289 & w12291 ) ;
  assign w12293 = ( w4143 & ~w12290 ) | ( w4143 & w12292 ) | ( ~w12290 & w12292 ) ;
  assign w12294 = \pi044 ^ w12293 ;
  assign w12295 = w12215 ^ w12286 ;
  assign w12296 = w12294 ^ w12295 ;
  assign w12297 = ~\pi105 & w3635 ;
  assign w12298 = \pi104 & w3817 ;
  assign w12299 = ( w3635 & ~w12297 ) | ( w3635 & w12298 ) | ( ~w12297 & w12298 ) ;
  assign w12300 = ~\pi106 & w3637 ;
  assign w12301 = w4068 | w12299 ;
  assign w12302 = ( w3638 & w12299 ) | ( w3638 & w12301 ) | ( w12299 & w12301 ) ;
  assign w12303 = ( w3637 & ~w12300 ) | ( w3637 & w12302 ) | ( ~w12300 & w12302 ) ;
  assign w12304 = \pi041 ^ w12303 ;
  assign w12305 = w12214 ^ w12296 ;
  assign w12306 = w12304 ^ w12305 ;
  assign w12307 = ~\pi108 & w3178 ;
  assign w12308 = \pi107 & w3340 ;
  assign w12309 = ( w3178 & ~w12307 ) | ( w3178 & w12308 ) | ( ~w12307 & w12308 ) ;
  assign w12310 = ~\pi109 & w3180 ;
  assign w12311 = w4599 | w12309 ;
  assign w12312 = ( w3181 & w12309 ) | ( w3181 & w12311 ) | ( w12309 & w12311 ) ;
  assign w12313 = ( w3180 & ~w12310 ) | ( w3180 & w12312 ) | ( ~w12310 & w12312 ) ;
  assign w12314 = \pi038 ^ w12313 ;
  assign w12315 = ( w12052 & w12053 ) | ( w12052 & w12158 ) | ( w12053 & w12158 ) ;
  assign w12316 = w12306 ^ w12315 ;
  assign w12317 = w12314 ^ w12316 ;
  assign w12318 = ~\pi111 & w2712 ;
  assign w12319 = \pi110 & w2872 ;
  assign w12320 = ( w2712 & ~w12318 ) | ( w2712 & w12319 ) | ( ~w12318 & w12319 ) ;
  assign w12321 = ~\pi112 & w2714 ;
  assign w12322 = w4999 | w12320 ;
  assign w12323 = ( w2715 & w12320 ) | ( w2715 & w12322 ) | ( w12320 & w12322 ) ;
  assign w12324 = ( w2714 & ~w12321 ) | ( w2714 & w12323 ) | ( ~w12321 & w12323 ) ;
  assign w12325 = \pi035 ^ w12324 ;
  assign w12326 = ( w12044 & w12160 ) | ( w12044 & w12168 ) | ( w12160 & w12168 ) ;
  assign w12327 = w12317 ^ w12326 ;
  assign w12328 = w12325 ^ w12327 ;
  assign w12329 = ~\pi114 & w2310 ;
  assign w12330 = \pi113 & w2443 ;
  assign w12331 = ( w2310 & ~w12329 ) | ( w2310 & w12330 ) | ( ~w12329 & w12330 ) ;
  assign w12332 = ~\pi115 & w2312 ;
  assign w12333 = w5585 | w12331 ;
  assign w12334 = ( w2313 & w12331 ) | ( w2313 & w12333 ) | ( w12331 & w12333 ) ;
  assign w12335 = ( w2312 & ~w12332 ) | ( w2312 & w12334 ) | ( ~w12332 & w12334 ) ;
  assign w12336 = \pi032 ^ w12335 ;
  assign w12337 = ( w12041 & w12042 ) | ( w12041 & w12170 ) | ( w12042 & w12170 ) ;
  assign w12338 = w12328 ^ w12337 ;
  assign w12339 = w12336 ^ w12338 ;
  assign w12340 = w12213 ^ w12339 ;
  assign w12341 = w12211 ^ w12340 ;
  assign w12342 = ~\pi120 & w1629 ;
  assign w12343 = \pi119 & w1722 ;
  assign w12344 = ( w1629 & ~w12342 ) | ( w1629 & w12343 ) | ( ~w12342 & w12343 ) ;
  assign w12345 = ~\pi121 & w1631 ;
  assign w12346 = w7050 | w12344 ;
  assign w12347 = ( w1632 & w12344 ) | ( w1632 & w12346 ) | ( w12344 & w12346 ) ;
  assign w12348 = ( w1631 & ~w12345 ) | ( w1631 & w12347 ) | ( ~w12345 & w12347 ) ;
  assign w12349 = \pi026 ^ w12348 ;
  assign w12350 = ( w12021 & w12023 ) | ( w12021 & w12173 ) | ( w12023 & w12173 ) ;
  assign w12351 = w12341 ^ w12350 ;
  assign w12352 = w12349 ^ w12351 ;
  assign w12353 = w12203 ^ w12352 ;
  assign w12354 = w12201 ^ w12353 ;
  assign w12355 = w12185 ^ w12354 ;
  assign w12356 = w12193 ^ w12355 ;
  assign w12357 = w12183 ^ w12184 ;
  assign w12358 = w12356 ^ w12357 ;
  assign w12359 = ( w12183 & w12184 ) | ( w12183 & w12356 ) | ( w12184 & w12356 ) ;
  assign w12360 = ( w12185 & w12193 ) | ( w12185 & w12354 ) | ( w12193 & w12354 ) ;
  assign w12361 = ~\pi124 & w1313 ;
  assign w12362 = \pi123 & w1417 ;
  assign w12363 = ( w1313 & ~w12361 ) | ( w1313 & w12362 ) | ( ~w12361 & w12362 ) ;
  assign w12364 = ~\pi125 & w1315 ;
  assign w12365 = w7988 | w12363 ;
  assign w12366 = ( w1316 & w12363 ) | ( w1316 & w12365 ) | ( w12363 & w12365 ) ;
  assign w12367 = ( w1315 & ~w12364 ) | ( w1315 & w12366 ) | ( ~w12364 & w12366 ) ;
  assign w12368 = \pi023 ^ w12367 ;
  assign w12369 = ( w12341 & w12349 ) | ( w12341 & w12350 ) | ( w12349 & w12350 ) ;
  assign w12370 = ~\pi121 & w1629 ;
  assign w12371 = \pi120 & w1722 ;
  assign w12372 = ( w1629 & ~w12370 ) | ( w1629 & w12371 ) | ( ~w12370 & w12371 ) ;
  assign w12373 = ~\pi122 & w1631 ;
  assign w12374 = w7069 | w12372 ;
  assign w12375 = ( w1632 & w12372 ) | ( w1632 & w12374 ) | ( w12372 & w12374 ) ;
  assign w12376 = ( w1631 & ~w12373 ) | ( w1631 & w12375 ) | ( ~w12373 & w12375 ) ;
  assign w12377 = \pi026 ^ w12376 ;
  assign w12378 = ( w12211 & w12213 ) | ( w12211 & w12339 ) | ( w12213 & w12339 ) ;
  assign w12379 = w12377 ^ w12378 ;
  assign w12380 = ~\pi118 & w1944 ;
  assign w12381 = \pi117 & w2072 ;
  assign w12382 = ( w1944 & ~w12380 ) | ( w1944 & w12381 ) | ( ~w12380 & w12381 ) ;
  assign w12383 = ~\pi119 & w1946 ;
  assign w12384 = w6616 | w12382 ;
  assign w12385 = ( w1947 & w12382 ) | ( w1947 & w12384 ) | ( w12382 & w12384 ) ;
  assign w12386 = ( w1946 & ~w12383 ) | ( w1946 & w12385 ) | ( ~w12383 & w12385 ) ;
  assign w12387 = \pi029 ^ w12386 ;
  assign w12388 = ( w12328 & w12336 ) | ( w12328 & w12337 ) | ( w12336 & w12337 ) ;
  assign w12389 = ~\pi115 & w2310 ;
  assign w12390 = \pi114 & w2443 ;
  assign w12391 = ( w2310 & ~w12389 ) | ( w2310 & w12390 ) | ( ~w12389 & w12390 ) ;
  assign w12392 = ~\pi116 & w2312 ;
  assign w12393 = w5976 | w12391 ;
  assign w12394 = ( w2313 & w12391 ) | ( w2313 & w12393 ) | ( w12391 & w12393 ) ;
  assign w12395 = ( w2312 & ~w12392 ) | ( w2312 & w12394 ) | ( ~w12392 & w12394 ) ;
  assign w12396 = \pi032 ^ w12395 ;
  assign w12397 = ( w12317 & w12325 ) | ( w12317 & w12326 ) | ( w12325 & w12326 ) ;
  assign w12398 = w12396 ^ w12397 ;
  assign w12399 = ~\pi106 & w3635 ;
  assign w12400 = \pi105 & w3817 ;
  assign w12401 = ( w3635 & ~w12399 ) | ( w3635 & w12400 ) | ( ~w12399 & w12400 ) ;
  assign w12402 = ~\pi107 & w3637 ;
  assign w12403 = w4087 | w12401 ;
  assign w12404 = ( w3638 & w12401 ) | ( w3638 & w12403 ) | ( w12401 & w12403 ) ;
  assign w12405 = ( w3637 & ~w12402 ) | ( w3637 & w12404 ) | ( ~w12402 & w12404 ) ;
  assign w12406 = \pi041 ^ w12405 ;
  assign w12407 = ( w12215 & w12286 ) | ( w12215 & ~w12294 ) | ( w12286 & ~w12294 ) ;
  assign w12408 = ~\pi103 & w4141 ;
  assign w12409 = \pi102 & w4334 ;
  assign w12410 = ( w4141 & ~w12408 ) | ( w4141 & w12409 ) | ( ~w12408 & w12409 ) ;
  assign w12411 = ~\pi104 & w4143 ;
  assign w12412 = w3740 | w12410 ;
  assign w12413 = ( w4144 & w12410 ) | ( w4144 & w12412 ) | ( w12410 & w12412 ) ;
  assign w12414 = ( w4143 & ~w12411 ) | ( w4143 & w12413 ) | ( ~w12411 & w12413 ) ;
  assign w12415 = \pi044 ^ w12414 ;
  assign w12416 = ( w12216 & ~w12276 ) | ( w12216 & w12284 ) | ( ~w12276 & w12284 ) ;
  assign w12417 = ~\pi094 & w5802 ;
  assign w12418 = \pi093 & w6052 ;
  assign w12419 = ( w5802 & ~w12417 ) | ( w5802 & w12418 ) | ( ~w12417 & w12418 ) ;
  assign w12420 = ~\pi095 & w5804 ;
  assign w12421 = w2409 | w12419 ;
  assign w12422 = ( w5805 & w12419 ) | ( w5805 & w12421 ) | ( w12419 & w12421 ) ;
  assign w12423 = ( w5804 & ~w12420 ) | ( w5804 & w12422 ) | ( ~w12420 & w12422 ) ;
  assign w12424 = \pi053 ^ w12423 ;
  assign w12425 = ( w12225 & ~w12241 ) | ( w12225 & w12249 ) | ( ~w12241 & w12249 ) ;
  assign w12426 = ~\pi088 & w7135 ;
  assign w12427 = \pi087 & w7359 ;
  assign w12428 = ( w7135 & ~w12426 ) | ( w7135 & w12427 ) | ( ~w12426 & w12427 ) ;
  assign w12429 = ~\pi089 & w7137 ;
  assign w12430 = w1595 | w12428 ;
  assign w12431 = ( w7138 & w12428 ) | ( w7138 & w12430 ) | ( w12428 & w12430 ) ;
  assign w12432 = ( w7137 & ~w12429 ) | ( w7137 & w12431 ) | ( ~w12429 & w12431 ) ;
  assign w12433 = \pi059 ^ w12432 ;
  assign w12434 = \pi062 ^ w11906 ;
  assign w12435 = ( \pi080 & \pi082 ) | ( \pi080 & w12434 ) | ( \pi082 & w12434 ) ;
  assign w12436 = ( ~\pi017 & \pi081 ) | ( ~\pi017 & w12435 ) | ( \pi081 & w12435 ) ;
  assign w12437 = w10655 & w12436 ;
  assign w12438 = ~\pi085 & w7811 ;
  assign w12439 = \pi084 & w8046 ;
  assign w12440 = ( w7811 & ~w12438 ) | ( w7811 & w12439 ) | ( ~w12438 & w12439 ) ;
  assign w12441 = ~\pi086 & w7813 ;
  assign w12442 = w1379 | w12440 ;
  assign w12443 = ( w7814 & w12440 ) | ( w7814 & w12442 ) | ( w12440 & w12442 ) ;
  assign w12444 = ( w7813 & ~w12441 ) | ( w7813 & w12443 ) | ( ~w12441 & w12443 ) ;
  assign w12445 = \pi062 ^ w12444 ;
  assign w12446 = w12437 ^ w12445 ;
  assign w12447 = ( \pi062 & \pi063 ) | ( \pi062 & \pi083 ) | ( \pi063 & \pi083 ) ;
  assign w12448 = \pi063 & ~\pi082 ;
  assign w12449 = \pi062 & w12448 ;
  assign w12450 = w12447 ^ w12449 ;
  assign w12451 = w12446 ^ w12450 ;
  assign w12452 = ( w12088 & w12233 ) | ( w12088 & ~w12239 ) | ( w12233 & ~w12239 ) ;
  assign w12453 = w12451 ^ w12452 ;
  assign w12454 = w12433 ^ w12453 ;
  assign w12455 = ~\pi091 & w6466 ;
  assign w12456 = \pi090 & w6702 ;
  assign w12457 = ( w6466 & ~w12455 ) | ( w6466 & w12456 ) | ( ~w12455 & w12456 ) ;
  assign w12458 = ~\pi092 & w6468 ;
  assign w12459 = w2033 | w12457 ;
  assign w12460 = ( w6469 & w12457 ) | ( w6469 & w12459 ) | ( w12457 & w12459 ) ;
  assign w12461 = ( w6468 & ~w12458 ) | ( w6468 & w12460 ) | ( ~w12458 & w12460 ) ;
  assign w12462 = \pi056 ^ w12461 ;
  assign w12463 = w12425 ^ w12454 ;
  assign w12464 = w12462 ^ w12463 ;
  assign w12465 = ( w12224 & ~w12251 ) | ( w12224 & w12252 ) | ( ~w12251 & w12252 ) ;
  assign w12466 = w12464 ^ w12465 ;
  assign w12467 = w12424 ^ w12466 ;
  assign w12468 = ( ~w12254 & w12262 ) | ( ~w12254 & w12263 ) | ( w12262 & w12263 ) ;
  assign w12469 = ~\pi097 & w5209 ;
  assign w12470 = \pi096 & w5433 ;
  assign w12471 = ( w5209 & ~w12469 ) | ( w5209 & w12470 ) | ( ~w12469 & w12470 ) ;
  assign w12472 = ~\pi098 & w5211 ;
  assign w12473 = w2824 | w12471 ;
  assign w12474 = ( w5212 & w12471 ) | ( w5212 & w12473 ) | ( w12471 & w12473 ) ;
  assign w12475 = ( w5211 & ~w12472 ) | ( w5211 & w12474 ) | ( ~w12472 & w12474 ) ;
  assign w12476 = \pi050 ^ w12475 ;
  assign w12477 = w12467 ^ w12468 ;
  assign w12478 = w12476 ^ w12477 ;
  assign w12479 = ( ~w12265 & w12273 ) | ( ~w12265 & w12274 ) | ( w12273 & w12274 ) ;
  assign w12480 = ~\pi100 & w4654 ;
  assign w12481 = \pi099 & w4876 ;
  assign w12482 = ( w4654 & ~w12480 ) | ( w4654 & w12481 ) | ( ~w12480 & w12481 ) ;
  assign w12483 = ~\pi101 & w4656 ;
  assign w12484 = w3264 | w12482 ;
  assign w12485 = ( w4657 & w12482 ) | ( w4657 & w12484 ) | ( w12482 & w12484 ) ;
  assign w12486 = ( w4656 & ~w12483 ) | ( w4656 & w12485 ) | ( ~w12483 & w12485 ) ;
  assign w12487 = \pi047 ^ w12486 ;
  assign w12488 = w12478 ^ w12479 ;
  assign w12489 = w12487 ^ w12488 ;
  assign w12490 = w12416 ^ w12489 ;
  assign w12491 = w12415 ^ w12490 ;
  assign w12492 = w12407 ^ w12491 ;
  assign w12493 = w12406 ^ w12492 ;
  assign w12494 = ( w12214 & w12296 ) | ( w12214 & w12304 ) | ( w12296 & w12304 ) ;
  assign w12495 = ~\pi109 & w3178 ;
  assign w12496 = \pi108 & w3340 ;
  assign w12497 = ( w3178 & ~w12495 ) | ( w3178 & w12496 ) | ( ~w12495 & w12496 ) ;
  assign w12498 = ~\pi110 & w3180 ;
  assign w12499 = w4792 | w12497 ;
  assign w12500 = ( w3181 & w12497 ) | ( w3181 & w12499 ) | ( w12497 & w12499 ) ;
  assign w12501 = ( w3180 & ~w12498 ) | ( w3180 & w12500 ) | ( ~w12498 & w12500 ) ;
  assign w12502 = \pi038 ^ w12501 ;
  assign w12503 = w12493 ^ w12494 ;
  assign w12504 = w12502 ^ w12503 ;
  assign w12505 = ( w12306 & w12314 ) | ( w12306 & w12315 ) | ( w12314 & w12315 ) ;
  assign w12506 = ~\pi112 & w2712 ;
  assign w12507 = \pi111 & w2872 ;
  assign w12508 = ( w2712 & ~w12506 ) | ( w2712 & w12507 ) | ( ~w12506 & w12507 ) ;
  assign w12509 = ~\pi113 & w2714 ;
  assign w12510 = w5366 | w12508 ;
  assign w12511 = ( w2715 & w12508 ) | ( w2715 & w12510 ) | ( w12508 & w12510 ) ;
  assign w12512 = ( w2714 & ~w12509 ) | ( w2714 & w12511 ) | ( ~w12509 & w12511 ) ;
  assign w12513 = \pi035 ^ w12512 ;
  assign w12514 = w12504 ^ w12505 ;
  assign w12515 = w12513 ^ w12514 ;
  assign w12516 = w12387 ^ w12515 ;
  assign w12517 = w12388 ^ w12516 ;
  assign w12518 = w12398 ^ w12517 ;
  assign w12519 = w12368 ^ w12518 ;
  assign w12520 = w12369 ^ w12519 ;
  assign w12521 = w12379 ^ w12520 ;
  assign w12522 = ( w12201 & w12203 ) | ( w12201 & w12352 ) | ( w12203 & w12352 ) ;
  assign w12523 = \pi127 & w1044 ;
  assign w12524 = ( \pi126 & ~w1047 ) | ( \pi126 & w8490 ) | ( ~w1047 & w8490 ) ;
  assign w12525 = \pi126 & ~w1138 ;
  assign w12526 = ( ~\pi126 & w12524 ) | ( ~\pi126 & w12525 ) | ( w12524 & w12525 ) ;
  assign w12527 = ( w9420 & w12523 ) | ( w9420 & ~w12526 ) | ( w12523 & ~w12526 ) ;
  assign w12528 = \pi020 ^ w12527 ;
  assign w12529 = w12522 ^ w12528 ;
  assign w12530 = w12521 ^ w12529 ;
  assign w12531 = w12359 ^ w12360 ;
  assign w12532 = w12530 ^ w12531 ;
  assign w12533 = ( w12359 & w12360 ) | ( w12359 & w12530 ) | ( w12360 & w12530 ) ;
  assign w12534 = ( w12521 & w12522 ) | ( w12521 & w12528 ) | ( w12522 & w12528 ) ;
  assign w12535 = w12379 ^ w12518 ;
  assign w12536 = ( w12368 & w12369 ) | ( w12368 & w12535 ) | ( w12369 & w12535 ) ;
  assign w12537 = w1047 & w8481 ;
  assign w12538 = w1138 | w12537 ;
  assign w12539 = ( \pi127 & w12537 ) | ( \pi127 & w12538 ) | ( w12537 & w12538 ) ;
  assign w12540 = \pi020 ^ w12539 ;
  assign w12541 = ~\pi125 & w1313 ;
  assign w12542 = \pi124 & w1417 ;
  assign w12543 = ( w1313 & ~w12541 ) | ( w1313 & w12542 ) | ( ~w12541 & w12542 ) ;
  assign w12544 = ~\pi126 & w1315 ;
  assign w12545 = w8231 | w12543 ;
  assign w12546 = ( w1316 & w12543 ) | ( w1316 & w12545 ) | ( w12543 & w12545 ) ;
  assign w12547 = ( w1315 & ~w12544 ) | ( w1315 & w12546 ) | ( ~w12544 & w12546 ) ;
  assign w12548 = \pi023 ^ w12547 ;
  assign w12549 = ( w12377 & w12378 ) | ( w12377 & w12518 ) | ( w12378 & w12518 ) ;
  assign w12550 = ~\pi122 & w1629 ;
  assign w12551 = \pi121 & w1722 ;
  assign w12552 = ( w1629 & ~w12550 ) | ( w1629 & w12551 ) | ( ~w12550 & w12551 ) ;
  assign w12553 = ~\pi123 & w1631 ;
  assign w12554 = w7516 | w12552 ;
  assign w12555 = ( w1632 & w12552 ) | ( w1632 & w12554 ) | ( w12552 & w12554 ) ;
  assign w12556 = ( w1631 & ~w12553 ) | ( w1631 & w12555 ) | ( ~w12553 & w12555 ) ;
  assign w12557 = \pi026 ^ w12556 ;
  assign w12558 = w12398 ^ w12515 ;
  assign w12559 = ( w12387 & w12388 ) | ( w12387 & w12558 ) | ( w12388 & w12558 ) ;
  assign w12560 = ~\pi119 & w1944 ;
  assign w12561 = \pi118 & w2072 ;
  assign w12562 = ( w1944 & ~w12560 ) | ( w1944 & w12561 ) | ( ~w12560 & w12561 ) ;
  assign w12563 = ~\pi120 & w1946 ;
  assign w12564 = w6634 | w12562 ;
  assign w12565 = ( w1947 & w12562 ) | ( w1947 & w12564 ) | ( w12562 & w12564 ) ;
  assign w12566 = ( w1946 & ~w12563 ) | ( w1946 & w12565 ) | ( ~w12563 & w12565 ) ;
  assign w12567 = \pi029 ^ w12566 ;
  assign w12568 = ( w12396 & w12397 ) | ( w12396 & w12515 ) | ( w12397 & w12515 ) ;
  assign w12569 = ~\pi116 & w2310 ;
  assign w12570 = \pi115 & w2443 ;
  assign w12571 = ( w2310 & ~w12569 ) | ( w2310 & w12570 ) | ( ~w12569 & w12570 ) ;
  assign w12572 = ~\pi117 & w2312 ;
  assign w12573 = w6185 | w12571 ;
  assign w12574 = ( w2313 & w12571 ) | ( w2313 & w12573 ) | ( w12571 & w12573 ) ;
  assign w12575 = ( w2312 & ~w12572 ) | ( w2312 & w12574 ) | ( ~w12572 & w12574 ) ;
  assign w12576 = \pi032 ^ w12575 ;
  assign w12577 = ( w12504 & w12505 ) | ( w12504 & w12513 ) | ( w12505 & w12513 ) ;
  assign w12578 = ( ~w12406 & w12407 ) | ( ~w12406 & w12491 ) | ( w12407 & w12491 ) ;
  assign w12579 = ~\pi107 & w3635 ;
  assign w12580 = \pi106 & w3817 ;
  assign w12581 = ( w3635 & ~w12579 ) | ( w3635 & w12580 ) | ( ~w12579 & w12580 ) ;
  assign w12582 = ~\pi108 & w3637 ;
  assign w12583 = w4425 | w12581 ;
  assign w12584 = ( w3638 & w12581 ) | ( w3638 & w12583 ) | ( w12581 & w12583 ) ;
  assign w12585 = ( w3637 & ~w12582 ) | ( w3637 & w12584 ) | ( ~w12582 & w12584 ) ;
  assign w12586 = \pi041 ^ w12585 ;
  assign w12587 = ( w12415 & w12416 ) | ( w12415 & ~w12489 ) | ( w12416 & ~w12489 ) ;
  assign w12588 = ~\pi104 & w4141 ;
  assign w12589 = \pi103 & w4334 ;
  assign w12590 = ( w4141 & ~w12588 ) | ( w4141 & w12589 ) | ( ~w12588 & w12589 ) ;
  assign w12591 = ~\pi105 & w4143 ;
  assign w12592 = w3905 | w12590 ;
  assign w12593 = ( w4144 & w12590 ) | ( w4144 & w12592 ) | ( w12590 & w12592 ) ;
  assign w12594 = ( w4143 & ~w12591 ) | ( w4143 & w12593 ) | ( ~w12591 & w12593 ) ;
  assign w12595 = \pi044 ^ w12594 ;
  assign w12596 = ( ~w12478 & w12479 ) | ( ~w12478 & w12487 ) | ( w12479 & w12487 ) ;
  assign w12597 = ~\pi101 & w4654 ;
  assign w12598 = \pi100 & w4876 ;
  assign w12599 = ( w4654 & ~w12597 ) | ( w4654 & w12598 ) | ( ~w12597 & w12598 ) ;
  assign w12600 = ~\pi102 & w4656 ;
  assign w12601 = w3284 | w12599 ;
  assign w12602 = ( w4657 & w12599 ) | ( w4657 & w12601 ) | ( w12599 & w12601 ) ;
  assign w12603 = ( w4656 & ~w12600 ) | ( w4656 & w12602 ) | ( ~w12600 & w12602 ) ;
  assign w12604 = \pi047 ^ w12603 ;
  assign w12605 = ( ~w12467 & w12468 ) | ( ~w12467 & w12476 ) | ( w12468 & w12476 ) ;
  assign w12606 = ~\pi098 & w5209 ;
  assign w12607 = \pi097 & w5433 ;
  assign w12608 = ( w5209 & ~w12606 ) | ( w5209 & w12607 ) | ( ~w12606 & w12607 ) ;
  assign w12609 = ~\pi099 & w5211 ;
  assign w12610 = w2966 | w12608 ;
  assign w12611 = ( w5212 & w12608 ) | ( w5212 & w12610 ) | ( w12608 & w12610 ) ;
  assign w12612 = ( w5211 & ~w12609 ) | ( w5211 & w12611 ) | ( ~w12609 & w12611 ) ;
  assign w12613 = \pi050 ^ w12612 ;
  assign w12614 = ( w12424 & ~w12464 ) | ( w12424 & w12465 ) | ( ~w12464 & w12465 ) ;
  assign w12615 = ( w12433 & ~w12451 ) | ( w12433 & w12452 ) | ( ~w12451 & w12452 ) ;
  assign w12616 = ~\pi089 & w7135 ;
  assign w12617 = \pi088 & w7359 ;
  assign w12618 = ( w7135 & ~w12616 ) | ( w7135 & w12617 ) | ( ~w12616 & w12617 ) ;
  assign w12619 = ~\pi090 & w7137 ;
  assign w12620 = w1801 | w12618 ;
  assign w12621 = ( w7138 & w12618 ) | ( w7138 & w12620 ) | ( w12618 & w12620 ) ;
  assign w12622 = ( w7137 & ~w12619 ) | ( w7137 & w12621 ) | ( ~w12619 & w12621 ) ;
  assign w12623 = \pi059 ^ w12622 ;
  assign w12624 = \pi063 & \pi082 ;
  assign w12625 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w12624 ) | ( \pi063 & w12624 ) ;
  assign w12626 = ( \pi062 & ~\pi063 ) | ( \pi062 & w12624 ) | ( ~\pi063 & w12624 ) ;
  assign w12627 = ( \pi083 & w12625 ) | ( \pi083 & w12626 ) | ( w12625 & w12626 ) ;
  assign w12628 = ( w12437 & w12445 ) | ( w12437 & ~w12627 ) | ( w12445 & ~w12627 ) ;
  assign w12629 = ~\pi086 & w7811 ;
  assign w12630 = \pi085 & w8046 ;
  assign w12631 = ( w7811 & ~w12629 ) | ( w7811 & w12630 ) | ( ~w12629 & w12630 ) ;
  assign w12632 = ~\pi087 & w7813 ;
  assign w12633 = ~w1477 & w7814 ;
  assign w12634 = ( w7814 & w12631 ) | ( w7814 & ~w12633 ) | ( w12631 & ~w12633 ) ;
  assign w12635 = ( w7813 & ~w12632 ) | ( w7813 & w12634 ) | ( ~w12632 & w12634 ) ;
  assign w12636 = ~\pi063 & \pi083 ;
  assign w12637 = ( \pi062 & ~w12448 ) | ( \pi062 & w12636 ) | ( ~w12448 & w12636 ) ;
  assign w12638 = w12635 ^ w12637 ;
  assign w12639 = \pi083 ^ w12638 ;
  assign w12640 = ( \pi063 & w12635 ) | ( \pi063 & ~w12636 ) | ( w12635 & ~w12636 ) ;
  assign w12641 = ( \pi062 & ~\pi063 ) | ( \pi062 & w12640 ) | ( ~\pi063 & w12640 ) ;
  assign w12642 = ( \pi062 & ~w12639 ) | ( \pi062 & w12641 ) | ( ~w12639 & w12641 ) ;
  assign w12643 = ( \pi063 & \pi084 ) | ( \pi063 & w12642 ) | ( \pi084 & w12642 ) ;
  assign w12644 = w12639 ^ w12643 ;
  assign w12645 = w12623 ^ w12628 ;
  assign w12646 = w12644 ^ w12645 ;
  assign w12647 = ~\pi092 & w6466 ;
  assign w12648 = \pi091 & w6702 ;
  assign w12649 = ( w6466 & ~w12647 ) | ( w6466 & w12648 ) | ( ~w12647 & w12648 ) ;
  assign w12650 = ~\pi093 & w6468 ;
  assign w12651 = w2155 | w12649 ;
  assign w12652 = ( w6469 & w12649 ) | ( w6469 & w12651 ) | ( w12649 & w12651 ) ;
  assign w12653 = ( w6468 & ~w12650 ) | ( w6468 & w12652 ) | ( ~w12650 & w12652 ) ;
  assign w12654 = \pi056 ^ w12653 ;
  assign w12655 = w12615 ^ w12646 ;
  assign w12656 = w12654 ^ w12655 ;
  assign w12657 = ( w12425 & ~w12454 ) | ( w12425 & w12462 ) | ( ~w12454 & w12462 ) ;
  assign w12658 = ~\pi095 & w5802 ;
  assign w12659 = \pi094 & w6052 ;
  assign w12660 = ( w5802 & ~w12658 ) | ( w5802 & w12659 ) | ( ~w12658 & w12659 ) ;
  assign w12661 = ~\pi096 & w5804 ;
  assign w12662 = w2546 | w12660 ;
  assign w12663 = ( w5805 & w12660 ) | ( w5805 & w12662 ) | ( w12660 & w12662 ) ;
  assign w12664 = ( w5804 & ~w12661 ) | ( w5804 & w12663 ) | ( ~w12661 & w12663 ) ;
  assign w12665 = \pi053 ^ w12664 ;
  assign w12666 = w12656 ^ w12657 ;
  assign w12667 = w12665 ^ w12666 ;
  assign w12668 = w12614 ^ w12667 ;
  assign w12669 = w12613 ^ w12668 ;
  assign w12670 = w12605 ^ w12669 ;
  assign w12671 = w12604 ^ w12670 ;
  assign w12672 = w12596 ^ w12671 ;
  assign w12673 = w12595 ^ w12672 ;
  assign w12674 = w12587 ^ w12673 ;
  assign w12675 = w12586 ^ w12674 ;
  assign w12676 = ~\pi110 & w3178 ;
  assign w12677 = \pi109 & w3340 ;
  assign w12678 = ( w3178 & ~w12676 ) | ( w3178 & w12677 ) | ( ~w12676 & w12677 ) ;
  assign w12679 = ~\pi111 & w3180 ;
  assign w12680 = w4811 | w12678 ;
  assign w12681 = ( w3181 & w12678 ) | ( w3181 & w12680 ) | ( w12678 & w12680 ) ;
  assign w12682 = ( w3180 & ~w12679 ) | ( w3180 & w12681 ) | ( ~w12679 & w12681 ) ;
  assign w12683 = \pi038 ^ w12682 ;
  assign w12684 = w12578 ^ w12675 ;
  assign w12685 = w12683 ^ w12684 ;
  assign w12686 = ( w12493 & w12494 ) | ( w12493 & w12502 ) | ( w12494 & w12502 ) ;
  assign w12687 = w12685 ^ w12686 ;
  assign w12688 = ~\pi113 & w2712 ;
  assign w12689 = \pi112 & w2872 ;
  assign w12690 = ( w2712 & ~w12688 ) | ( w2712 & w12689 ) | ( ~w12688 & w12689 ) ;
  assign w12691 = ~\pi114 & w2714 ;
  assign w12692 = w5565 | w12690 ;
  assign w12693 = ( w2715 & w12690 ) | ( w2715 & w12692 ) | ( w12690 & w12692 ) ;
  assign w12694 = ( w2714 & ~w12691 ) | ( w2714 & w12693 ) | ( ~w12691 & w12693 ) ;
  assign w12695 = \pi035 ^ w12694 ;
  assign w12696 = w12576 ^ w12695 ;
  assign w12697 = w12577 ^ w12696 ;
  assign w12698 = w12687 ^ w12697 ;
  assign w12699 = w12568 ^ w12698 ;
  assign w12700 = w12567 ^ w12699 ;
  assign w12701 = w12559 ^ w12700 ;
  assign w12702 = w12557 ^ w12701 ;
  assign w12703 = w12548 ^ w12549 ;
  assign w12704 = w12702 ^ w12703 ;
  assign w12705 = w12536 ^ w12704 ;
  assign w12706 = w12540 ^ w12705 ;
  assign w12707 = w12533 ^ w12534 ;
  assign w12708 = w12706 ^ w12707 ;
  assign w12709 = ( w12548 & w12549 ) | ( w12548 & w12702 ) | ( w12549 & w12702 ) ;
  assign w12710 = ~\pi126 & w1313 ;
  assign w12711 = \pi125 & w1417 ;
  assign w12712 = ( w1313 & ~w12710 ) | ( w1313 & w12711 ) | ( ~w12710 & w12711 ) ;
  assign w12713 = ~\pi127 & w1315 ;
  assign w12714 = w8466 | w12712 ;
  assign w12715 = ( w1316 & w12712 ) | ( w1316 & w12714 ) | ( w12712 & w12714 ) ;
  assign w12716 = ( w1315 & ~w12713 ) | ( w1315 & w12715 ) | ( ~w12713 & w12715 ) ;
  assign w12717 = \pi023 ^ w12716 ;
  assign w12718 = ~\pi123 & w1629 ;
  assign w12719 = \pi122 & w1722 ;
  assign w12720 = ( w1629 & ~w12718 ) | ( w1629 & w12719 ) | ( ~w12718 & w12719 ) ;
  assign w12721 = ~\pi124 & w1631 ;
  assign w12722 = w7538 | w12720 ;
  assign w12723 = ( w1632 & w12720 ) | ( w1632 & w12722 ) | ( w12720 & w12722 ) ;
  assign w12724 = ( w1631 & ~w12721 ) | ( w1631 & w12723 ) | ( ~w12721 & w12723 ) ;
  assign w12725 = \pi026 ^ w12724 ;
  assign w12726 = ( w12557 & w12559 ) | ( w12557 & w12700 ) | ( w12559 & w12700 ) ;
  assign w12727 = w12725 ^ w12726 ;
  assign w12728 = ( w12567 & w12568 ) | ( w12567 & w12698 ) | ( w12568 & w12698 ) ;
  assign w12729 = ~\pi120 & w1944 ;
  assign w12730 = \pi119 & w2072 ;
  assign w12731 = ( w1944 & ~w12729 ) | ( w1944 & w12730 ) | ( ~w12729 & w12730 ) ;
  assign w12732 = ~\pi121 & w1946 ;
  assign w12733 = w7050 | w12731 ;
  assign w12734 = ( w1947 & w12731 ) | ( w1947 & w12733 ) | ( w12731 & w12733 ) ;
  assign w12735 = ( w1946 & ~w12732 ) | ( w1946 & w12734 ) | ( ~w12732 & w12734 ) ;
  assign w12736 = \pi029 ^ w12735 ;
  assign w12737 = ~\pi117 & w2310 ;
  assign w12738 = \pi116 & w2443 ;
  assign w12739 = ( w2310 & ~w12737 ) | ( w2310 & w12738 ) | ( ~w12737 & w12738 ) ;
  assign w12740 = ~\pi118 & w2312 ;
  assign w12741 = w6206 | w12739 ;
  assign w12742 = ( w2313 & w12739 ) | ( w2313 & w12741 ) | ( w12739 & w12741 ) ;
  assign w12743 = ( w2312 & ~w12740 ) | ( w2312 & w12742 ) | ( ~w12740 & w12742 ) ;
  assign w12744 = \pi032 ^ w12743 ;
  assign w12745 = w12687 ^ w12695 ;
  assign w12746 = ( w12576 & w12577 ) | ( w12576 & w12745 ) | ( w12577 & w12745 ) ;
  assign w12747 = w12744 ^ w12746 ;
  assign w12748 = ( w12685 & w12686 ) | ( w12685 & w12695 ) | ( w12686 & w12695 ) ;
  assign w12749 = ( w12613 & w12614 ) | ( w12613 & ~w12667 ) | ( w12614 & ~w12667 ) ;
  assign w12750 = \pi083 ^ \pi085 ;
  assign w12751 = ( \pi062 & \pi063 ) | ( \pi062 & ~w12750 ) | ( \pi063 & ~w12750 ) ;
  assign w12752 = \pi083 ^ \pi084 ;
  assign w12753 = \pi062 & ~w12752 ;
  assign w12754 = ( \pi063 & ~w12752 ) | ( \pi063 & w12753 ) | ( ~w12752 & w12753 ) ;
  assign w12755 = \pi020 ^ w12754 ;
  assign w12756 = w12751 ^ w12755 ;
  assign w12757 = ~\pi087 & w7811 ;
  assign w12758 = \pi086 & w8046 ;
  assign w12759 = ( w7811 & ~w12757 ) | ( w7811 & w12758 ) | ( ~w12757 & w12758 ) ;
  assign w12760 = ~\pi088 & w7813 ;
  assign w12761 = w1574 | w12759 ;
  assign w12762 = ( w7814 & w12759 ) | ( w7814 & w12761 ) | ( w12759 & w12761 ) ;
  assign w12763 = ( w7813 & ~w12760 ) | ( w7813 & w12762 ) | ( ~w12760 & w12762 ) ;
  assign w12764 = \pi062 ^ w12763 ;
  assign w12765 = \pi063 ^ w12635 ;
  assign w12766 = ( ~\pi083 & \pi084 ) | ( ~\pi083 & w12765 ) | ( \pi084 & w12765 ) ;
  assign w12767 = w8323 ^ w12766 ;
  assign w12768 = ( \pi082 & \pi083 ) | ( \pi082 & w12635 ) | ( \pi083 & w12635 ) ;
  assign w12769 = ( ~\pi083 & w12765 ) | ( ~\pi083 & w12768 ) | ( w12765 & w12768 ) ;
  assign w12770 = ( ~w12766 & w12767 ) | ( ~w12766 & w12769 ) | ( w12767 & w12769 ) ;
  assign w12771 = w12764 ^ w12770 ;
  assign w12772 = w12756 ^ w12771 ;
  assign w12773 = ~\pi090 & w7135 ;
  assign w12774 = \pi089 & w7359 ;
  assign w12775 = ( w7135 & ~w12773 ) | ( w7135 & w12774 ) | ( ~w12773 & w12774 ) ;
  assign w12776 = ~\pi091 & w7137 ;
  assign w12777 = w1908 | w12775 ;
  assign w12778 = ( w7138 & w12775 ) | ( w7138 & w12777 ) | ( w12775 & w12777 ) ;
  assign w12779 = ( w7137 & ~w12776 ) | ( w7137 & w12778 ) | ( ~w12776 & w12778 ) ;
  assign w12780 = \pi059 ^ w12779 ;
  assign w12781 = ( w12623 & w12628 ) | ( w12623 & ~w12644 ) | ( w12628 & ~w12644 ) ;
  assign w12782 = w12772 ^ w12781 ;
  assign w12783 = w12780 ^ w12782 ;
  assign w12784 = ~\pi093 & w6466 ;
  assign w12785 = \pi092 & w6702 ;
  assign w12786 = ( w6466 & ~w12784 ) | ( w6466 & w12785 ) | ( ~w12784 & w12785 ) ;
  assign w12787 = ~\pi094 & w6468 ;
  assign w12788 = w2274 | w12786 ;
  assign w12789 = ( w6469 & w12786 ) | ( w6469 & w12788 ) | ( w12786 & w12788 ) ;
  assign w12790 = ( w6468 & ~w12787 ) | ( w6468 & w12789 ) | ( ~w12787 & w12789 ) ;
  assign w12791 = \pi056 ^ w12790 ;
  assign w12792 = ( w12615 & ~w12646 ) | ( w12615 & w12654 ) | ( ~w12646 & w12654 ) ;
  assign w12793 = w12783 ^ w12792 ;
  assign w12794 = w12791 ^ w12793 ;
  assign w12795 = ~\pi096 & w5802 ;
  assign w12796 = \pi095 & w6052 ;
  assign w12797 = ( w5802 & ~w12795 ) | ( w5802 & w12796 ) | ( ~w12795 & w12796 ) ;
  assign w12798 = ~\pi097 & w5804 ;
  assign w12799 = w2673 | w12797 ;
  assign w12800 = ( w5805 & w12797 ) | ( w5805 & w12799 ) | ( w12797 & w12799 ) ;
  assign w12801 = ( w5804 & ~w12798 ) | ( w5804 & w12800 ) | ( ~w12798 & w12800 ) ;
  assign w12802 = \pi053 ^ w12801 ;
  assign w12803 = ( ~w12656 & w12657 ) | ( ~w12656 & w12665 ) | ( w12657 & w12665 ) ;
  assign w12804 = w12794 ^ w12803 ;
  assign w12805 = w12802 ^ w12804 ;
  assign w12806 = ~\pi099 & w5209 ;
  assign w12807 = \pi098 & w5433 ;
  assign w12808 = ( w5209 & ~w12806 ) | ( w5209 & w12807 ) | ( ~w12806 & w12807 ) ;
  assign w12809 = ~\pi100 & w5211 ;
  assign w12810 = w3104 | w12808 ;
  assign w12811 = ( w5212 & w12808 ) | ( w5212 & w12810 ) | ( w12808 & w12810 ) ;
  assign w12812 = ( w5211 & ~w12809 ) | ( w5211 & w12811 ) | ( ~w12809 & w12811 ) ;
  assign w12813 = \pi050 ^ w12812 ;
  assign w12814 = w12749 ^ w12805 ;
  assign w12815 = w12813 ^ w12814 ;
  assign w12816 = ~\pi102 & w4654 ;
  assign w12817 = \pi101 & w4876 ;
  assign w12818 = ( w4654 & ~w12816 ) | ( w4654 & w12817 ) | ( ~w12816 & w12817 ) ;
  assign w12819 = ~\pi103 & w4656 ;
  assign w12820 = w3437 | w12818 ;
  assign w12821 = ( w4657 & w12818 ) | ( w4657 & w12820 ) | ( w12818 & w12820 ) ;
  assign w12822 = ( w4656 & ~w12819 ) | ( w4656 & w12821 ) | ( ~w12819 & w12821 ) ;
  assign w12823 = \pi047 ^ w12822 ;
  assign w12824 = ( w12604 & w12605 ) | ( w12604 & ~w12669 ) | ( w12605 & ~w12669 ) ;
  assign w12825 = w12815 ^ w12824 ;
  assign w12826 = w12823 ^ w12825 ;
  assign w12827 = ~\pi105 & w4141 ;
  assign w12828 = \pi104 & w4334 ;
  assign w12829 = ( w4141 & ~w12827 ) | ( w4141 & w12828 ) | ( ~w12827 & w12828 ) ;
  assign w12830 = ~\pi106 & w4143 ;
  assign w12831 = w4068 | w12829 ;
  assign w12832 = ( w4144 & w12829 ) | ( w4144 & w12831 ) | ( w12829 & w12831 ) ;
  assign w12833 = ( w4143 & ~w12830 ) | ( w4143 & w12832 ) | ( ~w12830 & w12832 ) ;
  assign w12834 = \pi044 ^ w12833 ;
  assign w12835 = ( w12595 & w12596 ) | ( w12595 & ~w12671 ) | ( w12596 & ~w12671 ) ;
  assign w12836 = w12826 ^ w12835 ;
  assign w12837 = w12834 ^ w12836 ;
  assign w12838 = ~\pi108 & w3635 ;
  assign w12839 = \pi107 & w3817 ;
  assign w12840 = ( w3635 & ~w12838 ) | ( w3635 & w12839 ) | ( ~w12838 & w12839 ) ;
  assign w12841 = ~\pi109 & w3637 ;
  assign w12842 = w4599 | w12840 ;
  assign w12843 = ( w3638 & w12840 ) | ( w3638 & w12842 ) | ( w12840 & w12842 ) ;
  assign w12844 = ( w3637 & ~w12841 ) | ( w3637 & w12843 ) | ( ~w12841 & w12843 ) ;
  assign w12845 = \pi041 ^ w12844 ;
  assign w12846 = ( w12586 & w12587 ) | ( w12586 & ~w12673 ) | ( w12587 & ~w12673 ) ;
  assign w12847 = w12837 ^ w12846 ;
  assign w12848 = w12845 ^ w12847 ;
  assign w12849 = ~\pi111 & w3178 ;
  assign w12850 = \pi110 & w3340 ;
  assign w12851 = ( w3178 & ~w12849 ) | ( w3178 & w12850 ) | ( ~w12849 & w12850 ) ;
  assign w12852 = ~\pi112 & w3180 ;
  assign w12853 = w4999 | w12851 ;
  assign w12854 = ( w3181 & w12851 ) | ( w3181 & w12853 ) | ( w12851 & w12853 ) ;
  assign w12855 = ( w3180 & ~w12852 ) | ( w3180 & w12854 ) | ( ~w12852 & w12854 ) ;
  assign w12856 = \pi038 ^ w12855 ;
  assign w12857 = ( w12578 & w12675 ) | ( w12578 & ~w12683 ) | ( w12675 & ~w12683 ) ;
  assign w12858 = w12848 ^ w12857 ;
  assign w12859 = w12856 ^ w12858 ;
  assign w12860 = ~\pi114 & w2712 ;
  assign w12861 = \pi113 & w2872 ;
  assign w12862 = ( w2712 & ~w12860 ) | ( w2712 & w12861 ) | ( ~w12860 & w12861 ) ;
  assign w12863 = ~\pi115 & w2714 ;
  assign w12864 = w5585 | w12862 ;
  assign w12865 = ( w2715 & w12862 ) | ( w2715 & w12864 ) | ( w12862 & w12864 ) ;
  assign w12866 = ( w2714 & ~w12863 ) | ( w2714 & w12865 ) | ( ~w12863 & w12865 ) ;
  assign w12867 = \pi035 ^ w12866 ;
  assign w12868 = ( w12748 & w12859 ) | ( w12748 & w12867 ) | ( w12859 & w12867 ) ;
  assign w12869 = w12748 ^ w12859 ;
  assign w12870 = w12867 ^ w12869 ;
  assign w12871 = w12736 ^ w12870 ;
  assign w12872 = w12728 ^ w12871 ;
  assign w12873 = w12747 ^ w12872 ;
  assign w12874 = w12727 ^ w12873 ;
  assign w12875 = w12709 ^ w12874 ;
  assign w12876 = w12717 ^ w12875 ;
  assign w12877 = ( w12536 & w12540 ) | ( w12536 & w12704 ) | ( w12540 & w12704 ) ;
  assign w12878 = ( w12533 & w12534 ) | ( w12533 & w12706 ) | ( w12534 & w12706 ) ;
  assign w12879 = w12877 ^ w12878 ;
  assign w12880 = w12876 ^ w12879 ;
  assign w12881 = ( w12725 & w12726 ) | ( w12725 & w12873 ) | ( w12726 & w12873 ) ;
  assign w12882 = \pi127 & w1313 ;
  assign w12883 = ( \pi126 & ~w1316 ) | ( \pi126 & w8490 ) | ( ~w1316 & w8490 ) ;
  assign w12884 = \pi126 & ~w1417 ;
  assign w12885 = ( ~\pi126 & w12883 ) | ( ~\pi126 & w12884 ) | ( w12883 & w12884 ) ;
  assign w12886 = ( w9420 & w12882 ) | ( w9420 & ~w12885 ) | ( w12882 & ~w12885 ) ;
  assign w12887 = ~\pi124 & w1629 ;
  assign w12888 = \pi123 & w1722 ;
  assign w12889 = ( w1629 & ~w12887 ) | ( w1629 & w12888 ) | ( ~w12887 & w12888 ) ;
  assign w12890 = ~\pi125 & w1631 ;
  assign w12891 = w7988 | w12889 ;
  assign w12892 = ( w1632 & w12889 ) | ( w1632 & w12891 ) | ( w12889 & w12891 ) ;
  assign w12893 = ( w1631 & ~w12890 ) | ( w1631 & w12892 ) | ( ~w12890 & w12892 ) ;
  assign w12894 = \pi026 ^ w12893 ;
  assign w12895 = w12747 ^ w12870 ;
  assign w12896 = ( w12728 & w12736 ) | ( w12728 & w12895 ) | ( w12736 & w12895 ) ;
  assign w12897 = w12894 ^ w12896 ;
  assign w12898 = ( w12744 & w12746 ) | ( w12744 & w12870 ) | ( w12746 & w12870 ) ;
  assign w12899 = \pi120 & w2072 ;
  assign w12900 = ( \pi122 & w1946 ) | ( \pi122 & w12899 ) | ( w1946 & w12899 ) ;
  assign w12901 = \pi121 | w12900 ;
  assign w12902 = ( w1944 & w12900 ) | ( w1944 & w12901 ) | ( w12900 & w12901 ) ;
  assign w12903 = w12899 | w12902 ;
  assign w12904 = ~w1947 & w7069 ;
  assign w12905 = ( w7069 & w12903 ) | ( w7069 & ~w12904 ) | ( w12903 & ~w12904 ) ;
  assign w12906 = \pi029 ^ w12905 ;
  assign w12907 = ~\pi118 & w2310 ;
  assign w12908 = \pi117 & w2443 ;
  assign w12909 = ( w2310 & ~w12907 ) | ( w2310 & w12908 ) | ( ~w12907 & w12908 ) ;
  assign w12910 = ~\pi119 & w2312 ;
  assign w12911 = w6616 | w12909 ;
  assign w12912 = ( w2313 & w12909 ) | ( w2313 & w12911 ) | ( w12909 & w12911 ) ;
  assign w12913 = ( w2312 & ~w12910 ) | ( w2312 & w12912 ) | ( ~w12910 & w12912 ) ;
  assign w12914 = \pi032 ^ w12913 ;
  assign w12915 = w12868 ^ w12914 ;
  assign w12916 = ~\pi106 & w4141 ;
  assign w12917 = \pi105 & w4334 ;
  assign w12918 = ( w4141 & ~w12916 ) | ( w4141 & w12917 ) | ( ~w12916 & w12917 ) ;
  assign w12919 = ~\pi107 & w4143 ;
  assign w12920 = w4087 | w12918 ;
  assign w12921 = ( w4144 & w12918 ) | ( w4144 & w12920 ) | ( w12918 & w12920 ) ;
  assign w12922 = ( w4143 & ~w12919 ) | ( w4143 & w12921 ) | ( ~w12919 & w12921 ) ;
  assign w12923 = \pi044 ^ w12922 ;
  assign w12924 = ( ~w12815 & w12823 ) | ( ~w12815 & w12824 ) | ( w12823 & w12824 ) ;
  assign w12925 = ~\pi103 & w4654 ;
  assign w12926 = \pi102 & w4876 ;
  assign w12927 = ( w4654 & ~w12925 ) | ( w4654 & w12926 ) | ( ~w12925 & w12926 ) ;
  assign w12928 = ~\pi104 & w4656 ;
  assign w12929 = w3740 | w12927 ;
  assign w12930 = ( w4657 & w12927 ) | ( w4657 & w12929 ) | ( w12927 & w12929 ) ;
  assign w12931 = ( w4656 & ~w12928 ) | ( w4656 & w12930 ) | ( ~w12928 & w12930 ) ;
  assign w12932 = \pi047 ^ w12931 ;
  assign w12933 = ( w12749 & ~w12805 ) | ( w12749 & w12813 ) | ( ~w12805 & w12813 ) ;
  assign w12934 = ( ~w12772 & w12780 ) | ( ~w12772 & w12781 ) | ( w12780 & w12781 ) ;
  assign w12935 = ~\pi091 & w7135 ;
  assign w12936 = \pi090 & w7359 ;
  assign w12937 = ( w7135 & ~w12935 ) | ( w7135 & w12936 ) | ( ~w12935 & w12936 ) ;
  assign w12938 = ~\pi092 & w7137 ;
  assign w12939 = w2033 | w12937 ;
  assign w12940 = ( w7138 & w12937 ) | ( w7138 & w12939 ) | ( w12937 & w12939 ) ;
  assign w12941 = ( w7137 & ~w12938 ) | ( w7137 & w12940 ) | ( ~w12938 & w12940 ) ;
  assign w12942 = \pi059 ^ w12941 ;
  assign w12943 = ( ~w12756 & w12764 ) | ( ~w12756 & w12770 ) | ( w12764 & w12770 ) ;
  assign w12944 = \pi063 ^ \pi083 ;
  assign w12945 = \pi062 ^ w12944 ;
  assign w12946 = ( \pi083 & \pi085 ) | ( \pi083 & w12945 ) | ( \pi085 & w12945 ) ;
  assign w12947 = ( ~\pi020 & \pi084 ) | ( ~\pi020 & w12946 ) | ( \pi084 & w12946 ) ;
  assign w12948 = w10655 & w12947 ;
  assign w12949 = ~\pi088 & w7811 ;
  assign w12950 = \pi087 & w8046 ;
  assign w12951 = ( w7811 & ~w12949 ) | ( w7811 & w12950 ) | ( ~w12949 & w12950 ) ;
  assign w12952 = ~\pi089 & w7813 ;
  assign w12953 = ~w1595 & w7814 ;
  assign w12954 = ( w7814 & w12951 ) | ( w7814 & ~w12953 ) | ( w12951 & ~w12953 ) ;
  assign w12955 = ( w7813 & ~w12952 ) | ( w7813 & w12954 ) | ( ~w12952 & w12954 ) ;
  assign w12956 = w12948 ^ w12955 ;
  assign w12957 = \pi062 ^ \pi086 ;
  assign w12958 = \pi063 ^ \pi086 ;
  assign w12959 = \pi062 & ~\pi085 ;
  assign w12960 = ( w12957 & ~w12958 ) | ( w12957 & w12959 ) | ( ~w12958 & w12959 ) ;
  assign w12961 = w12956 ^ w12960 ;
  assign w12962 = w12942 ^ w12943 ;
  assign w12963 = w12961 ^ w12962 ;
  assign w12964 = ~\pi094 & w6466 ;
  assign w12965 = \pi093 & w6702 ;
  assign w12966 = ( w6466 & ~w12964 ) | ( w6466 & w12965 ) | ( ~w12964 & w12965 ) ;
  assign w12967 = ~\pi095 & w6468 ;
  assign w12968 = w2409 | w12966 ;
  assign w12969 = ( w6469 & w12966 ) | ( w6469 & w12968 ) | ( w12966 & w12968 ) ;
  assign w12970 = ( w6468 & ~w12967 ) | ( w6468 & w12969 ) | ( ~w12967 & w12969 ) ;
  assign w12971 = \pi056 ^ w12970 ;
  assign w12972 = w12934 ^ w12963 ;
  assign w12973 = w12971 ^ w12972 ;
  assign w12974 = ( ~w12783 & w12791 ) | ( ~w12783 & w12792 ) | ( w12791 & w12792 ) ;
  assign w12975 = ~\pi097 & w5802 ;
  assign w12976 = \pi096 & w6052 ;
  assign w12977 = ( w5802 & ~w12975 ) | ( w5802 & w12976 ) | ( ~w12975 & w12976 ) ;
  assign w12978 = ~\pi098 & w5804 ;
  assign w12979 = w2824 | w12977 ;
  assign w12980 = ( w5805 & w12977 ) | ( w5805 & w12979 ) | ( w12977 & w12979 ) ;
  assign w12981 = ( w5804 & ~w12978 ) | ( w5804 & w12980 ) | ( ~w12978 & w12980 ) ;
  assign w12982 = \pi053 ^ w12981 ;
  assign w12983 = w12973 ^ w12974 ;
  assign w12984 = w12982 ^ w12983 ;
  assign w12985 = ( ~w12794 & w12802 ) | ( ~w12794 & w12803 ) | ( w12802 & w12803 ) ;
  assign w12986 = ~\pi100 & w5209 ;
  assign w12987 = \pi099 & w5433 ;
  assign w12988 = ( w5209 & ~w12986 ) | ( w5209 & w12987 ) | ( ~w12986 & w12987 ) ;
  assign w12989 = ~\pi101 & w5211 ;
  assign w12990 = w3264 | w12988 ;
  assign w12991 = ( w5212 & w12988 ) | ( w5212 & w12990 ) | ( w12988 & w12990 ) ;
  assign w12992 = ( w5211 & ~w12989 ) | ( w5211 & w12991 ) | ( ~w12989 & w12991 ) ;
  assign w12993 = \pi050 ^ w12992 ;
  assign w12994 = w12984 ^ w12985 ;
  assign w12995 = w12993 ^ w12994 ;
  assign w12996 = w12933 ^ w12995 ;
  assign w12997 = w12932 ^ w12996 ;
  assign w12998 = w12924 ^ w12997 ;
  assign w12999 = w12923 ^ w12998 ;
  assign w13000 = ( ~w12826 & w12834 ) | ( ~w12826 & w12835 ) | ( w12834 & w12835 ) ;
  assign w13001 = ~\pi109 & w3635 ;
  assign w13002 = \pi108 & w3817 ;
  assign w13003 = ( w3635 & ~w13001 ) | ( w3635 & w13002 ) | ( ~w13001 & w13002 ) ;
  assign w13004 = ~\pi110 & w3637 ;
  assign w13005 = w4792 | w13003 ;
  assign w13006 = ( w3638 & w13003 ) | ( w3638 & w13005 ) | ( w13003 & w13005 ) ;
  assign w13007 = ( w3637 & ~w13004 ) | ( w3637 & w13006 ) | ( ~w13004 & w13006 ) ;
  assign w13008 = \pi041 ^ w13007 ;
  assign w13009 = w12999 ^ w13000 ;
  assign w13010 = w13008 ^ w13009 ;
  assign w13011 = ( ~w12837 & w12845 ) | ( ~w12837 & w12846 ) | ( w12845 & w12846 ) ;
  assign w13012 = ~\pi112 & w3178 ;
  assign w13013 = \pi111 & w3340 ;
  assign w13014 = ( w3178 & ~w13012 ) | ( w3178 & w13013 ) | ( ~w13012 & w13013 ) ;
  assign w13015 = ~\pi113 & w3180 ;
  assign w13016 = w5366 | w13014 ;
  assign w13017 = ( w3181 & w13014 ) | ( w3181 & w13016 ) | ( w13014 & w13016 ) ;
  assign w13018 = ( w3180 & ~w13015 ) | ( w3180 & w13017 ) | ( ~w13015 & w13017 ) ;
  assign w13019 = \pi038 ^ w13018 ;
  assign w13020 = w13010 ^ w13011 ;
  assign w13021 = w13019 ^ w13020 ;
  assign w13022 = ( w12848 & ~w12856 ) | ( w12848 & w12857 ) | ( ~w12856 & w12857 ) ;
  assign w13023 = ~\pi115 & w2712 ;
  assign w13024 = \pi114 & w2872 ;
  assign w13025 = ( w2712 & ~w13023 ) | ( w2712 & w13024 ) | ( ~w13023 & w13024 ) ;
  assign w13026 = ~\pi116 & w2714 ;
  assign w13027 = w5976 | w13025 ;
  assign w13028 = ( w2715 & w13025 ) | ( w2715 & w13027 ) | ( w13025 & w13027 ) ;
  assign w13029 = ( w2714 & ~w13026 ) | ( w2714 & w13028 ) | ( ~w13026 & w13028 ) ;
  assign w13030 = \pi035 ^ w13029 ;
  assign w13031 = w13021 ^ w13022 ;
  assign w13032 = w13030 ^ w13031 ;
  assign w13033 = w12906 ^ w13032 ;
  assign w13034 = w12898 ^ w13033 ;
  assign w13035 = w12915 ^ w13034 ;
  assign w13036 = w12886 ^ w12897 ;
  assign w13037 = w12881 ^ w13035 ;
  assign w13038 = \pi023 ^ w13037 ;
  assign w13039 = w13036 ^ w13038 ;
  assign w13040 = ( w12709 & w12717 ) | ( w12709 & w12874 ) | ( w12717 & w12874 ) ;
  assign w13041 = ( w12876 & w12877 ) | ( w12876 & w12878 ) | ( w12877 & w12878 ) ;
  assign w13042 = w13040 ^ w13041 ;
  assign w13043 = w13039 ^ w13042 ;
  assign w13044 = ( w13039 & w13040 ) | ( w13039 & w13041 ) | ( w13040 & w13041 ) ;
  assign w13045 = w12897 ^ w13035 ;
  assign w13046 = \pi023 ^ w12886 ;
  assign w13047 = ( w12881 & w13045 ) | ( w12881 & w13046 ) | ( w13045 & w13046 ) ;
  assign w13048 = ( w12894 & w12896 ) | ( w12894 & w13035 ) | ( w12896 & w13035 ) ;
  assign w13049 = w1316 & w8481 ;
  assign w13050 = w1417 | w13049 ;
  assign w13051 = ( \pi127 & w13049 ) | ( \pi127 & w13050 ) | ( w13049 & w13050 ) ;
  assign w13052 = \pi023 ^ w13051 ;
  assign w13053 = ~\pi125 & w1629 ;
  assign w13054 = \pi124 & w1722 ;
  assign w13055 = ( w1629 & ~w13053 ) | ( w1629 & w13054 ) | ( ~w13053 & w13054 ) ;
  assign w13056 = ~\pi126 & w1631 ;
  assign w13057 = w8231 | w13055 ;
  assign w13058 = ( w1632 & w13055 ) | ( w1632 & w13057 ) | ( w13055 & w13057 ) ;
  assign w13059 = ( w1631 & ~w13056 ) | ( w1631 & w13058 ) | ( ~w13056 & w13058 ) ;
  assign w13060 = \pi026 ^ w13059 ;
  assign w13061 = w12915 ^ w13032 ;
  assign w13062 = ( w12898 & w12906 ) | ( w12898 & w13061 ) | ( w12906 & w13061 ) ;
  assign w13063 = ~\pi122 & w1944 ;
  assign w13064 = \pi121 & w2072 ;
  assign w13065 = ( w1944 & ~w13063 ) | ( w1944 & w13064 ) | ( ~w13063 & w13064 ) ;
  assign w13066 = ~\pi123 & w1946 ;
  assign w13067 = w7516 | w13065 ;
  assign w13068 = ( w1947 & w13065 ) | ( w1947 & w13067 ) | ( w13065 & w13067 ) ;
  assign w13069 = ( w1946 & ~w13066 ) | ( w1946 & w13068 ) | ( ~w13066 & w13068 ) ;
  assign w13070 = \pi029 ^ w13069 ;
  assign w13071 = ( w12868 & w12914 ) | ( w12868 & w13032 ) | ( w12914 & w13032 ) ;
  assign w13072 = ~\pi119 & w2310 ;
  assign w13073 = \pi118 & w2443 ;
  assign w13074 = ( w2310 & ~w13072 ) | ( w2310 & w13073 ) | ( ~w13072 & w13073 ) ;
  assign w13075 = ~\pi120 & w2312 ;
  assign w13076 = w6634 | w13074 ;
  assign w13077 = ( w2313 & w13074 ) | ( w2313 & w13076 ) | ( w13074 & w13076 ) ;
  assign w13078 = ( w2312 & ~w13075 ) | ( w2312 & w13077 ) | ( ~w13075 & w13077 ) ;
  assign w13079 = \pi032 ^ w13078 ;
  assign w13080 = ( w13021 & w13022 ) | ( w13021 & ~w13030 ) | ( w13022 & ~w13030 ) ;
  assign w13081 = ~\pi116 & w2712 ;
  assign w13082 = \pi115 & w2872 ;
  assign w13083 = ( w2712 & ~w13081 ) | ( w2712 & w13082 ) | ( ~w13081 & w13082 ) ;
  assign w13084 = ~\pi117 & w2714 ;
  assign w13085 = w6185 | w13083 ;
  assign w13086 = ( w2715 & w13083 ) | ( w2715 & w13085 ) | ( w13083 & w13085 ) ;
  assign w13087 = ( w2714 & ~w13084 ) | ( w2714 & w13086 ) | ( ~w13084 & w13086 ) ;
  assign w13088 = \pi035 ^ w13087 ;
  assign w13089 = ( ~w13010 & w13011 ) | ( ~w13010 & w13019 ) | ( w13011 & w13019 ) ;
  assign w13090 = ( w12923 & w12924 ) | ( w12923 & ~w12997 ) | ( w12924 & ~w12997 ) ;
  assign w13091 = ~\pi107 & w4141 ;
  assign w13092 = \pi106 & w4334 ;
  assign w13093 = ( w4141 & ~w13091 ) | ( w4141 & w13092 ) | ( ~w13091 & w13092 ) ;
  assign w13094 = ~\pi108 & w4143 ;
  assign w13095 = w4425 | w13093 ;
  assign w13096 = ( w4144 & w13093 ) | ( w4144 & w13095 ) | ( w13093 & w13095 ) ;
  assign w13097 = ( w4143 & ~w13094 ) | ( w4143 & w13096 ) | ( ~w13094 & w13096 ) ;
  assign w13098 = \pi044 ^ w13097 ;
  assign w13099 = ( w12932 & w12933 ) | ( w12932 & ~w12995 ) | ( w12933 & ~w12995 ) ;
  assign w13100 = ( ~w12973 & w12974 ) | ( ~w12973 & w12982 ) | ( w12974 & w12982 ) ;
  assign w13101 = ~\pi098 & w5802 ;
  assign w13102 = \pi097 & w6052 ;
  assign w13103 = ( w5802 & ~w13101 ) | ( w5802 & w13102 ) | ( ~w13101 & w13102 ) ;
  assign w13104 = ~\pi099 & w5804 ;
  assign w13105 = w2966 | w13103 ;
  assign w13106 = ( w5805 & w13103 ) | ( w5805 & w13105 ) | ( w13103 & w13105 ) ;
  assign w13107 = ( w5804 & ~w13104 ) | ( w5804 & w13106 ) | ( ~w13104 & w13106 ) ;
  assign w13108 = \pi053 ^ w13107 ;
  assign w13109 = ( w12934 & ~w12963 ) | ( w12934 & w12971 ) | ( ~w12963 & w12971 ) ;
  assign w13110 = \pi062 ^ w12955 ;
  assign w13111 = ( \pi062 & \pi063 ) | ( \pi062 & \pi086 ) | ( \pi063 & \pi086 ) ;
  assign w13112 = \pi062 & \pi085 ;
  assign w13113 = ( ~\pi062 & w13111 ) | ( ~\pi062 & w13112 ) | ( w13111 & w13112 ) ;
  assign w13114 = ( ~\pi063 & w13111 ) | ( ~\pi063 & w13113 ) | ( w13111 & w13113 ) ;
  assign w13115 = ( w12948 & w13110 ) | ( w12948 & ~w13114 ) | ( w13110 & ~w13114 ) ;
  assign w13116 = ~\pi089 & w7811 ;
  assign w13117 = \pi088 & w8046 ;
  assign w13118 = ( w7811 & ~w13116 ) | ( w7811 & w13117 ) | ( ~w13116 & w13117 ) ;
  assign w13119 = ~\pi090 & w7813 ;
  assign w13120 = ~w1801 & w7814 ;
  assign w13121 = ( w7814 & w13118 ) | ( w7814 & ~w13120 ) | ( w13118 & ~w13120 ) ;
  assign w13122 = ( w7813 & ~w13119 ) | ( w7813 & w13121 ) | ( ~w13119 & w13121 ) ;
  assign w13123 = \pi063 & ~\pi085 ;
  assign w13124 = ~\pi063 & \pi086 ;
  assign w13125 = ( \pi062 & ~w13123 ) | ( \pi062 & w13124 ) | ( ~w13123 & w13124 ) ;
  assign w13126 = w13122 ^ w13125 ;
  assign w13127 = \pi086 ^ w13126 ;
  assign w13128 = ( \pi063 & w13122 ) | ( \pi063 & ~w13124 ) | ( w13122 & ~w13124 ) ;
  assign w13129 = ( \pi062 & ~\pi063 ) | ( \pi062 & w13128 ) | ( ~\pi063 & w13128 ) ;
  assign w13130 = ( \pi062 & ~w13127 ) | ( \pi062 & w13129 ) | ( ~w13127 & w13129 ) ;
  assign w13131 = ( \pi063 & \pi087 ) | ( \pi063 & w13130 ) | ( \pi087 & w13130 ) ;
  assign w13132 = w13127 ^ w13131 ;
  assign w13133 = ~\pi092 & w7135 ;
  assign w13134 = \pi091 & w7359 ;
  assign w13135 = ( w7135 & ~w13133 ) | ( w7135 & w13134 ) | ( ~w13133 & w13134 ) ;
  assign w13136 = ~\pi093 & w7137 ;
  assign w13137 = w2155 | w13135 ;
  assign w13138 = ( w7138 & w13135 ) | ( w7138 & w13137 ) | ( w13135 & w13137 ) ;
  assign w13139 = ( w7137 & ~w13136 ) | ( w7137 & w13138 ) | ( ~w13136 & w13138 ) ;
  assign w13140 = \pi059 ^ w13139 ;
  assign w13141 = w13115 ^ w13132 ;
  assign w13142 = w13140 ^ w13141 ;
  assign w13143 = ( w12942 & w12943 ) | ( w12942 & ~w12961 ) | ( w12943 & ~w12961 ) ;
  assign w13144 = ~\pi095 & w6466 ;
  assign w13145 = \pi094 & w6702 ;
  assign w13146 = ( w6466 & ~w13144 ) | ( w6466 & w13145 ) | ( ~w13144 & w13145 ) ;
  assign w13147 = ~\pi096 & w6468 ;
  assign w13148 = w2546 | w13146 ;
  assign w13149 = ( w6469 & w13146 ) | ( w6469 & w13148 ) | ( w13146 & w13148 ) ;
  assign w13150 = ( w6468 & ~w13147 ) | ( w6468 & w13149 ) | ( ~w13147 & w13149 ) ;
  assign w13151 = \pi056 ^ w13150 ;
  assign w13152 = w13142 ^ w13143 ;
  assign w13153 = w13151 ^ w13152 ;
  assign w13154 = w13109 ^ w13153 ;
  assign w13155 = w13108 ^ w13154 ;
  assign w13156 = ~\pi101 & w5209 ;
  assign w13157 = \pi100 & w5433 ;
  assign w13158 = ( w5209 & ~w13156 ) | ( w5209 & w13157 ) | ( ~w13156 & w13157 ) ;
  assign w13159 = ~\pi102 & w5211 ;
  assign w13160 = w3284 | w13158 ;
  assign w13161 = ( w5212 & w13158 ) | ( w5212 & w13160 ) | ( w13158 & w13160 ) ;
  assign w13162 = ( w5211 & ~w13159 ) | ( w5211 & w13161 ) | ( ~w13159 & w13161 ) ;
  assign w13163 = \pi050 ^ w13162 ;
  assign w13164 = w13100 ^ w13155 ;
  assign w13165 = w13163 ^ w13164 ;
  assign w13166 = ( ~w12984 & w12985 ) | ( ~w12984 & w12993 ) | ( w12985 & w12993 ) ;
  assign w13167 = ~\pi104 & w4654 ;
  assign w13168 = \pi103 & w4876 ;
  assign w13169 = ( w4654 & ~w13167 ) | ( w4654 & w13168 ) | ( ~w13167 & w13168 ) ;
  assign w13170 = ~\pi105 & w4656 ;
  assign w13171 = w3905 | w13169 ;
  assign w13172 = ( w4657 & w13169 ) | ( w4657 & w13171 ) | ( w13169 & w13171 ) ;
  assign w13173 = ( w4656 & ~w13170 ) | ( w4656 & w13172 ) | ( ~w13170 & w13172 ) ;
  assign w13174 = \pi047 ^ w13173 ;
  assign w13175 = w13165 ^ w13166 ;
  assign w13176 = w13174 ^ w13175 ;
  assign w13177 = w13099 ^ w13176 ;
  assign w13178 = w13098 ^ w13177 ;
  assign w13179 = ~\pi110 & w3635 ;
  assign w13180 = \pi109 & w3817 ;
  assign w13181 = ( w3635 & ~w13179 ) | ( w3635 & w13180 ) | ( ~w13179 & w13180 ) ;
  assign w13182 = ~\pi111 & w3637 ;
  assign w13183 = w4811 | w13181 ;
  assign w13184 = ( w3638 & w13181 ) | ( w3638 & w13183 ) | ( w13181 & w13183 ) ;
  assign w13185 = ( w3637 & ~w13182 ) | ( w3637 & w13184 ) | ( ~w13182 & w13184 ) ;
  assign w13186 = \pi041 ^ w13185 ;
  assign w13187 = w13090 ^ w13178 ;
  assign w13188 = w13186 ^ w13187 ;
  assign w13189 = ( ~w12999 & w13000 ) | ( ~w12999 & w13008 ) | ( w13000 & w13008 ) ;
  assign w13190 = ~\pi113 & w3178 ;
  assign w13191 = \pi112 & w3340 ;
  assign w13192 = ( w3178 & ~w13190 ) | ( w3178 & w13191 ) | ( ~w13190 & w13191 ) ;
  assign w13193 = ~\pi114 & w3180 ;
  assign w13194 = w5565 | w13192 ;
  assign w13195 = ( w3181 & w13192 ) | ( w3181 & w13194 ) | ( w13192 & w13194 ) ;
  assign w13196 = ( w3180 & ~w13193 ) | ( w3180 & w13195 ) | ( ~w13193 & w13195 ) ;
  assign w13197 = \pi038 ^ w13196 ;
  assign w13198 = w13188 ^ w13189 ;
  assign w13199 = w13197 ^ w13198 ;
  assign w13200 = w13089 ^ w13199 ;
  assign w13201 = w13088 ^ w13200 ;
  assign w13202 = w13080 ^ w13201 ;
  assign w13203 = w13079 ^ w13202 ;
  assign w13204 = w13071 ^ w13203 ;
  assign w13205 = w13070 ^ w13204 ;
  assign w13206 = w13060 ^ w13062 ;
  assign w13207 = w13205 ^ w13206 ;
  assign w13208 = w13052 ^ w13207 ;
  assign w13209 = w13048 ^ w13208 ;
  assign w13210 = w13044 ^ w13209 ;
  assign w13211 = w13047 ^ w13210 ;
  assign w13212 = ( w13044 & w13047 ) | ( w13044 & w13209 ) | ( w13047 & w13209 ) ;
  assign w13213 = ( w13048 & w13052 ) | ( w13048 & w13207 ) | ( w13052 & w13207 ) ;
  assign w13214 = ( w13060 & w13062 ) | ( w13060 & w13205 ) | ( w13062 & w13205 ) ;
  assign w13215 = ~\pi126 & w1629 ;
  assign w13216 = \pi125 & w1722 ;
  assign w13217 = ( w1629 & ~w13215 ) | ( w1629 & w13216 ) | ( ~w13215 & w13216 ) ;
  assign w13218 = ~\pi127 & w1631 ;
  assign w13219 = w8466 | w13217 ;
  assign w13220 = ( w1632 & w13217 ) | ( w1632 & w13219 ) | ( w13217 & w13219 ) ;
  assign w13221 = ( w1631 & ~w13218 ) | ( w1631 & w13220 ) | ( ~w13218 & w13220 ) ;
  assign w13222 = \pi026 ^ w13221 ;
  assign w13223 = ( w13070 & w13071 ) | ( w13070 & w13203 ) | ( w13071 & w13203 ) ;
  assign w13224 = ~\pi123 & w1944 ;
  assign w13225 = \pi122 & w2072 ;
  assign w13226 = ( w1944 & ~w13224 ) | ( w1944 & w13225 ) | ( ~w13224 & w13225 ) ;
  assign w13227 = ~\pi124 & w1946 ;
  assign w13228 = w7538 | w13226 ;
  assign w13229 = ( w1947 & w13226 ) | ( w1947 & w13228 ) | ( w13226 & w13228 ) ;
  assign w13230 = ( w1946 & ~w13227 ) | ( w1946 & w13229 ) | ( ~w13227 & w13229 ) ;
  assign w13231 = \pi029 ^ w13230 ;
  assign w13232 = ~\pi120 & w2310 ;
  assign w13233 = \pi119 & w2443 ;
  assign w13234 = ( w2310 & ~w13232 ) | ( w2310 & w13233 ) | ( ~w13232 & w13233 ) ;
  assign w13235 = ~\pi121 & w2312 ;
  assign w13236 = w7050 | w13234 ;
  assign w13237 = ( w2313 & w13234 ) | ( w2313 & w13236 ) | ( w13234 & w13236 ) ;
  assign w13238 = ( w2312 & ~w13235 ) | ( w2312 & w13237 ) | ( ~w13235 & w13237 ) ;
  assign w13239 = \pi032 ^ w13238 ;
  assign w13240 = ( ~w13079 & w13080 ) | ( ~w13079 & w13201 ) | ( w13080 & w13201 ) ;
  assign w13241 = w13239 ^ w13240 ;
  assign w13242 = ( w13088 & w13089 ) | ( w13088 & ~w13199 ) | ( w13089 & ~w13199 ) ;
  assign w13243 = ( ~w13188 & w13189 ) | ( ~w13188 & w13197 ) | ( w13189 & w13197 ) ;
  assign w13244 = ( w13098 & w13099 ) | ( w13098 & ~w13176 ) | ( w13099 & ~w13176 ) ;
  assign w13245 = ( ~w13165 & w13166 ) | ( ~w13165 & w13174 ) | ( w13166 & w13174 ) ;
  assign w13246 = ~\pi099 & w5802 ;
  assign w13247 = \pi098 & w6052 ;
  assign w13248 = ( w5802 & ~w13246 ) | ( w5802 & w13247 ) | ( ~w13246 & w13247 ) ;
  assign w13249 = ~\pi100 & w5804 ;
  assign w13250 = w3104 | w13248 ;
  assign w13251 = ( w5805 & w13248 ) | ( w5805 & w13250 ) | ( w13248 & w13250 ) ;
  assign w13252 = ( w5804 & ~w13249 ) | ( w5804 & w13251 ) | ( ~w13249 & w13251 ) ;
  assign w13253 = \pi053 ^ w13252 ;
  assign w13254 = ( w13115 & ~w13132 ) | ( w13115 & w13140 ) | ( ~w13132 & w13140 ) ;
  assign w13255 = \pi063 ^ w13122 ;
  assign w13256 = ( ~\pi086 & \pi087 ) | ( ~\pi086 & w13255 ) | ( \pi087 & w13255 ) ;
  assign w13257 = w8323 ^ w13256 ;
  assign w13258 = ( \pi085 & \pi086 ) | ( \pi085 & w13122 ) | ( \pi086 & w13122 ) ;
  assign w13259 = ( ~\pi086 & w13255 ) | ( ~\pi086 & w13258 ) | ( w13255 & w13258 ) ;
  assign w13260 = ( ~w13256 & w13257 ) | ( ~w13256 & w13259 ) | ( w13257 & w13259 ) ;
  assign w13261 = \pi086 ^ \pi088 ;
  assign w13262 = ( \pi062 & \pi063 ) | ( \pi062 & ~w13261 ) | ( \pi063 & ~w13261 ) ;
  assign w13263 = \pi086 ^ \pi087 ;
  assign w13264 = \pi062 & ~w13263 ;
  assign w13265 = ( \pi063 & ~w13263 ) | ( \pi063 & w13264 ) | ( ~w13263 & w13264 ) ;
  assign w13266 = \pi023 ^ w13265 ;
  assign w13267 = w13262 ^ w13266 ;
  assign w13268 = ~\pi090 & w7811 ;
  assign w13269 = \pi089 & w8046 ;
  assign w13270 = ( w7811 & ~w13268 ) | ( w7811 & w13269 ) | ( ~w13268 & w13269 ) ;
  assign w13271 = ~\pi091 & w7813 ;
  assign w13272 = w1908 | w13270 ;
  assign w13273 = ( w7814 & w13270 ) | ( w7814 & w13272 ) | ( w13270 & w13272 ) ;
  assign w13274 = ( w7813 & ~w13271 ) | ( w7813 & w13273 ) | ( ~w13271 & w13273 ) ;
  assign w13275 = \pi062 ^ w13274 ;
  assign w13276 = w13260 ^ w13275 ;
  assign w13277 = w13267 ^ w13276 ;
  assign w13278 = ~\pi093 & w7135 ;
  assign w13279 = \pi092 & w7359 ;
  assign w13280 = ( w7135 & ~w13278 ) | ( w7135 & w13279 ) | ( ~w13278 & w13279 ) ;
  assign w13281 = ~\pi094 & w7137 ;
  assign w13282 = w2274 | w13280 ;
  assign w13283 = ( w7138 & w13280 ) | ( w7138 & w13282 ) | ( w13280 & w13282 ) ;
  assign w13284 = ( w7137 & ~w13281 ) | ( w7137 & w13283 ) | ( ~w13281 & w13283 ) ;
  assign w13285 = \pi059 ^ w13284 ;
  assign w13286 = w13254 ^ w13277 ;
  assign w13287 = w13285 ^ w13286 ;
  assign w13288 = ~\pi096 & w6466 ;
  assign w13289 = \pi095 & w6702 ;
  assign w13290 = ( w6466 & ~w13288 ) | ( w6466 & w13289 ) | ( ~w13288 & w13289 ) ;
  assign w13291 = ~\pi097 & w6468 ;
  assign w13292 = w2673 | w13290 ;
  assign w13293 = ( w6469 & w13290 ) | ( w6469 & w13292 ) | ( w13290 & w13292 ) ;
  assign w13294 = ( w6468 & ~w13291 ) | ( w6468 & w13293 ) | ( ~w13291 & w13293 ) ;
  assign w13295 = \pi056 ^ w13294 ;
  assign w13296 = ( ~w13142 & w13143 ) | ( ~w13142 & w13151 ) | ( w13143 & w13151 ) ;
  assign w13297 = w13287 ^ w13296 ;
  assign w13298 = w13295 ^ w13297 ;
  assign w13299 = ( w13108 & w13109 ) | ( w13108 & ~w13153 ) | ( w13109 & ~w13153 ) ;
  assign w13300 = w13298 ^ w13299 ;
  assign w13301 = w13253 ^ w13300 ;
  assign w13302 = ~\pi102 & w5209 ;
  assign w13303 = \pi101 & w5433 ;
  assign w13304 = ( w5209 & ~w13302 ) | ( w5209 & w13303 ) | ( ~w13302 & w13303 ) ;
  assign w13305 = ~\pi103 & w5211 ;
  assign w13306 = w3437 | w13304 ;
  assign w13307 = ( w5212 & w13304 ) | ( w5212 & w13306 ) | ( w13304 & w13306 ) ;
  assign w13308 = ( w5211 & ~w13305 ) | ( w5211 & w13307 ) | ( ~w13305 & w13307 ) ;
  assign w13309 = \pi050 ^ w13308 ;
  assign w13310 = ( w13100 & ~w13155 ) | ( w13100 & w13163 ) | ( ~w13155 & w13163 ) ;
  assign w13311 = w13301 ^ w13310 ;
  assign w13312 = w13309 ^ w13311 ;
  assign w13313 = ~\pi105 & w4654 ;
  assign w13314 = \pi104 & w4876 ;
  assign w13315 = ( w4654 & ~w13313 ) | ( w4654 & w13314 ) | ( ~w13313 & w13314 ) ;
  assign w13316 = ~\pi106 & w4656 ;
  assign w13317 = w4068 | w13315 ;
  assign w13318 = ( w4657 & w13315 ) | ( w4657 & w13317 ) | ( w13315 & w13317 ) ;
  assign w13319 = ( w4656 & ~w13316 ) | ( w4656 & w13318 ) | ( ~w13316 & w13318 ) ;
  assign w13320 = \pi047 ^ w13319 ;
  assign w13321 = w13245 ^ w13312 ;
  assign w13322 = w13320 ^ w13321 ;
  assign w13323 = ~\pi108 & w4141 ;
  assign w13324 = \pi107 & w4334 ;
  assign w13325 = ( w4141 & ~w13323 ) | ( w4141 & w13324 ) | ( ~w13323 & w13324 ) ;
  assign w13326 = ~\pi109 & w4143 ;
  assign w13327 = w4599 | w13325 ;
  assign w13328 = ( w4144 & w13325 ) | ( w4144 & w13327 ) | ( w13325 & w13327 ) ;
  assign w13329 = ( w4143 & ~w13326 ) | ( w4143 & w13328 ) | ( ~w13326 & w13328 ) ;
  assign w13330 = \pi044 ^ w13329 ;
  assign w13331 = w13244 ^ w13322 ;
  assign w13332 = w13330 ^ w13331 ;
  assign w13333 = ~\pi111 & w3635 ;
  assign w13334 = \pi110 & w3817 ;
  assign w13335 = ( w3635 & ~w13333 ) | ( w3635 & w13334 ) | ( ~w13333 & w13334 ) ;
  assign w13336 = ~\pi112 & w3637 ;
  assign w13337 = w4999 | w13335 ;
  assign w13338 = ( w3638 & w13335 ) | ( w3638 & w13337 ) | ( w13335 & w13337 ) ;
  assign w13339 = ( w3637 & ~w13336 ) | ( w3637 & w13338 ) | ( ~w13336 & w13338 ) ;
  assign w13340 = \pi041 ^ w13339 ;
  assign w13341 = ( w13090 & ~w13178 ) | ( w13090 & w13186 ) | ( ~w13178 & w13186 ) ;
  assign w13342 = w13332 ^ w13341 ;
  assign w13343 = w13340 ^ w13342 ;
  assign w13344 = ~\pi114 & w3178 ;
  assign w13345 = \pi113 & w3340 ;
  assign w13346 = ( w3178 & ~w13344 ) | ( w3178 & w13345 ) | ( ~w13344 & w13345 ) ;
  assign w13347 = ~\pi115 & w3180 ;
  assign w13348 = w5585 | w13346 ;
  assign w13349 = ( w3181 & w13346 ) | ( w3181 & w13348 ) | ( w13346 & w13348 ) ;
  assign w13350 = ( w3180 & ~w13347 ) | ( w3180 & w13349 ) | ( ~w13347 & w13349 ) ;
  assign w13351 = \pi038 ^ w13350 ;
  assign w13352 = ( w13243 & ~w13343 ) | ( w13243 & w13351 ) | ( ~w13343 & w13351 ) ;
  assign w13353 = w13243 ^ w13343 ;
  assign w13354 = w13351 ^ w13353 ;
  assign w13355 = ~\pi117 & w2712 ;
  assign w13356 = \pi116 & w2872 ;
  assign w13357 = ( w2712 & ~w13355 ) | ( w2712 & w13356 ) | ( ~w13355 & w13356 ) ;
  assign w13358 = ~\pi118 & w2714 ;
  assign w13359 = w6206 | w13357 ;
  assign w13360 = ( w2715 & w13357 ) | ( w2715 & w13359 ) | ( w13357 & w13359 ) ;
  assign w13361 = ( w2714 & ~w13358 ) | ( w2714 & w13360 ) | ( ~w13358 & w13360 ) ;
  assign w13362 = \pi035 ^ w13361 ;
  assign w13363 = w13242 ^ w13354 ;
  assign w13364 = w13362 ^ w13363 ;
  assign w13365 = w13231 ^ w13364 ;
  assign w13366 = w13223 ^ w13365 ;
  assign w13367 = w13241 ^ w13366 ;
  assign w13368 = w13214 ^ w13222 ;
  assign w13369 = w13367 ^ w13368 ;
  assign w13370 = w13212 ^ w13213 ;
  assign w13371 = w13369 ^ w13370 ;
  assign w13372 = ( w13212 & w13213 ) | ( w13212 & w13369 ) | ( w13213 & w13369 ) ;
  assign w13373 = ( w13214 & w13222 ) | ( w13214 & w13367 ) | ( w13222 & w13367 ) ;
  assign w13374 = ~\pi124 & w1944 ;
  assign w13375 = \pi123 & w2072 ;
  assign w13376 = ( w1944 & ~w13374 ) | ( w1944 & w13375 ) | ( ~w13374 & w13375 ) ;
  assign w13377 = ~\pi125 & w1946 ;
  assign w13378 = w7988 | w13376 ;
  assign w13379 = ( w1947 & w13376 ) | ( w1947 & w13378 ) | ( w13376 & w13378 ) ;
  assign w13380 = ( w1946 & ~w13377 ) | ( w1946 & w13379 ) | ( ~w13377 & w13379 ) ;
  assign w13381 = \pi029 ^ w13380 ;
  assign w13382 = ( ~w13239 & w13240 ) | ( ~w13239 & w13364 ) | ( w13240 & w13364 ) ;
  assign w13383 = ( w13242 & ~w13354 ) | ( w13242 & w13362 ) | ( ~w13354 & w13362 ) ;
  assign w13384 = \pi120 & w2443 ;
  assign w13385 = ( \pi122 & w2312 ) | ( \pi122 & w13384 ) | ( w2312 & w13384 ) ;
  assign w13386 = \pi121 | w13385 ;
  assign w13387 = ( w2310 & w13385 ) | ( w2310 & w13386 ) | ( w13385 & w13386 ) ;
  assign w13388 = w13384 | w13387 ;
  assign w13389 = ~\pi106 & w4654 ;
  assign w13390 = \pi105 & w4876 ;
  assign w13391 = ( w4654 & ~w13389 ) | ( w4654 & w13390 ) | ( ~w13389 & w13390 ) ;
  assign w13392 = ~\pi107 & w4656 ;
  assign w13393 = w4087 | w13391 ;
  assign w13394 = ( w4657 & w13391 ) | ( w4657 & w13393 ) | ( w13391 & w13393 ) ;
  assign w13395 = ( w4656 & ~w13392 ) | ( w4656 & w13394 ) | ( ~w13392 & w13394 ) ;
  assign w13396 = \pi047 ^ w13395 ;
  assign w13397 = ( ~w13301 & w13309 ) | ( ~w13301 & w13310 ) | ( w13309 & w13310 ) ;
  assign w13398 = ~\pi103 & w5209 ;
  assign w13399 = \pi102 & w5433 ;
  assign w13400 = ( w5209 & ~w13398 ) | ( w5209 & w13399 ) | ( ~w13398 & w13399 ) ;
  assign w13401 = ~\pi104 & w5211 ;
  assign w13402 = w3740 | w13400 ;
  assign w13403 = ( w5212 & w13400 ) | ( w5212 & w13402 ) | ( w13400 & w13402 ) ;
  assign w13404 = ( w5211 & ~w13401 ) | ( w5211 & w13403 ) | ( ~w13401 & w13403 ) ;
  assign w13405 = \pi050 ^ w13404 ;
  assign w13406 = ( w13253 & ~w13298 ) | ( w13253 & w13299 ) | ( ~w13298 & w13299 ) ;
  assign w13407 = ( w13260 & ~w13267 ) | ( w13260 & w13275 ) | ( ~w13267 & w13275 ) ;
  assign w13408 = \pi062 ^ w12958 ;
  assign w13409 = ( \pi086 & \pi088 ) | ( \pi086 & w13408 ) | ( \pi088 & w13408 ) ;
  assign w13410 = ( ~\pi023 & \pi087 ) | ( ~\pi023 & w13409 ) | ( \pi087 & w13409 ) ;
  assign w13411 = w10655 & w13410 ;
  assign w13412 = ~\pi091 & w7811 ;
  assign w13413 = \pi090 & w8046 ;
  assign w13414 = ( w7811 & ~w13412 ) | ( w7811 & w13413 ) | ( ~w13412 & w13413 ) ;
  assign w13415 = ~\pi092 & w7813 ;
  assign w13416 = ~w2033 & w7814 ;
  assign w13417 = ( w7814 & w13414 ) | ( w7814 & ~w13416 ) | ( w13414 & ~w13416 ) ;
  assign w13418 = ( w7813 & ~w13415 ) | ( w7813 & w13417 ) | ( ~w13415 & w13417 ) ;
  assign w13419 = w13411 ^ w13418 ;
  assign w13420 = \pi062 ^ \pi089 ;
  assign w13421 = \pi063 ^ \pi089 ;
  assign w13422 = \pi062 & ~\pi088 ;
  assign w13423 = ( w13420 & ~w13421 ) | ( w13420 & w13422 ) | ( ~w13421 & w13422 ) ;
  assign w13424 = w13419 ^ w13423 ;
  assign w13425 = ~\pi094 & w7135 ;
  assign w13426 = \pi093 & w7359 ;
  assign w13427 = ( w7135 & ~w13425 ) | ( w7135 & w13426 ) | ( ~w13425 & w13426 ) ;
  assign w13428 = ~\pi095 & w7137 ;
  assign w13429 = w2409 | w13427 ;
  assign w13430 = ( w7138 & w13427 ) | ( w7138 & w13429 ) | ( w13427 & w13429 ) ;
  assign w13431 = ( w7137 & ~w13428 ) | ( w7137 & w13430 ) | ( ~w13428 & w13430 ) ;
  assign w13432 = \pi059 ^ w13431 ;
  assign w13433 = w13407 ^ w13424 ;
  assign w13434 = w13432 ^ w13433 ;
  assign w13435 = ( w13254 & ~w13277 ) | ( w13254 & w13285 ) | ( ~w13277 & w13285 ) ;
  assign w13436 = ~\pi097 & w6466 ;
  assign w13437 = \pi096 & w6702 ;
  assign w13438 = ( w6466 & ~w13436 ) | ( w6466 & w13437 ) | ( ~w13436 & w13437 ) ;
  assign w13439 = ~\pi098 & w6468 ;
  assign w13440 = w2824 | w13438 ;
  assign w13441 = ( w6469 & w13438 ) | ( w6469 & w13440 ) | ( w13438 & w13440 ) ;
  assign w13442 = ( w6468 & ~w13439 ) | ( w6468 & w13441 ) | ( ~w13439 & w13441 ) ;
  assign w13443 = \pi056 ^ w13442 ;
  assign w13444 = w13434 ^ w13435 ;
  assign w13445 = w13443 ^ w13444 ;
  assign w13446 = ( ~w13287 & w13295 ) | ( ~w13287 & w13296 ) | ( w13295 & w13296 ) ;
  assign w13447 = ~\pi100 & w5802 ;
  assign w13448 = \pi099 & w6052 ;
  assign w13449 = ( w5802 & ~w13447 ) | ( w5802 & w13448 ) | ( ~w13447 & w13448 ) ;
  assign w13450 = ~\pi101 & w5804 ;
  assign w13451 = w3264 | w13449 ;
  assign w13452 = ( w5805 & w13449 ) | ( w5805 & w13451 ) | ( w13449 & w13451 ) ;
  assign w13453 = ( w5804 & ~w13450 ) | ( w5804 & w13452 ) | ( ~w13450 & w13452 ) ;
  assign w13454 = \pi053 ^ w13453 ;
  assign w13455 = w13445 ^ w13446 ;
  assign w13456 = w13454 ^ w13455 ;
  assign w13457 = w13406 ^ w13456 ;
  assign w13458 = w13405 ^ w13457 ;
  assign w13459 = w13397 ^ w13458 ;
  assign w13460 = w13396 ^ w13459 ;
  assign w13461 = ( w13245 & ~w13312 ) | ( w13245 & w13320 ) | ( ~w13312 & w13320 ) ;
  assign w13462 = ~\pi109 & w4141 ;
  assign w13463 = \pi108 & w4334 ;
  assign w13464 = ( w4141 & ~w13462 ) | ( w4141 & w13463 ) | ( ~w13462 & w13463 ) ;
  assign w13465 = ~\pi110 & w4143 ;
  assign w13466 = w4792 | w13464 ;
  assign w13467 = ( w4144 & w13464 ) | ( w4144 & w13466 ) | ( w13464 & w13466 ) ;
  assign w13468 = ( w4143 & ~w13465 ) | ( w4143 & w13467 ) | ( ~w13465 & w13467 ) ;
  assign w13469 = \pi044 ^ w13468 ;
  assign w13470 = w13460 ^ w13461 ;
  assign w13471 = w13469 ^ w13470 ;
  assign w13472 = ( w13244 & ~w13322 ) | ( w13244 & w13330 ) | ( ~w13322 & w13330 ) ;
  assign w13473 = ~\pi112 & w3635 ;
  assign w13474 = \pi111 & w3817 ;
  assign w13475 = ( w3635 & ~w13473 ) | ( w3635 & w13474 ) | ( ~w13473 & w13474 ) ;
  assign w13476 = ~\pi113 & w3637 ;
  assign w13477 = w5366 | w13475 ;
  assign w13478 = ( w3638 & w13475 ) | ( w3638 & w13477 ) | ( w13475 & w13477 ) ;
  assign w13479 = ( w3637 & ~w13476 ) | ( w3637 & w13478 ) | ( ~w13476 & w13478 ) ;
  assign w13480 = \pi041 ^ w13479 ;
  assign w13481 = w13471 ^ w13472 ;
  assign w13482 = w13480 ^ w13481 ;
  assign w13483 = ( ~w13332 & w13340 ) | ( ~w13332 & w13341 ) | ( w13340 & w13341 ) ;
  assign w13484 = ~\pi115 & w3178 ;
  assign w13485 = \pi114 & w3340 ;
  assign w13486 = ( w3178 & ~w13484 ) | ( w3178 & w13485 ) | ( ~w13484 & w13485 ) ;
  assign w13487 = ~\pi116 & w3180 ;
  assign w13488 = w5976 | w13486 ;
  assign w13489 = ( w3181 & w13486 ) | ( w3181 & w13488 ) | ( w13486 & w13488 ) ;
  assign w13490 = ( w3180 & ~w13487 ) | ( w3180 & w13489 ) | ( ~w13487 & w13489 ) ;
  assign w13491 = \pi038 ^ w13490 ;
  assign w13492 = w13482 ^ w13483 ;
  assign w13493 = w13491 ^ w13492 ;
  assign w13494 = ~\pi118 & w2712 ;
  assign w13495 = \pi117 & w2872 ;
  assign w13496 = ( w2712 & ~w13494 ) | ( w2712 & w13495 ) | ( ~w13494 & w13495 ) ;
  assign w13497 = ~\pi119 & w2714 ;
  assign w13498 = w6616 | w13496 ;
  assign w13499 = ( w2715 & w13496 ) | ( w2715 & w13498 ) | ( w13496 & w13498 ) ;
  assign w13500 = ( w2714 & ~w13497 ) | ( w2714 & w13499 ) | ( ~w13497 & w13499 ) ;
  assign w13501 = \pi035 ^ w13500 ;
  assign w13502 = w13352 ^ w13493 ;
  assign w13503 = w13501 ^ w13502 ;
  assign w13504 = w2313 & ~w7069 ;
  assign w13505 = ( w2313 & w13388 ) | ( w2313 & ~w13504 ) | ( w13388 & ~w13504 ) ;
  assign w13506 = w13383 ^ w13505 ;
  assign w13507 = \pi032 ^ w13503 ;
  assign w13508 = w13506 ^ w13507 ;
  assign w13509 = w13381 ^ w13382 ;
  assign w13510 = w13508 ^ w13509 ;
  assign w13511 = w13241 ^ w13364 ;
  assign w13512 = ( w13223 & w13231 ) | ( w13223 & w13511 ) | ( w13231 & w13511 ) ;
  assign w13513 = \pi127 & w1629 ;
  assign w13514 = ( \pi126 & ~w1632 ) | ( \pi126 & w8490 ) | ( ~w1632 & w8490 ) ;
  assign w13515 = \pi126 & ~w1722 ;
  assign w13516 = ( ~\pi126 & w13514 ) | ( ~\pi126 & w13515 ) | ( w13514 & w13515 ) ;
  assign w13517 = ( w9420 & w13513 ) | ( w9420 & ~w13516 ) | ( w13513 & ~w13516 ) ;
  assign w13518 = \pi026 ^ w13517 ;
  assign w13519 = w13510 ^ w13518 ;
  assign w13520 = w13512 ^ w13519 ;
  assign w13521 = w13372 ^ w13373 ;
  assign w13522 = w13520 ^ w13521 ;
  assign w13523 = ( w13372 & w13373 ) | ( w13372 & w13520 ) | ( w13373 & w13520 ) ;
  assign w13524 = ( w13510 & w13512 ) | ( w13510 & w13518 ) | ( w13512 & w13518 ) ;
  assign w13525 = ( ~w13381 & w13382 ) | ( ~w13381 & w13508 ) | ( w13382 & w13508 ) ;
  assign w13526 = w1632 & w8481 ;
  assign w13527 = w1722 | w13526 ;
  assign w13528 = ( \pi127 & w13526 ) | ( \pi127 & w13527 ) | ( w13526 & w13527 ) ;
  assign w13529 = \pi026 ^ w13528 ;
  assign w13530 = ~\pi125 & w1944 ;
  assign w13531 = \pi124 & w2072 ;
  assign w13532 = ( w1944 & ~w13530 ) | ( w1944 & w13531 ) | ( ~w13530 & w13531 ) ;
  assign w13533 = ~\pi126 & w1946 ;
  assign w13534 = w8231 | w13532 ;
  assign w13535 = ( w1947 & w13532 ) | ( w1947 & w13534 ) | ( w13532 & w13534 ) ;
  assign w13536 = ( w1946 & ~w13533 ) | ( w1946 & w13535 ) | ( ~w13533 & w13535 ) ;
  assign w13537 = \pi029 ^ w13536 ;
  assign w13538 = w7069 | w13388 ;
  assign w13539 = ( w2313 & w13388 ) | ( w2313 & w13538 ) | ( w13388 & w13538 ) ;
  assign w13540 = \pi032 ^ w13539 ;
  assign w13541 = ( w13383 & ~w13503 ) | ( w13383 & w13540 ) | ( ~w13503 & w13540 ) ;
  assign w13542 = ~\pi122 & w2310 ;
  assign w13543 = \pi121 & w2443 ;
  assign w13544 = ( w2310 & ~w13542 ) | ( w2310 & w13543 ) | ( ~w13542 & w13543 ) ;
  assign w13545 = ~\pi123 & w2312 ;
  assign w13546 = w7516 | w13544 ;
  assign w13547 = ( w2313 & w13544 ) | ( w2313 & w13546 ) | ( w13544 & w13546 ) ;
  assign w13548 = ( w2312 & ~w13545 ) | ( w2312 & w13547 ) | ( ~w13545 & w13547 ) ;
  assign w13549 = \pi032 ^ w13548 ;
  assign w13550 = ( w13352 & ~w13493 ) | ( w13352 & w13501 ) | ( ~w13493 & w13501 ) ;
  assign w13551 = ~\pi119 & w2712 ;
  assign w13552 = \pi118 & w2872 ;
  assign w13553 = ( w2712 & ~w13551 ) | ( w2712 & w13552 ) | ( ~w13551 & w13552 ) ;
  assign w13554 = ~\pi120 & w2714 ;
  assign w13555 = w6634 | w13553 ;
  assign w13556 = ( w2715 & w13553 ) | ( w2715 & w13555 ) | ( w13553 & w13555 ) ;
  assign w13557 = ( w2714 & ~w13554 ) | ( w2714 & w13556 ) | ( ~w13554 & w13556 ) ;
  assign w13558 = \pi035 ^ w13557 ;
  assign w13559 = ( ~w13482 & w13483 ) | ( ~w13482 & w13491 ) | ( w13483 & w13491 ) ;
  assign w13560 = ~\pi116 & w3178 ;
  assign w13561 = \pi115 & w3340 ;
  assign w13562 = ( w3178 & ~w13560 ) | ( w3178 & w13561 ) | ( ~w13560 & w13561 ) ;
  assign w13563 = ~\pi117 & w3180 ;
  assign w13564 = w6185 | w13562 ;
  assign w13565 = ( w3181 & w13562 ) | ( w3181 & w13564 ) | ( w13562 & w13564 ) ;
  assign w13566 = ( w3180 & ~w13563 ) | ( w3180 & w13565 ) | ( ~w13563 & w13565 ) ;
  assign w13567 = \pi038 ^ w13566 ;
  assign w13568 = ( ~w13471 & w13472 ) | ( ~w13471 & w13480 ) | ( w13472 & w13480 ) ;
  assign w13569 = ( w13396 & w13397 ) | ( w13396 & ~w13458 ) | ( w13397 & ~w13458 ) ;
  assign w13570 = ~\pi107 & w4654 ;
  assign w13571 = \pi106 & w4876 ;
  assign w13572 = ( w4654 & ~w13570 ) | ( w4654 & w13571 ) | ( ~w13570 & w13571 ) ;
  assign w13573 = ~\pi108 & w4656 ;
  assign w13574 = w4425 | w13572 ;
  assign w13575 = ( w4657 & w13572 ) | ( w4657 & w13574 ) | ( w13572 & w13574 ) ;
  assign w13576 = ( w4656 & ~w13573 ) | ( w4656 & w13575 ) | ( ~w13573 & w13575 ) ;
  assign w13577 = \pi047 ^ w13576 ;
  assign w13578 = ( w13405 & w13406 ) | ( w13405 & ~w13456 ) | ( w13406 & ~w13456 ) ;
  assign w13579 = ( ~w13434 & w13435 ) | ( ~w13434 & w13443 ) | ( w13435 & w13443 ) ;
  assign w13580 = ~\pi098 & w6466 ;
  assign w13581 = \pi097 & w6702 ;
  assign w13582 = ( w6466 & ~w13580 ) | ( w6466 & w13581 ) | ( ~w13580 & w13581 ) ;
  assign w13583 = ~\pi099 & w6468 ;
  assign w13584 = w2966 | w13582 ;
  assign w13585 = ( w6469 & w13582 ) | ( w6469 & w13584 ) | ( w13582 & w13584 ) ;
  assign w13586 = ( w6468 & ~w13583 ) | ( w6468 & w13585 ) | ( ~w13583 & w13585 ) ;
  assign w13587 = \pi056 ^ w13586 ;
  assign w13588 = ( w13407 & ~w13424 ) | ( w13407 & w13432 ) | ( ~w13424 & w13432 ) ;
  assign w13589 = ~\pi095 & w7135 ;
  assign w13590 = \pi094 & w7359 ;
  assign w13591 = ( w7135 & ~w13589 ) | ( w7135 & w13590 ) | ( ~w13589 & w13590 ) ;
  assign w13592 = ~\pi096 & w7137 ;
  assign w13593 = w2546 | w13591 ;
  assign w13594 = ( w7138 & w13591 ) | ( w7138 & w13593 ) | ( w13591 & w13593 ) ;
  assign w13595 = ( w7137 & ~w13592 ) | ( w7137 & w13594 ) | ( ~w13592 & w13594 ) ;
  assign w13596 = \pi059 ^ w13595 ;
  assign w13597 = \pi062 ^ w13418 ;
  assign w13598 = ( \pi062 & \pi063 ) | ( \pi062 & \pi089 ) | ( \pi063 & \pi089 ) ;
  assign w13599 = \pi062 & \pi088 ;
  assign w13600 = ( ~\pi062 & w13598 ) | ( ~\pi062 & w13599 ) | ( w13598 & w13599 ) ;
  assign w13601 = ( ~\pi063 & w13598 ) | ( ~\pi063 & w13600 ) | ( w13598 & w13600 ) ;
  assign w13602 = ( w13411 & w13597 ) | ( w13411 & ~w13601 ) | ( w13597 & ~w13601 ) ;
  assign w13603 = ~\pi092 & w7811 ;
  assign w13604 = \pi091 & w8046 ;
  assign w13605 = ( w7811 & ~w13603 ) | ( w7811 & w13604 ) | ( ~w13603 & w13604 ) ;
  assign w13606 = ~\pi093 & w7813 ;
  assign w13607 = ~w2155 & w7814 ;
  assign w13608 = ( w7814 & w13605 ) | ( w7814 & ~w13607 ) | ( w13605 & ~w13607 ) ;
  assign w13609 = ( w7813 & ~w13606 ) | ( w7813 & w13608 ) | ( ~w13606 & w13608 ) ;
  assign w13610 = \pi063 & ~\pi088 ;
  assign w13611 = ~\pi063 & \pi089 ;
  assign w13612 = ( \pi062 & ~w13610 ) | ( \pi062 & w13611 ) | ( ~w13610 & w13611 ) ;
  assign w13613 = w13609 ^ w13612 ;
  assign w13614 = \pi089 ^ w13613 ;
  assign w13615 = ( \pi063 & w13609 ) | ( \pi063 & ~w13611 ) | ( w13609 & ~w13611 ) ;
  assign w13616 = ( \pi062 & ~\pi063 ) | ( \pi062 & w13615 ) | ( ~\pi063 & w13615 ) ;
  assign w13617 = ( \pi062 & ~w13614 ) | ( \pi062 & w13616 ) | ( ~w13614 & w13616 ) ;
  assign w13618 = ( \pi063 & \pi090 ) | ( \pi063 & w13617 ) | ( \pi090 & w13617 ) ;
  assign w13619 = w13614 ^ w13618 ;
  assign w13620 = w13596 ^ w13602 ;
  assign w13621 = w13619 ^ w13620 ;
  assign w13622 = w13587 ^ w13588 ;
  assign w13623 = w13621 ^ w13622 ;
  assign w13624 = ~\pi101 & w5802 ;
  assign w13625 = \pi100 & w6052 ;
  assign w13626 = ( w5802 & ~w13624 ) | ( w5802 & w13625 ) | ( ~w13624 & w13625 ) ;
  assign w13627 = ~\pi102 & w5804 ;
  assign w13628 = w3284 | w13626 ;
  assign w13629 = ( w5805 & w13626 ) | ( w5805 & w13628 ) | ( w13626 & w13628 ) ;
  assign w13630 = ( w5804 & ~w13627 ) | ( w5804 & w13629 ) | ( ~w13627 & w13629 ) ;
  assign w13631 = \pi053 ^ w13630 ;
  assign w13632 = w13579 ^ w13623 ;
  assign w13633 = w13631 ^ w13632 ;
  assign w13634 = ( ~w13445 & w13446 ) | ( ~w13445 & w13454 ) | ( w13446 & w13454 ) ;
  assign w13635 = ~\pi104 & w5209 ;
  assign w13636 = \pi103 & w5433 ;
  assign w13637 = ( w5209 & ~w13635 ) | ( w5209 & w13636 ) | ( ~w13635 & w13636 ) ;
  assign w13638 = ~\pi105 & w5211 ;
  assign w13639 = w3905 | w13637 ;
  assign w13640 = ( w5212 & w13637 ) | ( w5212 & w13639 ) | ( w13637 & w13639 ) ;
  assign w13641 = ( w5211 & ~w13638 ) | ( w5211 & w13640 ) | ( ~w13638 & w13640 ) ;
  assign w13642 = \pi050 ^ w13641 ;
  assign w13643 = w13633 ^ w13634 ;
  assign w13644 = w13642 ^ w13643 ;
  assign w13645 = w13578 ^ w13644 ;
  assign w13646 = w13577 ^ w13645 ;
  assign w13647 = ~\pi110 & w4141 ;
  assign w13648 = \pi109 & w4334 ;
  assign w13649 = ( w4141 & ~w13647 ) | ( w4141 & w13648 ) | ( ~w13647 & w13648 ) ;
  assign w13650 = ~\pi111 & w4143 ;
  assign w13651 = w4811 | w13649 ;
  assign w13652 = ( w4144 & w13649 ) | ( w4144 & w13651 ) | ( w13649 & w13651 ) ;
  assign w13653 = ( w4143 & ~w13650 ) | ( w4143 & w13652 ) | ( ~w13650 & w13652 ) ;
  assign w13654 = \pi044 ^ w13653 ;
  assign w13655 = w13569 ^ w13646 ;
  assign w13656 = w13654 ^ w13655 ;
  assign w13657 = ( ~w13460 & w13461 ) | ( ~w13460 & w13469 ) | ( w13461 & w13469 ) ;
  assign w13658 = ~\pi113 & w3635 ;
  assign w13659 = \pi112 & w3817 ;
  assign w13660 = ( w3635 & ~w13658 ) | ( w3635 & w13659 ) | ( ~w13658 & w13659 ) ;
  assign w13661 = ~\pi114 & w3637 ;
  assign w13662 = w5565 | w13660 ;
  assign w13663 = ( w3638 & w13660 ) | ( w3638 & w13662 ) | ( w13660 & w13662 ) ;
  assign w13664 = ( w3637 & ~w13661 ) | ( w3637 & w13663 ) | ( ~w13661 & w13663 ) ;
  assign w13665 = \pi041 ^ w13664 ;
  assign w13666 = w13656 ^ w13657 ;
  assign w13667 = w13665 ^ w13666 ;
  assign w13668 = w13568 ^ w13667 ;
  assign w13669 = w13567 ^ w13668 ;
  assign w13670 = w13559 ^ w13669 ;
  assign w13671 = w13558 ^ w13670 ;
  assign w13672 = w13549 ^ w13550 ;
  assign w13673 = w13671 ^ w13672 ;
  assign w13674 = w13537 ^ w13541 ;
  assign w13675 = w13673 ^ w13674 ;
  assign w13676 = w13529 ^ w13675 ;
  assign w13677 = w13525 ^ w13676 ;
  assign w13678 = w13523 ^ w13677 ;
  assign w13679 = w13524 ^ w13678 ;
  assign w13680 = ( w13525 & ~w13529 ) | ( w13525 & w13675 ) | ( ~w13529 & w13675 ) ;
  assign w13681 = ( w13537 & w13541 ) | ( w13537 & ~w13673 ) | ( w13541 & ~w13673 ) ;
  assign w13682 = ~\pi126 & w1944 ;
  assign w13683 = \pi125 & w2072 ;
  assign w13684 = ( w1944 & ~w13682 ) | ( w1944 & w13683 ) | ( ~w13682 & w13683 ) ;
  assign w13685 = ~\pi127 & w1946 ;
  assign w13686 = w8466 | w13684 ;
  assign w13687 = ( w1947 & w13684 ) | ( w1947 & w13686 ) | ( w13684 & w13686 ) ;
  assign w13688 = ( w1946 & ~w13685 ) | ( w1946 & w13687 ) | ( ~w13685 & w13687 ) ;
  assign w13689 = \pi029 ^ w13688 ;
  assign w13690 = ~\pi120 & w2712 ;
  assign w13691 = \pi119 & w2872 ;
  assign w13692 = ( w2712 & ~w13690 ) | ( w2712 & w13691 ) | ( ~w13690 & w13691 ) ;
  assign w13693 = ~\pi121 & w2714 ;
  assign w13694 = w7050 | w13692 ;
  assign w13695 = ( w2715 & w13692 ) | ( w2715 & w13694 ) | ( w13692 & w13694 ) ;
  assign w13696 = ( w2714 & ~w13693 ) | ( w2714 & w13695 ) | ( ~w13693 & w13695 ) ;
  assign w13697 = \pi035 ^ w13696 ;
  assign w13698 = ( w13567 & w13568 ) | ( w13567 & ~w13667 ) | ( w13568 & ~w13667 ) ;
  assign w13699 = ( ~w13656 & w13657 ) | ( ~w13656 & w13665 ) | ( w13657 & w13665 ) ;
  assign w13700 = ( w13577 & w13578 ) | ( w13577 & ~w13644 ) | ( w13578 & ~w13644 ) ;
  assign w13701 = ( ~w13633 & w13634 ) | ( ~w13633 & w13642 ) | ( w13634 & w13642 ) ;
  assign w13702 = ~\pi096 & w7135 ;
  assign w13703 = \pi095 & w7359 ;
  assign w13704 = ( w7135 & ~w13702 ) | ( w7135 & w13703 ) | ( ~w13702 & w13703 ) ;
  assign w13705 = ~\pi097 & w7137 ;
  assign w13706 = w2673 | w13704 ;
  assign w13707 = ( w7138 & w13704 ) | ( w7138 & w13706 ) | ( w13704 & w13706 ) ;
  assign w13708 = ( w7137 & ~w13705 ) | ( w7137 & w13707 ) | ( ~w13705 & w13707 ) ;
  assign w13709 = \pi059 ^ w13708 ;
  assign w13710 = ( w13596 & w13602 ) | ( w13596 & ~w13619 ) | ( w13602 & ~w13619 ) ;
  assign w13711 = \pi063 ^ w13609 ;
  assign w13712 = ( ~\pi089 & \pi090 ) | ( ~\pi089 & w13711 ) | ( \pi090 & w13711 ) ;
  assign w13713 = w8323 ^ w13712 ;
  assign w13714 = ( \pi088 & \pi089 ) | ( \pi088 & w13609 ) | ( \pi089 & w13609 ) ;
  assign w13715 = ( ~\pi089 & w13711 ) | ( ~\pi089 & w13714 ) | ( w13711 & w13714 ) ;
  assign w13716 = ( ~w13712 & w13713 ) | ( ~w13712 & w13715 ) | ( w13713 & w13715 ) ;
  assign w13717 = \pi089 ^ \pi091 ;
  assign w13718 = ( \pi062 & \pi063 ) | ( \pi062 & ~w13717 ) | ( \pi063 & ~w13717 ) ;
  assign w13719 = \pi089 ^ \pi090 ;
  assign w13720 = \pi062 & ~w13719 ;
  assign w13721 = ( \pi063 & ~w13719 ) | ( \pi063 & w13720 ) | ( ~w13719 & w13720 ) ;
  assign w13722 = \pi026 ^ w13721 ;
  assign w13723 = w13718 ^ w13722 ;
  assign w13724 = ~\pi093 & w7811 ;
  assign w13725 = \pi092 & w8046 ;
  assign w13726 = ( w7811 & ~w13724 ) | ( w7811 & w13725 ) | ( ~w13724 & w13725 ) ;
  assign w13727 = ~\pi094 & w7813 ;
  assign w13728 = w2274 | w13726 ;
  assign w13729 = ( w7814 & w13726 ) | ( w7814 & w13728 ) | ( w13726 & w13728 ) ;
  assign w13730 = ( w7813 & ~w13727 ) | ( w7813 & w13729 ) | ( ~w13727 & w13729 ) ;
  assign w13731 = \pi062 ^ w13730 ;
  assign w13732 = w13716 ^ w13731 ;
  assign w13733 = w13723 ^ w13732 ;
  assign w13734 = w13710 ^ w13733 ;
  assign w13735 = w13709 ^ w13734 ;
  assign w13736 = ~\pi099 & w6466 ;
  assign w13737 = \pi098 & w6702 ;
  assign w13738 = ( w6466 & ~w13736 ) | ( w6466 & w13737 ) | ( ~w13736 & w13737 ) ;
  assign w13739 = ~\pi100 & w6468 ;
  assign w13740 = w3104 | w13738 ;
  assign w13741 = ( w6469 & w13738 ) | ( w6469 & w13740 ) | ( w13738 & w13740 ) ;
  assign w13742 = ( w6468 & ~w13739 ) | ( w6468 & w13741 ) | ( ~w13739 & w13741 ) ;
  assign w13743 = \pi056 ^ w13742 ;
  assign w13744 = ( w13587 & w13588 ) | ( w13587 & ~w13621 ) | ( w13588 & ~w13621 ) ;
  assign w13745 = w13735 ^ w13744 ;
  assign w13746 = w13743 ^ w13745 ;
  assign w13747 = ~\pi102 & w5802 ;
  assign w13748 = \pi101 & w6052 ;
  assign w13749 = ( w5802 & ~w13747 ) | ( w5802 & w13748 ) | ( ~w13747 & w13748 ) ;
  assign w13750 = ~\pi103 & w5804 ;
  assign w13751 = w3437 | w13749 ;
  assign w13752 = ( w5805 & w13749 ) | ( w5805 & w13751 ) | ( w13749 & w13751 ) ;
  assign w13753 = ( w5804 & ~w13750 ) | ( w5804 & w13752 ) | ( ~w13750 & w13752 ) ;
  assign w13754 = \pi053 ^ w13753 ;
  assign w13755 = ( w13579 & ~w13623 ) | ( w13579 & w13631 ) | ( ~w13623 & w13631 ) ;
  assign w13756 = w13746 ^ w13755 ;
  assign w13757 = w13754 ^ w13756 ;
  assign w13758 = ~\pi105 & w5209 ;
  assign w13759 = \pi104 & w5433 ;
  assign w13760 = ( w5209 & ~w13758 ) | ( w5209 & w13759 ) | ( ~w13758 & w13759 ) ;
  assign w13761 = ~\pi106 & w5211 ;
  assign w13762 = w4068 | w13760 ;
  assign w13763 = ( w5212 & w13760 ) | ( w5212 & w13762 ) | ( w13760 & w13762 ) ;
  assign w13764 = ( w5211 & ~w13761 ) | ( w5211 & w13763 ) | ( ~w13761 & w13763 ) ;
  assign w13765 = \pi050 ^ w13764 ;
  assign w13766 = w13701 ^ w13757 ;
  assign w13767 = w13765 ^ w13766 ;
  assign w13768 = ~\pi108 & w4654 ;
  assign w13769 = \pi107 & w4876 ;
  assign w13770 = ( w4654 & ~w13768 ) | ( w4654 & w13769 ) | ( ~w13768 & w13769 ) ;
  assign w13771 = ~\pi109 & w4656 ;
  assign w13772 = w4599 | w13770 ;
  assign w13773 = ( w4657 & w13770 ) | ( w4657 & w13772 ) | ( w13770 & w13772 ) ;
  assign w13774 = ( w4656 & ~w13771 ) | ( w4656 & w13773 ) | ( ~w13771 & w13773 ) ;
  assign w13775 = \pi047 ^ w13774 ;
  assign w13776 = w13700 ^ w13767 ;
  assign w13777 = w13775 ^ w13776 ;
  assign w13778 = ~\pi111 & w4141 ;
  assign w13779 = \pi110 & w4334 ;
  assign w13780 = ( w4141 & ~w13778 ) | ( w4141 & w13779 ) | ( ~w13778 & w13779 ) ;
  assign w13781 = ~\pi112 & w4143 ;
  assign w13782 = w4999 | w13780 ;
  assign w13783 = ( w4144 & w13780 ) | ( w4144 & w13782 ) | ( w13780 & w13782 ) ;
  assign w13784 = ( w4143 & ~w13781 ) | ( w4143 & w13783 ) | ( ~w13781 & w13783 ) ;
  assign w13785 = \pi044 ^ w13784 ;
  assign w13786 = ( w13569 & ~w13646 ) | ( w13569 & w13654 ) | ( ~w13646 & w13654 ) ;
  assign w13787 = w13777 ^ w13786 ;
  assign w13788 = w13785 ^ w13787 ;
  assign w13789 = ~\pi114 & w3635 ;
  assign w13790 = \pi113 & w3817 ;
  assign w13791 = ( w3635 & ~w13789 ) | ( w3635 & w13790 ) | ( ~w13789 & w13790 ) ;
  assign w13792 = ~\pi115 & w3637 ;
  assign w13793 = w5585 | w13791 ;
  assign w13794 = ( w3638 & w13791 ) | ( w3638 & w13793 ) | ( w13791 & w13793 ) ;
  assign w13795 = ( w3637 & ~w13792 ) | ( w3637 & w13794 ) | ( ~w13792 & w13794 ) ;
  assign w13796 = \pi041 ^ w13795 ;
  assign w13797 = ( w13699 & ~w13788 ) | ( w13699 & w13796 ) | ( ~w13788 & w13796 ) ;
  assign w13798 = w13699 ^ w13788 ;
  assign w13799 = w13796 ^ w13798 ;
  assign w13800 = ~\pi117 & w3178 ;
  assign w13801 = \pi116 & w3340 ;
  assign w13802 = ( w3178 & ~w13800 ) | ( w3178 & w13801 ) | ( ~w13800 & w13801 ) ;
  assign w13803 = ~\pi118 & w3180 ;
  assign w13804 = w6206 | w13802 ;
  assign w13805 = ( w3181 & w13802 ) | ( w3181 & w13804 ) | ( w13802 & w13804 ) ;
  assign w13806 = ( w3180 & ~w13803 ) | ( w3180 & w13805 ) | ( ~w13803 & w13805 ) ;
  assign w13807 = \pi038 ^ w13806 ;
  assign w13808 = w13698 ^ w13799 ;
  assign w13809 = w13807 ^ w13808 ;
  assign w13810 = ( w13558 & w13559 ) | ( w13558 & ~w13669 ) | ( w13559 & ~w13669 ) ;
  assign w13811 = w13809 ^ w13810 ;
  assign w13812 = w13697 ^ w13811 ;
  assign w13813 = ~\pi123 & w2310 ;
  assign w13814 = \pi122 & w2443 ;
  assign w13815 = ( w2310 & ~w13813 ) | ( w2310 & w13814 ) | ( ~w13813 & w13814 ) ;
  assign w13816 = ~\pi124 & w2312 ;
  assign w13817 = w7538 | w13815 ;
  assign w13818 = ( w2313 & w13815 ) | ( w2313 & w13817 ) | ( w13815 & w13817 ) ;
  assign w13819 = ( w2312 & ~w13816 ) | ( w2312 & w13818 ) | ( ~w13816 & w13818 ) ;
  assign w13820 = \pi032 ^ w13819 ;
  assign w13821 = ( w13549 & w13550 ) | ( w13549 & ~w13671 ) | ( w13550 & ~w13671 ) ;
  assign w13822 = w13820 ^ w13821 ;
  assign w13823 = w13812 ^ w13822 ;
  assign w13824 = w13681 ^ w13689 ;
  assign w13825 = w13823 ^ w13824 ;
  assign w13826 = ( w13523 & w13524 ) | ( w13523 & w13677 ) | ( w13524 & w13677 ) ;
  assign w13827 = w13680 ^ w13826 ;
  assign w13828 = w13825 ^ w13827 ;
  assign w13829 = ( ~w13812 & w13820 ) | ( ~w13812 & w13821 ) | ( w13820 & w13821 ) ;
  assign w13830 = \pi127 & w1944 ;
  assign w13831 = ( \pi126 & ~w1947 ) | ( \pi126 & w8490 ) | ( ~w1947 & w8490 ) ;
  assign w13832 = \pi126 & ~w2072 ;
  assign w13833 = ( ~\pi126 & w13831 ) | ( ~\pi126 & w13832 ) | ( w13831 & w13832 ) ;
  assign w13834 = ( w9420 & w13830 ) | ( w9420 & ~w13833 ) | ( w13830 & ~w13833 ) ;
  assign w13835 = ~\pi124 & w2310 ;
  assign w13836 = \pi123 & w2443 ;
  assign w13837 = ( w2310 & ~w13835 ) | ( w2310 & w13836 ) | ( ~w13835 & w13836 ) ;
  assign w13838 = ~\pi125 & w2312 ;
  assign w13839 = w7988 | w13837 ;
  assign w13840 = ( w2313 & w13837 ) | ( w2313 & w13839 ) | ( w13837 & w13839 ) ;
  assign w13841 = ( w2312 & ~w13838 ) | ( w2312 & w13840 ) | ( ~w13838 & w13840 ) ;
  assign w13842 = \pi032 ^ w13841 ;
  assign w13843 = ( w13697 & ~w13809 ) | ( w13697 & w13810 ) | ( ~w13809 & w13810 ) ;
  assign w13844 = w13842 ^ w13843 ;
  assign w13845 = ~\pi121 & w2712 ;
  assign w13846 = \pi120 & w2872 ;
  assign w13847 = ( w2712 & ~w13845 ) | ( w2712 & w13846 ) | ( ~w13845 & w13846 ) ;
  assign w13848 = ~\pi122 & w2714 ;
  assign w13849 = w7069 | w13847 ;
  assign w13850 = ( w2715 & w13847 ) | ( w2715 & w13849 ) | ( w13847 & w13849 ) ;
  assign w13851 = ( w2714 & ~w13848 ) | ( w2714 & w13850 ) | ( ~w13848 & w13850 ) ;
  assign w13852 = \pi035 ^ w13851 ;
  assign w13853 = ( w13698 & ~w13799 ) | ( w13698 & w13807 ) | ( ~w13799 & w13807 ) ;
  assign w13854 = ~\pi106 & w5209 ;
  assign w13855 = \pi105 & w5433 ;
  assign w13856 = ( w5209 & ~w13854 ) | ( w5209 & w13855 ) | ( ~w13854 & w13855 ) ;
  assign w13857 = ~\pi107 & w5211 ;
  assign w13858 = w4087 | w13856 ;
  assign w13859 = ( w5212 & w13856 ) | ( w5212 & w13858 ) | ( w13856 & w13858 ) ;
  assign w13860 = ( w5211 & ~w13857 ) | ( w5211 & w13859 ) | ( ~w13857 & w13859 ) ;
  assign w13861 = \pi050 ^ w13860 ;
  assign w13862 = ( ~w13746 & w13754 ) | ( ~w13746 & w13755 ) | ( w13754 & w13755 ) ;
  assign w13863 = ~\pi103 & w5802 ;
  assign w13864 = \pi102 & w6052 ;
  assign w13865 = ( w5802 & ~w13863 ) | ( w5802 & w13864 ) | ( ~w13863 & w13864 ) ;
  assign w13866 = ~\pi104 & w5804 ;
  assign w13867 = w3740 | w13865 ;
  assign w13868 = ( w5805 & w13865 ) | ( w5805 & w13867 ) | ( w13865 & w13867 ) ;
  assign w13869 = ( w5804 & ~w13866 ) | ( w5804 & w13868 ) | ( ~w13866 & w13868 ) ;
  assign w13870 = \pi053 ^ w13869 ;
  assign w13871 = ( ~w13735 & w13743 ) | ( ~w13735 & w13744 ) | ( w13743 & w13744 ) ;
  assign w13872 = ~\pi097 & w7135 ;
  assign w13873 = \pi096 & w7359 ;
  assign w13874 = ( w7135 & ~w13872 ) | ( w7135 & w13873 ) | ( ~w13872 & w13873 ) ;
  assign w13875 = ~\pi098 & w7137 ;
  assign w13876 = w2824 | w13874 ;
  assign w13877 = ( w7138 & w13874 ) | ( w7138 & w13876 ) | ( w13874 & w13876 ) ;
  assign w13878 = ( w7137 & ~w13875 ) | ( w7137 & w13877 ) | ( ~w13875 & w13877 ) ;
  assign w13879 = \pi059 ^ w13878 ;
  assign w13880 = \pi062 ^ w13421 ;
  assign w13881 = ( \pi089 & \pi091 ) | ( \pi089 & w13880 ) | ( \pi091 & w13880 ) ;
  assign w13882 = ( ~\pi026 & \pi090 ) | ( ~\pi026 & w13881 ) | ( \pi090 & w13881 ) ;
  assign w13883 = w10655 & w13882 ;
  assign w13884 = ~\pi094 & w7811 ;
  assign w13885 = \pi093 & w8046 ;
  assign w13886 = ( w7811 & ~w13884 ) | ( w7811 & w13885 ) | ( ~w13884 & w13885 ) ;
  assign w13887 = ~\pi095 & w7813 ;
  assign w13888 = w2409 | w13886 ;
  assign w13889 = ( w7814 & w13886 ) | ( w7814 & w13888 ) | ( w13886 & w13888 ) ;
  assign w13890 = ( w7813 & ~w13887 ) | ( w7813 & w13889 ) | ( ~w13887 & w13889 ) ;
  assign w13891 = \pi062 ^ w13890 ;
  assign w13892 = w13883 ^ w13891 ;
  assign w13893 = ( \pi062 & \pi063 ) | ( \pi062 & \pi092 ) | ( \pi063 & \pi092 ) ;
  assign w13894 = \pi063 & ~\pi091 ;
  assign w13895 = \pi062 & w13894 ;
  assign w13896 = w13893 ^ w13895 ;
  assign w13897 = w13892 ^ w13896 ;
  assign w13898 = ( w13716 & ~w13723 ) | ( w13716 & w13731 ) | ( ~w13723 & w13731 ) ;
  assign w13899 = w13879 ^ w13897 ;
  assign w13900 = w13898 ^ w13899 ;
  assign w13901 = ( w13709 & w13710 ) | ( w13709 & ~w13733 ) | ( w13710 & ~w13733 ) ;
  assign w13902 = ~\pi100 & w6466 ;
  assign w13903 = \pi099 & w6702 ;
  assign w13904 = ( w6466 & ~w13902 ) | ( w6466 & w13903 ) | ( ~w13902 & w13903 ) ;
  assign w13905 = ~\pi101 & w6468 ;
  assign w13906 = w3264 | w13904 ;
  assign w13907 = ( w6469 & w13904 ) | ( w6469 & w13906 ) | ( w13904 & w13906 ) ;
  assign w13908 = ( w6468 & ~w13905 ) | ( w6468 & w13907 ) | ( ~w13905 & w13907 ) ;
  assign w13909 = \pi056 ^ w13908 ;
  assign w13910 = w13900 ^ w13901 ;
  assign w13911 = w13909 ^ w13910 ;
  assign w13912 = w13871 ^ w13911 ;
  assign w13913 = w13870 ^ w13912 ;
  assign w13914 = w13862 ^ w13913 ;
  assign w13915 = w13861 ^ w13914 ;
  assign w13916 = ( w13701 & ~w13757 ) | ( w13701 & w13765 ) | ( ~w13757 & w13765 ) ;
  assign w13917 = ~\pi109 & w4654 ;
  assign w13918 = \pi108 & w4876 ;
  assign w13919 = ( w4654 & ~w13917 ) | ( w4654 & w13918 ) | ( ~w13917 & w13918 ) ;
  assign w13920 = ~\pi110 & w4656 ;
  assign w13921 = w4792 | w13919 ;
  assign w13922 = ( w4657 & w13919 ) | ( w4657 & w13921 ) | ( w13919 & w13921 ) ;
  assign w13923 = ( w4656 & ~w13920 ) | ( w4656 & w13922 ) | ( ~w13920 & w13922 ) ;
  assign w13924 = \pi047 ^ w13923 ;
  assign w13925 = w13915 ^ w13916 ;
  assign w13926 = w13924 ^ w13925 ;
  assign w13927 = ( w13700 & ~w13767 ) | ( w13700 & w13775 ) | ( ~w13767 & w13775 ) ;
  assign w13928 = ~\pi112 & w4141 ;
  assign w13929 = \pi111 & w4334 ;
  assign w13930 = ( w4141 & ~w13928 ) | ( w4141 & w13929 ) | ( ~w13928 & w13929 ) ;
  assign w13931 = ~\pi113 & w4143 ;
  assign w13932 = w5366 | w13930 ;
  assign w13933 = ( w4144 & w13930 ) | ( w4144 & w13932 ) | ( w13930 & w13932 ) ;
  assign w13934 = ( w4143 & ~w13931 ) | ( w4143 & w13933 ) | ( ~w13931 & w13933 ) ;
  assign w13935 = \pi044 ^ w13934 ;
  assign w13936 = w13926 ^ w13927 ;
  assign w13937 = w13935 ^ w13936 ;
  assign w13938 = ( ~w13777 & w13785 ) | ( ~w13777 & w13786 ) | ( w13785 & w13786 ) ;
  assign w13939 = ~\pi115 & w3635 ;
  assign w13940 = \pi114 & w3817 ;
  assign w13941 = ( w3635 & ~w13939 ) | ( w3635 & w13940 ) | ( ~w13939 & w13940 ) ;
  assign w13942 = ~\pi116 & w3637 ;
  assign w13943 = w5976 | w13941 ;
  assign w13944 = ( w3638 & w13941 ) | ( w3638 & w13943 ) | ( w13941 & w13943 ) ;
  assign w13945 = ( w3637 & ~w13942 ) | ( w3637 & w13944 ) | ( ~w13942 & w13944 ) ;
  assign w13946 = \pi041 ^ w13945 ;
  assign w13947 = w13937 ^ w13938 ;
  assign w13948 = w13946 ^ w13947 ;
  assign w13949 = ~\pi118 & w3178 ;
  assign w13950 = \pi117 & w3340 ;
  assign w13951 = ( w3178 & ~w13949 ) | ( w3178 & w13950 ) | ( ~w13949 & w13950 ) ;
  assign w13952 = ~\pi119 & w3180 ;
  assign w13953 = w6616 | w13951 ;
  assign w13954 = ( w3181 & w13951 ) | ( w3181 & w13953 ) | ( w13951 & w13953 ) ;
  assign w13955 = ( w3180 & ~w13952 ) | ( w3180 & w13954 ) | ( ~w13952 & w13954 ) ;
  assign w13956 = \pi038 ^ w13955 ;
  assign w13957 = w13797 ^ w13948 ;
  assign w13958 = w13956 ^ w13957 ;
  assign w13959 = w13852 ^ w13853 ;
  assign w13960 = w13958 ^ w13959 ;
  assign w13961 = w13829 ^ w13844 ;
  assign w13962 = w13834 ^ w13960 ;
  assign w13963 = \pi029 ^ w13962 ;
  assign w13964 = w13961 ^ w13963 ;
  assign w13965 = ( w13681 & w13689 ) | ( w13681 & ~w13823 ) | ( w13689 & ~w13823 ) ;
  assign w13966 = ( w13680 & w13825 ) | ( w13680 & ~w13826 ) | ( w13825 & ~w13826 ) ;
  assign w13967 = w13965 ^ w13966 ;
  assign w13968 = w13964 ^ w13967 ;
  assign w13969 = ( w13964 & ~w13965 ) | ( w13964 & w13966 ) | ( ~w13965 & w13966 ) ;
  assign w13970 = \pi029 ^ w13834 ;
  assign w13971 = w13844 ^ w13960 ;
  assign w13972 = ( w13829 & w13970 ) | ( w13829 & ~w13971 ) | ( w13970 & ~w13971 ) ;
  assign w13973 = ( w13842 & w13843 ) | ( w13842 & ~w13960 ) | ( w13843 & ~w13960 ) ;
  assign w13974 = w1947 & w8481 ;
  assign w13975 = w2072 | w13974 ;
  assign w13976 = ( \pi127 & w13974 ) | ( \pi127 & w13975 ) | ( w13974 & w13975 ) ;
  assign w13977 = \pi029 ^ w13976 ;
  assign w13978 = ~\pi125 & w2310 ;
  assign w13979 = \pi124 & w2443 ;
  assign w13980 = ( w2310 & ~w13978 ) | ( w2310 & w13979 ) | ( ~w13978 & w13979 ) ;
  assign w13981 = ~\pi126 & w2312 ;
  assign w13982 = w8231 | w13980 ;
  assign w13983 = ( w2313 & w13980 ) | ( w2313 & w13982 ) | ( w13980 & w13982 ) ;
  assign w13984 = ( w2312 & ~w13981 ) | ( w2312 & w13983 ) | ( ~w13981 & w13983 ) ;
  assign w13985 = \pi032 ^ w13984 ;
  assign w13986 = ( w13852 & w13853 ) | ( w13852 & ~w13958 ) | ( w13853 & ~w13958 ) ;
  assign w13987 = ( w13797 & ~w13948 ) | ( w13797 & w13956 ) | ( ~w13948 & w13956 ) ;
  assign w13988 = ~\pi119 & w3178 ;
  assign w13989 = \pi118 & w3340 ;
  assign w13990 = ( w3178 & ~w13988 ) | ( w3178 & w13989 ) | ( ~w13988 & w13989 ) ;
  assign w13991 = ~\pi120 & w3180 ;
  assign w13992 = w6634 | w13990 ;
  assign w13993 = ( w3181 & w13990 ) | ( w3181 & w13992 ) | ( w13990 & w13992 ) ;
  assign w13994 = ( w3180 & ~w13991 ) | ( w3180 & w13993 ) | ( ~w13991 & w13993 ) ;
  assign w13995 = \pi038 ^ w13994 ;
  assign w13996 = ( ~w13937 & w13938 ) | ( ~w13937 & w13946 ) | ( w13938 & w13946 ) ;
  assign w13997 = ~\pi116 & w3635 ;
  assign w13998 = \pi115 & w3817 ;
  assign w13999 = ( w3635 & ~w13997 ) | ( w3635 & w13998 ) | ( ~w13997 & w13998 ) ;
  assign w14000 = ~\pi117 & w3637 ;
  assign w14001 = w6185 | w13999 ;
  assign w14002 = ( w3638 & w13999 ) | ( w3638 & w14001 ) | ( w13999 & w14001 ) ;
  assign w14003 = ( w3637 & ~w14000 ) | ( w3637 & w14002 ) | ( ~w14000 & w14002 ) ;
  assign w14004 = \pi041 ^ w14003 ;
  assign w14005 = ( ~w13926 & w13927 ) | ( ~w13926 & w13935 ) | ( w13927 & w13935 ) ;
  assign w14006 = ( w13861 & w13862 ) | ( w13861 & ~w13913 ) | ( w13862 & ~w13913 ) ;
  assign w14007 = ~\pi107 & w5209 ;
  assign w14008 = \pi106 & w5433 ;
  assign w14009 = ( w5209 & ~w14007 ) | ( w5209 & w14008 ) | ( ~w14007 & w14008 ) ;
  assign w14010 = ~\pi108 & w5211 ;
  assign w14011 = w4425 | w14009 ;
  assign w14012 = ( w5212 & w14009 ) | ( w5212 & w14011 ) | ( w14009 & w14011 ) ;
  assign w14013 = ( w5211 & ~w14010 ) | ( w5211 & w14012 ) | ( ~w14010 & w14012 ) ;
  assign w14014 = \pi050 ^ w14013 ;
  assign w14015 = ( w13870 & w13871 ) | ( w13870 & ~w13911 ) | ( w13871 & ~w13911 ) ;
  assign w14016 = ( w13879 & ~w13897 ) | ( w13879 & w13898 ) | ( ~w13897 & w13898 ) ;
  assign w14017 = ~\pi098 & w7135 ;
  assign w14018 = \pi097 & w7359 ;
  assign w14019 = ( w7135 & ~w14017 ) | ( w7135 & w14018 ) | ( ~w14017 & w14018 ) ;
  assign w14020 = ~\pi099 & w7137 ;
  assign w14021 = w2966 | w14019 ;
  assign w14022 = ( w7138 & w14019 ) | ( w7138 & w14021 ) | ( w14019 & w14021 ) ;
  assign w14023 = ( w7137 & ~w14020 ) | ( w7137 & w14022 ) | ( ~w14020 & w14022 ) ;
  assign w14024 = \pi059 ^ w14023 ;
  assign w14025 = \pi063 & \pi091 ;
  assign w14026 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w14025 ) | ( \pi063 & w14025 ) ;
  assign w14027 = ( \pi062 & ~\pi063 ) | ( \pi062 & w14025 ) | ( ~\pi063 & w14025 ) ;
  assign w14028 = ( \pi092 & w14026 ) | ( \pi092 & w14027 ) | ( w14026 & w14027 ) ;
  assign w14029 = ( w13883 & w13891 ) | ( w13883 & ~w14028 ) | ( w13891 & ~w14028 ) ;
  assign w14030 = \pi092 & ~w14029 ;
  assign w14031 = ( \pi063 & ~\pi091 ) | ( \pi063 & w14030 ) | ( ~\pi091 & w14030 ) ;
  assign w14032 = ( \pi062 & ~\pi063 ) | ( \pi062 & w14031 ) | ( ~\pi063 & w14031 ) ;
  assign w14033 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi093 ) | ( \pi063 & ~\pi093 ) ;
  assign w14034 = ( \pi092 & w14029 ) | ( \pi092 & w14033 ) | ( w14029 & w14033 ) ;
  assign w14035 = ( ~\pi063 & w14029 ) | ( ~\pi063 & w14030 ) | ( w14029 & w14030 ) ;
  assign w14036 = ( \pi062 & ~\pi092 ) | ( \pi062 & w14035 ) | ( ~\pi092 & w14035 ) ;
  assign w14037 = ( ~w14032 & w14034 ) | ( ~w14032 & w14036 ) | ( w14034 & w14036 ) ;
  assign w14038 = \pi091 ^ \pi093 ;
  assign w14039 = ( \pi062 & \pi063 ) | ( \pi062 & ~w14038 ) | ( \pi063 & ~w14038 ) ;
  assign w14040 = \pi091 ^ \pi092 ;
  assign w14041 = \pi062 & ~w14040 ;
  assign w14042 = ( \pi063 & ~w14040 ) | ( \pi063 & w14041 ) | ( ~w14040 & w14041 ) ;
  assign w14043 = w14029 ^ w14042 ;
  assign w14044 = w14039 ^ w14043 ;
  assign w14045 = ~\pi095 & w7811 ;
  assign w14046 = \pi094 & w8046 ;
  assign w14047 = ( w7811 & ~w14045 ) | ( w7811 & w14046 ) | ( ~w14045 & w14046 ) ;
  assign w14048 = ~\pi096 & w7813 ;
  assign w14049 = w2546 | w14047 ;
  assign w14050 = ( w7814 & w14047 ) | ( w7814 & w14049 ) | ( w14047 & w14049 ) ;
  assign w14051 = ( w7813 & ~w14048 ) | ( w7813 & w14050 ) | ( ~w14048 & w14050 ) ;
  assign w14052 = \pi062 ^ w14051 ;
  assign w14053 = w14024 ^ w14044 ;
  assign w14054 = w14052 ^ w14053 ;
  assign w14055 = ~\pi101 & w6466 ;
  assign w14056 = \pi100 & w6702 ;
  assign w14057 = ( w6466 & ~w14055 ) | ( w6466 & w14056 ) | ( ~w14055 & w14056 ) ;
  assign w14058 = ~\pi102 & w6468 ;
  assign w14059 = w3284 | w14057 ;
  assign w14060 = ( w6469 & w14057 ) | ( w6469 & w14059 ) | ( w14057 & w14059 ) ;
  assign w14061 = ( w6468 & ~w14058 ) | ( w6468 & w14060 ) | ( ~w14058 & w14060 ) ;
  assign w14062 = \pi056 ^ w14061 ;
  assign w14063 = w14016 ^ w14054 ;
  assign w14064 = w14062 ^ w14063 ;
  assign w14065 = ( ~w13900 & w13901 ) | ( ~w13900 & w13909 ) | ( w13901 & w13909 ) ;
  assign w14066 = ~\pi104 & w5802 ;
  assign w14067 = \pi103 & w6052 ;
  assign w14068 = ( w5802 & ~w14066 ) | ( w5802 & w14067 ) | ( ~w14066 & w14067 ) ;
  assign w14069 = ~\pi105 & w5804 ;
  assign w14070 = w3905 | w14068 ;
  assign w14071 = ( w5805 & w14068 ) | ( w5805 & w14070 ) | ( w14068 & w14070 ) ;
  assign w14072 = ( w5804 & ~w14069 ) | ( w5804 & w14071 ) | ( ~w14069 & w14071 ) ;
  assign w14073 = \pi053 ^ w14072 ;
  assign w14074 = w14064 ^ w14065 ;
  assign w14075 = w14073 ^ w14074 ;
  assign w14076 = w14015 ^ w14075 ;
  assign w14077 = w14014 ^ w14076 ;
  assign w14078 = ~\pi110 & w4654 ;
  assign w14079 = \pi109 & w4876 ;
  assign w14080 = ( w4654 & ~w14078 ) | ( w4654 & w14079 ) | ( ~w14078 & w14079 ) ;
  assign w14081 = ~\pi111 & w4656 ;
  assign w14082 = w4811 | w14080 ;
  assign w14083 = ( w4657 & w14080 ) | ( w4657 & w14082 ) | ( w14080 & w14082 ) ;
  assign w14084 = ( w4656 & ~w14081 ) | ( w4656 & w14083 ) | ( ~w14081 & w14083 ) ;
  assign w14085 = \pi047 ^ w14084 ;
  assign w14086 = w14006 ^ w14077 ;
  assign w14087 = w14085 ^ w14086 ;
  assign w14088 = ( ~w13915 & w13916 ) | ( ~w13915 & w13924 ) | ( w13916 & w13924 ) ;
  assign w14089 = ~\pi113 & w4141 ;
  assign w14090 = \pi112 & w4334 ;
  assign w14091 = ( w4141 & ~w14089 ) | ( w4141 & w14090 ) | ( ~w14089 & w14090 ) ;
  assign w14092 = ~\pi114 & w4143 ;
  assign w14093 = w5565 | w14091 ;
  assign w14094 = ( w4144 & w14091 ) | ( w4144 & w14093 ) | ( w14091 & w14093 ) ;
  assign w14095 = ( w4143 & ~w14092 ) | ( w4143 & w14094 ) | ( ~w14092 & w14094 ) ;
  assign w14096 = \pi044 ^ w14095 ;
  assign w14097 = w14087 ^ w14088 ;
  assign w14098 = w14096 ^ w14097 ;
  assign w14099 = w14005 ^ w14098 ;
  assign w14100 = w14004 ^ w14099 ;
  assign w14101 = w13996 ^ w14100 ;
  assign w14102 = w13995 ^ w14101 ;
  assign w14103 = ~\pi122 & w2712 ;
  assign w14104 = \pi121 & w2872 ;
  assign w14105 = ( w2712 & ~w14103 ) | ( w2712 & w14104 ) | ( ~w14103 & w14104 ) ;
  assign w14106 = ~\pi123 & w2714 ;
  assign w14107 = w7516 | w14105 ;
  assign w14108 = ( w2715 & w14105 ) | ( w2715 & w14107 ) | ( w14105 & w14107 ) ;
  assign w14109 = ( w2714 & ~w14106 ) | ( w2714 & w14108 ) | ( ~w14106 & w14108 ) ;
  assign w14110 = \pi035 ^ w14109 ;
  assign w14111 = w13987 ^ w14110 ;
  assign w14112 = w14102 ^ w14111 ;
  assign w14113 = w13985 ^ w14112 ;
  assign w14114 = w13986 ^ w14113 ;
  assign w14115 = w13977 ^ w14114 ;
  assign w14116 = w13973 ^ w14115 ;
  assign w14117 = w13969 ^ w14116 ;
  assign w14118 = w13972 ^ w14117 ;
  assign w14119 = ( w13969 & ~w13972 ) | ( w13969 & w14116 ) | ( ~w13972 & w14116 ) ;
  assign w14120 = ( w13973 & w13977 ) | ( w13973 & ~w14114 ) | ( w13977 & ~w14114 ) ;
  assign w14121 = ~\pi120 & w3178 ;
  assign w14122 = \pi119 & w3340 ;
  assign w14123 = ( w3178 & ~w14121 ) | ( w3178 & w14122 ) | ( ~w14121 & w14122 ) ;
  assign w14124 = ~\pi121 & w3180 ;
  assign w14125 = w7050 | w14123 ;
  assign w14126 = ( w3181 & w14123 ) | ( w3181 & w14125 ) | ( w14123 & w14125 ) ;
  assign w14127 = ( w3180 & ~w14124 ) | ( w3180 & w14126 ) | ( ~w14124 & w14126 ) ;
  assign w14128 = \pi038 ^ w14127 ;
  assign w14129 = ( w14004 & w14005 ) | ( w14004 & ~w14098 ) | ( w14005 & ~w14098 ) ;
  assign w14130 = ( ~w14087 & w14088 ) | ( ~w14087 & w14096 ) | ( w14088 & w14096 ) ;
  assign w14131 = ( w14014 & w14015 ) | ( w14014 & ~w14075 ) | ( w14015 & ~w14075 ) ;
  assign w14132 = ( ~w14064 & w14065 ) | ( ~w14064 & w14073 ) | ( w14065 & w14073 ) ;
  assign w14133 = ~\pi102 & w6466 ;
  assign w14134 = \pi101 & w6702 ;
  assign w14135 = ( w6466 & ~w14133 ) | ( w6466 & w14134 ) | ( ~w14133 & w14134 ) ;
  assign w14136 = ~\pi103 & w6468 ;
  assign w14137 = w3437 | w14135 ;
  assign w14138 = ( w6469 & w14135 ) | ( w6469 & w14137 ) | ( w14135 & w14137 ) ;
  assign w14139 = ( w6468 & ~w14136 ) | ( w6468 & w14138 ) | ( ~w14136 & w14138 ) ;
  assign w14140 = \pi056 ^ w14139 ;
  assign w14141 = ( w14024 & ~w14044 ) | ( w14024 & w14052 ) | ( ~w14044 & w14052 ) ;
  assign w14142 = \pi092 ^ \pi094 ;
  assign w14143 = ( \pi062 & \pi063 ) | ( \pi062 & ~w14142 ) | ( \pi063 & ~w14142 ) ;
  assign w14144 = \pi062 & ~w2154 ;
  assign w14145 = ( \pi063 & ~w2154 ) | ( \pi063 & w14144 ) | ( ~w2154 & w14144 ) ;
  assign w14146 = \pi029 ^ w14145 ;
  assign w14147 = w14143 ^ w14146 ;
  assign w14148 = ~\pi096 & w7811 ;
  assign w14149 = \pi095 & w8046 ;
  assign w14150 = ( w7811 & ~w14148 ) | ( w7811 & w14149 ) | ( ~w14148 & w14149 ) ;
  assign w14151 = ~\pi097 & w7813 ;
  assign w14152 = w2673 | w14150 ;
  assign w14153 = ( w7814 & w14150 ) | ( w7814 & w14152 ) | ( w14150 & w14152 ) ;
  assign w14154 = ( w7813 & ~w14151 ) | ( w7813 & w14153 ) | ( ~w14151 & w14153 ) ;
  assign w14155 = \pi062 ^ w14154 ;
  assign w14156 = w14037 ^ w14155 ;
  assign w14157 = w14147 ^ w14156 ;
  assign w14158 = ~\pi099 & w7135 ;
  assign w14159 = \pi098 & w7359 ;
  assign w14160 = ( w7135 & ~w14158 ) | ( w7135 & w14159 ) | ( ~w14158 & w14159 ) ;
  assign w14161 = ~\pi100 & w7137 ;
  assign w14162 = w3104 | w14160 ;
  assign w14163 = ( w7138 & w14160 ) | ( w7138 & w14162 ) | ( w14160 & w14162 ) ;
  assign w14164 = ( w7137 & ~w14161 ) | ( w7137 & w14163 ) | ( ~w14161 & w14163 ) ;
  assign w14165 = \pi059 ^ w14164 ;
  assign w14166 = w14141 ^ w14157 ;
  assign w14167 = w14165 ^ w14166 ;
  assign w14168 = ( w14016 & ~w14054 ) | ( w14016 & w14062 ) | ( ~w14054 & w14062 ) ;
  assign w14169 = w14167 ^ w14168 ;
  assign w14170 = w14140 ^ w14169 ;
  assign w14171 = ~\pi105 & w5802 ;
  assign w14172 = \pi104 & w6052 ;
  assign w14173 = ( w5802 & ~w14171 ) | ( w5802 & w14172 ) | ( ~w14171 & w14172 ) ;
  assign w14174 = ~\pi106 & w5804 ;
  assign w14175 = w4068 | w14173 ;
  assign w14176 = ( w5805 & w14173 ) | ( w5805 & w14175 ) | ( w14173 & w14175 ) ;
  assign w14177 = ( w5804 & ~w14174 ) | ( w5804 & w14176 ) | ( ~w14174 & w14176 ) ;
  assign w14178 = \pi053 ^ w14177 ;
  assign w14179 = w14132 ^ w14170 ;
  assign w14180 = w14178 ^ w14179 ;
  assign w14181 = ~\pi108 & w5209 ;
  assign w14182 = \pi107 & w5433 ;
  assign w14183 = ( w5209 & ~w14181 ) | ( w5209 & w14182 ) | ( ~w14181 & w14182 ) ;
  assign w14184 = ~\pi109 & w5211 ;
  assign w14185 = w4599 | w14183 ;
  assign w14186 = ( w5212 & w14183 ) | ( w5212 & w14185 ) | ( w14183 & w14185 ) ;
  assign w14187 = ( w5211 & ~w14184 ) | ( w5211 & w14186 ) | ( ~w14184 & w14186 ) ;
  assign w14188 = \pi050 ^ w14187 ;
  assign w14189 = w14131 ^ w14180 ;
  assign w14190 = w14188 ^ w14189 ;
  assign w14191 = ~\pi111 & w4654 ;
  assign w14192 = \pi110 & w4876 ;
  assign w14193 = ( w4654 & ~w14191 ) | ( w4654 & w14192 ) | ( ~w14191 & w14192 ) ;
  assign w14194 = ~\pi112 & w4656 ;
  assign w14195 = w4999 | w14193 ;
  assign w14196 = ( w4657 & w14193 ) | ( w4657 & w14195 ) | ( w14193 & w14195 ) ;
  assign w14197 = ( w4656 & ~w14194 ) | ( w4656 & w14196 ) | ( ~w14194 & w14196 ) ;
  assign w14198 = \pi047 ^ w14197 ;
  assign w14199 = ( w14006 & ~w14077 ) | ( w14006 & w14085 ) | ( ~w14077 & w14085 ) ;
  assign w14200 = w14190 ^ w14199 ;
  assign w14201 = w14198 ^ w14200 ;
  assign w14202 = ~\pi114 & w4141 ;
  assign w14203 = \pi113 & w4334 ;
  assign w14204 = ( w4141 & ~w14202 ) | ( w4141 & w14203 ) | ( ~w14202 & w14203 ) ;
  assign w14205 = ~\pi115 & w4143 ;
  assign w14206 = w5585 | w14204 ;
  assign w14207 = ( w4144 & w14204 ) | ( w4144 & w14206 ) | ( w14204 & w14206 ) ;
  assign w14208 = ( w4143 & ~w14205 ) | ( w4143 & w14207 ) | ( ~w14205 & w14207 ) ;
  assign w14209 = \pi044 ^ w14208 ;
  assign w14210 = ( w14130 & ~w14201 ) | ( w14130 & w14209 ) | ( ~w14201 & w14209 ) ;
  assign w14211 = w14130 ^ w14201 ;
  assign w14212 = w14209 ^ w14211 ;
  assign w14213 = ~\pi117 & w3635 ;
  assign w14214 = \pi116 & w3817 ;
  assign w14215 = ( w3635 & ~w14213 ) | ( w3635 & w14214 ) | ( ~w14213 & w14214 ) ;
  assign w14216 = ~\pi118 & w3637 ;
  assign w14217 = w6206 | w14215 ;
  assign w14218 = ( w3638 & w14215 ) | ( w3638 & w14217 ) | ( w14215 & w14217 ) ;
  assign w14219 = ( w3637 & ~w14216 ) | ( w3637 & w14218 ) | ( ~w14216 & w14218 ) ;
  assign w14220 = \pi041 ^ w14219 ;
  assign w14221 = w14129 ^ w14212 ;
  assign w14222 = w14220 ^ w14221 ;
  assign w14223 = ( w13995 & w13996 ) | ( w13995 & ~w14100 ) | ( w13996 & ~w14100 ) ;
  assign w14224 = w14222 ^ w14223 ;
  assign w14225 = w14128 ^ w14224 ;
  assign w14226 = ~\pi123 & w2712 ;
  assign w14227 = \pi122 & w2872 ;
  assign w14228 = ( w2712 & ~w14226 ) | ( w2712 & w14227 ) | ( ~w14226 & w14227 ) ;
  assign w14229 = ~\pi124 & w2714 ;
  assign w14230 = w7538 | w14228 ;
  assign w14231 = ( w2715 & w14228 ) | ( w2715 & w14230 ) | ( w14228 & w14230 ) ;
  assign w14232 = ( w2714 & ~w14229 ) | ( w2714 & w14231 ) | ( ~w14229 & w14231 ) ;
  assign w14233 = \pi035 ^ w14232 ;
  assign w14234 = ( w13987 & ~w14102 ) | ( w13987 & w14110 ) | ( ~w14102 & w14110 ) ;
  assign w14235 = w14233 ^ w14234 ;
  assign w14236 = w14225 ^ w14235 ;
  assign w14237 = ( w13985 & w13986 ) | ( w13985 & ~w14112 ) | ( w13986 & ~w14112 ) ;
  assign w14238 = ~\pi126 & w2310 ;
  assign w14239 = \pi125 & w2443 ;
  assign w14240 = ( w2310 & ~w14238 ) | ( w2310 & w14239 ) | ( ~w14238 & w14239 ) ;
  assign w14241 = ~\pi127 & w2312 ;
  assign w14242 = w8466 | w14240 ;
  assign w14243 = ( w2313 & w14240 ) | ( w2313 & w14242 ) | ( w14240 & w14242 ) ;
  assign w14244 = ( w2312 & ~w14241 ) | ( w2312 & w14243 ) | ( ~w14241 & w14243 ) ;
  assign w14245 = \pi032 ^ w14244 ;
  assign w14246 = w14237 ^ w14245 ;
  assign w14247 = w14236 ^ w14246 ;
  assign w14248 = w14119 ^ w14120 ;
  assign w14249 = w14247 ^ w14248 ;
  assign w14250 = ( ~w14225 & w14233 ) | ( ~w14225 & w14234 ) | ( w14233 & w14234 ) ;
  assign w14251 = \pi127 & w2310 ;
  assign w14252 = ( \pi126 & ~w2313 ) | ( \pi126 & w8490 ) | ( ~w2313 & w8490 ) ;
  assign w14253 = \pi126 & ~w2443 ;
  assign w14254 = ( ~\pi126 & w14252 ) | ( ~\pi126 & w14253 ) | ( w14252 & w14253 ) ;
  assign w14255 = ( w9420 & w14251 ) | ( w9420 & ~w14254 ) | ( w14251 & ~w14254 ) ;
  assign w14256 = ~\pi121 & w3178 ;
  assign w14257 = \pi120 & w3340 ;
  assign w14258 = ( w3178 & ~w14256 ) | ( w3178 & w14257 ) | ( ~w14256 & w14257 ) ;
  assign w14259 = ~\pi122 & w3180 ;
  assign w14260 = w7069 | w14258 ;
  assign w14261 = ( w3181 & w14258 ) | ( w3181 & w14260 ) | ( w14258 & w14260 ) ;
  assign w14262 = ( w3180 & ~w14259 ) | ( w3180 & w14261 ) | ( ~w14259 & w14261 ) ;
  assign w14263 = \pi038 ^ w14262 ;
  assign w14264 = ( w14129 & ~w14212 ) | ( w14129 & w14220 ) | ( ~w14212 & w14220 ) ;
  assign w14265 = ~\pi106 & w5802 ;
  assign w14266 = \pi105 & w6052 ;
  assign w14267 = ( w5802 & ~w14265 ) | ( w5802 & w14266 ) | ( ~w14265 & w14266 ) ;
  assign w14268 = ~\pi107 & w5804 ;
  assign w14269 = w4087 | w14267 ;
  assign w14270 = ( w5805 & w14267 ) | ( w5805 & w14269 ) | ( w14267 & w14269 ) ;
  assign w14271 = ( w5804 & ~w14268 ) | ( w5804 & w14270 ) | ( ~w14268 & w14270 ) ;
  assign w14272 = \pi053 ^ w14271 ;
  assign w14273 = ( w14140 & ~w14167 ) | ( w14140 & w14168 ) | ( ~w14167 & w14168 ) ;
  assign w14274 = ~\pi103 & w6466 ;
  assign w14275 = \pi102 & w6702 ;
  assign w14276 = ( w6466 & ~w14274 ) | ( w6466 & w14275 ) | ( ~w14274 & w14275 ) ;
  assign w14277 = ~\pi104 & w6468 ;
  assign w14278 = w3740 | w14276 ;
  assign w14279 = ( w6469 & w14276 ) | ( w6469 & w14278 ) | ( w14276 & w14278 ) ;
  assign w14280 = ( w6468 & ~w14277 ) | ( w6468 & w14279 ) | ( ~w14277 & w14279 ) ;
  assign w14281 = \pi056 ^ w14280 ;
  assign w14282 = ( w14141 & ~w14157 ) | ( w14141 & w14165 ) | ( ~w14157 & w14165 ) ;
  assign w14283 = ~\pi100 & w7135 ;
  assign w14284 = \pi099 & w7359 ;
  assign w14285 = ( w7135 & ~w14283 ) | ( w7135 & w14284 ) | ( ~w14283 & w14284 ) ;
  assign w14286 = ~\pi101 & w7137 ;
  assign w14287 = w3264 | w14285 ;
  assign w14288 = ( w7138 & w14285 ) | ( w7138 & w14287 ) | ( w14285 & w14287 ) ;
  assign w14289 = ( w7137 & ~w14286 ) | ( w7137 & w14288 ) | ( ~w14286 & w14288 ) ;
  assign w14290 = \pi059 ^ w14289 ;
  assign w14291 = ( w14037 & ~w14147 ) | ( w14037 & w14155 ) | ( ~w14147 & w14155 ) ;
  assign w14292 = \pi063 ^ \pi092 ;
  assign w14293 = \pi062 ^ w14292 ;
  assign w14294 = ( \pi092 & \pi094 ) | ( \pi092 & w14293 ) | ( \pi094 & w14293 ) ;
  assign w14295 = ( ~\pi029 & \pi093 ) | ( ~\pi029 & w14294 ) | ( \pi093 & w14294 ) ;
  assign w14296 = w10655 & w14295 ;
  assign w14297 = ~\pi097 & w7811 ;
  assign w14298 = \pi096 & w8046 ;
  assign w14299 = ( w7811 & ~w14297 ) | ( w7811 & w14298 ) | ( ~w14297 & w14298 ) ;
  assign w14300 = ~\pi098 & w7813 ;
  assign w14301 = w2824 | w14299 ;
  assign w14302 = ( w7814 & w14299 ) | ( w7814 & w14301 ) | ( w14299 & w14301 ) ;
  assign w14303 = ( w7813 & ~w14300 ) | ( w7813 & w14302 ) | ( ~w14300 & w14302 ) ;
  assign w14304 = \pi062 ^ w14303 ;
  assign w14305 = w14296 ^ w14304 ;
  assign w14306 = ( \pi062 & \pi063 ) | ( \pi062 & \pi095 ) | ( \pi063 & \pi095 ) ;
  assign w14307 = \pi063 & ~\pi094 ;
  assign w14308 = \pi062 & w14307 ;
  assign w14309 = w14306 ^ w14308 ;
  assign w14310 = w14305 ^ w14309 ;
  assign w14311 = w14291 ^ w14310 ;
  assign w14312 = w14290 ^ w14311 ;
  assign w14313 = w14282 ^ w14312 ;
  assign w14314 = w14281 ^ w14313 ;
  assign w14315 = w14273 ^ w14314 ;
  assign w14316 = w14272 ^ w14315 ;
  assign w14317 = ( w14132 & ~w14170 ) | ( w14132 & w14178 ) | ( ~w14170 & w14178 ) ;
  assign w14318 = ~\pi109 & w5209 ;
  assign w14319 = \pi108 & w5433 ;
  assign w14320 = ( w5209 & ~w14318 ) | ( w5209 & w14319 ) | ( ~w14318 & w14319 ) ;
  assign w14321 = ~\pi110 & w5211 ;
  assign w14322 = w4792 | w14320 ;
  assign w14323 = ( w5212 & w14320 ) | ( w5212 & w14322 ) | ( w14320 & w14322 ) ;
  assign w14324 = ( w5211 & ~w14321 ) | ( w5211 & w14323 ) | ( ~w14321 & w14323 ) ;
  assign w14325 = \pi050 ^ w14324 ;
  assign w14326 = w14316 ^ w14317 ;
  assign w14327 = w14325 ^ w14326 ;
  assign w14328 = ( w14131 & ~w14180 ) | ( w14131 & w14188 ) | ( ~w14180 & w14188 ) ;
  assign w14329 = ~\pi112 & w4654 ;
  assign w14330 = \pi111 & w4876 ;
  assign w14331 = ( w4654 & ~w14329 ) | ( w4654 & w14330 ) | ( ~w14329 & w14330 ) ;
  assign w14332 = ~\pi113 & w4656 ;
  assign w14333 = w5366 | w14331 ;
  assign w14334 = ( w4657 & w14331 ) | ( w4657 & w14333 ) | ( w14331 & w14333 ) ;
  assign w14335 = ( w4656 & ~w14332 ) | ( w4656 & w14334 ) | ( ~w14332 & w14334 ) ;
  assign w14336 = \pi047 ^ w14335 ;
  assign w14337 = w14327 ^ w14328 ;
  assign w14338 = w14336 ^ w14337 ;
  assign w14339 = ( ~w14190 & w14198 ) | ( ~w14190 & w14199 ) | ( w14198 & w14199 ) ;
  assign w14340 = ~\pi115 & w4141 ;
  assign w14341 = \pi114 & w4334 ;
  assign w14342 = ( w4141 & ~w14340 ) | ( w4141 & w14341 ) | ( ~w14340 & w14341 ) ;
  assign w14343 = ~\pi116 & w4143 ;
  assign w14344 = w5976 | w14342 ;
  assign w14345 = ( w4144 & w14342 ) | ( w4144 & w14344 ) | ( w14342 & w14344 ) ;
  assign w14346 = ( w4143 & ~w14343 ) | ( w4143 & w14345 ) | ( ~w14343 & w14345 ) ;
  assign w14347 = \pi044 ^ w14346 ;
  assign w14348 = w14338 ^ w14339 ;
  assign w14349 = w14347 ^ w14348 ;
  assign w14350 = ~\pi118 & w3635 ;
  assign w14351 = \pi117 & w3817 ;
  assign w14352 = ( w3635 & ~w14350 ) | ( w3635 & w14351 ) | ( ~w14350 & w14351 ) ;
  assign w14353 = ~\pi119 & w3637 ;
  assign w14354 = w6616 | w14352 ;
  assign w14355 = ( w3638 & w14352 ) | ( w3638 & w14354 ) | ( w14352 & w14354 ) ;
  assign w14356 = ( w3637 & ~w14353 ) | ( w3637 & w14355 ) | ( ~w14353 & w14355 ) ;
  assign w14357 = \pi041 ^ w14356 ;
  assign w14358 = w14210 ^ w14349 ;
  assign w14359 = w14357 ^ w14358 ;
  assign w14360 = w14263 ^ w14264 ;
  assign w14361 = w14359 ^ w14360 ;
  assign w14362 = ( w14128 & ~w14222 ) | ( w14128 & w14223 ) | ( ~w14222 & w14223 ) ;
  assign w14363 = w14361 ^ w14362 ;
  assign w14364 = ~\pi124 & w2712 ;
  assign w14365 = \pi123 & w2872 ;
  assign w14366 = ( w2712 & ~w14364 ) | ( w2712 & w14365 ) | ( ~w14364 & w14365 ) ;
  assign w14367 = ~\pi125 & w2714 ;
  assign w14368 = w7988 | w14366 ;
  assign w14369 = ( w2715 & w14366 ) | ( w2715 & w14368 ) | ( w14366 & w14368 ) ;
  assign w14370 = ( w2714 & ~w14367 ) | ( w2714 & w14369 ) | ( ~w14367 & w14369 ) ;
  assign w14371 = \pi035 ^ w14370 ;
  assign w14372 = w14250 ^ w14371 ;
  assign w14373 = w14255 ^ w14363 ;
  assign w14374 = \pi032 ^ w14373 ;
  assign w14375 = w14372 ^ w14374 ;
  assign w14376 = ( ~w14236 & w14237 ) | ( ~w14236 & w14245 ) | ( w14237 & w14245 ) ;
  assign w14377 = ( w14119 & ~w14120 ) | ( w14119 & w14247 ) | ( ~w14120 & w14247 ) ;
  assign w14378 = w14376 ^ w14377 ;
  assign w14379 = w14375 ^ w14378 ;
  assign w14380 = ( w14375 & ~w14376 ) | ( w14375 & w14377 ) | ( ~w14376 & w14377 ) ;
  assign w14381 = \pi032 ^ w14255 ;
  assign w14382 = w14363 ^ w14371 ;
  assign w14383 = ( w14250 & w14381 ) | ( w14250 & ~w14382 ) | ( w14381 & ~w14382 ) ;
  assign w14384 = ( ~w14361 & w14362 ) | ( ~w14361 & w14371 ) | ( w14362 & w14371 ) ;
  assign w14385 = w2313 & w8481 ;
  assign w14386 = w2443 | w14385 ;
  assign w14387 = ( \pi127 & w14385 ) | ( \pi127 & w14386 ) | ( w14385 & w14386 ) ;
  assign w14388 = \pi032 ^ w14387 ;
  assign w14389 = ( w14210 & ~w14349 ) | ( w14210 & w14357 ) | ( ~w14349 & w14357 ) ;
  assign w14390 = ~\pi119 & w3635 ;
  assign w14391 = \pi118 & w3817 ;
  assign w14392 = ( w3635 & ~w14390 ) | ( w3635 & w14391 ) | ( ~w14390 & w14391 ) ;
  assign w14393 = ~\pi120 & w3637 ;
  assign w14394 = w6634 | w14392 ;
  assign w14395 = ( w3638 & w14392 ) | ( w3638 & w14394 ) | ( w14392 & w14394 ) ;
  assign w14396 = ( w3637 & ~w14393 ) | ( w3637 & w14395 ) | ( ~w14393 & w14395 ) ;
  assign w14397 = \pi041 ^ w14396 ;
  assign w14398 = ( ~w14338 & w14339 ) | ( ~w14338 & w14347 ) | ( w14339 & w14347 ) ;
  assign w14399 = ~\pi116 & w4141 ;
  assign w14400 = \pi115 & w4334 ;
  assign w14401 = ( w4141 & ~w14399 ) | ( w4141 & w14400 ) | ( ~w14399 & w14400 ) ;
  assign w14402 = ~\pi117 & w4143 ;
  assign w14403 = w6185 | w14401 ;
  assign w14404 = ( w4144 & w14401 ) | ( w4144 & w14403 ) | ( w14401 & w14403 ) ;
  assign w14405 = ( w4143 & ~w14402 ) | ( w4143 & w14404 ) | ( ~w14402 & w14404 ) ;
  assign w14406 = \pi044 ^ w14405 ;
  assign w14407 = ( ~w14327 & w14328 ) | ( ~w14327 & w14336 ) | ( w14328 & w14336 ) ;
  assign w14408 = ( w14272 & w14273 ) | ( w14272 & ~w14314 ) | ( w14273 & ~w14314 ) ;
  assign w14409 = ~\pi107 & w5802 ;
  assign w14410 = \pi106 & w6052 ;
  assign w14411 = ( w5802 & ~w14409 ) | ( w5802 & w14410 ) | ( ~w14409 & w14410 ) ;
  assign w14412 = ~\pi108 & w5804 ;
  assign w14413 = w4425 | w14411 ;
  assign w14414 = ( w5805 & w14411 ) | ( w5805 & w14413 ) | ( w14411 & w14413 ) ;
  assign w14415 = ( w5804 & ~w14412 ) | ( w5804 & w14414 ) | ( ~w14412 & w14414 ) ;
  assign w14416 = \pi053 ^ w14415 ;
  assign w14417 = ( w14281 & w14282 ) | ( w14281 & ~w14312 ) | ( w14282 & ~w14312 ) ;
  assign w14418 = ~\pi104 & w6466 ;
  assign w14419 = \pi103 & w6702 ;
  assign w14420 = ( w6466 & ~w14418 ) | ( w6466 & w14419 ) | ( ~w14418 & w14419 ) ;
  assign w14421 = ~\pi105 & w6468 ;
  assign w14422 = w3905 | w14420 ;
  assign w14423 = ( w6469 & w14420 ) | ( w6469 & w14422 ) | ( w14420 & w14422 ) ;
  assign w14424 = ( w6468 & ~w14421 ) | ( w6468 & w14423 ) | ( ~w14421 & w14423 ) ;
  assign w14425 = \pi056 ^ w14424 ;
  assign w14426 = ( w14290 & w14291 ) | ( w14290 & ~w14310 ) | ( w14291 & ~w14310 ) ;
  assign w14427 = \pi063 & \pi094 ;
  assign w14428 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w14427 ) | ( \pi063 & w14427 ) ;
  assign w14429 = ( \pi062 & ~\pi063 ) | ( \pi062 & w14427 ) | ( ~\pi063 & w14427 ) ;
  assign w14430 = ( \pi095 & w14428 ) | ( \pi095 & w14429 ) | ( w14428 & w14429 ) ;
  assign w14431 = ( w14296 & w14304 ) | ( w14296 & ~w14430 ) | ( w14304 & ~w14430 ) ;
  assign w14432 = \pi095 & ~w14431 ;
  assign w14433 = ( \pi063 & ~\pi094 ) | ( \pi063 & w14432 ) | ( ~\pi094 & w14432 ) ;
  assign w14434 = ( \pi062 & ~\pi063 ) | ( \pi062 & w14433 ) | ( ~\pi063 & w14433 ) ;
  assign w14435 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi096 ) | ( \pi063 & ~\pi096 ) ;
  assign w14436 = ( \pi095 & w14431 ) | ( \pi095 & w14435 ) | ( w14431 & w14435 ) ;
  assign w14437 = ( ~\pi063 & w14431 ) | ( ~\pi063 & w14432 ) | ( w14431 & w14432 ) ;
  assign w14438 = ( \pi062 & ~\pi095 ) | ( \pi062 & w14437 ) | ( ~\pi095 & w14437 ) ;
  assign w14439 = ( ~w14434 & w14436 ) | ( ~w14434 & w14438 ) | ( w14436 & w14438 ) ;
  assign w14440 = \pi094 ^ \pi096 ;
  assign w14441 = ( \pi062 & \pi063 ) | ( \pi062 & ~w14440 ) | ( \pi063 & ~w14440 ) ;
  assign w14442 = \pi094 ^ \pi095 ;
  assign w14443 = \pi062 & ~w14442 ;
  assign w14444 = ( \pi063 & ~w14442 ) | ( \pi063 & w14443 ) | ( ~w14442 & w14443 ) ;
  assign w14445 = w14431 ^ w14444 ;
  assign w14446 = w14441 ^ w14445 ;
  assign w14447 = ~\pi098 & w7811 ;
  assign w14448 = \pi097 & w8046 ;
  assign w14449 = ( w7811 & ~w14447 ) | ( w7811 & w14448 ) | ( ~w14447 & w14448 ) ;
  assign w14450 = ~\pi099 & w7813 ;
  assign w14451 = w2966 | w14449 ;
  assign w14452 = ( w7814 & w14449 ) | ( w7814 & w14451 ) | ( w14449 & w14451 ) ;
  assign w14453 = ( w7813 & ~w14450 ) | ( w7813 & w14452 ) | ( ~w14450 & w14452 ) ;
  assign w14454 = \pi062 ^ w14453 ;
  assign w14455 = ~\pi101 & w7135 ;
  assign w14456 = \pi100 & w7359 ;
  assign w14457 = ( w7135 & ~w14455 ) | ( w7135 & w14456 ) | ( ~w14455 & w14456 ) ;
  assign w14458 = ~\pi102 & w7137 ;
  assign w14459 = w3284 | w14457 ;
  assign w14460 = ( w7138 & w14457 ) | ( w7138 & w14459 ) | ( w14457 & w14459 ) ;
  assign w14461 = ( w7137 & ~w14458 ) | ( w7137 & w14460 ) | ( ~w14458 & w14460 ) ;
  assign w14462 = \pi059 ^ w14461 ;
  assign w14463 = w14446 ^ w14462 ;
  assign w14464 = w14454 ^ w14463 ;
  assign w14465 = w14426 ^ w14464 ;
  assign w14466 = w14425 ^ w14465 ;
  assign w14467 = w14417 ^ w14466 ;
  assign w14468 = w14416 ^ w14467 ;
  assign w14469 = ~\pi110 & w5209 ;
  assign w14470 = \pi109 & w5433 ;
  assign w14471 = ( w5209 & ~w14469 ) | ( w5209 & w14470 ) | ( ~w14469 & w14470 ) ;
  assign w14472 = ~\pi111 & w5211 ;
  assign w14473 = w4811 | w14471 ;
  assign w14474 = ( w5212 & w14471 ) | ( w5212 & w14473 ) | ( w14471 & w14473 ) ;
  assign w14475 = ( w5211 & ~w14472 ) | ( w5211 & w14474 ) | ( ~w14472 & w14474 ) ;
  assign w14476 = \pi050 ^ w14475 ;
  assign w14477 = w14408 ^ w14468 ;
  assign w14478 = w14476 ^ w14477 ;
  assign w14479 = ( ~w14316 & w14317 ) | ( ~w14316 & w14325 ) | ( w14317 & w14325 ) ;
  assign w14480 = ~\pi113 & w4654 ;
  assign w14481 = \pi112 & w4876 ;
  assign w14482 = ( w4654 & ~w14480 ) | ( w4654 & w14481 ) | ( ~w14480 & w14481 ) ;
  assign w14483 = ~\pi114 & w4656 ;
  assign w14484 = w5565 | w14482 ;
  assign w14485 = ( w4657 & w14482 ) | ( w4657 & w14484 ) | ( w14482 & w14484 ) ;
  assign w14486 = ( w4656 & ~w14483 ) | ( w4656 & w14485 ) | ( ~w14483 & w14485 ) ;
  assign w14487 = \pi047 ^ w14486 ;
  assign w14488 = w14478 ^ w14479 ;
  assign w14489 = w14487 ^ w14488 ;
  assign w14490 = w14407 ^ w14489 ;
  assign w14491 = w14406 ^ w14490 ;
  assign w14492 = w14398 ^ w14491 ;
  assign w14493 = w14397 ^ w14492 ;
  assign w14494 = ~\pi122 & w3178 ;
  assign w14495 = \pi121 & w3340 ;
  assign w14496 = ( w3178 & ~w14494 ) | ( w3178 & w14495 ) | ( ~w14494 & w14495 ) ;
  assign w14497 = ~\pi123 & w3180 ;
  assign w14498 = w7516 | w14496 ;
  assign w14499 = ( w3181 & w14496 ) | ( w3181 & w14498 ) | ( w14496 & w14498 ) ;
  assign w14500 = ( w3180 & ~w14497 ) | ( w3180 & w14499 ) | ( ~w14497 & w14499 ) ;
  assign w14501 = \pi038 ^ w14500 ;
  assign w14502 = w14389 ^ w14501 ;
  assign w14503 = w14493 ^ w14502 ;
  assign w14504 = ( w14263 & w14264 ) | ( w14263 & ~w14359 ) | ( w14264 & ~w14359 ) ;
  assign w14505 = ~\pi125 & w2712 ;
  assign w14506 = \pi124 & w2872 ;
  assign w14507 = ( w2712 & ~w14505 ) | ( w2712 & w14506 ) | ( ~w14505 & w14506 ) ;
  assign w14508 = ~\pi126 & w2714 ;
  assign w14509 = w8231 | w14507 ;
  assign w14510 = ( w2715 & w14507 ) | ( w2715 & w14509 ) | ( w14507 & w14509 ) ;
  assign w14511 = ( w2714 & ~w14508 ) | ( w2714 & w14510 ) | ( ~w14508 & w14510 ) ;
  assign w14512 = \pi035 ^ w14511 ;
  assign w14513 = w14503 ^ w14512 ;
  assign w14514 = w14504 ^ w14513 ;
  assign w14515 = w14388 ^ w14514 ;
  assign w14516 = w14384 ^ w14515 ;
  assign w14517 = w14380 ^ w14516 ;
  assign w14518 = w14383 ^ w14517 ;
  assign w14519 = ( w14380 & ~w14383 ) | ( w14380 & w14516 ) | ( ~w14383 & w14516 ) ;
  assign w14520 = ( w14384 & w14388 ) | ( w14384 & ~w14514 ) | ( w14388 & ~w14514 ) ;
  assign w14521 = ~\pi120 & w3635 ;
  assign w14522 = \pi119 & w3817 ;
  assign w14523 = ( w3635 & ~w14521 ) | ( w3635 & w14522 ) | ( ~w14521 & w14522 ) ;
  assign w14524 = ~\pi121 & w3637 ;
  assign w14525 = w7050 | w14523 ;
  assign w14526 = ( w3638 & w14523 ) | ( w3638 & w14525 ) | ( w14523 & w14525 ) ;
  assign w14527 = ( w3637 & ~w14524 ) | ( w3637 & w14526 ) | ( ~w14524 & w14526 ) ;
  assign w14528 = \pi041 ^ w14527 ;
  assign w14529 = ( w14406 & w14407 ) | ( w14406 & ~w14489 ) | ( w14407 & ~w14489 ) ;
  assign w14530 = ( ~w14478 & w14479 ) | ( ~w14478 & w14487 ) | ( w14479 & w14487 ) ;
  assign w14531 = ~\pi105 & w6466 ;
  assign w14532 = \pi104 & w6702 ;
  assign w14533 = ( w6466 & ~w14531 ) | ( w6466 & w14532 ) | ( ~w14531 & w14532 ) ;
  assign w14534 = ~\pi106 & w6468 ;
  assign w14535 = w4068 | w14533 ;
  assign w14536 = ( w6469 & w14533 ) | ( w6469 & w14535 ) | ( w14533 & w14535 ) ;
  assign w14537 = ( w6468 & ~w14534 ) | ( w6468 & w14536 ) | ( ~w14534 & w14536 ) ;
  assign w14538 = \pi056 ^ w14537 ;
  assign w14539 = ( ~w14446 & w14454 ) | ( ~w14446 & w14462 ) | ( w14454 & w14462 ) ;
  assign w14540 = \pi095 ^ \pi097 ;
  assign w14541 = ( \pi062 & \pi063 ) | ( \pi062 & ~w14540 ) | ( \pi063 & ~w14540 ) ;
  assign w14542 = \pi095 ^ \pi096 ;
  assign w14543 = \pi062 & ~w14542 ;
  assign w14544 = ( \pi063 & ~w14542 ) | ( \pi063 & w14543 ) | ( ~w14542 & w14543 ) ;
  assign w14545 = \pi032 ^ w14544 ;
  assign w14546 = w14541 ^ w14545 ;
  assign w14547 = ~\pi099 & w7811 ;
  assign w14548 = \pi098 & w8046 ;
  assign w14549 = ( w7811 & ~w14547 ) | ( w7811 & w14548 ) | ( ~w14547 & w14548 ) ;
  assign w14550 = ~\pi100 & w7813 ;
  assign w14551 = w3104 | w14549 ;
  assign w14552 = ( w7814 & w14549 ) | ( w7814 & w14551 ) | ( w14549 & w14551 ) ;
  assign w14553 = ( w7813 & ~w14550 ) | ( w7813 & w14552 ) | ( ~w14550 & w14552 ) ;
  assign w14554 = \pi062 ^ w14553 ;
  assign w14555 = w14439 ^ w14554 ;
  assign w14556 = w14546 ^ w14555 ;
  assign w14557 = ~\pi102 & w7135 ;
  assign w14558 = \pi101 & w7359 ;
  assign w14559 = ( w7135 & ~w14557 ) | ( w7135 & w14558 ) | ( ~w14557 & w14558 ) ;
  assign w14560 = ~\pi103 & w7137 ;
  assign w14561 = w3437 | w14559 ;
  assign w14562 = ( w7138 & w14559 ) | ( w7138 & w14561 ) | ( w14559 & w14561 ) ;
  assign w14563 = ( w7137 & ~w14560 ) | ( w7137 & w14562 ) | ( ~w14560 & w14562 ) ;
  assign w14564 = \pi059 ^ w14563 ;
  assign w14565 = w14539 ^ w14556 ;
  assign w14566 = w14564 ^ w14565 ;
  assign w14567 = ( w14425 & w14426 ) | ( w14425 & ~w14464 ) | ( w14426 & ~w14464 ) ;
  assign w14568 = w14566 ^ w14567 ;
  assign w14569 = w14538 ^ w14568 ;
  assign w14570 = ~\pi108 & w5802 ;
  assign w14571 = \pi107 & w6052 ;
  assign w14572 = ( w5802 & ~w14570 ) | ( w5802 & w14571 ) | ( ~w14570 & w14571 ) ;
  assign w14573 = ~\pi109 & w5804 ;
  assign w14574 = w4599 | w14572 ;
  assign w14575 = ( w5805 & w14572 ) | ( w5805 & w14574 ) | ( w14572 & w14574 ) ;
  assign w14576 = ( w5804 & ~w14573 ) | ( w5804 & w14575 ) | ( ~w14573 & w14575 ) ;
  assign w14577 = \pi053 ^ w14576 ;
  assign w14578 = ( w14416 & w14417 ) | ( w14416 & ~w14466 ) | ( w14417 & ~w14466 ) ;
  assign w14579 = w14569 ^ w14578 ;
  assign w14580 = w14577 ^ w14579 ;
  assign w14581 = ~\pi111 & w5209 ;
  assign w14582 = \pi110 & w5433 ;
  assign w14583 = ( w5209 & ~w14581 ) | ( w5209 & w14582 ) | ( ~w14581 & w14582 ) ;
  assign w14584 = ~\pi112 & w5211 ;
  assign w14585 = w4999 | w14583 ;
  assign w14586 = ( w5212 & w14583 ) | ( w5212 & w14585 ) | ( w14583 & w14585 ) ;
  assign w14587 = ( w5211 & ~w14584 ) | ( w5211 & w14586 ) | ( ~w14584 & w14586 ) ;
  assign w14588 = \pi050 ^ w14587 ;
  assign w14589 = ( w14408 & ~w14468 ) | ( w14408 & w14476 ) | ( ~w14468 & w14476 ) ;
  assign w14590 = w14580 ^ w14589 ;
  assign w14591 = w14588 ^ w14590 ;
  assign w14592 = ~\pi114 & w4654 ;
  assign w14593 = \pi113 & w4876 ;
  assign w14594 = ( w4654 & ~w14592 ) | ( w4654 & w14593 ) | ( ~w14592 & w14593 ) ;
  assign w14595 = ~\pi115 & w4656 ;
  assign w14596 = w5585 | w14594 ;
  assign w14597 = ( w4657 & w14594 ) | ( w4657 & w14596 ) | ( w14594 & w14596 ) ;
  assign w14598 = ( w4656 & ~w14595 ) | ( w4656 & w14597 ) | ( ~w14595 & w14597 ) ;
  assign w14599 = \pi047 ^ w14598 ;
  assign w14600 = ( w14530 & ~w14591 ) | ( w14530 & w14599 ) | ( ~w14591 & w14599 ) ;
  assign w14601 = w14530 ^ w14591 ;
  assign w14602 = w14599 ^ w14601 ;
  assign w14603 = ~\pi117 & w4141 ;
  assign w14604 = \pi116 & w4334 ;
  assign w14605 = ( w4141 & ~w14603 ) | ( w4141 & w14604 ) | ( ~w14603 & w14604 ) ;
  assign w14606 = ~\pi118 & w4143 ;
  assign w14607 = w6206 | w14605 ;
  assign w14608 = ( w4144 & w14605 ) | ( w4144 & w14607 ) | ( w14605 & w14607 ) ;
  assign w14609 = ( w4143 & ~w14606 ) | ( w4143 & w14608 ) | ( ~w14606 & w14608 ) ;
  assign w14610 = \pi044 ^ w14609 ;
  assign w14611 = w14529 ^ w14602 ;
  assign w14612 = w14610 ^ w14611 ;
  assign w14613 = ( w14397 & w14398 ) | ( w14397 & ~w14491 ) | ( w14398 & ~w14491 ) ;
  assign w14614 = w14612 ^ w14613 ;
  assign w14615 = w14528 ^ w14614 ;
  assign w14616 = ~\pi123 & w3178 ;
  assign w14617 = \pi122 & w3340 ;
  assign w14618 = ( w3178 & ~w14616 ) | ( w3178 & w14617 ) | ( ~w14616 & w14617 ) ;
  assign w14619 = ~\pi124 & w3180 ;
  assign w14620 = w7538 | w14618 ;
  assign w14621 = ( w3181 & w14618 ) | ( w3181 & w14620 ) | ( w14618 & w14620 ) ;
  assign w14622 = ( w3180 & ~w14619 ) | ( w3180 & w14621 ) | ( ~w14619 & w14621 ) ;
  assign w14623 = \pi038 ^ w14622 ;
  assign w14624 = ( w14389 & ~w14493 ) | ( w14389 & w14501 ) | ( ~w14493 & w14501 ) ;
  assign w14625 = w14623 ^ w14624 ;
  assign w14626 = w14615 ^ w14625 ;
  assign w14627 = ( ~w14503 & w14504 ) | ( ~w14503 & w14512 ) | ( w14504 & w14512 ) ;
  assign w14628 = ~\pi126 & w2712 ;
  assign w14629 = \pi125 & w2872 ;
  assign w14630 = ( w2712 & ~w14628 ) | ( w2712 & w14629 ) | ( ~w14628 & w14629 ) ;
  assign w14631 = ~\pi127 & w2714 ;
  assign w14632 = w8466 | w14630 ;
  assign w14633 = ( w2715 & w14630 ) | ( w2715 & w14632 ) | ( w14630 & w14632 ) ;
  assign w14634 = ( w2714 & ~w14631 ) | ( w2714 & w14633 ) | ( ~w14631 & w14633 ) ;
  assign w14635 = \pi035 ^ w14634 ;
  assign w14636 = w14627 ^ w14635 ;
  assign w14637 = w14626 ^ w14636 ;
  assign w14638 = w14519 ^ w14520 ;
  assign w14639 = w14637 ^ w14638 ;
  assign w14640 = ( ~w14615 & w14623 ) | ( ~w14615 & w14624 ) | ( w14623 & w14624 ) ;
  assign w14641 = \pi127 & w2712 ;
  assign w14642 = ( \pi126 & ~w2715 ) | ( \pi126 & w8490 ) | ( ~w2715 & w8490 ) ;
  assign w14643 = \pi126 & ~w2872 ;
  assign w14644 = ( ~\pi126 & w14642 ) | ( ~\pi126 & w14643 ) | ( w14642 & w14643 ) ;
  assign w14645 = ( w9420 & w14641 ) | ( w9420 & ~w14644 ) | ( w14641 & ~w14644 ) ;
  assign w14646 = ~\pi121 & w3635 ;
  assign w14647 = \pi120 & w3817 ;
  assign w14648 = ( w3635 & ~w14646 ) | ( w3635 & w14647 ) | ( ~w14646 & w14647 ) ;
  assign w14649 = ~\pi122 & w3637 ;
  assign w14650 = w7069 | w14648 ;
  assign w14651 = ( w3638 & w14648 ) | ( w3638 & w14650 ) | ( w14648 & w14650 ) ;
  assign w14652 = ( w3637 & ~w14649 ) | ( w3637 & w14651 ) | ( ~w14649 & w14651 ) ;
  assign w14653 = \pi041 ^ w14652 ;
  assign w14654 = ( w14529 & ~w14602 ) | ( w14529 & w14610 ) | ( ~w14602 & w14610 ) ;
  assign w14655 = ~\pi106 & w6466 ;
  assign w14656 = \pi105 & w6702 ;
  assign w14657 = ( w6466 & ~w14655 ) | ( w6466 & w14656 ) | ( ~w14655 & w14656 ) ;
  assign w14658 = ~\pi107 & w6468 ;
  assign w14659 = w4087 | w14657 ;
  assign w14660 = ( w6469 & w14657 ) | ( w6469 & w14659 ) | ( w14657 & w14659 ) ;
  assign w14661 = ( w6468 & ~w14658 ) | ( w6468 & w14660 ) | ( ~w14658 & w14660 ) ;
  assign w14662 = \pi056 ^ w14661 ;
  assign w14663 = ( w14539 & ~w14556 ) | ( w14539 & w14564 ) | ( ~w14556 & w14564 ) ;
  assign w14664 = ~\pi103 & w7135 ;
  assign w14665 = \pi102 & w7359 ;
  assign w14666 = ( w7135 & ~w14664 ) | ( w7135 & w14665 ) | ( ~w14664 & w14665 ) ;
  assign w14667 = ~\pi104 & w7137 ;
  assign w14668 = w3740 | w14666 ;
  assign w14669 = ( w7138 & w14666 ) | ( w7138 & w14668 ) | ( w14666 & w14668 ) ;
  assign w14670 = ( w7137 & ~w14667 ) | ( w7137 & w14669 ) | ( ~w14667 & w14669 ) ;
  assign w14671 = \pi059 ^ w14670 ;
  assign w14672 = ( w14439 & ~w14546 ) | ( w14439 & w14554 ) | ( ~w14546 & w14554 ) ;
  assign w14673 = \pi063 ^ \pi095 ;
  assign w14674 = \pi062 ^ w14673 ;
  assign w14675 = ( \pi095 & \pi097 ) | ( \pi095 & w14674 ) | ( \pi097 & w14674 ) ;
  assign w14676 = ( ~\pi032 & \pi096 ) | ( ~\pi032 & w14675 ) | ( \pi096 & w14675 ) ;
  assign w14677 = w10655 & w14676 ;
  assign w14678 = ~\pi100 & w7811 ;
  assign w14679 = \pi099 & w8046 ;
  assign w14680 = ( w7811 & ~w14678 ) | ( w7811 & w14679 ) | ( ~w14678 & w14679 ) ;
  assign w14681 = ~\pi101 & w7813 ;
  assign w14682 = w3264 | w14680 ;
  assign w14683 = ( w7814 & w14680 ) | ( w7814 & w14682 ) | ( w14680 & w14682 ) ;
  assign w14684 = ( w7813 & ~w14681 ) | ( w7813 & w14683 ) | ( ~w14681 & w14683 ) ;
  assign w14685 = \pi062 ^ w14684 ;
  assign w14686 = w14677 ^ w14685 ;
  assign w14687 = ( \pi062 & \pi063 ) | ( \pi062 & \pi098 ) | ( \pi063 & \pi098 ) ;
  assign w14688 = \pi063 & ~\pi097 ;
  assign w14689 = \pi062 & w14688 ;
  assign w14690 = w14687 ^ w14689 ;
  assign w14691 = w14686 ^ w14690 ;
  assign w14692 = w14671 ^ w14672 ;
  assign w14693 = w14691 ^ w14692 ;
  assign w14694 = w14663 ^ w14693 ;
  assign w14695 = w14662 ^ w14694 ;
  assign w14696 = ( w14538 & ~w14566 ) | ( w14538 & w14567 ) | ( ~w14566 & w14567 ) ;
  assign w14697 = ~\pi109 & w5802 ;
  assign w14698 = \pi108 & w6052 ;
  assign w14699 = ( w5802 & ~w14697 ) | ( w5802 & w14698 ) | ( ~w14697 & w14698 ) ;
  assign w14700 = ~\pi110 & w5804 ;
  assign w14701 = w4792 | w14699 ;
  assign w14702 = ( w5805 & w14699 ) | ( w5805 & w14701 ) | ( w14699 & w14701 ) ;
  assign w14703 = ( w5804 & ~w14700 ) | ( w5804 & w14702 ) | ( ~w14700 & w14702 ) ;
  assign w14704 = \pi053 ^ w14703 ;
  assign w14705 = w14695 ^ w14696 ;
  assign w14706 = w14704 ^ w14705 ;
  assign w14707 = ( ~w14569 & w14577 ) | ( ~w14569 & w14578 ) | ( w14577 & w14578 ) ;
  assign w14708 = ~\pi112 & w5209 ;
  assign w14709 = \pi111 & w5433 ;
  assign w14710 = ( w5209 & ~w14708 ) | ( w5209 & w14709 ) | ( ~w14708 & w14709 ) ;
  assign w14711 = ~\pi113 & w5211 ;
  assign w14712 = w5366 | w14710 ;
  assign w14713 = ( w5212 & w14710 ) | ( w5212 & w14712 ) | ( w14710 & w14712 ) ;
  assign w14714 = ( w5211 & ~w14711 ) | ( w5211 & w14713 ) | ( ~w14711 & w14713 ) ;
  assign w14715 = \pi050 ^ w14714 ;
  assign w14716 = w14706 ^ w14707 ;
  assign w14717 = w14715 ^ w14716 ;
  assign w14718 = ( ~w14580 & w14588 ) | ( ~w14580 & w14589 ) | ( w14588 & w14589 ) ;
  assign w14719 = ~\pi115 & w4654 ;
  assign w14720 = \pi114 & w4876 ;
  assign w14721 = ( w4654 & ~w14719 ) | ( w4654 & w14720 ) | ( ~w14719 & w14720 ) ;
  assign w14722 = ~\pi116 & w4656 ;
  assign w14723 = w5976 | w14721 ;
  assign w14724 = ( w4657 & w14721 ) | ( w4657 & w14723 ) | ( w14721 & w14723 ) ;
  assign w14725 = ( w4656 & ~w14722 ) | ( w4656 & w14724 ) | ( ~w14722 & w14724 ) ;
  assign w14726 = \pi047 ^ w14725 ;
  assign w14727 = w14717 ^ w14718 ;
  assign w14728 = w14726 ^ w14727 ;
  assign w14729 = ~\pi118 & w4141 ;
  assign w14730 = \pi117 & w4334 ;
  assign w14731 = ( w4141 & ~w14729 ) | ( w4141 & w14730 ) | ( ~w14729 & w14730 ) ;
  assign w14732 = ~\pi119 & w4143 ;
  assign w14733 = w6616 | w14731 ;
  assign w14734 = ( w4144 & w14731 ) | ( w4144 & w14733 ) | ( w14731 & w14733 ) ;
  assign w14735 = ( w4143 & ~w14732 ) | ( w4143 & w14734 ) | ( ~w14732 & w14734 ) ;
  assign w14736 = \pi044 ^ w14735 ;
  assign w14737 = w14600 ^ w14728 ;
  assign w14738 = w14736 ^ w14737 ;
  assign w14739 = w14653 ^ w14654 ;
  assign w14740 = w14738 ^ w14739 ;
  assign w14741 = ( w14528 & ~w14612 ) | ( w14528 & w14613 ) | ( ~w14612 & w14613 ) ;
  assign w14742 = w14740 ^ w14741 ;
  assign w14743 = ~\pi124 & w3178 ;
  assign w14744 = \pi123 & w3340 ;
  assign w14745 = ( w3178 & ~w14743 ) | ( w3178 & w14744 ) | ( ~w14743 & w14744 ) ;
  assign w14746 = ~\pi125 & w3180 ;
  assign w14747 = w7988 | w14745 ;
  assign w14748 = ( w3181 & w14745 ) | ( w3181 & w14747 ) | ( w14745 & w14747 ) ;
  assign w14749 = ( w3180 & ~w14746 ) | ( w3180 & w14748 ) | ( ~w14746 & w14748 ) ;
  assign w14750 = \pi038 ^ w14749 ;
  assign w14751 = w14640 ^ w14750 ;
  assign w14752 = w14645 ^ w14742 ;
  assign w14753 = \pi035 ^ w14752 ;
  assign w14754 = w14751 ^ w14753 ;
  assign w14755 = ( ~w14626 & w14627 ) | ( ~w14626 & w14635 ) | ( w14627 & w14635 ) ;
  assign w14756 = ( w14519 & ~w14520 ) | ( w14519 & w14637 ) | ( ~w14520 & w14637 ) ;
  assign w14757 = w14755 ^ w14756 ;
  assign w14758 = w14754 ^ w14757 ;
  assign w14759 = ( w14754 & ~w14755 ) | ( w14754 & w14756 ) | ( ~w14755 & w14756 ) ;
  assign w14760 = \pi035 ^ w14645 ;
  assign w14761 = w14742 ^ w14750 ;
  assign w14762 = ( w14640 & w14760 ) | ( w14640 & ~w14761 ) | ( w14760 & ~w14761 ) ;
  assign w14763 = ( ~w14740 & w14741 ) | ( ~w14740 & w14750 ) | ( w14741 & w14750 ) ;
  assign w14764 = w2715 & w8481 ;
  assign w14765 = w2872 | w14764 ;
  assign w14766 = ( \pi127 & w14764 ) | ( \pi127 & w14765 ) | ( w14764 & w14765 ) ;
  assign w14767 = \pi035 ^ w14766 ;
  assign w14768 = ( w14600 & ~w14728 ) | ( w14600 & w14736 ) | ( ~w14728 & w14736 ) ;
  assign w14769 = ~\pi119 & w4141 ;
  assign w14770 = \pi118 & w4334 ;
  assign w14771 = ( w4141 & ~w14769 ) | ( w4141 & w14770 ) | ( ~w14769 & w14770 ) ;
  assign w14772 = ~\pi120 & w4143 ;
  assign w14773 = w6634 | w14771 ;
  assign w14774 = ( w4144 & w14771 ) | ( w4144 & w14773 ) | ( w14771 & w14773 ) ;
  assign w14775 = ( w4143 & ~w14772 ) | ( w4143 & w14774 ) | ( ~w14772 & w14774 ) ;
  assign w14776 = \pi044 ^ w14775 ;
  assign w14777 = ( ~w14717 & w14718 ) | ( ~w14717 & w14726 ) | ( w14718 & w14726 ) ;
  assign w14778 = ~\pi116 & w4654 ;
  assign w14779 = \pi115 & w4876 ;
  assign w14780 = ( w4654 & ~w14778 ) | ( w4654 & w14779 ) | ( ~w14778 & w14779 ) ;
  assign w14781 = ~\pi117 & w4656 ;
  assign w14782 = w6185 | w14780 ;
  assign w14783 = ( w4657 & w14780 ) | ( w4657 & w14782 ) | ( w14780 & w14782 ) ;
  assign w14784 = ( w4656 & ~w14781 ) | ( w4656 & w14783 ) | ( ~w14781 & w14783 ) ;
  assign w14785 = \pi047 ^ w14784 ;
  assign w14786 = ( ~w14706 & w14707 ) | ( ~w14706 & w14715 ) | ( w14707 & w14715 ) ;
  assign w14787 = ( w14662 & w14663 ) | ( w14662 & ~w14693 ) | ( w14663 & ~w14693 ) ;
  assign w14788 = ~\pi107 & w6466 ;
  assign w14789 = \pi106 & w6702 ;
  assign w14790 = ( w6466 & ~w14788 ) | ( w6466 & w14789 ) | ( ~w14788 & w14789 ) ;
  assign w14791 = ~\pi108 & w6468 ;
  assign w14792 = w4425 | w14790 ;
  assign w14793 = ( w6469 & w14790 ) | ( w6469 & w14792 ) | ( w14790 & w14792 ) ;
  assign w14794 = ( w6468 & ~w14791 ) | ( w6468 & w14793 ) | ( ~w14791 & w14793 ) ;
  assign w14795 = \pi056 ^ w14794 ;
  assign w14796 = ( w14671 & w14672 ) | ( w14671 & ~w14691 ) | ( w14672 & ~w14691 ) ;
  assign w14797 = \pi063 & \pi097 ;
  assign w14798 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w14797 ) | ( \pi063 & w14797 ) ;
  assign w14799 = ( \pi062 & ~\pi063 ) | ( \pi062 & w14797 ) | ( ~\pi063 & w14797 ) ;
  assign w14800 = ( \pi098 & w14798 ) | ( \pi098 & w14799 ) | ( w14798 & w14799 ) ;
  assign w14801 = ( w14677 & w14685 ) | ( w14677 & ~w14800 ) | ( w14685 & ~w14800 ) ;
  assign w14802 = \pi098 & ~w14801 ;
  assign w14803 = ( \pi063 & ~\pi097 ) | ( \pi063 & w14802 ) | ( ~\pi097 & w14802 ) ;
  assign w14804 = ( \pi062 & ~\pi063 ) | ( \pi062 & w14803 ) | ( ~\pi063 & w14803 ) ;
  assign w14805 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi099 ) | ( \pi063 & ~\pi099 ) ;
  assign w14806 = ( \pi098 & w14801 ) | ( \pi098 & w14805 ) | ( w14801 & w14805 ) ;
  assign w14807 = ( ~\pi063 & w14801 ) | ( ~\pi063 & w14802 ) | ( w14801 & w14802 ) ;
  assign w14808 = ( \pi062 & ~\pi098 ) | ( \pi062 & w14807 ) | ( ~\pi098 & w14807 ) ;
  assign w14809 = ( ~w14804 & w14806 ) | ( ~w14804 & w14808 ) | ( w14806 & w14808 ) ;
  assign w14810 = \pi097 ^ \pi099 ;
  assign w14811 = ( \pi062 & \pi063 ) | ( \pi062 & ~w14810 ) | ( \pi063 & ~w14810 ) ;
  assign w14812 = \pi097 ^ \pi098 ;
  assign w14813 = \pi062 & ~w14812 ;
  assign w14814 = ( \pi063 & ~w14812 ) | ( \pi063 & w14813 ) | ( ~w14812 & w14813 ) ;
  assign w14815 = w14801 ^ w14814 ;
  assign w14816 = w14811 ^ w14815 ;
  assign w14817 = ~\pi101 & w7811 ;
  assign w14818 = \pi100 & w8046 ;
  assign w14819 = ( w7811 & ~w14817 ) | ( w7811 & w14818 ) | ( ~w14817 & w14818 ) ;
  assign w14820 = ~\pi102 & w7813 ;
  assign w14821 = w3284 | w14819 ;
  assign w14822 = ( w7814 & w14819 ) | ( w7814 & w14821 ) | ( w14819 & w14821 ) ;
  assign w14823 = ( w7813 & ~w14820 ) | ( w7813 & w14822 ) | ( ~w14820 & w14822 ) ;
  assign w14824 = \pi062 ^ w14823 ;
  assign w14825 = ~\pi104 & w7135 ;
  assign w14826 = \pi103 & w7359 ;
  assign w14827 = ( w7135 & ~w14825 ) | ( w7135 & w14826 ) | ( ~w14825 & w14826 ) ;
  assign w14828 = ~\pi105 & w7137 ;
  assign w14829 = w3905 | w14827 ;
  assign w14830 = ( w7138 & w14827 ) | ( w7138 & w14829 ) | ( w14827 & w14829 ) ;
  assign w14831 = ( w7137 & ~w14828 ) | ( w7137 & w14830 ) | ( ~w14828 & w14830 ) ;
  assign w14832 = \pi059 ^ w14831 ;
  assign w14833 = w14816 ^ w14824 ;
  assign w14834 = w14832 ^ w14833 ;
  assign w14835 = w14796 ^ w14834 ;
  assign w14836 = w14795 ^ w14835 ;
  assign w14837 = ~\pi110 & w5802 ;
  assign w14838 = \pi109 & w6052 ;
  assign w14839 = ( w5802 & ~w14837 ) | ( w5802 & w14838 ) | ( ~w14837 & w14838 ) ;
  assign w14840 = ~\pi111 & w5804 ;
  assign w14841 = w4811 | w14839 ;
  assign w14842 = ( w5805 & w14839 ) | ( w5805 & w14841 ) | ( w14839 & w14841 ) ;
  assign w14843 = ( w5804 & ~w14840 ) | ( w5804 & w14842 ) | ( ~w14840 & w14842 ) ;
  assign w14844 = \pi053 ^ w14843 ;
  assign w14845 = w14787 ^ w14836 ;
  assign w14846 = w14844 ^ w14845 ;
  assign w14847 = ( ~w14695 & w14696 ) | ( ~w14695 & w14704 ) | ( w14696 & w14704 ) ;
  assign w14848 = ~\pi113 & w5209 ;
  assign w14849 = \pi112 & w5433 ;
  assign w14850 = ( w5209 & ~w14848 ) | ( w5209 & w14849 ) | ( ~w14848 & w14849 ) ;
  assign w14851 = ~\pi114 & w5211 ;
  assign w14852 = w5565 | w14850 ;
  assign w14853 = ( w5212 & w14850 ) | ( w5212 & w14852 ) | ( w14850 & w14852 ) ;
  assign w14854 = ( w5211 & ~w14851 ) | ( w5211 & w14853 ) | ( ~w14851 & w14853 ) ;
  assign w14855 = \pi050 ^ w14854 ;
  assign w14856 = w14846 ^ w14847 ;
  assign w14857 = w14855 ^ w14856 ;
  assign w14858 = w14786 ^ w14857 ;
  assign w14859 = w14785 ^ w14858 ;
  assign w14860 = w14777 ^ w14859 ;
  assign w14861 = w14776 ^ w14860 ;
  assign w14862 = ~\pi122 & w3635 ;
  assign w14863 = \pi121 & w3817 ;
  assign w14864 = ( w3635 & ~w14862 ) | ( w3635 & w14863 ) | ( ~w14862 & w14863 ) ;
  assign w14865 = ~\pi123 & w3637 ;
  assign w14866 = w7516 | w14864 ;
  assign w14867 = ( w3638 & w14864 ) | ( w3638 & w14866 ) | ( w14864 & w14866 ) ;
  assign w14868 = ( w3637 & ~w14865 ) | ( w3637 & w14867 ) | ( ~w14865 & w14867 ) ;
  assign w14869 = \pi041 ^ w14868 ;
  assign w14870 = w14768 ^ w14869 ;
  assign w14871 = w14861 ^ w14870 ;
  assign w14872 = ( w14653 & w14654 ) | ( w14653 & ~w14738 ) | ( w14654 & ~w14738 ) ;
  assign w14873 = ~\pi125 & w3178 ;
  assign w14874 = \pi124 & w3340 ;
  assign w14875 = ( w3178 & ~w14873 ) | ( w3178 & w14874 ) | ( ~w14873 & w14874 ) ;
  assign w14876 = ~\pi126 & w3180 ;
  assign w14877 = w8231 | w14875 ;
  assign w14878 = ( w3181 & w14875 ) | ( w3181 & w14877 ) | ( w14875 & w14877 ) ;
  assign w14879 = ( w3180 & ~w14876 ) | ( w3180 & w14878 ) | ( ~w14876 & w14878 ) ;
  assign w14880 = \pi038 ^ w14879 ;
  assign w14881 = w14871 ^ w14880 ;
  assign w14882 = w14872 ^ w14881 ;
  assign w14883 = w14767 ^ w14882 ;
  assign w14884 = w14763 ^ w14883 ;
  assign w14885 = w14759 ^ w14884 ;
  assign w14886 = w14762 ^ w14885 ;
  assign w14887 = ( w14759 & ~w14762 ) | ( w14759 & w14884 ) | ( ~w14762 & w14884 ) ;
  assign w14888 = ( w14785 & w14786 ) | ( w14785 & ~w14857 ) | ( w14786 & ~w14857 ) ;
  assign w14889 = ~\pi117 & w4654 ;
  assign w14890 = \pi116 & w4876 ;
  assign w14891 = ( w4654 & ~w14889 ) | ( w4654 & w14890 ) | ( ~w14889 & w14890 ) ;
  assign w14892 = ~\pi118 & w4656 ;
  assign w14893 = w6206 | w14891 ;
  assign w14894 = ( w4657 & w14891 ) | ( w4657 & w14893 ) | ( w14891 & w14893 ) ;
  assign w14895 = ( w4656 & ~w14892 ) | ( w4656 & w14894 ) | ( ~w14892 & w14894 ) ;
  assign w14896 = \pi047 ^ w14895 ;
  assign w14897 = ( ~w14846 & w14847 ) | ( ~w14846 & w14855 ) | ( w14847 & w14855 ) ;
  assign w14898 = \pi098 ^ \pi100 ;
  assign w14899 = ( \pi062 & \pi063 ) | ( \pi062 & ~w14898 ) | ( \pi063 & ~w14898 ) ;
  assign w14900 = \pi098 ^ \pi099 ;
  assign w14901 = \pi062 & ~w14900 ;
  assign w14902 = ( \pi063 & ~w14900 ) | ( \pi063 & w14901 ) | ( ~w14900 & w14901 ) ;
  assign w14903 = \pi035 ^ w14902 ;
  assign w14904 = w14899 ^ w14903 ;
  assign w14905 = ~\pi102 & w7811 ;
  assign w14906 = \pi101 & w8046 ;
  assign w14907 = ( w7811 & ~w14905 ) | ( w7811 & w14906 ) | ( ~w14905 & w14906 ) ;
  assign w14908 = ~\pi103 & w7813 ;
  assign w14909 = w3437 | w14907 ;
  assign w14910 = ( w7814 & w14907 ) | ( w7814 & w14909 ) | ( w14907 & w14909 ) ;
  assign w14911 = ( w7813 & ~w14908 ) | ( w7813 & w14910 ) | ( ~w14908 & w14910 ) ;
  assign w14912 = \pi062 ^ w14911 ;
  assign w14913 = w14809 ^ w14912 ;
  assign w14914 = w14904 ^ w14913 ;
  assign w14915 = ~\pi105 & w7135 ;
  assign w14916 = \pi104 & w7359 ;
  assign w14917 = ( w7135 & ~w14915 ) | ( w7135 & w14916 ) | ( ~w14915 & w14916 ) ;
  assign w14918 = ~\pi106 & w7137 ;
  assign w14919 = w4068 | w14917 ;
  assign w14920 = ( w7138 & w14917 ) | ( w7138 & w14919 ) | ( w14917 & w14919 ) ;
  assign w14921 = ( w7137 & ~w14918 ) | ( w7137 & w14920 ) | ( ~w14918 & w14920 ) ;
  assign w14922 = \pi059 ^ w14921 ;
  assign w14923 = ( ~w14816 & w14824 ) | ( ~w14816 & w14832 ) | ( w14824 & w14832 ) ;
  assign w14924 = w14914 ^ w14923 ;
  assign w14925 = w14922 ^ w14924 ;
  assign w14926 = ~\pi108 & w6466 ;
  assign w14927 = \pi107 & w6702 ;
  assign w14928 = ( w6466 & ~w14926 ) | ( w6466 & w14927 ) | ( ~w14926 & w14927 ) ;
  assign w14929 = ~\pi109 & w6468 ;
  assign w14930 = w4599 | w14928 ;
  assign w14931 = ( w6469 & w14928 ) | ( w6469 & w14930 ) | ( w14928 & w14930 ) ;
  assign w14932 = ( w6468 & ~w14929 ) | ( w6468 & w14931 ) | ( ~w14929 & w14931 ) ;
  assign w14933 = \pi056 ^ w14932 ;
  assign w14934 = ( w14795 & w14796 ) | ( w14795 & ~w14834 ) | ( w14796 & ~w14834 ) ;
  assign w14935 = w14925 ^ w14934 ;
  assign w14936 = w14933 ^ w14935 ;
  assign w14937 = ~\pi111 & w5802 ;
  assign w14938 = \pi110 & w6052 ;
  assign w14939 = ( w5802 & ~w14937 ) | ( w5802 & w14938 ) | ( ~w14937 & w14938 ) ;
  assign w14940 = ~\pi112 & w5804 ;
  assign w14941 = w4999 | w14939 ;
  assign w14942 = ( w5805 & w14939 ) | ( w5805 & w14941 ) | ( w14939 & w14941 ) ;
  assign w14943 = ( w5804 & ~w14940 ) | ( w5804 & w14942 ) | ( ~w14940 & w14942 ) ;
  assign w14944 = \pi053 ^ w14943 ;
  assign w14945 = ( w14787 & ~w14836 ) | ( w14787 & w14844 ) | ( ~w14836 & w14844 ) ;
  assign w14946 = w14936 ^ w14945 ;
  assign w14947 = w14944 ^ w14946 ;
  assign w14948 = ~\pi114 & w5209 ;
  assign w14949 = \pi113 & w5433 ;
  assign w14950 = ( w5209 & ~w14948 ) | ( w5209 & w14949 ) | ( ~w14948 & w14949 ) ;
  assign w14951 = ~\pi115 & w5211 ;
  assign w14952 = w5585 | w14950 ;
  assign w14953 = ( w5212 & w14950 ) | ( w5212 & w14952 ) | ( w14950 & w14952 ) ;
  assign w14954 = ( w5211 & ~w14951 ) | ( w5211 & w14953 ) | ( ~w14951 & w14953 ) ;
  assign w14955 = \pi050 ^ w14954 ;
  assign w14956 = w14897 ^ w14947 ;
  assign w14957 = w14955 ^ w14956 ;
  assign w14958 = w14888 ^ w14957 ;
  assign w14959 = w14896 ^ w14958 ;
  assign w14960 = ~\pi120 & w4141 ;
  assign w14961 = \pi119 & w4334 ;
  assign w14962 = ( w4141 & ~w14960 ) | ( w4141 & w14961 ) | ( ~w14960 & w14961 ) ;
  assign w14963 = ~\pi121 & w4143 ;
  assign w14964 = w7050 | w14962 ;
  assign w14965 = ( w4144 & w14962 ) | ( w4144 & w14964 ) | ( w14962 & w14964 ) ;
  assign w14966 = ( w4143 & ~w14963 ) | ( w4143 & w14965 ) | ( ~w14963 & w14965 ) ;
  assign w14967 = \pi044 ^ w14966 ;
  assign w14968 = ( w14776 & w14777 ) | ( w14776 & ~w14859 ) | ( w14777 & ~w14859 ) ;
  assign w14969 = w14959 ^ w14968 ;
  assign w14970 = w14967 ^ w14969 ;
  assign w14971 = ~\pi123 & w3635 ;
  assign w14972 = \pi122 & w3817 ;
  assign w14973 = ( w3635 & ~w14971 ) | ( w3635 & w14972 ) | ( ~w14971 & w14972 ) ;
  assign w14974 = ~\pi124 & w3637 ;
  assign w14975 = w7538 | w14973 ;
  assign w14976 = ( w3638 & w14973 ) | ( w3638 & w14975 ) | ( w14973 & w14975 ) ;
  assign w14977 = ( w3637 & ~w14974 ) | ( w3637 & w14976 ) | ( ~w14974 & w14976 ) ;
  assign w14978 = \pi041 ^ w14977 ;
  assign w14979 = ( w14768 & ~w14861 ) | ( w14768 & w14869 ) | ( ~w14861 & w14869 ) ;
  assign w14980 = w14978 ^ w14979 ;
  assign w14981 = w14970 ^ w14980 ;
  assign w14982 = ~\pi126 & w3178 ;
  assign w14983 = \pi125 & w3340 ;
  assign w14984 = ( w3178 & ~w14982 ) | ( w3178 & w14983 ) | ( ~w14982 & w14983 ) ;
  assign w14985 = ~\pi127 & w3180 ;
  assign w14986 = w8466 | w14984 ;
  assign w14987 = ( w3181 & w14984 ) | ( w3181 & w14986 ) | ( w14984 & w14986 ) ;
  assign w14988 = ( w3180 & ~w14985 ) | ( w3180 & w14987 ) | ( ~w14985 & w14987 ) ;
  assign w14989 = \pi038 ^ w14988 ;
  assign w14990 = ( ~w14871 & w14872 ) | ( ~w14871 & w14880 ) | ( w14872 & w14880 ) ;
  assign w14991 = w14989 ^ w14990 ;
  assign w14992 = w14981 ^ w14991 ;
  assign w14993 = ( w14763 & w14767 ) | ( w14763 & ~w14882 ) | ( w14767 & ~w14882 ) ;
  assign w14994 = w14887 ^ w14992 ;
  assign w14995 = w14993 ^ w14994 ;
  assign w14996 = ( ~w14970 & w14978 ) | ( ~w14970 & w14979 ) | ( w14978 & w14979 ) ;
  assign w14997 = \pi127 & w3178 ;
  assign w14998 = ( \pi126 & ~w3181 ) | ( \pi126 & w8490 ) | ( ~w3181 & w8490 ) ;
  assign w14999 = \pi126 & ~w3340 ;
  assign w15000 = ( ~\pi126 & w14998 ) | ( ~\pi126 & w14999 ) | ( w14998 & w14999 ) ;
  assign w15001 = ( w9420 & w14997 ) | ( w9420 & ~w15000 ) | ( w14997 & ~w15000 ) ;
  assign w15002 = ~\pi103 & w7811 ;
  assign w15003 = \pi102 & w8046 ;
  assign w15004 = ( w7811 & ~w15002 ) | ( w7811 & w15003 ) | ( ~w15002 & w15003 ) ;
  assign w15005 = ~\pi104 & w7813 ;
  assign w15006 = w3740 | w15004 ;
  assign w15007 = ( w7814 & w15004 ) | ( w7814 & w15006 ) | ( w15004 & w15006 ) ;
  assign w15008 = ( w7813 & ~w15005 ) | ( w7813 & w15007 ) | ( ~w15005 & w15007 ) ;
  assign w15009 = \pi062 ^ w15008 ;
  assign w15010 = ( \pi062 & \pi063 ) | ( \pi062 & \pi101 ) | ( \pi063 & \pi101 ) ;
  assign w15011 = \pi063 & ~\pi100 ;
  assign w15012 = w15010 & ~w15011 ;
  assign w15013 = ( ~\pi062 & w15010 ) | ( ~\pi062 & w15012 ) | ( w15010 & w15012 ) ;
  assign w15014 = \pi063 ^ \pi098 ;
  assign w15015 = \pi062 ^ w15014 ;
  assign w15016 = ( \pi098 & \pi100 ) | ( \pi098 & w15015 ) | ( \pi100 & w15015 ) ;
  assign w15017 = ( ~\pi035 & \pi099 ) | ( ~\pi035 & w15016 ) | ( \pi099 & w15016 ) ;
  assign w15018 = w10655 & w15017 ;
  assign w15019 = w15009 ^ w15013 ;
  assign w15020 = w15018 ^ w15019 ;
  assign w15021 = ( w14809 & ~w14904 ) | ( w14809 & w14912 ) | ( ~w14904 & w14912 ) ;
  assign w15022 = ~\pi106 & w7135 ;
  assign w15023 = \pi105 & w7359 ;
  assign w15024 = ( w7135 & ~w15022 ) | ( w7135 & w15023 ) | ( ~w15022 & w15023 ) ;
  assign w15025 = ~\pi107 & w7137 ;
  assign w15026 = w4087 | w15024 ;
  assign w15027 = ( w7138 & w15024 ) | ( w7138 & w15026 ) | ( w15024 & w15026 ) ;
  assign w15028 = ( w7137 & ~w15025 ) | ( w7137 & w15027 ) | ( ~w15025 & w15027 ) ;
  assign w15029 = \pi059 ^ w15028 ;
  assign w15030 = w15020 ^ w15021 ;
  assign w15031 = w15029 ^ w15030 ;
  assign w15032 = ( ~w14914 & w14922 ) | ( ~w14914 & w14923 ) | ( w14922 & w14923 ) ;
  assign w15033 = ~\pi109 & w6466 ;
  assign w15034 = \pi108 & w6702 ;
  assign w15035 = ( w6466 & ~w15033 ) | ( w6466 & w15034 ) | ( ~w15033 & w15034 ) ;
  assign w15036 = ~\pi110 & w6468 ;
  assign w15037 = w4792 | w15035 ;
  assign w15038 = ( w6469 & w15035 ) | ( w6469 & w15037 ) | ( w15035 & w15037 ) ;
  assign w15039 = ( w6468 & ~w15036 ) | ( w6468 & w15038 ) | ( ~w15036 & w15038 ) ;
  assign w15040 = \pi056 ^ w15039 ;
  assign w15041 = w15031 ^ w15032 ;
  assign w15042 = w15040 ^ w15041 ;
  assign w15043 = ( ~w14925 & w14933 ) | ( ~w14925 & w14934 ) | ( w14933 & w14934 ) ;
  assign w15044 = ~\pi112 & w5802 ;
  assign w15045 = \pi111 & w6052 ;
  assign w15046 = ( w5802 & ~w15044 ) | ( w5802 & w15045 ) | ( ~w15044 & w15045 ) ;
  assign w15047 = ~\pi113 & w5804 ;
  assign w15048 = w5366 | w15046 ;
  assign w15049 = ( w5805 & w15046 ) | ( w5805 & w15048 ) | ( w15046 & w15048 ) ;
  assign w15050 = ( w5804 & ~w15047 ) | ( w5804 & w15049 ) | ( ~w15047 & w15049 ) ;
  assign w15051 = \pi053 ^ w15050 ;
  assign w15052 = w15042 ^ w15043 ;
  assign w15053 = w15051 ^ w15052 ;
  assign w15054 = ( ~w14936 & w14944 ) | ( ~w14936 & w14945 ) | ( w14944 & w14945 ) ;
  assign w15055 = ~\pi115 & w5209 ;
  assign w15056 = \pi114 & w5433 ;
  assign w15057 = ( w5209 & ~w15055 ) | ( w5209 & w15056 ) | ( ~w15055 & w15056 ) ;
  assign w15058 = ~\pi116 & w5211 ;
  assign w15059 = w5976 | w15057 ;
  assign w15060 = ( w5212 & w15057 ) | ( w5212 & w15059 ) | ( w15057 & w15059 ) ;
  assign w15061 = ( w5211 & ~w15058 ) | ( w5211 & w15060 ) | ( ~w15058 & w15060 ) ;
  assign w15062 = \pi050 ^ w15061 ;
  assign w15063 = w15053 ^ w15054 ;
  assign w15064 = w15062 ^ w15063 ;
  assign w15065 = ( w14897 & ~w14947 ) | ( w14897 & w14955 ) | ( ~w14947 & w14955 ) ;
  assign w15066 = ~\pi118 & w4654 ;
  assign w15067 = \pi117 & w4876 ;
  assign w15068 = ( w4654 & ~w15066 ) | ( w4654 & w15067 ) | ( ~w15066 & w15067 ) ;
  assign w15069 = ~\pi119 & w4656 ;
  assign w15070 = w6616 | w15068 ;
  assign w15071 = ( w4657 & w15068 ) | ( w4657 & w15070 ) | ( w15068 & w15070 ) ;
  assign w15072 = ( w4656 & ~w15069 ) | ( w4656 & w15071 ) | ( ~w15069 & w15071 ) ;
  assign w15073 = \pi047 ^ w15072 ;
  assign w15074 = w15064 ^ w15065 ;
  assign w15075 = w15073 ^ w15074 ;
  assign w15076 = ( w14888 & w14896 ) | ( w14888 & ~w14957 ) | ( w14896 & ~w14957 ) ;
  assign w15077 = ~\pi121 & w4141 ;
  assign w15078 = \pi120 & w4334 ;
  assign w15079 = ( w4141 & ~w15077 ) | ( w4141 & w15078 ) | ( ~w15077 & w15078 ) ;
  assign w15080 = ~\pi122 & w4143 ;
  assign w15081 = w7069 | w15079 ;
  assign w15082 = ( w4144 & w15079 ) | ( w4144 & w15081 ) | ( w15079 & w15081 ) ;
  assign w15083 = ( w4143 & ~w15080 ) | ( w4143 & w15082 ) | ( ~w15080 & w15082 ) ;
  assign w15084 = \pi044 ^ w15083 ;
  assign w15085 = w15075 ^ w15076 ;
  assign w15086 = w15084 ^ w15085 ;
  assign w15087 = ( ~w14959 & w14967 ) | ( ~w14959 & w14968 ) | ( w14967 & w14968 ) ;
  assign w15088 = w15086 ^ w15087 ;
  assign w15089 = ~\pi124 & w3635 ;
  assign w15090 = \pi123 & w3817 ;
  assign w15091 = ( w3635 & ~w15089 ) | ( w3635 & w15090 ) | ( ~w15089 & w15090 ) ;
  assign w15092 = ~\pi125 & w3637 ;
  assign w15093 = w7988 | w15091 ;
  assign w15094 = ( w3638 & w15091 ) | ( w3638 & w15093 ) | ( w15091 & w15093 ) ;
  assign w15095 = ( w3637 & ~w15092 ) | ( w3637 & w15094 ) | ( ~w15092 & w15094 ) ;
  assign w15096 = \pi041 ^ w15095 ;
  assign w15097 = w14996 ^ w15096 ;
  assign w15098 = w15001 ^ w15088 ;
  assign w15099 = \pi038 ^ w15098 ;
  assign w15100 = w15097 ^ w15099 ;
  assign w15101 = ( ~w14981 & w14989 ) | ( ~w14981 & w14990 ) | ( w14989 & w14990 ) ;
  assign w15102 = ( w14887 & w14992 ) | ( w14887 & ~w14993 ) | ( w14992 & ~w14993 ) ;
  assign w15103 = w15101 ^ w15102 ;
  assign w15104 = w15100 ^ w15103 ;
  assign w15105 = ( w15100 & ~w15101 ) | ( w15100 & w15102 ) | ( ~w15101 & w15102 ) ;
  assign w15106 = \pi038 ^ w15001 ;
  assign w15107 = w15088 ^ w15096 ;
  assign w15108 = ( w14996 & w15106 ) | ( w14996 & ~w15107 ) | ( w15106 & ~w15107 ) ;
  assign w15109 = ( ~w15086 & w15087 ) | ( ~w15086 & w15096 ) | ( w15087 & w15096 ) ;
  assign w15110 = w3181 & w8481 ;
  assign w15111 = w3340 | w15110 ;
  assign w15112 = ( \pi127 & w15110 ) | ( \pi127 & w15111 ) | ( w15110 & w15111 ) ;
  assign w15113 = \pi038 ^ w15112 ;
  assign w15114 = ( ~w15064 & w15065 ) | ( ~w15064 & w15073 ) | ( w15065 & w15073 ) ;
  assign w15115 = ~\pi119 & w4654 ;
  assign w15116 = \pi118 & w4876 ;
  assign w15117 = ( w4654 & ~w15115 ) | ( w4654 & w15116 ) | ( ~w15115 & w15116 ) ;
  assign w15118 = ~\pi120 & w4656 ;
  assign w15119 = w6634 | w15117 ;
  assign w15120 = ( w4657 & w15117 ) | ( w4657 & w15119 ) | ( w15117 & w15119 ) ;
  assign w15121 = ( w4656 & ~w15118 ) | ( w4656 & w15120 ) | ( ~w15118 & w15120 ) ;
  assign w15122 = \pi047 ^ w15121 ;
  assign w15123 = ( ~w15053 & w15054 ) | ( ~w15053 & w15062 ) | ( w15054 & w15062 ) ;
  assign w15124 = ~\pi116 & w5209 ;
  assign w15125 = \pi115 & w5433 ;
  assign w15126 = ( w5209 & ~w15124 ) | ( w5209 & w15125 ) | ( ~w15124 & w15125 ) ;
  assign w15127 = ~\pi117 & w5211 ;
  assign w15128 = w6185 | w15126 ;
  assign w15129 = ( w5212 & w15126 ) | ( w5212 & w15128 ) | ( w15126 & w15128 ) ;
  assign w15130 = ( w5211 & ~w15127 ) | ( w5211 & w15129 ) | ( ~w15127 & w15129 ) ;
  assign w15131 = \pi050 ^ w15130 ;
  assign w15132 = ( ~w15042 & w15043 ) | ( ~w15042 & w15051 ) | ( w15043 & w15051 ) ;
  assign w15133 = ( w15009 & ~w15013 ) | ( w15009 & w15018 ) | ( ~w15013 & w15018 ) ;
  assign w15134 = \pi100 ^ \pi102 ;
  assign w15135 = ( \pi062 & \pi063 ) | ( \pi062 & ~w15134 ) | ( \pi063 & ~w15134 ) ;
  assign w15136 = \pi062 & ~w3263 ;
  assign w15137 = ( \pi063 & ~w3263 ) | ( \pi063 & w15136 ) | ( ~w3263 & w15136 ) ;
  assign w15138 = w15133 ^ w15137 ;
  assign w15139 = w15135 ^ w15138 ;
  assign w15140 = ~\pi104 & w7811 ;
  assign w15141 = \pi103 & w8046 ;
  assign w15142 = ( w7811 & ~w15140 ) | ( w7811 & w15141 ) | ( ~w15140 & w15141 ) ;
  assign w15143 = ~\pi105 & w7813 ;
  assign w15144 = w3905 | w15142 ;
  assign w15145 = ( w7814 & w15142 ) | ( w7814 & w15144 ) | ( w15142 & w15144 ) ;
  assign w15146 = ( w7813 & ~w15143 ) | ( w7813 & w15145 ) | ( ~w15143 & w15145 ) ;
  assign w15147 = \pi062 ^ w15146 ;
  assign w15148 = ~\pi107 & w7135 ;
  assign w15149 = \pi106 & w7359 ;
  assign w15150 = ( w7135 & ~w15148 ) | ( w7135 & w15149 ) | ( ~w15148 & w15149 ) ;
  assign w15151 = ~\pi108 & w7137 ;
  assign w15152 = w4425 | w15150 ;
  assign w15153 = ( w7138 & w15150 ) | ( w7138 & w15152 ) | ( w15150 & w15152 ) ;
  assign w15154 = ( w7137 & ~w15151 ) | ( w7137 & w15153 ) | ( ~w15151 & w15153 ) ;
  assign w15155 = \pi059 ^ w15154 ;
  assign w15156 = w15139 ^ w15155 ;
  assign w15157 = w15147 ^ w15156 ;
  assign w15158 = ( ~w15020 & w15021 ) | ( ~w15020 & w15029 ) | ( w15021 & w15029 ) ;
  assign w15159 = ~\pi110 & w6466 ;
  assign w15160 = \pi109 & w6702 ;
  assign w15161 = ( w6466 & ~w15159 ) | ( w6466 & w15160 ) | ( ~w15159 & w15160 ) ;
  assign w15162 = ~\pi111 & w6468 ;
  assign w15163 = w4811 | w15161 ;
  assign w15164 = ( w6469 & w15161 ) | ( w6469 & w15163 ) | ( w15161 & w15163 ) ;
  assign w15165 = ( w6468 & ~w15162 ) | ( w6468 & w15164 ) | ( ~w15162 & w15164 ) ;
  assign w15166 = \pi056 ^ w15165 ;
  assign w15167 = w15157 ^ w15158 ;
  assign w15168 = w15166 ^ w15167 ;
  assign w15169 = ( ~w15031 & w15032 ) | ( ~w15031 & w15040 ) | ( w15032 & w15040 ) ;
  assign w15170 = ~\pi113 & w5802 ;
  assign w15171 = \pi112 & w6052 ;
  assign w15172 = ( w5802 & ~w15170 ) | ( w5802 & w15171 ) | ( ~w15170 & w15171 ) ;
  assign w15173 = ~\pi114 & w5804 ;
  assign w15174 = w5565 | w15172 ;
  assign w15175 = ( w5805 & w15172 ) | ( w5805 & w15174 ) | ( w15172 & w15174 ) ;
  assign w15176 = ( w5804 & ~w15173 ) | ( w5804 & w15175 ) | ( ~w15173 & w15175 ) ;
  assign w15177 = \pi053 ^ w15176 ;
  assign w15178 = w15168 ^ w15169 ;
  assign w15179 = w15177 ^ w15178 ;
  assign w15180 = w15132 ^ w15179 ;
  assign w15181 = w15131 ^ w15180 ;
  assign w15182 = w15123 ^ w15181 ;
  assign w15183 = w15122 ^ w15182 ;
  assign w15184 = ~\pi122 & w4141 ;
  assign w15185 = \pi121 & w4334 ;
  assign w15186 = ( w4141 & ~w15184 ) | ( w4141 & w15185 ) | ( ~w15184 & w15185 ) ;
  assign w15187 = ~\pi123 & w4143 ;
  assign w15188 = w7516 | w15186 ;
  assign w15189 = ( w4144 & w15186 ) | ( w4144 & w15188 ) | ( w15186 & w15188 ) ;
  assign w15190 = ( w4143 & ~w15187 ) | ( w4143 & w15189 ) | ( ~w15187 & w15189 ) ;
  assign w15191 = \pi044 ^ w15190 ;
  assign w15192 = w15114 ^ w15191 ;
  assign w15193 = w15183 ^ w15192 ;
  assign w15194 = ( ~w15075 & w15076 ) | ( ~w15075 & w15084 ) | ( w15076 & w15084 ) ;
  assign w15195 = ~\pi125 & w3635 ;
  assign w15196 = \pi124 & w3817 ;
  assign w15197 = ( w3635 & ~w15195 ) | ( w3635 & w15196 ) | ( ~w15195 & w15196 ) ;
  assign w15198 = ~\pi126 & w3637 ;
  assign w15199 = w8231 | w15197 ;
  assign w15200 = ( w3638 & w15197 ) | ( w3638 & w15199 ) | ( w15197 & w15199 ) ;
  assign w15201 = ( w3637 & ~w15198 ) | ( w3637 & w15200 ) | ( ~w15198 & w15200 ) ;
  assign w15202 = \pi041 ^ w15201 ;
  assign w15203 = w15193 ^ w15202 ;
  assign w15204 = w15194 ^ w15203 ;
  assign w15205 = w15113 ^ w15204 ;
  assign w15206 = w15109 ^ w15205 ;
  assign w15207 = w15105 ^ w15206 ;
  assign w15208 = w15108 ^ w15207 ;
  assign w15209 = ( w15105 & ~w15108 ) | ( w15105 & w15206 ) | ( ~w15108 & w15206 ) ;
  assign w15210 = ( w15131 & w15132 ) | ( w15131 & ~w15179 ) | ( w15132 & ~w15179 ) ;
  assign w15211 = ~\pi117 & w5209 ;
  assign w15212 = \pi116 & w5433 ;
  assign w15213 = ( w5209 & ~w15211 ) | ( w5209 & w15212 ) | ( ~w15211 & w15212 ) ;
  assign w15214 = ~\pi118 & w5211 ;
  assign w15215 = w6206 | w15213 ;
  assign w15216 = ( w5212 & w15213 ) | ( w5212 & w15215 ) | ( w15213 & w15215 ) ;
  assign w15217 = ( w5211 & ~w15214 ) | ( w5211 & w15216 ) | ( ~w15214 & w15216 ) ;
  assign w15218 = \pi050 ^ w15217 ;
  assign w15219 = ( ~w15168 & w15169 ) | ( ~w15168 & w15177 ) | ( w15169 & w15177 ) ;
  assign w15220 = \pi101 | w15133 ;
  assign w15221 = ( \pi063 & \pi100 ) | ( \pi063 & ~w15220 ) | ( \pi100 & ~w15220 ) ;
  assign w15222 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15221 ) | ( ~\pi063 & w15221 ) ;
  assign w15223 = ( \pi062 & \pi063 ) | ( \pi062 & \pi102 ) | ( \pi063 & \pi102 ) ;
  assign w15224 = ( ~\pi101 & w15133 ) | ( ~\pi101 & w15223 ) | ( w15133 & w15223 ) ;
  assign w15225 = ( \pi063 & ~w15133 ) | ( \pi063 & w15220 ) | ( ~w15133 & w15220 ) ;
  assign w15226 = ( \pi062 & \pi101 ) | ( \pi062 & ~w15225 ) | ( \pi101 & ~w15225 ) ;
  assign w15227 = ( ~w15222 & w15224 ) | ( ~w15222 & w15226 ) | ( w15224 & w15226 ) ;
  assign w15228 = \pi038 ^ w15013 ;
  assign w15229 = ( \pi062 & \pi063 ) | ( \pi062 & \pi103 ) | ( \pi063 & \pi103 ) ;
  assign w15230 = \pi063 & ~\pi102 ;
  assign w15231 = \pi062 & w15230 ;
  assign w15232 = w15229 ^ w15231 ;
  assign w15233 = w15228 ^ w15232 ;
  assign w15234 = ~\pi105 & w7811 ;
  assign w15235 = \pi104 & w8046 ;
  assign w15236 = ( w7811 & ~w15234 ) | ( w7811 & w15235 ) | ( ~w15234 & w15235 ) ;
  assign w15237 = ~\pi106 & w7813 ;
  assign w15238 = w4068 | w15236 ;
  assign w15239 = ( w7814 & w15236 ) | ( w7814 & w15238 ) | ( w15236 & w15238 ) ;
  assign w15240 = ( w7813 & ~w15237 ) | ( w7813 & w15239 ) | ( ~w15237 & w15239 ) ;
  assign w15241 = \pi062 ^ w15240 ;
  assign w15242 = w15227 ^ w15241 ;
  assign w15243 = w15233 ^ w15242 ;
  assign w15244 = ~\pi108 & w7135 ;
  assign w15245 = \pi107 & w7359 ;
  assign w15246 = ( w7135 & ~w15244 ) | ( w7135 & w15245 ) | ( ~w15244 & w15245 ) ;
  assign w15247 = ~\pi109 & w7137 ;
  assign w15248 = w4599 | w15246 ;
  assign w15249 = ( w7138 & w15246 ) | ( w7138 & w15248 ) | ( w15246 & w15248 ) ;
  assign w15250 = ( w7137 & ~w15247 ) | ( w7137 & w15249 ) | ( ~w15247 & w15249 ) ;
  assign w15251 = \pi059 ^ w15250 ;
  assign w15252 = ( ~w15139 & w15147 ) | ( ~w15139 & w15155 ) | ( w15147 & w15155 ) ;
  assign w15253 = w15243 ^ w15252 ;
  assign w15254 = w15251 ^ w15253 ;
  assign w15255 = ~\pi111 & w6466 ;
  assign w15256 = \pi110 & w6702 ;
  assign w15257 = ( w6466 & ~w15255 ) | ( w6466 & w15256 ) | ( ~w15255 & w15256 ) ;
  assign w15258 = ~\pi112 & w6468 ;
  assign w15259 = w4999 | w15257 ;
  assign w15260 = ( w6469 & w15257 ) | ( w6469 & w15259 ) | ( w15257 & w15259 ) ;
  assign w15261 = ( w6468 & ~w15258 ) | ( w6468 & w15260 ) | ( ~w15258 & w15260 ) ;
  assign w15262 = \pi056 ^ w15261 ;
  assign w15263 = ( ~w15157 & w15158 ) | ( ~w15157 & w15166 ) | ( w15158 & w15166 ) ;
  assign w15264 = w15254 ^ w15263 ;
  assign w15265 = w15262 ^ w15264 ;
  assign w15266 = ~\pi114 & w5802 ;
  assign w15267 = \pi113 & w6052 ;
  assign w15268 = ( w5802 & ~w15266 ) | ( w5802 & w15267 ) | ( ~w15266 & w15267 ) ;
  assign w15269 = ~\pi115 & w5804 ;
  assign w15270 = w5585 | w15268 ;
  assign w15271 = ( w5805 & w15268 ) | ( w5805 & w15270 ) | ( w15268 & w15270 ) ;
  assign w15272 = ( w5804 & ~w15269 ) | ( w5804 & w15271 ) | ( ~w15269 & w15271 ) ;
  assign w15273 = \pi053 ^ w15272 ;
  assign w15274 = w15219 ^ w15265 ;
  assign w15275 = w15273 ^ w15274 ;
  assign w15276 = w15210 ^ w15275 ;
  assign w15277 = w15218 ^ w15276 ;
  assign w15278 = ~\pi120 & w4654 ;
  assign w15279 = \pi119 & w4876 ;
  assign w15280 = ( w4654 & ~w15278 ) | ( w4654 & w15279 ) | ( ~w15278 & w15279 ) ;
  assign w15281 = ~\pi121 & w4656 ;
  assign w15282 = w7050 | w15280 ;
  assign w15283 = ( w4657 & w15280 ) | ( w4657 & w15282 ) | ( w15280 & w15282 ) ;
  assign w15284 = ( w4656 & ~w15281 ) | ( w4656 & w15283 ) | ( ~w15281 & w15283 ) ;
  assign w15285 = \pi047 ^ w15284 ;
  assign w15286 = ( w15122 & w15123 ) | ( w15122 & ~w15181 ) | ( w15123 & ~w15181 ) ;
  assign w15287 = w15277 ^ w15286 ;
  assign w15288 = w15285 ^ w15287 ;
  assign w15289 = ~\pi123 & w4141 ;
  assign w15290 = \pi122 & w4334 ;
  assign w15291 = ( w4141 & ~w15289 ) | ( w4141 & w15290 ) | ( ~w15289 & w15290 ) ;
  assign w15292 = ~\pi124 & w4143 ;
  assign w15293 = w7538 | w15291 ;
  assign w15294 = ( w4144 & w15291 ) | ( w4144 & w15293 ) | ( w15291 & w15293 ) ;
  assign w15295 = ( w4143 & ~w15292 ) | ( w4143 & w15294 ) | ( ~w15292 & w15294 ) ;
  assign w15296 = \pi044 ^ w15295 ;
  assign w15297 = ( w15114 & ~w15183 ) | ( w15114 & w15191 ) | ( ~w15183 & w15191 ) ;
  assign w15298 = w15296 ^ w15297 ;
  assign w15299 = w15288 ^ w15298 ;
  assign w15300 = ~\pi126 & w3635 ;
  assign w15301 = \pi125 & w3817 ;
  assign w15302 = ( w3635 & ~w15300 ) | ( w3635 & w15301 ) | ( ~w15300 & w15301 ) ;
  assign w15303 = ~\pi127 & w3637 ;
  assign w15304 = w8466 | w15302 ;
  assign w15305 = ( w3638 & w15302 ) | ( w3638 & w15304 ) | ( w15302 & w15304 ) ;
  assign w15306 = ( w3637 & ~w15303 ) | ( w3637 & w15305 ) | ( ~w15303 & w15305 ) ;
  assign w15307 = \pi041 ^ w15306 ;
  assign w15308 = ( ~w15193 & w15194 ) | ( ~w15193 & w15202 ) | ( w15194 & w15202 ) ;
  assign w15309 = w15307 ^ w15308 ;
  assign w15310 = w15299 ^ w15309 ;
  assign w15311 = ( w15109 & w15113 ) | ( w15109 & ~w15204 ) | ( w15113 & ~w15204 ) ;
  assign w15312 = w15209 ^ w15310 ;
  assign w15313 = w15311 ^ w15312 ;
  assign w15314 = ( ~w15288 & w15296 ) | ( ~w15288 & w15297 ) | ( w15296 & w15297 ) ;
  assign w15315 = \pi127 & w3635 ;
  assign w15316 = ( \pi126 & ~w3638 ) | ( \pi126 & w8490 ) | ( ~w3638 & w8490 ) ;
  assign w15317 = \pi126 & ~w3817 ;
  assign w15318 = ( ~\pi126 & w15316 ) | ( ~\pi126 & w15317 ) | ( w15316 & w15317 ) ;
  assign w15319 = ( w9420 & w15315 ) | ( w9420 & ~w15318 ) | ( w15315 & ~w15318 ) ;
  assign w15320 = ( w15227 & ~w15233 ) | ( w15227 & w15241 ) | ( ~w15233 & w15241 ) ;
  assign w15321 = ( \pi062 & \pi063 ) | ( \pi062 & \pi104 ) | ( \pi063 & \pi104 ) ;
  assign w15322 = \pi063 & ~\pi103 ;
  assign w15323 = w15321 & ~w15322 ;
  assign w15324 = ( ~\pi062 & w15321 ) | ( ~\pi062 & w15323 ) | ( w15321 & w15323 ) ;
  assign w15325 = \pi063 & \pi102 ;
  assign w15326 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w15325 ) | ( \pi063 & w15325 ) ;
  assign w15327 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15325 ) | ( ~\pi063 & w15325 ) ;
  assign w15328 = ( \pi103 & w15326 ) | ( \pi103 & w15327 ) | ( w15326 & w15327 ) ;
  assign w15329 = ( ~\pi038 & w15013 ) | ( ~\pi038 & w15328 ) | ( w15013 & w15328 ) ;
  assign w15330 = \pi105 & w8046 ;
  assign w15331 = ( \pi107 & w7813 ) | ( \pi107 & w15330 ) | ( w7813 & w15330 ) ;
  assign w15332 = \pi106 | w15331 ;
  assign w15333 = ( w7811 & w15331 ) | ( w7811 & w15332 ) | ( w15331 & w15332 ) ;
  assign w15334 = w15330 | w15333 ;
  assign w15335 = ~w4087 & w7814 ;
  assign w15336 = ( w7814 & w15334 ) | ( w7814 & ~w15335 ) | ( w15334 & ~w15335 ) ;
  assign w15337 = w15329 ^ w15336 ;
  assign w15338 = \pi062 ^ w15324 ;
  assign w15339 = w15337 ^ w15338 ;
  assign w15340 = ~\pi109 & w7135 ;
  assign w15341 = \pi108 & w7359 ;
  assign w15342 = ( w7135 & ~w15340 ) | ( w7135 & w15341 ) | ( ~w15340 & w15341 ) ;
  assign w15343 = ~\pi110 & w7137 ;
  assign w15344 = w4792 | w15342 ;
  assign w15345 = ( w7138 & w15342 ) | ( w7138 & w15344 ) | ( w15342 & w15344 ) ;
  assign w15346 = ( w7137 & ~w15343 ) | ( w7137 & w15345 ) | ( ~w15343 & w15345 ) ;
  assign w15347 = \pi059 ^ w15346 ;
  assign w15348 = w15320 ^ w15347 ;
  assign w15349 = w15339 ^ w15348 ;
  assign w15350 = ( ~w15243 & w15251 ) | ( ~w15243 & w15252 ) | ( w15251 & w15252 ) ;
  assign w15351 = ~\pi112 & w6466 ;
  assign w15352 = \pi111 & w6702 ;
  assign w15353 = ( w6466 & ~w15351 ) | ( w6466 & w15352 ) | ( ~w15351 & w15352 ) ;
  assign w15354 = ~\pi113 & w6468 ;
  assign w15355 = w5366 | w15353 ;
  assign w15356 = ( w6469 & w15353 ) | ( w6469 & w15355 ) | ( w15353 & w15355 ) ;
  assign w15357 = ( w6468 & ~w15354 ) | ( w6468 & w15356 ) | ( ~w15354 & w15356 ) ;
  assign w15358 = \pi056 ^ w15357 ;
  assign w15359 = w15349 ^ w15350 ;
  assign w15360 = w15358 ^ w15359 ;
  assign w15361 = ( ~w15254 & w15262 ) | ( ~w15254 & w15263 ) | ( w15262 & w15263 ) ;
  assign w15362 = ~\pi115 & w5802 ;
  assign w15363 = \pi114 & w6052 ;
  assign w15364 = ( w5802 & ~w15362 ) | ( w5802 & w15363 ) | ( ~w15362 & w15363 ) ;
  assign w15365 = ~\pi116 & w5804 ;
  assign w15366 = w5976 | w15364 ;
  assign w15367 = ( w5805 & w15364 ) | ( w5805 & w15366 ) | ( w15364 & w15366 ) ;
  assign w15368 = ( w5804 & ~w15365 ) | ( w5804 & w15367 ) | ( ~w15365 & w15367 ) ;
  assign w15369 = \pi053 ^ w15368 ;
  assign w15370 = w15360 ^ w15361 ;
  assign w15371 = w15369 ^ w15370 ;
  assign w15372 = ( w15219 & ~w15265 ) | ( w15219 & w15273 ) | ( ~w15265 & w15273 ) ;
  assign w15373 = ~\pi118 & w5209 ;
  assign w15374 = \pi117 & w5433 ;
  assign w15375 = ( w5209 & ~w15373 ) | ( w5209 & w15374 ) | ( ~w15373 & w15374 ) ;
  assign w15376 = ~\pi119 & w5211 ;
  assign w15377 = w6616 | w15375 ;
  assign w15378 = ( w5212 & w15375 ) | ( w5212 & w15377 ) | ( w15375 & w15377 ) ;
  assign w15379 = ( w5211 & ~w15376 ) | ( w5211 & w15378 ) | ( ~w15376 & w15378 ) ;
  assign w15380 = \pi050 ^ w15379 ;
  assign w15381 = w15371 ^ w15372 ;
  assign w15382 = w15380 ^ w15381 ;
  assign w15383 = ( w15210 & w15218 ) | ( w15210 & ~w15275 ) | ( w15218 & ~w15275 ) ;
  assign w15384 = ~\pi121 & w4654 ;
  assign w15385 = \pi120 & w4876 ;
  assign w15386 = ( w4654 & ~w15384 ) | ( w4654 & w15385 ) | ( ~w15384 & w15385 ) ;
  assign w15387 = ~\pi122 & w4656 ;
  assign w15388 = w7069 | w15386 ;
  assign w15389 = ( w4657 & w15386 ) | ( w4657 & w15388 ) | ( w15386 & w15388 ) ;
  assign w15390 = ( w4656 & ~w15387 ) | ( w4656 & w15389 ) | ( ~w15387 & w15389 ) ;
  assign w15391 = \pi047 ^ w15390 ;
  assign w15392 = w15383 ^ w15391 ;
  assign w15393 = w15382 ^ w15392 ;
  assign w15394 = ( ~w15277 & w15285 ) | ( ~w15277 & w15286 ) | ( w15285 & w15286 ) ;
  assign w15395 = w15393 ^ w15394 ;
  assign w15396 = ~\pi124 & w4141 ;
  assign w15397 = \pi123 & w4334 ;
  assign w15398 = ( w4141 & ~w15396 ) | ( w4141 & w15397 ) | ( ~w15396 & w15397 ) ;
  assign w15399 = ~\pi125 & w4143 ;
  assign w15400 = w7988 | w15398 ;
  assign w15401 = ( w4144 & w15398 ) | ( w4144 & w15400 ) | ( w15398 & w15400 ) ;
  assign w15402 = ( w4143 & ~w15399 ) | ( w4143 & w15401 ) | ( ~w15399 & w15401 ) ;
  assign w15403 = \pi044 ^ w15402 ;
  assign w15404 = w15314 ^ w15403 ;
  assign w15405 = w15319 ^ w15395 ;
  assign w15406 = \pi041 ^ w15405 ;
  assign w15407 = w15404 ^ w15406 ;
  assign w15408 = ( ~w15299 & w15307 ) | ( ~w15299 & w15308 ) | ( w15307 & w15308 ) ;
  assign w15409 = ( w15209 & w15310 ) | ( w15209 & ~w15311 ) | ( w15310 & ~w15311 ) ;
  assign w15410 = w15408 ^ w15409 ;
  assign w15411 = w15407 ^ w15410 ;
  assign w15412 = ( w15407 & ~w15408 ) | ( w15407 & w15409 ) | ( ~w15408 & w15409 ) ;
  assign w15413 = \pi041 ^ w15319 ;
  assign w15414 = w15395 ^ w15403 ;
  assign w15415 = ( w15314 & w15413 ) | ( w15314 & ~w15414 ) | ( w15413 & ~w15414 ) ;
  assign w15416 = ( ~w15393 & w15394 ) | ( ~w15393 & w15403 ) | ( w15394 & w15403 ) ;
  assign w15417 = w3638 & w8481 ;
  assign w15418 = w3817 | w15417 ;
  assign w15419 = ( \pi127 & w15417 ) | ( \pi127 & w15418 ) | ( w15417 & w15418 ) ;
  assign w15420 = \pi041 ^ w15419 ;
  assign w15421 = ~\pi122 & w4654 ;
  assign w15422 = \pi121 & w4876 ;
  assign w15423 = ( w4654 & ~w15421 ) | ( w4654 & w15422 ) | ( ~w15421 & w15422 ) ;
  assign w15424 = ~\pi123 & w4656 ;
  assign w15425 = w7516 | w15423 ;
  assign w15426 = ( w4657 & w15423 ) | ( w4657 & w15425 ) | ( w15423 & w15425 ) ;
  assign w15427 = ( w4656 & ~w15424 ) | ( w4656 & w15426 ) | ( ~w15424 & w15426 ) ;
  assign w15428 = \pi047 ^ w15427 ;
  assign w15429 = ( ~w15371 & w15372 ) | ( ~w15371 & w15380 ) | ( w15372 & w15380 ) ;
  assign w15430 = ~\pi119 & w5209 ;
  assign w15431 = \pi118 & w5433 ;
  assign w15432 = ( w5209 & ~w15430 ) | ( w5209 & w15431 ) | ( ~w15430 & w15431 ) ;
  assign w15433 = ~\pi120 & w5211 ;
  assign w15434 = w6634 | w15432 ;
  assign w15435 = ( w5212 & w15432 ) | ( w5212 & w15434 ) | ( w15432 & w15434 ) ;
  assign w15436 = ( w5211 & ~w15433 ) | ( w5211 & w15435 ) | ( ~w15433 & w15435 ) ;
  assign w15437 = \pi050 ^ w15436 ;
  assign w15438 = ( ~w15360 & w15361 ) | ( ~w15360 & w15369 ) | ( w15361 & w15369 ) ;
  assign w15439 = ~\pi116 & w5802 ;
  assign w15440 = \pi115 & w6052 ;
  assign w15441 = ( w5802 & ~w15439 ) | ( w5802 & w15440 ) | ( ~w15439 & w15440 ) ;
  assign w15442 = ~\pi117 & w5804 ;
  assign w15443 = w6185 | w15441 ;
  assign w15444 = ( w5805 & w15441 ) | ( w5805 & w15443 ) | ( w15441 & w15443 ) ;
  assign w15445 = ( w5804 & ~w15442 ) | ( w5804 & w15444 ) | ( ~w15442 & w15444 ) ;
  assign w15446 = \pi053 ^ w15445 ;
  assign w15447 = ( ~w15349 & w15350 ) | ( ~w15349 & w15358 ) | ( w15350 & w15358 ) ;
  assign w15448 = ( w15320 & ~w15339 ) | ( w15320 & w15347 ) | ( ~w15339 & w15347 ) ;
  assign w15449 = w4087 | w15334 ;
  assign w15450 = ( w7814 & w15334 ) | ( w7814 & w15449 ) | ( w15334 & w15449 ) ;
  assign w15451 = \pi062 ^ w15450 ;
  assign w15452 = ( ~w15324 & w15329 ) | ( ~w15324 & w15451 ) | ( w15329 & w15451 ) ;
  assign w15453 = \pi103 ^ \pi105 ;
  assign w15454 = ( \pi062 & \pi063 ) | ( \pi062 & ~w15453 ) | ( \pi063 & ~w15453 ) ;
  assign w15455 = \pi103 ^ \pi104 ;
  assign w15456 = \pi062 & ~w15455 ;
  assign w15457 = ( \pi063 & ~w15455 ) | ( \pi063 & w15456 ) | ( ~w15455 & w15456 ) ;
  assign w15458 = w15452 ^ w15457 ;
  assign w15459 = w15454 ^ w15458 ;
  assign w15460 = ~\pi107 & w7811 ;
  assign w15461 = \pi106 & w8046 ;
  assign w15462 = ( w7811 & ~w15460 ) | ( w7811 & w15461 ) | ( ~w15460 & w15461 ) ;
  assign w15463 = ~\pi108 & w7813 ;
  assign w15464 = w4425 | w15462 ;
  assign w15465 = ( w7814 & w15462 ) | ( w7814 & w15464 ) | ( w15462 & w15464 ) ;
  assign w15466 = ( w7813 & ~w15463 ) | ( w7813 & w15465 ) | ( ~w15463 & w15465 ) ;
  assign w15467 = \pi062 ^ w15466 ;
  assign w15468 = ~\pi110 & w7135 ;
  assign w15469 = \pi109 & w7359 ;
  assign w15470 = ( w7135 & ~w15468 ) | ( w7135 & w15469 ) | ( ~w15468 & w15469 ) ;
  assign w15471 = ~\pi111 & w7137 ;
  assign w15472 = w4811 | w15470 ;
  assign w15473 = ( w7138 & w15470 ) | ( w7138 & w15472 ) | ( w15470 & w15472 ) ;
  assign w15474 = ( w7137 & ~w15471 ) | ( w7137 & w15473 ) | ( ~w15471 & w15473 ) ;
  assign w15475 = \pi059 ^ w15474 ;
  assign w15476 = w15459 ^ w15475 ;
  assign w15477 = w15467 ^ w15476 ;
  assign w15478 = ~\pi113 & w6466 ;
  assign w15479 = \pi112 & w6702 ;
  assign w15480 = ( w6466 & ~w15478 ) | ( w6466 & w15479 ) | ( ~w15478 & w15479 ) ;
  assign w15481 = ~\pi114 & w6468 ;
  assign w15482 = w5565 | w15480 ;
  assign w15483 = ( w6469 & w15480 ) | ( w6469 & w15482 ) | ( w15480 & w15482 ) ;
  assign w15484 = ( w6468 & ~w15481 ) | ( w6468 & w15483 ) | ( ~w15481 & w15483 ) ;
  assign w15485 = \pi056 ^ w15484 ;
  assign w15486 = w15448 ^ w15477 ;
  assign w15487 = w15485 ^ w15486 ;
  assign w15488 = w15447 ^ w15487 ;
  assign w15489 = w15446 ^ w15488 ;
  assign w15490 = w15437 ^ w15438 ;
  assign w15491 = w15489 ^ w15490 ;
  assign w15492 = w15428 ^ w15429 ;
  assign w15493 = w15491 ^ w15492 ;
  assign w15494 = ( ~w15382 & w15383 ) | ( ~w15382 & w15391 ) | ( w15383 & w15391 ) ;
  assign w15495 = ~\pi125 & w4141 ;
  assign w15496 = \pi124 & w4334 ;
  assign w15497 = ( w4141 & ~w15495 ) | ( w4141 & w15496 ) | ( ~w15495 & w15496 ) ;
  assign w15498 = ~\pi126 & w4143 ;
  assign w15499 = w8231 | w15497 ;
  assign w15500 = ( w4144 & w15497 ) | ( w4144 & w15499 ) | ( w15497 & w15499 ) ;
  assign w15501 = ( w4143 & ~w15498 ) | ( w4143 & w15500 ) | ( ~w15498 & w15500 ) ;
  assign w15502 = \pi044 ^ w15501 ;
  assign w15503 = w15493 ^ w15502 ;
  assign w15504 = w15494 ^ w15503 ;
  assign w15505 = w15420 ^ w15504 ;
  assign w15506 = w15416 ^ w15505 ;
  assign w15507 = w15412 ^ w15506 ;
  assign w15508 = w15415 ^ w15507 ;
  assign w15509 = ( w15412 & ~w15415 ) | ( w15412 & w15506 ) | ( ~w15415 & w15506 ) ;
  assign w15510 = ~\pi123 & w4654 ;
  assign w15511 = \pi122 & w4876 ;
  assign w15512 = ( w4654 & ~w15510 ) | ( w4654 & w15511 ) | ( ~w15510 & w15511 ) ;
  assign w15513 = ~\pi124 & w4656 ;
  assign w15514 = w7538 | w15512 ;
  assign w15515 = ( w4657 & w15512 ) | ( w4657 & w15514 ) | ( w15512 & w15514 ) ;
  assign w15516 = ( w4656 & ~w15513 ) | ( w4656 & w15515 ) | ( ~w15513 & w15515 ) ;
  assign w15517 = \pi047 ^ w15516 ;
  assign w15518 = ( w15437 & w15438 ) | ( w15437 & ~w15489 ) | ( w15438 & ~w15489 ) ;
  assign w15519 = ~\pi120 & w5209 ;
  assign w15520 = \pi119 & w5433 ;
  assign w15521 = ( w5209 & ~w15519 ) | ( w5209 & w15520 ) | ( ~w15519 & w15520 ) ;
  assign w15522 = ~\pi121 & w5211 ;
  assign w15523 = w7050 | w15521 ;
  assign w15524 = ( w5212 & w15521 ) | ( w5212 & w15523 ) | ( w15521 & w15523 ) ;
  assign w15525 = ( w5211 & ~w15522 ) | ( w5211 & w15524 ) | ( ~w15522 & w15524 ) ;
  assign w15526 = \pi050 ^ w15525 ;
  assign w15527 = ( w15446 & w15447 ) | ( w15446 & ~w15487 ) | ( w15447 & ~w15487 ) ;
  assign w15528 = ( w15448 & ~w15477 ) | ( w15448 & w15485 ) | ( ~w15477 & w15485 ) ;
  assign w15529 = ~\pi114 & w6466 ;
  assign w15530 = \pi113 & w6702 ;
  assign w15531 = ( w6466 & ~w15529 ) | ( w6466 & w15530 ) | ( ~w15529 & w15530 ) ;
  assign w15532 = ~\pi115 & w6468 ;
  assign w15533 = w5585 | w15531 ;
  assign w15534 = ( w6469 & w15531 ) | ( w6469 & w15533 ) | ( w15531 & w15533 ) ;
  assign w15535 = ( w6468 & ~w15532 ) | ( w6468 & w15534 ) | ( ~w15532 & w15534 ) ;
  assign w15536 = \pi056 ^ w15535 ;
  assign w15537 = \pi041 ^ w15324 ;
  assign w15538 = ( \pi062 & \pi063 ) | ( \pi062 & \pi106 ) | ( \pi063 & \pi106 ) ;
  assign w15539 = \pi063 & ~\pi105 ;
  assign w15540 = \pi062 & w15539 ;
  assign w15541 = w15538 ^ w15540 ;
  assign w15542 = w15537 ^ w15541 ;
  assign w15543 = ~\pi108 & w7811 ;
  assign w15544 = \pi107 & w8046 ;
  assign w15545 = ( w7811 & ~w15543 ) | ( w7811 & w15544 ) | ( ~w15543 & w15544 ) ;
  assign w15546 = ~\pi109 & w7813 ;
  assign w15547 = w4599 | w15545 ;
  assign w15548 = ( w7814 & w15545 ) | ( w7814 & w15547 ) | ( w15545 & w15547 ) ;
  assign w15549 = ( w7813 & ~w15546 ) | ( w7813 & w15548 ) | ( ~w15546 & w15548 ) ;
  assign w15550 = \pi062 ^ w15549 ;
  assign w15551 = \pi104 | w15452 ;
  assign w15552 = ( \pi063 & \pi103 ) | ( \pi063 & ~w15551 ) | ( \pi103 & ~w15551 ) ;
  assign w15553 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15552 ) | ( ~\pi063 & w15552 ) ;
  assign w15554 = ( \pi062 & \pi063 ) | ( \pi062 & \pi105 ) | ( \pi063 & \pi105 ) ;
  assign w15555 = ( ~\pi104 & w15452 ) | ( ~\pi104 & w15554 ) | ( w15452 & w15554 ) ;
  assign w15556 = ( \pi063 & ~w15452 ) | ( \pi063 & w15551 ) | ( ~w15452 & w15551 ) ;
  assign w15557 = ( \pi062 & \pi104 ) | ( \pi062 & ~w15556 ) | ( \pi104 & ~w15556 ) ;
  assign w15558 = ( ~w15553 & w15555 ) | ( ~w15553 & w15557 ) | ( w15555 & w15557 ) ;
  assign w15559 = w15550 ^ w15558 ;
  assign w15560 = w15542 ^ w15559 ;
  assign w15561 = ~\pi111 & w7135 ;
  assign w15562 = \pi110 & w7359 ;
  assign w15563 = ( w7135 & ~w15561 ) | ( w7135 & w15562 ) | ( ~w15561 & w15562 ) ;
  assign w15564 = ~\pi112 & w7137 ;
  assign w15565 = w4999 | w15563 ;
  assign w15566 = ( w7138 & w15563 ) | ( w7138 & w15565 ) | ( w15563 & w15565 ) ;
  assign w15567 = ( w7137 & ~w15564 ) | ( w7137 & w15566 ) | ( ~w15564 & w15566 ) ;
  assign w15568 = \pi059 ^ w15567 ;
  assign w15569 = ( ~w15459 & w15467 ) | ( ~w15459 & w15475 ) | ( w15467 & w15475 ) ;
  assign w15570 = w15560 ^ w15569 ;
  assign w15571 = w15568 ^ w15570 ;
  assign w15572 = w15528 ^ w15571 ;
  assign w15573 = w15536 ^ w15572 ;
  assign w15574 = ~\pi117 & w5802 ;
  assign w15575 = \pi116 & w6052 ;
  assign w15576 = ( w5802 & ~w15574 ) | ( w5802 & w15575 ) | ( ~w15574 & w15575 ) ;
  assign w15577 = ~\pi118 & w5804 ;
  assign w15578 = w6206 | w15576 ;
  assign w15579 = ( w5805 & w15576 ) | ( w5805 & w15578 ) | ( w15576 & w15578 ) ;
  assign w15580 = ( w5804 & ~w15577 ) | ( w5804 & w15579 ) | ( ~w15577 & w15579 ) ;
  assign w15581 = \pi053 ^ w15580 ;
  assign w15582 = w15527 ^ w15573 ;
  assign w15583 = w15581 ^ w15582 ;
  assign w15584 = w15518 ^ w15526 ;
  assign w15585 = w15583 ^ w15584 ;
  assign w15586 = ( w15428 & w15429 ) | ( w15428 & ~w15491 ) | ( w15429 & ~w15491 ) ;
  assign w15587 = w15517 ^ w15586 ;
  assign w15588 = w15585 ^ w15587 ;
  assign w15589 = ~\pi126 & w4141 ;
  assign w15590 = \pi125 & w4334 ;
  assign w15591 = ( w4141 & ~w15589 ) | ( w4141 & w15590 ) | ( ~w15589 & w15590 ) ;
  assign w15592 = ~\pi127 & w4143 ;
  assign w15593 = w8466 | w15591 ;
  assign w15594 = ( w4144 & w15591 ) | ( w4144 & w15593 ) | ( w15591 & w15593 ) ;
  assign w15595 = ( w4143 & ~w15592 ) | ( w4143 & w15594 ) | ( ~w15592 & w15594 ) ;
  assign w15596 = \pi044 ^ w15595 ;
  assign w15597 = ( ~w15493 & w15494 ) | ( ~w15493 & w15502 ) | ( w15494 & w15502 ) ;
  assign w15598 = w15596 ^ w15597 ;
  assign w15599 = w15588 ^ w15598 ;
  assign w15600 = ( w15416 & w15420 ) | ( w15416 & ~w15504 ) | ( w15420 & ~w15504 ) ;
  assign w15601 = w15509 ^ w15599 ;
  assign w15602 = w15600 ^ w15601 ;
  assign w15603 = ( w15517 & ~w15585 ) | ( w15517 & w15586 ) | ( ~w15585 & w15586 ) ;
  assign w15604 = \pi127 & w4141 ;
  assign w15605 = ( \pi126 & ~w4144 ) | ( \pi126 & w8490 ) | ( ~w4144 & w8490 ) ;
  assign w15606 = \pi126 & ~w4334 ;
  assign w15607 = ( ~\pi126 & w15605 ) | ( ~\pi126 & w15606 ) | ( w15605 & w15606 ) ;
  assign w15608 = ( w9420 & w15604 ) | ( w9420 & ~w15607 ) | ( w15604 & ~w15607 ) ;
  assign w15609 = ~\pi124 & w4654 ;
  assign w15610 = \pi123 & w4876 ;
  assign w15611 = ( w4654 & ~w15609 ) | ( w4654 & w15610 ) | ( ~w15609 & w15610 ) ;
  assign w15612 = ~\pi125 & w4656 ;
  assign w15613 = w7988 | w15611 ;
  assign w15614 = ( w4657 & w15611 ) | ( w4657 & w15613 ) | ( w15611 & w15613 ) ;
  assign w15615 = ( w4656 & ~w15612 ) | ( w4656 & w15614 ) | ( ~w15612 & w15614 ) ;
  assign w15616 = \pi047 ^ w15615 ;
  assign w15617 = ( w15518 & w15526 ) | ( w15518 & ~w15583 ) | ( w15526 & ~w15583 ) ;
  assign w15618 = ( w15527 & ~w15573 ) | ( w15527 & w15581 ) | ( ~w15573 & w15581 ) ;
  assign w15619 = ( ~w15542 & w15550 ) | ( ~w15542 & w15558 ) | ( w15550 & w15558 ) ;
  assign w15620 = ( \pi062 & \pi063 ) | ( \pi062 & \pi107 ) | ( \pi063 & \pi107 ) ;
  assign w15621 = \pi063 & ~\pi106 ;
  assign w15622 = w15620 & ~w15621 ;
  assign w15623 = ( ~\pi062 & w15620 ) | ( ~\pi062 & w15622 ) | ( w15620 & w15622 ) ;
  assign w15624 = \pi063 & \pi105 ;
  assign w15625 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w15624 ) | ( \pi063 & w15624 ) ;
  assign w15626 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15624 ) | ( ~\pi063 & w15624 ) ;
  assign w15627 = ( \pi106 & w15625 ) | ( \pi106 & w15626 ) | ( w15625 & w15626 ) ;
  assign w15628 = ( ~\pi041 & w15324 ) | ( ~\pi041 & w15627 ) | ( w15324 & w15627 ) ;
  assign w15629 = \pi108 & w8046 ;
  assign w15630 = ( \pi110 & w7813 ) | ( \pi110 & w15629 ) | ( w7813 & w15629 ) ;
  assign w15631 = \pi109 | w15630 ;
  assign w15632 = ( w7811 & w15630 ) | ( w7811 & w15631 ) | ( w15630 & w15631 ) ;
  assign w15633 = w15629 | w15632 ;
  assign w15634 = ~w4792 & w7814 ;
  assign w15635 = ( w7814 & w15633 ) | ( w7814 & ~w15634 ) | ( w15633 & ~w15634 ) ;
  assign w15636 = w15628 ^ w15635 ;
  assign w15637 = \pi062 ^ w15623 ;
  assign w15638 = w15636 ^ w15637 ;
  assign w15639 = ~\pi112 & w7135 ;
  assign w15640 = \pi111 & w7359 ;
  assign w15641 = ( w7135 & ~w15639 ) | ( w7135 & w15640 ) | ( ~w15639 & w15640 ) ;
  assign w15642 = ~\pi113 & w7137 ;
  assign w15643 = w5366 | w15641 ;
  assign w15644 = ( w7138 & w15641 ) | ( w7138 & w15643 ) | ( w15641 & w15643 ) ;
  assign w15645 = ( w7137 & ~w15642 ) | ( w7137 & w15644 ) | ( ~w15642 & w15644 ) ;
  assign w15646 = \pi059 ^ w15645 ;
  assign w15647 = w15619 ^ w15638 ;
  assign w15648 = w15646 ^ w15647 ;
  assign w15649 = ( ~w15560 & w15568 ) | ( ~w15560 & w15569 ) | ( w15568 & w15569 ) ;
  assign w15650 = ~\pi115 & w6466 ;
  assign w15651 = \pi114 & w6702 ;
  assign w15652 = ( w6466 & ~w15650 ) | ( w6466 & w15651 ) | ( ~w15650 & w15651 ) ;
  assign w15653 = ~\pi116 & w6468 ;
  assign w15654 = w5976 | w15652 ;
  assign w15655 = ( w6469 & w15652 ) | ( w6469 & w15654 ) | ( w15652 & w15654 ) ;
  assign w15656 = ( w6468 & ~w15653 ) | ( w6468 & w15655 ) | ( ~w15653 & w15655 ) ;
  assign w15657 = \pi056 ^ w15656 ;
  assign w15658 = w15648 ^ w15649 ;
  assign w15659 = w15657 ^ w15658 ;
  assign w15660 = ( w15528 & w15536 ) | ( w15528 & ~w15571 ) | ( w15536 & ~w15571 ) ;
  assign w15661 = ~\pi118 & w5802 ;
  assign w15662 = \pi117 & w6052 ;
  assign w15663 = ( w5802 & ~w15661 ) | ( w5802 & w15662 ) | ( ~w15661 & w15662 ) ;
  assign w15664 = ~\pi119 & w5804 ;
  assign w15665 = w6616 | w15663 ;
  assign w15666 = ( w5805 & w15663 ) | ( w5805 & w15665 ) | ( w15663 & w15665 ) ;
  assign w15667 = ( w5804 & ~w15664 ) | ( w5804 & w15666 ) | ( ~w15664 & w15666 ) ;
  assign w15668 = \pi053 ^ w15667 ;
  assign w15669 = w15659 ^ w15660 ;
  assign w15670 = w15668 ^ w15669 ;
  assign w15671 = ~\pi121 & w5209 ;
  assign w15672 = \pi120 & w5433 ;
  assign w15673 = ( w5209 & ~w15671 ) | ( w5209 & w15672 ) | ( ~w15671 & w15672 ) ;
  assign w15674 = ~\pi122 & w5211 ;
  assign w15675 = w7069 | w15673 ;
  assign w15676 = ( w5212 & w15673 ) | ( w5212 & w15675 ) | ( w15673 & w15675 ) ;
  assign w15677 = ( w5211 & ~w15674 ) | ( w5211 & w15676 ) | ( ~w15674 & w15676 ) ;
  assign w15678 = \pi050 ^ w15677 ;
  assign w15679 = w15618 ^ w15678 ;
  assign w15680 = w15670 ^ w15679 ;
  assign w15681 = w15616 ^ w15680 ;
  assign w15682 = w15617 ^ w15681 ;
  assign w15683 = \pi044 ^ w15603 ;
  assign w15684 = w15608 ^ w15683 ;
  assign w15685 = w15682 ^ w15684 ;
  assign w15686 = ( ~w15588 & w15596 ) | ( ~w15588 & w15597 ) | ( w15596 & w15597 ) ;
  assign w15687 = ( w15509 & w15599 ) | ( w15509 & ~w15600 ) | ( w15599 & ~w15600 ) ;
  assign w15688 = w15686 ^ w15687 ;
  assign w15689 = w15685 ^ w15688 ;
  assign w15690 = ( w15685 & ~w15686 ) | ( w15685 & w15687 ) | ( ~w15686 & w15687 ) ;
  assign w15691 = \pi044 ^ w15608 ;
  assign w15692 = ( w15603 & ~w15682 ) | ( w15603 & w15691 ) | ( ~w15682 & w15691 ) ;
  assign w15693 = ( w15616 & w15617 ) | ( w15616 & ~w15680 ) | ( w15617 & ~w15680 ) ;
  assign w15694 = w4144 & w8481 ;
  assign w15695 = w4334 | w15694 ;
  assign w15696 = ( \pi127 & w15694 ) | ( \pi127 & w15695 ) | ( w15694 & w15695 ) ;
  assign w15697 = \pi044 ^ w15696 ;
  assign w15698 = ~\pi122 & w5209 ;
  assign w15699 = \pi121 & w5433 ;
  assign w15700 = ( w5209 & ~w15698 ) | ( w5209 & w15699 ) | ( ~w15698 & w15699 ) ;
  assign w15701 = ~\pi123 & w5211 ;
  assign w15702 = w7516 | w15700 ;
  assign w15703 = ( w5212 & w15700 ) | ( w5212 & w15702 ) | ( w15700 & w15702 ) ;
  assign w15704 = ( w5211 & ~w15701 ) | ( w5211 & w15703 ) | ( ~w15701 & w15703 ) ;
  assign w15705 = \pi050 ^ w15704 ;
  assign w15706 = ( ~w15659 & w15660 ) | ( ~w15659 & w15668 ) | ( w15660 & w15668 ) ;
  assign w15707 = ~\pi119 & w5802 ;
  assign w15708 = \pi118 & w6052 ;
  assign w15709 = ( w5802 & ~w15707 ) | ( w5802 & w15708 ) | ( ~w15707 & w15708 ) ;
  assign w15710 = ~\pi120 & w5804 ;
  assign w15711 = w6634 | w15709 ;
  assign w15712 = ( w5805 & w15709 ) | ( w5805 & w15711 ) | ( w15709 & w15711 ) ;
  assign w15713 = ( w5804 & ~w15710 ) | ( w5804 & w15712 ) | ( ~w15710 & w15712 ) ;
  assign w15714 = \pi053 ^ w15713 ;
  assign w15715 = ( ~w15648 & w15649 ) | ( ~w15648 & w15657 ) | ( w15649 & w15657 ) ;
  assign w15716 = ~\pi116 & w6466 ;
  assign w15717 = \pi115 & w6702 ;
  assign w15718 = ( w6466 & ~w15716 ) | ( w6466 & w15717 ) | ( ~w15716 & w15717 ) ;
  assign w15719 = ~\pi117 & w6468 ;
  assign w15720 = w6185 | w15718 ;
  assign w15721 = ( w6469 & w15718 ) | ( w6469 & w15720 ) | ( w15718 & w15720 ) ;
  assign w15722 = ( w6468 & ~w15719 ) | ( w6468 & w15721 ) | ( ~w15719 & w15721 ) ;
  assign w15723 = \pi056 ^ w15722 ;
  assign w15724 = ( w15619 & ~w15638 ) | ( w15619 & w15646 ) | ( ~w15638 & w15646 ) ;
  assign w15725 = ~\pi113 & w7135 ;
  assign w15726 = \pi112 & w7359 ;
  assign w15727 = ( w7135 & ~w15725 ) | ( w7135 & w15726 ) | ( ~w15725 & w15726 ) ;
  assign w15728 = ~\pi114 & w7137 ;
  assign w15729 = w5565 | w15727 ;
  assign w15730 = ( w7138 & w15727 ) | ( w7138 & w15729 ) | ( w15727 & w15729 ) ;
  assign w15731 = ( w7137 & ~w15728 ) | ( w7137 & w15730 ) | ( ~w15728 & w15730 ) ;
  assign w15732 = \pi059 ^ w15731 ;
  assign w15733 = w4792 | w15633 ;
  assign w15734 = ( w7814 & w15633 ) | ( w7814 & w15733 ) | ( w15633 & w15733 ) ;
  assign w15735 = \pi062 ^ w15734 ;
  assign w15736 = ( ~w15623 & w15628 ) | ( ~w15623 & w15735 ) | ( w15628 & w15735 ) ;
  assign w15737 = ~\pi110 & w7811 ;
  assign w15738 = \pi109 & w8046 ;
  assign w15739 = ( w7811 & ~w15737 ) | ( w7811 & w15738 ) | ( ~w15737 & w15738 ) ;
  assign w15740 = ~\pi111 & w7813 ;
  assign w15741 = ~w4811 & w7814 ;
  assign w15742 = ( w7814 & w15739 ) | ( w7814 & ~w15741 ) | ( w15739 & ~w15741 ) ;
  assign w15743 = ( w7813 & ~w15740 ) | ( w7813 & w15742 ) | ( ~w15740 & w15742 ) ;
  assign w15744 = ~\pi063 & \pi107 ;
  assign w15745 = ( \pi062 & ~w15621 ) | ( \pi062 & w15744 ) | ( ~w15621 & w15744 ) ;
  assign w15746 = w15743 ^ w15745 ;
  assign w15747 = \pi107 ^ w15746 ;
  assign w15748 = ( \pi063 & w15743 ) | ( \pi063 & ~w15744 ) | ( w15743 & ~w15744 ) ;
  assign w15749 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15748 ) | ( ~\pi063 & w15748 ) ;
  assign w15750 = ( \pi062 & ~w15747 ) | ( \pi062 & w15749 ) | ( ~w15747 & w15749 ) ;
  assign w15751 = ( \pi063 & \pi108 ) | ( \pi063 & w15750 ) | ( \pi108 & w15750 ) ;
  assign w15752 = w15747 ^ w15751 ;
  assign w15753 = w15732 ^ w15752 ;
  assign w15754 = w15736 ^ w15753 ;
  assign w15755 = w15724 ^ w15754 ;
  assign w15756 = w15723 ^ w15755 ;
  assign w15757 = w15714 ^ w15715 ;
  assign w15758 = w15756 ^ w15757 ;
  assign w15759 = w15705 ^ w15706 ;
  assign w15760 = w15758 ^ w15759 ;
  assign w15761 = ( w15618 & ~w15670 ) | ( w15618 & w15678 ) | ( ~w15670 & w15678 ) ;
  assign w15762 = ~\pi125 & w4654 ;
  assign w15763 = \pi124 & w4876 ;
  assign w15764 = ( w4654 & ~w15762 ) | ( w4654 & w15763 ) | ( ~w15762 & w15763 ) ;
  assign w15765 = ~\pi126 & w4656 ;
  assign w15766 = w8231 | w15764 ;
  assign w15767 = ( w4657 & w15764 ) | ( w4657 & w15766 ) | ( w15764 & w15766 ) ;
  assign w15768 = ( w4656 & ~w15765 ) | ( w4656 & w15767 ) | ( ~w15765 & w15767 ) ;
  assign w15769 = \pi047 ^ w15768 ;
  assign w15770 = w15760 ^ w15769 ;
  assign w15771 = w15761 ^ w15770 ;
  assign w15772 = w15697 ^ w15771 ;
  assign w15773 = w15693 ^ w15772 ;
  assign w15774 = w15690 ^ w15773 ;
  assign w15775 = w15692 ^ w15774 ;
  assign w15776 = ( w15690 & ~w15692 ) | ( w15690 & w15773 ) | ( ~w15692 & w15773 ) ;
  assign w15777 = ~\pi126 & w4654 ;
  assign w15778 = \pi125 & w4876 ;
  assign w15779 = ( w4654 & ~w15777 ) | ( w4654 & w15778 ) | ( ~w15777 & w15778 ) ;
  assign w15780 = ~\pi127 & w4656 ;
  assign w15781 = w8466 | w15779 ;
  assign w15782 = ( w4657 & w15779 ) | ( w4657 & w15781 ) | ( w15779 & w15781 ) ;
  assign w15783 = ( w4656 & ~w15780 ) | ( w4656 & w15782 ) | ( ~w15780 & w15782 ) ;
  assign w15784 = \pi047 ^ w15783 ;
  assign w15785 = ( w15705 & w15706 ) | ( w15705 & ~w15758 ) | ( w15706 & ~w15758 ) ;
  assign w15786 = ~\pi123 & w5209 ;
  assign w15787 = \pi122 & w5433 ;
  assign w15788 = ( w5209 & ~w15786 ) | ( w5209 & w15787 ) | ( ~w15786 & w15787 ) ;
  assign w15789 = ~\pi124 & w5211 ;
  assign w15790 = w7538 | w15788 ;
  assign w15791 = ( w5212 & w15788 ) | ( w5212 & w15790 ) | ( w15788 & w15790 ) ;
  assign w15792 = ( w5211 & ~w15789 ) | ( w5211 & w15791 ) | ( ~w15789 & w15791 ) ;
  assign w15793 = \pi050 ^ w15792 ;
  assign w15794 = ( w15714 & w15715 ) | ( w15714 & ~w15756 ) | ( w15715 & ~w15756 ) ;
  assign w15795 = ~\pi120 & w5802 ;
  assign w15796 = \pi119 & w6052 ;
  assign w15797 = ( w5802 & ~w15795 ) | ( w5802 & w15796 ) | ( ~w15795 & w15796 ) ;
  assign w15798 = ~\pi121 & w5804 ;
  assign w15799 = w7050 | w15797 ;
  assign w15800 = ( w5805 & w15797 ) | ( w5805 & w15799 ) | ( w15797 & w15799 ) ;
  assign w15801 = ( w5804 & ~w15798 ) | ( w5804 & w15800 ) | ( ~w15798 & w15800 ) ;
  assign w15802 = \pi053 ^ w15801 ;
  assign w15803 = ( w15723 & w15724 ) | ( w15723 & ~w15754 ) | ( w15724 & ~w15754 ) ;
  assign w15804 = ~\pi117 & w6466 ;
  assign w15805 = \pi116 & w6702 ;
  assign w15806 = ( w6466 & ~w15804 ) | ( w6466 & w15805 ) | ( ~w15804 & w15805 ) ;
  assign w15807 = ~\pi118 & w6468 ;
  assign w15808 = w6206 | w15806 ;
  assign w15809 = ( w6469 & w15806 ) | ( w6469 & w15808 ) | ( w15806 & w15808 ) ;
  assign w15810 = ( w6468 & ~w15807 ) | ( w6468 & w15809 ) | ( ~w15807 & w15809 ) ;
  assign w15811 = \pi056 ^ w15810 ;
  assign w15812 = ( w15732 & w15736 ) | ( w15732 & ~w15752 ) | ( w15736 & ~w15752 ) ;
  assign w15813 = \pi063 ^ w15743 ;
  assign w15814 = ( \pi107 & ~\pi108 ) | ( \pi107 & w15813 ) | ( ~\pi108 & w15813 ) ;
  assign w15815 = w8323 ^ w15814 ;
  assign w15816 = ( \pi106 & \pi107 ) | ( \pi106 & ~w15743 ) | ( \pi107 & ~w15743 ) ;
  assign w15817 = ( \pi107 & w15813 ) | ( \pi107 & ~w15816 ) | ( w15813 & ~w15816 ) ;
  assign w15818 = ( ~w15814 & w15815 ) | ( ~w15814 & w15817 ) | ( w15815 & w15817 ) ;
  assign w15819 = ( \pi062 & \pi063 ) | ( \pi062 & \pi109 ) | ( \pi063 & \pi109 ) ;
  assign w15820 = \pi108 | w8323 ;
  assign w15821 = w15819 & w15820 ;
  assign w15822 = \pi044 ^ w15821 ;
  assign w15823 = ~\pi111 & w7811 ;
  assign w15824 = \pi110 & w8046 ;
  assign w15825 = ( w7811 & ~w15823 ) | ( w7811 & w15824 ) | ( ~w15823 & w15824 ) ;
  assign w15826 = ~\pi112 & w7813 ;
  assign w15827 = w4999 | w15825 ;
  assign w15828 = ( w7814 & w15825 ) | ( w7814 & w15827 ) | ( w15825 & w15827 ) ;
  assign w15829 = ( w7813 & ~w15826 ) | ( w7813 & w15828 ) | ( ~w15826 & w15828 ) ;
  assign w15830 = \pi062 ^ w15829 ;
  assign w15831 = w15623 ^ w15822 ;
  assign w15832 = w15818 ^ w15831 ;
  assign w15833 = w15830 ^ w15832 ;
  assign w15834 = ~\pi114 & w7135 ;
  assign w15835 = \pi113 & w7359 ;
  assign w15836 = ( w7135 & ~w15834 ) | ( w7135 & w15835 ) | ( ~w15834 & w15835 ) ;
  assign w15837 = ~\pi115 & w7137 ;
  assign w15838 = w5585 | w15836 ;
  assign w15839 = ( w7138 & w15836 ) | ( w7138 & w15838 ) | ( w15836 & w15838 ) ;
  assign w15840 = ( w7137 & ~w15837 ) | ( w7137 & w15839 ) | ( ~w15837 & w15839 ) ;
  assign w15841 = \pi059 ^ w15840 ;
  assign w15842 = w15812 ^ w15833 ;
  assign w15843 = w15841 ^ w15842 ;
  assign w15844 = w15803 ^ w15843 ;
  assign w15845 = w15811 ^ w15844 ;
  assign w15846 = w15794 ^ w15802 ;
  assign w15847 = w15845 ^ w15846 ;
  assign w15848 = w15785 ^ w15793 ;
  assign w15849 = w15847 ^ w15848 ;
  assign w15850 = ( ~w15760 & w15761 ) | ( ~w15760 & w15769 ) | ( w15761 & w15769 ) ;
  assign w15851 = w15784 ^ w15850 ;
  assign w15852 = w15849 ^ w15851 ;
  assign w15853 = ( w15693 & w15697 ) | ( w15693 & ~w15771 ) | ( w15697 & ~w15771 ) ;
  assign w15854 = w15776 ^ w15852 ;
  assign w15855 = w15853 ^ w15854 ;
  assign w15856 = ( w15785 & w15793 ) | ( w15785 & ~w15847 ) | ( w15793 & ~w15847 ) ;
  assign w15857 = \pi127 & w4654 ;
  assign w15858 = ( \pi126 & ~w4657 ) | ( \pi126 & w8490 ) | ( ~w4657 & w8490 ) ;
  assign w15859 = \pi126 & ~w4876 ;
  assign w15860 = ( ~\pi126 & w15858 ) | ( ~\pi126 & w15859 ) | ( w15858 & w15859 ) ;
  assign w15861 = ( w9420 & w15857 ) | ( w9420 & ~w15860 ) | ( w15857 & ~w15860 ) ;
  assign w15862 = ~\pi124 & w5209 ;
  assign w15863 = \pi123 & w5433 ;
  assign w15864 = ( w5209 & ~w15862 ) | ( w5209 & w15863 ) | ( ~w15862 & w15863 ) ;
  assign w15865 = ~\pi125 & w5211 ;
  assign w15866 = w7988 | w15864 ;
  assign w15867 = ( w5212 & w15864 ) | ( w5212 & w15866 ) | ( w15864 & w15866 ) ;
  assign w15868 = ( w5211 & ~w15865 ) | ( w5211 & w15867 ) | ( ~w15865 & w15867 ) ;
  assign w15869 = \pi050 ^ w15868 ;
  assign w15870 = ( w15794 & w15802 ) | ( w15794 & ~w15845 ) | ( w15802 & ~w15845 ) ;
  assign w15871 = ( w15803 & w15811 ) | ( w15803 & ~w15843 ) | ( w15811 & ~w15843 ) ;
  assign w15872 = ~\pi118 & w6466 ;
  assign w15873 = \pi117 & w6702 ;
  assign w15874 = ( w6466 & ~w15872 ) | ( w6466 & w15873 ) | ( ~w15872 & w15873 ) ;
  assign w15875 = ~\pi119 & w6468 ;
  assign w15876 = w6616 | w15874 ;
  assign w15877 = ( w6469 & w15874 ) | ( w6469 & w15876 ) | ( w15874 & w15876 ) ;
  assign w15878 = ( w6468 & ~w15875 ) | ( w6468 & w15877 ) | ( ~w15875 & w15877 ) ;
  assign w15879 = \pi056 ^ w15878 ;
  assign w15880 = ( w15812 & ~w15833 ) | ( w15812 & w15841 ) | ( ~w15833 & w15841 ) ;
  assign w15881 = ~\pi115 & w7135 ;
  assign w15882 = \pi114 & w7359 ;
  assign w15883 = ( w7135 & ~w15881 ) | ( w7135 & w15882 ) | ( ~w15881 & w15882 ) ;
  assign w15884 = ~\pi116 & w7137 ;
  assign w15885 = w5976 | w15883 ;
  assign w15886 = ( w7138 & w15883 ) | ( w7138 & w15885 ) | ( w15883 & w15885 ) ;
  assign w15887 = ( w7137 & ~w15884 ) | ( w7137 & w15886 ) | ( ~w15884 & w15886 ) ;
  assign w15888 = \pi059 ^ w15887 ;
  assign w15889 = ( w15818 & w15830 ) | ( w15818 & ~w15831 ) | ( w15830 & ~w15831 ) ;
  assign w15890 = \pi063 & \pi108 ;
  assign w15891 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w15890 ) | ( \pi063 & w15890 ) ;
  assign w15892 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15890 ) | ( ~\pi063 & w15890 ) ;
  assign w15893 = ( \pi109 & w15891 ) | ( \pi109 & w15892 ) | ( w15891 & w15892 ) ;
  assign w15894 = ( ~\pi044 & w15623 ) | ( ~\pi044 & w15893 ) | ( w15623 & w15893 ) ;
  assign w15895 = ~\pi112 & w7811 ;
  assign w15896 = \pi111 & w8046 ;
  assign w15897 = ( w7811 & ~w15895 ) | ( w7811 & w15896 ) | ( ~w15895 & w15896 ) ;
  assign w15898 = ~\pi113 & w7813 ;
  assign w15899 = w5366 | w15897 ;
  assign w15900 = ( w7814 & w15897 ) | ( w7814 & w15899 ) | ( w15897 & w15899 ) ;
  assign w15901 = ( w7813 & ~w15898 ) | ( w7813 & w15900 ) | ( ~w15898 & w15900 ) ;
  assign w15902 = \pi062 ^ w15901 ;
  assign w15903 = w15894 ^ w15902 ;
  assign w15904 = ( \pi062 & \pi063 ) | ( \pi062 & \pi110 ) | ( \pi063 & \pi110 ) ;
  assign w15905 = \pi063 & ~\pi109 ;
  assign w15906 = \pi062 & w15905 ;
  assign w15907 = w15904 ^ w15906 ;
  assign w15908 = w15903 ^ w15907 ;
  assign w15909 = w15888 ^ w15889 ;
  assign w15910 = w15908 ^ w15909 ;
  assign w15911 = w15879 ^ w15880 ;
  assign w15912 = w15910 ^ w15911 ;
  assign w15913 = ~\pi121 & w5802 ;
  assign w15914 = \pi120 & w6052 ;
  assign w15915 = ( w5802 & ~w15913 ) | ( w5802 & w15914 ) | ( ~w15913 & w15914 ) ;
  assign w15916 = ~\pi122 & w5804 ;
  assign w15917 = w7069 | w15915 ;
  assign w15918 = ( w5805 & w15915 ) | ( w5805 & w15917 ) | ( w15915 & w15917 ) ;
  assign w15919 = ( w5804 & ~w15916 ) | ( w5804 & w15918 ) | ( ~w15916 & w15918 ) ;
  assign w15920 = \pi053 ^ w15919 ;
  assign w15921 = w15871 ^ w15920 ;
  assign w15922 = w15912 ^ w15921 ;
  assign w15923 = w15869 ^ w15922 ;
  assign w15924 = w15870 ^ w15923 ;
  assign w15925 = \pi047 ^ w15856 ;
  assign w15926 = w15861 ^ w15925 ;
  assign w15927 = w15924 ^ w15926 ;
  assign w15928 = ( w15784 & ~w15849 ) | ( w15784 & w15850 ) | ( ~w15849 & w15850 ) ;
  assign w15929 = ( w15776 & w15852 ) | ( w15776 & ~w15853 ) | ( w15852 & ~w15853 ) ;
  assign w15930 = w15928 ^ w15929 ;
  assign w15931 = w15927 ^ w15930 ;
  assign w15932 = ~\pi122 & w5802 ;
  assign w15933 = \pi121 & w6052 ;
  assign w15934 = ( w5802 & ~w15932 ) | ( w5802 & w15933 ) | ( ~w15932 & w15933 ) ;
  assign w15935 = ~\pi123 & w5804 ;
  assign w15936 = w7516 | w15934 ;
  assign w15937 = ( w5805 & w15934 ) | ( w5805 & w15936 ) | ( w15934 & w15936 ) ;
  assign w15938 = ( w5804 & ~w15935 ) | ( w5804 & w15937 ) | ( ~w15935 & w15937 ) ;
  assign w15939 = \pi053 ^ w15938 ;
  assign w15940 = ( w15879 & w15880 ) | ( w15879 & ~w15910 ) | ( w15880 & ~w15910 ) ;
  assign w15941 = ~\pi119 & w6466 ;
  assign w15942 = \pi118 & w6702 ;
  assign w15943 = ( w6466 & ~w15941 ) | ( w6466 & w15942 ) | ( ~w15941 & w15942 ) ;
  assign w15944 = ~\pi120 & w6468 ;
  assign w15945 = w6634 | w15943 ;
  assign w15946 = ( w6469 & w15943 ) | ( w6469 & w15945 ) | ( w15943 & w15945 ) ;
  assign w15947 = ( w6468 & ~w15944 ) | ( w6468 & w15946 ) | ( ~w15944 & w15946 ) ;
  assign w15948 = \pi056 ^ w15947 ;
  assign w15949 = ( w15888 & w15889 ) | ( w15888 & ~w15908 ) | ( w15889 & ~w15908 ) ;
  assign w15950 = ~\pi116 & w7135 ;
  assign w15951 = \pi115 & w7359 ;
  assign w15952 = ( w7135 & ~w15950 ) | ( w7135 & w15951 ) | ( ~w15950 & w15951 ) ;
  assign w15953 = ~\pi117 & w7137 ;
  assign w15954 = w6185 | w15952 ;
  assign w15955 = ( w7138 & w15952 ) | ( w7138 & w15954 ) | ( w15952 & w15954 ) ;
  assign w15956 = ( w7137 & ~w15953 ) | ( w7137 & w15955 ) | ( ~w15953 & w15955 ) ;
  assign w15957 = \pi059 ^ w15956 ;
  assign w15958 = \pi063 & \pi109 ;
  assign w15959 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w15958 ) | ( \pi063 & w15958 ) ;
  assign w15960 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15958 ) | ( ~\pi063 & w15958 ) ;
  assign w15961 = ( \pi110 & w15959 ) | ( \pi110 & w15960 ) | ( w15959 & w15960 ) ;
  assign w15962 = ( w15894 & w15902 ) | ( w15894 & ~w15961 ) | ( w15902 & ~w15961 ) ;
  assign w15963 = \pi110 & ~w15962 ;
  assign w15964 = ( \pi063 & ~\pi109 ) | ( \pi063 & w15963 ) | ( ~\pi109 & w15963 ) ;
  assign w15965 = ( \pi062 & ~\pi063 ) | ( \pi062 & w15964 ) | ( ~\pi063 & w15964 ) ;
  assign w15966 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi111 ) | ( \pi063 & ~\pi111 ) ;
  assign w15967 = ( \pi110 & w15962 ) | ( \pi110 & w15966 ) | ( w15962 & w15966 ) ;
  assign w15968 = ( ~\pi063 & w15962 ) | ( ~\pi063 & w15963 ) | ( w15962 & w15963 ) ;
  assign w15969 = ( \pi062 & ~\pi110 ) | ( \pi062 & w15968 ) | ( ~\pi110 & w15968 ) ;
  assign w15970 = ( ~w15965 & w15967 ) | ( ~w15965 & w15969 ) | ( w15967 & w15969 ) ;
  assign w15971 = \pi109 ^ \pi111 ;
  assign w15972 = ( \pi062 & \pi063 ) | ( \pi062 & ~w15971 ) | ( \pi063 & ~w15971 ) ;
  assign w15973 = \pi109 ^ \pi110 ;
  assign w15974 = \pi062 & ~w15973 ;
  assign w15975 = ( \pi063 & ~w15973 ) | ( \pi063 & w15974 ) | ( ~w15973 & w15974 ) ;
  assign w15976 = w15962 ^ w15975 ;
  assign w15977 = w15972 ^ w15976 ;
  assign w15978 = ~\pi113 & w7811 ;
  assign w15979 = \pi112 & w8046 ;
  assign w15980 = ( w7811 & ~w15978 ) | ( w7811 & w15979 ) | ( ~w15978 & w15979 ) ;
  assign w15981 = ~\pi114 & w7813 ;
  assign w15982 = w5565 | w15980 ;
  assign w15983 = ( w7814 & w15980 ) | ( w7814 & w15982 ) | ( w15980 & w15982 ) ;
  assign w15984 = ( w7813 & ~w15981 ) | ( w7813 & w15983 ) | ( ~w15981 & w15983 ) ;
  assign w15985 = \pi062 ^ w15984 ;
  assign w15986 = w15957 ^ w15977 ;
  assign w15987 = w15985 ^ w15986 ;
  assign w15988 = w15948 ^ w15949 ;
  assign w15989 = w15987 ^ w15988 ;
  assign w15990 = w15939 ^ w15989 ;
  assign w15991 = w15940 ^ w15990 ;
  assign w15992 = ( w15871 & ~w15912 ) | ( w15871 & w15920 ) | ( ~w15912 & w15920 ) ;
  assign w15993 = ~\pi125 & w5209 ;
  assign w15994 = \pi124 & w5433 ;
  assign w15995 = ( w5209 & ~w15993 ) | ( w5209 & w15994 ) | ( ~w15993 & w15994 ) ;
  assign w15996 = ~\pi126 & w5211 ;
  assign w15997 = w8231 | w15995 ;
  assign w15998 = ( w5212 & w15995 ) | ( w5212 & w15997 ) | ( w15995 & w15997 ) ;
  assign w15999 = ( w5211 & ~w15996 ) | ( w5211 & w15998 ) | ( ~w15996 & w15998 ) ;
  assign w16000 = \pi050 ^ w15999 ;
  assign w16001 = w15991 ^ w16000 ;
  assign w16002 = w15992 ^ w16001 ;
  assign w16003 = ( w15869 & w15870 ) | ( w15869 & ~w15922 ) | ( w15870 & ~w15922 ) ;
  assign w16004 = w4657 & w8481 ;
  assign w16005 = w4876 | w16004 ;
  assign w16006 = ( \pi127 & w16004 ) | ( \pi127 & w16005 ) | ( w16004 & w16005 ) ;
  assign w16007 = \pi047 ^ w16006 ;
  assign w16008 = w16002 ^ w16007 ;
  assign w16009 = w16003 ^ w16008 ;
  assign w16010 = \pi047 ^ w15861 ;
  assign w16011 = ( w15856 & ~w15924 ) | ( w15856 & w16010 ) | ( ~w15924 & w16010 ) ;
  assign w16012 = ( w15927 & ~w15928 ) | ( w15927 & w15929 ) | ( ~w15928 & w15929 ) ;
  assign w16013 = w16009 ^ w16012 ;
  assign w16014 = w16011 ^ w16013 ;
  assign w16015 = ~\pi126 & w5209 ;
  assign w16016 = \pi125 & w5433 ;
  assign w16017 = ( w5209 & ~w16015 ) | ( w5209 & w16016 ) | ( ~w16015 & w16016 ) ;
  assign w16018 = ~\pi127 & w5211 ;
  assign w16019 = w8466 | w16017 ;
  assign w16020 = ( w5212 & w16017 ) | ( w5212 & w16019 ) | ( w16017 & w16019 ) ;
  assign w16021 = ( w5211 & ~w16018 ) | ( w5211 & w16020 ) | ( ~w16018 & w16020 ) ;
  assign w16022 = \pi050 ^ w16021 ;
  assign w16023 = ( w15939 & w15940 ) | ( w15939 & ~w15989 ) | ( w15940 & ~w15989 ) ;
  assign w16024 = ~\pi123 & w5802 ;
  assign w16025 = \pi122 & w6052 ;
  assign w16026 = ( w5802 & ~w16024 ) | ( w5802 & w16025 ) | ( ~w16024 & w16025 ) ;
  assign w16027 = ~\pi124 & w5804 ;
  assign w16028 = w7538 | w16026 ;
  assign w16029 = ( w5805 & w16026 ) | ( w5805 & w16028 ) | ( w16026 & w16028 ) ;
  assign w16030 = ( w5804 & ~w16027 ) | ( w5804 & w16029 ) | ( ~w16027 & w16029 ) ;
  assign w16031 = \pi053 ^ w16030 ;
  assign w16032 = ( w15948 & w15949 ) | ( w15948 & ~w15987 ) | ( w15949 & ~w15987 ) ;
  assign w16033 = ~\pi120 & w6466 ;
  assign w16034 = \pi119 & w6702 ;
  assign w16035 = ( w6466 & ~w16033 ) | ( w6466 & w16034 ) | ( ~w16033 & w16034 ) ;
  assign w16036 = ~\pi121 & w6468 ;
  assign w16037 = w7050 | w16035 ;
  assign w16038 = ( w6469 & w16035 ) | ( w6469 & w16037 ) | ( w16035 & w16037 ) ;
  assign w16039 = ( w6468 & ~w16036 ) | ( w6468 & w16038 ) | ( ~w16036 & w16038 ) ;
  assign w16040 = \pi056 ^ w16039 ;
  assign w16041 = ( w15957 & ~w15977 ) | ( w15957 & w15985 ) | ( ~w15977 & w15985 ) ;
  assign w16042 = ~\pi114 & w7811 ;
  assign w16043 = \pi113 & w8046 ;
  assign w16044 = ( w7811 & ~w16042 ) | ( w7811 & w16043 ) | ( ~w16042 & w16043 ) ;
  assign w16045 = ~\pi115 & w7813 ;
  assign w16046 = w5585 | w16044 ;
  assign w16047 = ( w7814 & w16044 ) | ( w7814 & w16046 ) | ( w16044 & w16046 ) ;
  assign w16048 = ( w7813 & ~w16045 ) | ( w7813 & w16047 ) | ( ~w16045 & w16047 ) ;
  assign w16049 = \pi062 ^ w16048 ;
  assign w16050 = \pi110 ^ \pi112 ;
  assign w16051 = ( \pi062 & \pi063 ) | ( \pi062 & ~w16050 ) | ( \pi063 & ~w16050 ) ;
  assign w16052 = \pi110 ^ \pi111 ;
  assign w16053 = \pi062 & ~w16052 ;
  assign w16054 = ( \pi063 & ~w16052 ) | ( \pi063 & w16053 ) | ( ~w16052 & w16053 ) ;
  assign w16055 = \pi047 ^ w16054 ;
  assign w16056 = w16051 ^ w16055 ;
  assign w16057 = w15970 ^ w16049 ;
  assign w16058 = w16056 ^ w16057 ;
  assign w16059 = ~\pi117 & w7135 ;
  assign w16060 = \pi116 & w7359 ;
  assign w16061 = ( w7135 & ~w16059 ) | ( w7135 & w16060 ) | ( ~w16059 & w16060 ) ;
  assign w16062 = ~\pi118 & w7137 ;
  assign w16063 = w6206 | w16061 ;
  assign w16064 = ( w7138 & w16061 ) | ( w7138 & w16063 ) | ( w16061 & w16063 ) ;
  assign w16065 = ( w7137 & ~w16062 ) | ( w7137 & w16064 ) | ( ~w16062 & w16064 ) ;
  assign w16066 = \pi059 ^ w16065 ;
  assign w16067 = w16041 ^ w16058 ;
  assign w16068 = w16066 ^ w16067 ;
  assign w16069 = w16032 ^ w16040 ;
  assign w16070 = w16068 ^ w16069 ;
  assign w16071 = w16023 ^ w16031 ;
  assign w16072 = w16070 ^ w16071 ;
  assign w16073 = ( ~w15991 & w15992 ) | ( ~w15991 & w16000 ) | ( w15992 & w16000 ) ;
  assign w16074 = w16022 ^ w16073 ;
  assign w16075 = w16072 ^ w16074 ;
  assign w16076 = ( ~w16002 & w16003 ) | ( ~w16002 & w16007 ) | ( w16003 & w16007 ) ;
  assign w16077 = ( w16009 & ~w16011 ) | ( w16009 & w16012 ) | ( ~w16011 & w16012 ) ;
  assign w16078 = w16075 ^ w16077 ;
  assign w16079 = w16076 ^ w16078 ;
  assign w16080 = \pi127 & w5209 ;
  assign w16081 = ( \pi126 & w5433 ) | ( \pi126 & w16080 ) | ( w5433 & w16080 ) ;
  assign w16082 = ( \pi126 & ~w8464 ) | ( \pi126 & w16081 ) | ( ~w8464 & w16081 ) ;
  assign w16083 = ( \pi127 & ~w5212 ) | ( \pi127 & w8464 ) | ( ~w5212 & w8464 ) ;
  assign w16084 = ( ~w16080 & w16082 ) | ( ~w16080 & w16083 ) | ( w16082 & w16083 ) ;
  assign w16085 = \pi126 | \pi127 ;
  assign w16086 = ( w16081 & ~w16084 ) | ( w16081 & w16085 ) | ( ~w16084 & w16085 ) ;
  assign w16087 = ( w16023 & w16031 ) | ( w16023 & ~w16070 ) | ( w16031 & ~w16070 ) ;
  assign w16088 = ~\pi124 & w5802 ;
  assign w16089 = \pi123 & w6052 ;
  assign w16090 = ( w5802 & ~w16088 ) | ( w5802 & w16089 ) | ( ~w16088 & w16089 ) ;
  assign w16091 = ~\pi125 & w5804 ;
  assign w16092 = w7988 | w16090 ;
  assign w16093 = ( w5805 & w16090 ) | ( w5805 & w16092 ) | ( w16090 & w16092 ) ;
  assign w16094 = ( w5804 & ~w16091 ) | ( w5804 & w16093 ) | ( ~w16091 & w16093 ) ;
  assign w16095 = \pi053 ^ w16094 ;
  assign w16096 = ( w16032 & w16040 ) | ( w16032 & ~w16068 ) | ( w16040 & ~w16068 ) ;
  assign w16097 = ~\pi121 & w6466 ;
  assign w16098 = \pi120 & w6702 ;
  assign w16099 = ( w6466 & ~w16097 ) | ( w6466 & w16098 ) | ( ~w16097 & w16098 ) ;
  assign w16100 = ~\pi122 & w6468 ;
  assign w16101 = w7069 | w16099 ;
  assign w16102 = ( w6469 & w16099 ) | ( w6469 & w16101 ) | ( w16099 & w16101 ) ;
  assign w16103 = ( w6468 & ~w16100 ) | ( w6468 & w16102 ) | ( ~w16100 & w16102 ) ;
  assign w16104 = \pi056 ^ w16103 ;
  assign w16105 = ( w16041 & ~w16058 ) | ( w16041 & w16066 ) | ( ~w16058 & w16066 ) ;
  assign w16106 = ~\pi118 & w7135 ;
  assign w16107 = \pi117 & w7359 ;
  assign w16108 = ( w7135 & ~w16106 ) | ( w7135 & w16107 ) | ( ~w16106 & w16107 ) ;
  assign w16109 = ~\pi119 & w7137 ;
  assign w16110 = w6616 | w16108 ;
  assign w16111 = ( w7138 & w16108 ) | ( w7138 & w16110 ) | ( w16108 & w16110 ) ;
  assign w16112 = ( w7137 & ~w16109 ) | ( w7137 & w16111 ) | ( ~w16109 & w16111 ) ;
  assign w16113 = \pi059 ^ w16112 ;
  assign w16114 = ( w15970 & w16049 ) | ( w15970 & ~w16056 ) | ( w16049 & ~w16056 ) ;
  assign w16115 = ( \pi062 & \pi063 ) | ( \pi062 & \pi113 ) | ( \pi063 & \pi113 ) ;
  assign w16116 = \pi063 & ~\pi112 ;
  assign w16117 = w16115 & ~w16116 ;
  assign w16118 = ( ~\pi062 & w16115 ) | ( ~\pi062 & w16117 ) | ( w16115 & w16117 ) ;
  assign w16119 = \pi063 ^ \pi110 ;
  assign w16120 = \pi062 ^ w16119 ;
  assign w16121 = ( \pi110 & \pi112 ) | ( \pi110 & w16120 ) | ( \pi112 & w16120 ) ;
  assign w16122 = ( ~\pi047 & \pi111 ) | ( ~\pi047 & w16121 ) | ( \pi111 & w16121 ) ;
  assign w16123 = w10655 & w16122 ;
  assign w16124 = \pi114 & w8046 ;
  assign w16125 = ( \pi116 & w7813 ) | ( \pi116 & w16124 ) | ( w7813 & w16124 ) ;
  assign w16126 = \pi115 | w16125 ;
  assign w16127 = ( w7811 & w16125 ) | ( w7811 & w16126 ) | ( w16125 & w16126 ) ;
  assign w16128 = w16124 | w16127 ;
  assign w16129 = ~w5976 & w7814 ;
  assign w16130 = ( w7814 & w16128 ) | ( w7814 & ~w16129 ) | ( w16128 & ~w16129 ) ;
  assign w16131 = w16118 ^ w16130 ;
  assign w16132 = \pi062 ^ w16123 ;
  assign w16133 = w16131 ^ w16132 ;
  assign w16134 = w16113 ^ w16114 ;
  assign w16135 = w16133 ^ w16134 ;
  assign w16136 = w16104 ^ w16105 ;
  assign w16137 = w16135 ^ w16136 ;
  assign w16138 = w16095 ^ w16137 ;
  assign w16139 = w16096 ^ w16138 ;
  assign w16140 = \pi050 ^ w16087 ;
  assign w16141 = w16086 ^ w16140 ;
  assign w16142 = w16139 ^ w16141 ;
  assign w16143 = ( w16022 & ~w16072 ) | ( w16022 & w16073 ) | ( ~w16072 & w16073 ) ;
  assign w16144 = ( w16075 & ~w16076 ) | ( w16075 & w16077 ) | ( ~w16076 & w16077 ) ;
  assign w16145 = w16143 ^ w16144 ;
  assign w16146 = w16142 ^ w16145 ;
  assign w16147 = ~\pi122 & w6466 ;
  assign w16148 = \pi121 & w6702 ;
  assign w16149 = ( w6466 & ~w16147 ) | ( w6466 & w16148 ) | ( ~w16147 & w16148 ) ;
  assign w16150 = ~\pi123 & w6468 ;
  assign w16151 = w7516 | w16149 ;
  assign w16152 = ( w6469 & w16149 ) | ( w6469 & w16151 ) | ( w16149 & w16151 ) ;
  assign w16153 = ( w6468 & ~w16150 ) | ( w6468 & w16152 ) | ( ~w16150 & w16152 ) ;
  assign w16154 = \pi056 ^ w16153 ;
  assign w16155 = ( w16113 & w16114 ) | ( w16113 & ~w16133 ) | ( w16114 & ~w16133 ) ;
  assign w16156 = ~\pi116 & w7811 ;
  assign w16157 = \pi115 & w8046 ;
  assign w16158 = ( w7811 & ~w16156 ) | ( w7811 & w16157 ) | ( ~w16156 & w16157 ) ;
  assign w16159 = ~\pi117 & w7813 ;
  assign w16160 = w6185 | w16158 ;
  assign w16161 = ( w7814 & w16158 ) | ( w7814 & w16160 ) | ( w16158 & w16160 ) ;
  assign w16162 = ( w7813 & ~w16159 ) | ( w7813 & w16161 ) | ( ~w16159 & w16161 ) ;
  assign w16163 = \pi062 ^ w16162 ;
  assign w16164 = \pi112 ^ \pi114 ;
  assign w16165 = ( \pi062 & \pi063 ) | ( \pi062 & ~w16164 ) | ( \pi063 & ~w16164 ) ;
  assign w16166 = \pi062 & ~w5365 ;
  assign w16167 = ( \pi063 & ~w5365 ) | ( \pi063 & w16166 ) | ( ~w5365 & w16166 ) ;
  assign w16168 = w16163 ^ w16167 ;
  assign w16169 = w16165 ^ w16168 ;
  assign w16170 = w5976 | w16128 ;
  assign w16171 = ( w7814 & w16128 ) | ( w7814 & w16170 ) | ( w16128 & w16170 ) ;
  assign w16172 = \pi062 ^ w16171 ;
  assign w16173 = ( ~w16118 & w16123 ) | ( ~w16118 & w16172 ) | ( w16123 & w16172 ) ;
  assign w16174 = ~\pi119 & w7135 ;
  assign w16175 = \pi118 & w7359 ;
  assign w16176 = ( w7135 & ~w16174 ) | ( w7135 & w16175 ) | ( ~w16174 & w16175 ) ;
  assign w16177 = ~\pi120 & w7137 ;
  assign w16178 = w6634 | w16176 ;
  assign w16179 = ( w7138 & w16176 ) | ( w7138 & w16178 ) | ( w16176 & w16178 ) ;
  assign w16180 = ( w7137 & ~w16177 ) | ( w7137 & w16179 ) | ( ~w16177 & w16179 ) ;
  assign w16181 = \pi059 ^ w16180 ;
  assign w16182 = w16169 ^ w16181 ;
  assign w16183 = w16173 ^ w16182 ;
  assign w16184 = w16154 ^ w16183 ;
  assign w16185 = w16155 ^ w16184 ;
  assign w16186 = ( w16104 & w16105 ) | ( w16104 & ~w16135 ) | ( w16105 & ~w16135 ) ;
  assign w16187 = ~\pi125 & w5802 ;
  assign w16188 = \pi124 & w6052 ;
  assign w16189 = ( w5802 & ~w16187 ) | ( w5802 & w16188 ) | ( ~w16187 & w16188 ) ;
  assign w16190 = ~\pi126 & w5804 ;
  assign w16191 = w8231 | w16189 ;
  assign w16192 = ( w5805 & w16189 ) | ( w5805 & w16191 ) | ( w16189 & w16191 ) ;
  assign w16193 = ( w5804 & ~w16190 ) | ( w5804 & w16192 ) | ( ~w16190 & w16192 ) ;
  assign w16194 = \pi053 ^ w16193 ;
  assign w16195 = w16185 ^ w16194 ;
  assign w16196 = w16186 ^ w16195 ;
  assign w16197 = ( w16095 & w16096 ) | ( w16095 & ~w16137 ) | ( w16096 & ~w16137 ) ;
  assign w16198 = w5212 & w8481 ;
  assign w16199 = w5433 | w16198 ;
  assign w16200 = ( \pi127 & w16198 ) | ( \pi127 & w16199 ) | ( w16198 & w16199 ) ;
  assign w16201 = \pi050 ^ w16200 ;
  assign w16202 = w16196 ^ w16201 ;
  assign w16203 = w16197 ^ w16202 ;
  assign w16204 = \pi050 ^ w16086 ;
  assign w16205 = ( w16087 & ~w16139 ) | ( w16087 & w16204 ) | ( ~w16139 & w16204 ) ;
  assign w16206 = ( w16142 & ~w16143 ) | ( w16142 & w16144 ) | ( ~w16143 & w16144 ) ;
  assign w16207 = w16203 ^ w16206 ;
  assign w16208 = w16205 ^ w16207 ;
  assign w16209 = ( w16154 & w16155 ) | ( w16154 & ~w16183 ) | ( w16155 & ~w16183 ) ;
  assign w16210 = ~\pi123 & w6466 ;
  assign w16211 = \pi122 & w6702 ;
  assign w16212 = ( w6466 & ~w16210 ) | ( w6466 & w16211 ) | ( ~w16210 & w16211 ) ;
  assign w16213 = ~\pi124 & w6468 ;
  assign w16214 = w7538 | w16212 ;
  assign w16215 = ( w6469 & w16212 ) | ( w6469 & w16214 ) | ( w16212 & w16214 ) ;
  assign w16216 = ( w6468 & ~w16213 ) | ( w6468 & w16215 ) | ( ~w16213 & w16215 ) ;
  assign w16217 = \pi056 ^ w16216 ;
  assign w16218 = ( ~w16169 & w16173 ) | ( ~w16169 & w16181 ) | ( w16173 & w16181 ) ;
  assign w16219 = ~\pi120 & w7135 ;
  assign w16220 = \pi119 & w7359 ;
  assign w16221 = ( w7135 & ~w16219 ) | ( w7135 & w16220 ) | ( ~w16219 & w16220 ) ;
  assign w16222 = ~\pi121 & w7137 ;
  assign w16223 = w7050 | w16221 ;
  assign w16224 = ( w7138 & w16221 ) | ( w7138 & w16223 ) | ( w16221 & w16223 ) ;
  assign w16225 = ( w7137 & ~w16222 ) | ( w7137 & w16224 ) | ( ~w16222 & w16224 ) ;
  assign w16226 = \pi059 ^ w16225 ;
  assign w16227 = ~\pi117 & w7811 ;
  assign w16228 = \pi116 & w8046 ;
  assign w16229 = ( w7811 & ~w16227 ) | ( w7811 & w16228 ) | ( ~w16227 & w16228 ) ;
  assign w16230 = ~\pi118 & w7813 ;
  assign w16231 = w6206 | w16229 ;
  assign w16232 = ( w7814 & w16229 ) | ( w7814 & w16231 ) | ( w16229 & w16231 ) ;
  assign w16233 = ( w7813 & ~w16230 ) | ( w7813 & w16232 ) | ( ~w16230 & w16232 ) ;
  assign w16234 = \pi062 ^ w16233 ;
  assign w16235 = \pi113 | w16163 ;
  assign w16236 = ( \pi063 & \pi112 ) | ( \pi063 & ~w16235 ) | ( \pi112 & ~w16235 ) ;
  assign w16237 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16236 ) | ( ~\pi063 & w16236 ) ;
  assign w16238 = ( \pi062 & \pi063 ) | ( \pi062 & \pi114 ) | ( \pi063 & \pi114 ) ;
  assign w16239 = ( ~\pi113 & w16163 ) | ( ~\pi113 & w16238 ) | ( w16163 & w16238 ) ;
  assign w16240 = ( \pi063 & ~w16163 ) | ( \pi063 & w16235 ) | ( ~w16163 & w16235 ) ;
  assign w16241 = ( \pi062 & \pi113 ) | ( \pi062 & ~w16240 ) | ( \pi113 & ~w16240 ) ;
  assign w16242 = ( ~w16237 & w16239 ) | ( ~w16237 & w16241 ) | ( w16239 & w16241 ) ;
  assign w16243 = \pi050 ^ w16118 ;
  assign w16244 = ( \pi062 & \pi063 ) | ( \pi062 & \pi115 ) | ( \pi063 & \pi115 ) ;
  assign w16245 = \pi063 & ~\pi114 ;
  assign w16246 = \pi062 & w16245 ;
  assign w16247 = w16244 ^ w16246 ;
  assign w16248 = w16243 ^ w16247 ;
  assign w16249 = w16234 ^ w16242 ;
  assign w16250 = w16248 ^ w16249 ;
  assign w16251 = w16218 ^ w16226 ;
  assign w16252 = w16250 ^ w16251 ;
  assign w16253 = w16209 ^ w16217 ;
  assign w16254 = w16252 ^ w16253 ;
  assign w16255 = ~\pi126 & w5802 ;
  assign w16256 = \pi125 & w6052 ;
  assign w16257 = ( w5802 & ~w16255 ) | ( w5802 & w16256 ) | ( ~w16255 & w16256 ) ;
  assign w16258 = ~\pi127 & w5804 ;
  assign w16259 = w8466 | w16257 ;
  assign w16260 = ( w5805 & w16257 ) | ( w5805 & w16259 ) | ( w16257 & w16259 ) ;
  assign w16261 = ( w5804 & ~w16258 ) | ( w5804 & w16260 ) | ( ~w16258 & w16260 ) ;
  assign w16262 = \pi053 ^ w16261 ;
  assign w16263 = ( ~w16185 & w16186 ) | ( ~w16185 & w16194 ) | ( w16186 & w16194 ) ;
  assign w16264 = w16262 ^ w16263 ;
  assign w16265 = w16254 ^ w16264 ;
  assign w16266 = ( ~w16196 & w16197 ) | ( ~w16196 & w16201 ) | ( w16197 & w16201 ) ;
  assign w16267 = ( w16203 & ~w16205 ) | ( w16203 & w16206 ) | ( ~w16205 & w16206 ) ;
  assign w16268 = w16265 ^ w16267 ;
  assign w16269 = w16266 ^ w16268 ;
  assign w16270 = \pi127 & w5802 ;
  assign w16271 = ( \pi126 & w6052 ) | ( \pi126 & w16270 ) | ( w6052 & w16270 ) ;
  assign w16272 = ( \pi126 & ~w8464 ) | ( \pi126 & w16271 ) | ( ~w8464 & w16271 ) ;
  assign w16273 = ( \pi127 & ~w5805 ) | ( \pi127 & w8464 ) | ( ~w5805 & w8464 ) ;
  assign w16274 = ( ~w16270 & w16272 ) | ( ~w16270 & w16273 ) | ( w16272 & w16273 ) ;
  assign w16275 = ( w16085 & w16271 ) | ( w16085 & ~w16274 ) | ( w16271 & ~w16274 ) ;
  assign w16276 = ( w16209 & w16217 ) | ( w16209 & ~w16252 ) | ( w16217 & ~w16252 ) ;
  assign w16277 = ~\pi124 & w6466 ;
  assign w16278 = \pi123 & w6702 ;
  assign w16279 = ( w6466 & ~w16277 ) | ( w6466 & w16278 ) | ( ~w16277 & w16278 ) ;
  assign w16280 = ~\pi125 & w6468 ;
  assign w16281 = w7988 | w16279 ;
  assign w16282 = ( w6469 & w16279 ) | ( w6469 & w16281 ) | ( w16279 & w16281 ) ;
  assign w16283 = ( w6468 & ~w16280 ) | ( w6468 & w16282 ) | ( ~w16280 & w16282 ) ;
  assign w16284 = \pi056 ^ w16283 ;
  assign w16285 = ( w16218 & w16226 ) | ( w16218 & ~w16250 ) | ( w16226 & ~w16250 ) ;
  assign w16286 = ~\pi121 & w7135 ;
  assign w16287 = \pi120 & w7359 ;
  assign w16288 = ( w7135 & ~w16286 ) | ( w7135 & w16287 ) | ( ~w16286 & w16287 ) ;
  assign w16289 = ~\pi122 & w7137 ;
  assign w16290 = w7069 | w16288 ;
  assign w16291 = ( w7138 & w16288 ) | ( w7138 & w16290 ) | ( w16288 & w16290 ) ;
  assign w16292 = ( w7137 & ~w16289 ) | ( w7137 & w16291 ) | ( ~w16289 & w16291 ) ;
  assign w16293 = \pi059 ^ w16292 ;
  assign w16294 = ( w16234 & w16242 ) | ( w16234 & ~w16248 ) | ( w16242 & ~w16248 ) ;
  assign w16295 = \pi063 & \pi114 ;
  assign w16296 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w16295 ) | ( \pi063 & w16295 ) ;
  assign w16297 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16295 ) | ( ~\pi063 & w16295 ) ;
  assign w16298 = ( \pi115 & w16296 ) | ( \pi115 & w16297 ) | ( w16296 & w16297 ) ;
  assign w16299 = ( ~\pi050 & w16118 ) | ( ~\pi050 & w16298 ) | ( w16118 & w16298 ) ;
  assign w16300 = ~\pi118 & w7811 ;
  assign w16301 = \pi117 & w8046 ;
  assign w16302 = ( w7811 & ~w16300 ) | ( w7811 & w16301 ) | ( ~w16300 & w16301 ) ;
  assign w16303 = ~\pi119 & w7813 ;
  assign w16304 = w6616 | w16302 ;
  assign w16305 = ( w7814 & w16302 ) | ( w7814 & w16304 ) | ( w16302 & w16304 ) ;
  assign w16306 = ( w7813 & ~w16303 ) | ( w7813 & w16305 ) | ( ~w16303 & w16305 ) ;
  assign w16307 = \pi062 ^ w16306 ;
  assign w16308 = w16299 ^ w16307 ;
  assign w16309 = ( \pi062 & \pi063 ) | ( \pi062 & \pi116 ) | ( \pi063 & \pi116 ) ;
  assign w16310 = \pi063 & ~\pi115 ;
  assign w16311 = \pi062 & w16310 ;
  assign w16312 = w16309 ^ w16311 ;
  assign w16313 = w16308 ^ w16312 ;
  assign w16314 = w16293 ^ w16313 ;
  assign w16315 = w16294 ^ w16314 ;
  assign w16316 = w16284 ^ w16315 ;
  assign w16317 = w16285 ^ w16316 ;
  assign w16318 = \pi053 ^ w16276 ;
  assign w16319 = w16275 ^ w16318 ;
  assign w16320 = w16317 ^ w16319 ;
  assign w16321 = ( ~w16254 & w16262 ) | ( ~w16254 & w16263 ) | ( w16262 & w16263 ) ;
  assign w16322 = ( w16265 & ~w16266 ) | ( w16265 & w16267 ) | ( ~w16266 & w16267 ) ;
  assign w16323 = w16321 ^ w16322 ;
  assign w16324 = w16320 ^ w16323 ;
  assign w16325 = ( w16293 & w16294 ) | ( w16293 & ~w16313 ) | ( w16294 & ~w16313 ) ;
  assign w16326 = \pi063 & \pi115 ;
  assign w16327 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w16326 ) | ( \pi063 & w16326 ) ;
  assign w16328 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16326 ) | ( ~\pi063 & w16326 ) ;
  assign w16329 = ( \pi116 & w16327 ) | ( \pi116 & w16328 ) | ( w16327 & w16328 ) ;
  assign w16330 = ( w16299 & w16307 ) | ( w16299 & ~w16329 ) | ( w16307 & ~w16329 ) ;
  assign w16331 = \pi116 & ~w16330 ;
  assign w16332 = ( \pi063 & ~\pi115 ) | ( \pi063 & w16331 ) | ( ~\pi115 & w16331 ) ;
  assign w16333 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16332 ) | ( ~\pi063 & w16332 ) ;
  assign w16334 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi117 ) | ( \pi063 & ~\pi117 ) ;
  assign w16335 = ( \pi116 & w16330 ) | ( \pi116 & w16334 ) | ( w16330 & w16334 ) ;
  assign w16336 = ( ~\pi063 & w16330 ) | ( ~\pi063 & w16331 ) | ( w16330 & w16331 ) ;
  assign w16337 = ( \pi062 & ~\pi116 ) | ( \pi062 & w16336 ) | ( ~\pi116 & w16336 ) ;
  assign w16338 = ( ~w16333 & w16335 ) | ( ~w16333 & w16337 ) | ( w16335 & w16337 ) ;
  assign w16339 = \pi115 ^ \pi117 ;
  assign w16340 = ( \pi062 & \pi063 ) | ( \pi062 & ~w16339 ) | ( \pi063 & ~w16339 ) ;
  assign w16341 = \pi115 ^ \pi116 ;
  assign w16342 = \pi062 & ~w16341 ;
  assign w16343 = ( \pi063 & ~w16341 ) | ( \pi063 & w16342 ) | ( ~w16341 & w16342 ) ;
  assign w16344 = w16330 ^ w16343 ;
  assign w16345 = w16340 ^ w16344 ;
  assign w16346 = ~\pi119 & w7811 ;
  assign w16347 = \pi118 & w8046 ;
  assign w16348 = ( w7811 & ~w16346 ) | ( w7811 & w16347 ) | ( ~w16346 & w16347 ) ;
  assign w16349 = ~\pi120 & w7813 ;
  assign w16350 = w6634 | w16348 ;
  assign w16351 = ( w7814 & w16348 ) | ( w7814 & w16350 ) | ( w16348 & w16350 ) ;
  assign w16352 = ( w7813 & ~w16349 ) | ( w7813 & w16351 ) | ( ~w16349 & w16351 ) ;
  assign w16353 = \pi062 ^ w16352 ;
  assign w16354 = ~\pi122 & w7135 ;
  assign w16355 = \pi121 & w7359 ;
  assign w16356 = ( w7135 & ~w16354 ) | ( w7135 & w16355 ) | ( ~w16354 & w16355 ) ;
  assign w16357 = ~\pi123 & w7137 ;
  assign w16358 = w7516 | w16356 ;
  assign w16359 = ( w7138 & w16356 ) | ( w7138 & w16358 ) | ( w16356 & w16358 ) ;
  assign w16360 = ( w7137 & ~w16357 ) | ( w7137 & w16359 ) | ( ~w16357 & w16359 ) ;
  assign w16361 = \pi059 ^ w16360 ;
  assign w16362 = w16345 ^ w16361 ;
  assign w16363 = w16353 ^ w16362 ;
  assign w16364 = ~\pi125 & w6466 ;
  assign w16365 = \pi124 & w6702 ;
  assign w16366 = ( w6466 & ~w16364 ) | ( w6466 & w16365 ) | ( ~w16364 & w16365 ) ;
  assign w16367 = ~\pi126 & w6468 ;
  assign w16368 = w8231 | w16366 ;
  assign w16369 = ( w6469 & w16366 ) | ( w6469 & w16368 ) | ( w16366 & w16368 ) ;
  assign w16370 = ( w6468 & ~w16367 ) | ( w6468 & w16369 ) | ( ~w16367 & w16369 ) ;
  assign w16371 = \pi056 ^ w16370 ;
  assign w16372 = w16363 ^ w16371 ;
  assign w16373 = w16325 ^ w16372 ;
  assign w16374 = ( w16284 & w16285 ) | ( w16284 & ~w16315 ) | ( w16285 & ~w16315 ) ;
  assign w16375 = w5805 & w8481 ;
  assign w16376 = w6052 | w16375 ;
  assign w16377 = ( \pi127 & w16375 ) | ( \pi127 & w16376 ) | ( w16375 & w16376 ) ;
  assign w16378 = \pi053 ^ w16377 ;
  assign w16379 = w16373 ^ w16378 ;
  assign w16380 = w16374 ^ w16379 ;
  assign w16381 = \pi053 ^ w16275 ;
  assign w16382 = ( w16276 & ~w16317 ) | ( w16276 & w16381 ) | ( ~w16317 & w16381 ) ;
  assign w16383 = ( w16320 & ~w16321 ) | ( w16320 & w16322 ) | ( ~w16321 & w16322 ) ;
  assign w16384 = w16380 ^ w16383 ;
  assign w16385 = w16382 ^ w16384 ;
  assign w16386 = ( w16380 & ~w16382 ) | ( w16380 & w16383 ) | ( ~w16382 & w16383 ) ;
  assign w16387 = ( ~w16373 & w16374 ) | ( ~w16373 & w16378 ) | ( w16374 & w16378 ) ;
  assign w16388 = ( w16325 & ~w16363 ) | ( w16325 & w16371 ) | ( ~w16363 & w16371 ) ;
  assign w16389 = ~\pi126 & w6466 ;
  assign w16390 = \pi125 & w6702 ;
  assign w16391 = ( w6466 & ~w16389 ) | ( w6466 & w16390 ) | ( ~w16389 & w16390 ) ;
  assign w16392 = ~\pi127 & w6468 ;
  assign w16393 = w8466 | w16391 ;
  assign w16394 = ( w6469 & w16391 ) | ( w6469 & w16393 ) | ( w16391 & w16393 ) ;
  assign w16395 = ( w6468 & ~w16392 ) | ( w6468 & w16394 ) | ( ~w16392 & w16394 ) ;
  assign w16396 = \pi056 ^ w16395 ;
  assign w16397 = ( ~w16345 & w16353 ) | ( ~w16345 & w16361 ) | ( w16353 & w16361 ) ;
  assign w16398 = ~\pi123 & w7135 ;
  assign w16399 = \pi122 & w7359 ;
  assign w16400 = ( w7135 & ~w16398 ) | ( w7135 & w16399 ) | ( ~w16398 & w16399 ) ;
  assign w16401 = ~\pi124 & w7137 ;
  assign w16402 = w7538 | w16400 ;
  assign w16403 = ( w7138 & w16400 ) | ( w7138 & w16402 ) | ( w16400 & w16402 ) ;
  assign w16404 = ( w7137 & ~w16401 ) | ( w7137 & w16403 ) | ( ~w16401 & w16403 ) ;
  assign w16405 = \pi059 ^ w16404 ;
  assign w16406 = \pi116 ^ \pi118 ;
  assign w16407 = ( \pi062 & \pi063 ) | ( \pi062 & ~w16406 ) | ( \pi063 & ~w16406 ) ;
  assign w16408 = \pi062 & ~w6184 ;
  assign w16409 = ( \pi063 & ~w6184 ) | ( \pi063 & w16408 ) | ( ~w6184 & w16408 ) ;
  assign w16410 = \pi053 ^ w16409 ;
  assign w16411 = w16407 ^ w16410 ;
  assign w16412 = ~\pi120 & w7811 ;
  assign w16413 = \pi119 & w8046 ;
  assign w16414 = ( w7811 & ~w16412 ) | ( w7811 & w16413 ) | ( ~w16412 & w16413 ) ;
  assign w16415 = ~\pi121 & w7813 ;
  assign w16416 = w7050 | w16414 ;
  assign w16417 = ( w7814 & w16414 ) | ( w7814 & w16416 ) | ( w16414 & w16416 ) ;
  assign w16418 = ( w7813 & ~w16415 ) | ( w7813 & w16417 ) | ( ~w16415 & w16417 ) ;
  assign w16419 = \pi062 ^ w16418 ;
  assign w16420 = w16338 ^ w16419 ;
  assign w16421 = w16411 ^ w16420 ;
  assign w16422 = w16397 ^ w16405 ;
  assign w16423 = w16421 ^ w16422 ;
  assign w16424 = w16388 ^ w16396 ;
  assign w16425 = w16423 ^ w16424 ;
  assign w16426 = w16386 ^ w16387 ;
  assign w16427 = w16425 ^ w16426 ;
  assign w16428 = \pi127 & w6466 ;
  assign w16429 = ( \pi126 & w6702 ) | ( \pi126 & w16428 ) | ( w6702 & w16428 ) ;
  assign w16430 = ( \pi126 & ~w8464 ) | ( \pi126 & w16429 ) | ( ~w8464 & w16429 ) ;
  assign w16431 = ( \pi127 & ~w6469 ) | ( \pi127 & w8464 ) | ( ~w6469 & w8464 ) ;
  assign w16432 = ( ~w16428 & w16430 ) | ( ~w16428 & w16431 ) | ( w16430 & w16431 ) ;
  assign w16433 = ( w16085 & w16429 ) | ( w16085 & ~w16432 ) | ( w16429 & ~w16432 ) ;
  assign w16434 = ( w16397 & w16405 ) | ( w16397 & ~w16421 ) | ( w16405 & ~w16421 ) ;
  assign w16435 = ~\pi124 & w7135 ;
  assign w16436 = \pi123 & w7359 ;
  assign w16437 = ( w7135 & ~w16435 ) | ( w7135 & w16436 ) | ( ~w16435 & w16436 ) ;
  assign w16438 = ~\pi125 & w7137 ;
  assign w16439 = w7988 | w16437 ;
  assign w16440 = ( w7138 & w16437 ) | ( w7138 & w16439 ) | ( w16437 & w16439 ) ;
  assign w16441 = ( w7137 & ~w16438 ) | ( w7137 & w16440 ) | ( ~w16438 & w16440 ) ;
  assign w16442 = \pi059 ^ w16441 ;
  assign w16443 = ( w16338 & ~w16411 ) | ( w16338 & w16419 ) | ( ~w16411 & w16419 ) ;
  assign w16444 = ( \pi062 & \pi063 ) | ( \pi062 & \pi119 ) | ( \pi063 & \pi119 ) ;
  assign w16445 = \pi063 & ~\pi118 ;
  assign w16446 = w16444 & ~w16445 ;
  assign w16447 = ( ~\pi062 & w16444 ) | ( ~\pi062 & w16446 ) | ( w16444 & w16446 ) ;
  assign w16448 = \pi063 ^ \pi116 ;
  assign w16449 = \pi062 ^ w16448 ;
  assign w16450 = ( \pi116 & \pi118 ) | ( \pi116 & w16449 ) | ( \pi118 & w16449 ) ;
  assign w16451 = ( ~\pi053 & \pi117 ) | ( ~\pi053 & w16450 ) | ( \pi117 & w16450 ) ;
  assign w16452 = w10655 & w16451 ;
  assign w16453 = \pi120 & w8046 ;
  assign w16454 = ( \pi122 & w7813 ) | ( \pi122 & w16453 ) | ( w7813 & w16453 ) ;
  assign w16455 = \pi121 | w16454 ;
  assign w16456 = ( w7811 & w16454 ) | ( w7811 & w16455 ) | ( w16454 & w16455 ) ;
  assign w16457 = w16453 | w16456 ;
  assign w16458 = ~w7069 & w7814 ;
  assign w16459 = ( w7814 & w16457 ) | ( w7814 & ~w16458 ) | ( w16457 & ~w16458 ) ;
  assign w16460 = w16447 ^ w16459 ;
  assign w16461 = \pi062 ^ w16452 ;
  assign w16462 = w16460 ^ w16461 ;
  assign w16463 = w16442 ^ w16443 ;
  assign w16464 = w16462 ^ w16463 ;
  assign w16465 = \pi056 ^ w16434 ;
  assign w16466 = w16433 ^ w16465 ;
  assign w16467 = w16464 ^ w16466 ;
  assign w16468 = ( w16388 & w16396 ) | ( w16388 & ~w16423 ) | ( w16396 & ~w16423 ) ;
  assign w16469 = ( w16386 & ~w16387 ) | ( w16386 & w16425 ) | ( ~w16387 & w16425 ) ;
  assign w16470 = w16468 ^ w16469 ;
  assign w16471 = w16467 ^ w16470 ;
  assign w16472 = ~\pi122 & w7811 ;
  assign w16473 = \pi121 & w8046 ;
  assign w16474 = ( w7811 & ~w16472 ) | ( w7811 & w16473 ) | ( ~w16472 & w16473 ) ;
  assign w16475 = ~\pi123 & w7813 ;
  assign w16476 = w7516 | w16474 ;
  assign w16477 = ( w7814 & w16474 ) | ( w7814 & w16476 ) | ( w16474 & w16476 ) ;
  assign w16478 = ( w7813 & ~w16475 ) | ( w7813 & w16477 ) | ( ~w16475 & w16477 ) ;
  assign w16479 = \pi062 ^ w16478 ;
  assign w16480 = \pi118 ^ \pi120 ;
  assign w16481 = ( \pi062 & \pi063 ) | ( \pi062 & ~w16480 ) | ( \pi063 & ~w16480 ) ;
  assign w16482 = \pi118 ^ \pi119 ;
  assign w16483 = \pi062 & ~w16482 ;
  assign w16484 = ( \pi063 & ~w16482 ) | ( \pi063 & w16483 ) | ( ~w16482 & w16483 ) ;
  assign w16485 = w16479 ^ w16484 ;
  assign w16486 = w16481 ^ w16485 ;
  assign w16487 = w7069 | w16457 ;
  assign w16488 = ( w7814 & w16457 ) | ( w7814 & w16487 ) | ( w16457 & w16487 ) ;
  assign w16489 = \pi062 ^ w16488 ;
  assign w16490 = ( ~w16447 & w16452 ) | ( ~w16447 & w16489 ) | ( w16452 & w16489 ) ;
  assign w16491 = ~\pi125 & w7135 ;
  assign w16492 = \pi124 & w7359 ;
  assign w16493 = ( w7135 & ~w16491 ) | ( w7135 & w16492 ) | ( ~w16491 & w16492 ) ;
  assign w16494 = ~\pi126 & w7137 ;
  assign w16495 = w8231 | w16493 ;
  assign w16496 = ( w7138 & w16493 ) | ( w7138 & w16495 ) | ( w16493 & w16495 ) ;
  assign w16497 = ( w7137 & ~w16494 ) | ( w7137 & w16496 ) | ( ~w16494 & w16496 ) ;
  assign w16498 = \pi059 ^ w16497 ;
  assign w16499 = w16486 ^ w16498 ;
  assign w16500 = w16490 ^ w16499 ;
  assign w16501 = ( w16442 & w16443 ) | ( w16442 & ~w16462 ) | ( w16443 & ~w16462 ) ;
  assign w16502 = w6469 & w8481 ;
  assign w16503 = w6702 | w16502 ;
  assign w16504 = ( \pi127 & w16502 ) | ( \pi127 & w16503 ) | ( w16502 & w16503 ) ;
  assign w16505 = \pi056 ^ w16504 ;
  assign w16506 = w16500 ^ w16505 ;
  assign w16507 = w16501 ^ w16506 ;
  assign w16508 = \pi056 ^ w16433 ;
  assign w16509 = ( w16434 & ~w16464 ) | ( w16434 & w16508 ) | ( ~w16464 & w16508 ) ;
  assign w16510 = ( w16467 & ~w16468 ) | ( w16467 & w16469 ) | ( ~w16468 & w16469 ) ;
  assign w16511 = w16507 ^ w16510 ;
  assign w16512 = w16509 ^ w16511 ;
  assign w16513 = ( ~w16486 & w16490 ) | ( ~w16486 & w16498 ) | ( w16490 & w16498 ) ;
  assign w16514 = ~\pi126 & w7135 ;
  assign w16515 = \pi125 & w7359 ;
  assign w16516 = ( w7135 & ~w16514 ) | ( w7135 & w16515 ) | ( ~w16514 & w16515 ) ;
  assign w16517 = ~\pi127 & w7137 ;
  assign w16518 = w8466 | w16516 ;
  assign w16519 = ( w7138 & w16516 ) | ( w7138 & w16518 ) | ( w16516 & w16518 ) ;
  assign w16520 = ( w7137 & ~w16517 ) | ( w7137 & w16519 ) | ( ~w16517 & w16519 ) ;
  assign w16521 = \pi059 ^ w16520 ;
  assign w16522 = ( \pi062 & \pi063 ) | ( \pi062 & \pi121 ) | ( \pi063 & \pi121 ) ;
  assign w16523 = \pi120 | w8323 ;
  assign w16524 = w16522 & w16523 ;
  assign w16525 = \pi056 ^ w16524 ;
  assign w16526 = \pi119 | w16479 ;
  assign w16527 = ( \pi063 & \pi118 ) | ( \pi063 & ~w16526 ) | ( \pi118 & ~w16526 ) ;
  assign w16528 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16527 ) | ( ~\pi063 & w16527 ) ;
  assign w16529 = ( \pi062 & \pi063 ) | ( \pi062 & \pi120 ) | ( \pi063 & \pi120 ) ;
  assign w16530 = ( ~\pi119 & w16479 ) | ( ~\pi119 & w16529 ) | ( w16479 & w16529 ) ;
  assign w16531 = ( \pi063 & ~w16479 ) | ( \pi063 & w16526 ) | ( ~w16479 & w16526 ) ;
  assign w16532 = ( \pi062 & \pi119 ) | ( \pi062 & ~w16531 ) | ( \pi119 & ~w16531 ) ;
  assign w16533 = ( ~w16528 & w16530 ) | ( ~w16528 & w16532 ) | ( w16530 & w16532 ) ;
  assign w16534 = w16447 ^ w16533 ;
  assign w16535 = w16525 ^ w16534 ;
  assign w16536 = ~\pi123 & w7811 ;
  assign w16537 = \pi122 & w8046 ;
  assign w16538 = ( w7811 & ~w16536 ) | ( w7811 & w16537 ) | ( ~w16536 & w16537 ) ;
  assign w16539 = ~\pi124 & w7813 ;
  assign w16540 = w7538 | w16538 ;
  assign w16541 = ( w7814 & w16538 ) | ( w7814 & w16540 ) | ( w16538 & w16540 ) ;
  assign w16542 = ( w7813 & ~w16539 ) | ( w7813 & w16541 ) | ( ~w16539 & w16541 ) ;
  assign w16543 = \pi062 ^ w16542 ;
  assign w16544 = w16535 ^ w16543 ;
  assign w16545 = w16513 ^ w16544 ;
  assign w16546 = w16521 ^ w16545 ;
  assign w16547 = ( ~w16500 & w16501 ) | ( ~w16500 & w16505 ) | ( w16501 & w16505 ) ;
  assign w16548 = ( w16507 & ~w16509 ) | ( w16507 & w16510 ) | ( ~w16509 & w16510 ) ;
  assign w16549 = w16546 ^ w16548 ;
  assign w16550 = w16547 ^ w16549 ;
  assign w16551 = w16447 ^ w16525 ;
  assign w16552 = ( w16533 & w16543 ) | ( w16533 & ~w16551 ) | ( w16543 & ~w16551 ) ;
  assign w16553 = \pi063 & \pi120 ;
  assign w16554 = ( ~\pi062 & \pi063 ) | ( ~\pi062 & w16553 ) | ( \pi063 & w16553 ) ;
  assign w16555 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16553 ) | ( ~\pi063 & w16553 ) ;
  assign w16556 = ( \pi121 & w16554 ) | ( \pi121 & w16555 ) | ( w16554 & w16555 ) ;
  assign w16557 = ( ~\pi056 & w16447 ) | ( ~\pi056 & w16556 ) | ( w16447 & w16556 ) ;
  assign w16558 = ~\pi124 & w7811 ;
  assign w16559 = \pi123 & w8046 ;
  assign w16560 = ( w7811 & ~w16558 ) | ( w7811 & w16559 ) | ( ~w16558 & w16559 ) ;
  assign w16561 = ~\pi125 & w7813 ;
  assign w16562 = w7814 & ~w7988 ;
  assign w16563 = ( w7814 & w16560 ) | ( w7814 & ~w16562 ) | ( w16560 & ~w16562 ) ;
  assign w16564 = ( w7813 & ~w16561 ) | ( w7813 & w16563 ) | ( ~w16561 & w16563 ) ;
  assign w16565 = w16557 ^ w16564 ;
  assign w16566 = \pi062 ^ \pi122 ;
  assign w16567 = \pi063 ^ \pi122 ;
  assign w16568 = \pi062 & ~\pi121 ;
  assign w16569 = ( w16566 & ~w16567 ) | ( w16566 & w16568 ) | ( ~w16567 & w16568 ) ;
  assign w16570 = w16565 ^ w16569 ;
  assign w16571 = \pi127 & w7135 ;
  assign w16572 = ( \pi126 & w7359 ) | ( \pi126 & w16571 ) | ( w7359 & w16571 ) ;
  assign w16573 = ( \pi126 & ~w8464 ) | ( \pi126 & w16572 ) | ( ~w8464 & w16572 ) ;
  assign w16574 = ( \pi127 & ~w7138 ) | ( \pi127 & w8464 ) | ( ~w7138 & w8464 ) ;
  assign w16575 = ( ~w16571 & w16573 ) | ( ~w16571 & w16574 ) | ( w16573 & w16574 ) ;
  assign w16576 = ( w16085 & w16572 ) | ( w16085 & ~w16575 ) | ( w16572 & ~w16575 ) ;
  assign w16577 = \pi059 ^ w16552 ;
  assign w16578 = w16570 ^ w16577 ;
  assign w16579 = w16576 ^ w16578 ;
  assign w16580 = ( w16513 & w16521 ) | ( w16513 & ~w16544 ) | ( w16521 & ~w16544 ) ;
  assign w16581 = ( w16546 & ~w16547 ) | ( w16546 & w16548 ) | ( ~w16547 & w16548 ) ;
  assign w16582 = w16580 ^ w16581 ;
  assign w16583 = w16579 ^ w16582 ;
  assign w16584 = ( w16579 & ~w16580 ) | ( w16579 & w16581 ) | ( ~w16580 & w16581 ) ;
  assign w16585 = \pi059 ^ w16576 ;
  assign w16586 = ( w16552 & ~w16570 ) | ( w16552 & w16585 ) | ( ~w16570 & w16585 ) ;
  assign w16587 = \pi062 ^ w16564 ;
  assign w16588 = ( \pi062 & \pi063 ) | ( \pi062 & \pi122 ) | ( \pi063 & \pi122 ) ;
  assign w16589 = \pi062 & \pi121 ;
  assign w16590 = ( ~\pi062 & w16588 ) | ( ~\pi062 & w16589 ) | ( w16588 & w16589 ) ;
  assign w16591 = ( ~\pi063 & w16588 ) | ( ~\pi063 & w16590 ) | ( w16588 & w16590 ) ;
  assign w16592 = ( w16557 & w16587 ) | ( w16557 & ~w16591 ) | ( w16587 & ~w16591 ) ;
  assign w16593 = \pi122 & ~w16592 ;
  assign w16594 = ( \pi063 & ~\pi121 ) | ( \pi063 & w16593 ) | ( ~\pi121 & w16593 ) ;
  assign w16595 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16594 ) | ( ~\pi063 & w16594 ) ;
  assign w16596 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi123 ) | ( \pi063 & ~\pi123 ) ;
  assign w16597 = ( \pi122 & w16592 ) | ( \pi122 & w16596 ) | ( w16592 & w16596 ) ;
  assign w16598 = ( ~\pi063 & w16592 ) | ( ~\pi063 & w16593 ) | ( w16592 & w16593 ) ;
  assign w16599 = ( \pi062 & ~\pi122 ) | ( \pi062 & w16598 ) | ( ~\pi122 & w16598 ) ;
  assign w16600 = ( ~w16595 & w16597 ) | ( ~w16595 & w16599 ) | ( w16597 & w16599 ) ;
  assign w16601 = \pi121 ^ \pi123 ;
  assign w16602 = ( \pi062 & \pi063 ) | ( \pi062 & ~w16601 ) | ( \pi063 & ~w16601 ) ;
  assign w16603 = \pi121 ^ \pi122 ;
  assign w16604 = \pi062 & ~w16603 ;
  assign w16605 = ( \pi063 & ~w16603 ) | ( \pi063 & w16604 ) | ( ~w16603 & w16604 ) ;
  assign w16606 = w16592 ^ w16605 ;
  assign w16607 = w16602 ^ w16606 ;
  assign w16608 = ~\pi125 & w7811 ;
  assign w16609 = \pi124 & w8046 ;
  assign w16610 = ( w7811 & ~w16608 ) | ( w7811 & w16609 ) | ( ~w16608 & w16609 ) ;
  assign w16611 = ~\pi126 & w7813 ;
  assign w16612 = w8231 | w16610 ;
  assign w16613 = ( w7814 & w16610 ) | ( w7814 & w16612 ) | ( w16610 & w16612 ) ;
  assign w16614 = ( w7813 & ~w16611 ) | ( w7813 & w16613 ) | ( ~w16611 & w16613 ) ;
  assign w16615 = \pi062 ^ w16614 ;
  assign w16616 = w7138 & w8481 ;
  assign w16617 = w7359 | w16616 ;
  assign w16618 = ( \pi127 & w16616 ) | ( \pi127 & w16617 ) | ( w16616 & w16617 ) ;
  assign w16619 = \pi059 ^ w16618 ;
  assign w16620 = w16607 ^ w16619 ;
  assign w16621 = w16615 ^ w16620 ;
  assign w16622 = w16584 ^ w16621 ;
  assign w16623 = w16586 ^ w16622 ;
  assign w16624 = ( w16584 & ~w16586 ) | ( w16584 & w16621 ) | ( ~w16586 & w16621 ) ;
  assign w16625 = ( ~w16607 & w16615 ) | ( ~w16607 & w16619 ) | ( w16615 & w16619 ) ;
  assign w16626 = \pi122 ^ \pi124 ;
  assign w16627 = ( \pi062 & \pi063 ) | ( \pi062 & ~w16626 ) | ( \pi063 & ~w16626 ) ;
  assign w16628 = \pi122 ^ \pi123 ;
  assign w16629 = \pi062 & ~w16628 ;
  assign w16630 = ( \pi063 & ~w16628 ) | ( \pi063 & w16629 ) | ( ~w16628 & w16629 ) ;
  assign w16631 = \pi059 ^ w16630 ;
  assign w16632 = w16627 ^ w16631 ;
  assign w16633 = ~\pi126 & w7811 ;
  assign w16634 = \pi125 & w8046 ;
  assign w16635 = ( w7811 & ~w16633 ) | ( w7811 & w16634 ) | ( ~w16633 & w16634 ) ;
  assign w16636 = ~\pi127 & w7813 ;
  assign w16637 = w8466 | w16635 ;
  assign w16638 = ( w7814 & w16635 ) | ( w7814 & w16637 ) | ( w16635 & w16637 ) ;
  assign w16639 = ( w7813 & ~w16636 ) | ( w7813 & w16638 ) | ( ~w16636 & w16638 ) ;
  assign w16640 = \pi062 ^ w16639 ;
  assign w16641 = w16600 ^ w16640 ;
  assign w16642 = w16632 ^ w16641 ;
  assign w16643 = w16624 ^ w16625 ;
  assign w16644 = w16642 ^ w16643 ;
  assign w16645 = ( w16624 & ~w16625 ) | ( w16624 & w16642 ) | ( ~w16625 & w16642 ) ;
  assign w16646 = ( w16600 & ~w16632 ) | ( w16600 & w16640 ) | ( ~w16632 & w16640 ) ;
  assign w16647 = ( \pi062 & \pi063 ) | ( \pi062 & \pi125 ) | ( \pi063 & \pi125 ) ;
  assign w16648 = \pi063 & ~\pi124 ;
  assign w16649 = w16647 & ~w16648 ;
  assign w16650 = ( ~\pi062 & w16647 ) | ( ~\pi062 & w16649 ) | ( w16647 & w16649 ) ;
  assign w16651 = \pi062 ^ w16567 ;
  assign w16652 = ( \pi122 & \pi124 ) | ( \pi122 & w16651 ) | ( \pi124 & w16651 ) ;
  assign w16653 = ( ~\pi059 & \pi123 ) | ( ~\pi059 & w16652 ) | ( \pi123 & w16652 ) ;
  assign w16654 = w10655 & w16653 ;
  assign w16655 = \pi127 & w7811 ;
  assign w16656 = ( \pi126 & ~w7814 ) | ( \pi126 & w8490 ) | ( ~w7814 & w8490 ) ;
  assign w16657 = \pi126 & ~w8046 ;
  assign w16658 = ( ~\pi126 & w16656 ) | ( ~\pi126 & w16657 ) | ( w16656 & w16657 ) ;
  assign w16659 = ( w9420 & w16655 ) | ( w9420 & ~w16658 ) | ( w16655 & ~w16658 ) ;
  assign w16660 = \pi062 ^ w16654 ;
  assign w16661 = w16659 ^ w16660 ;
  assign w16662 = w16650 ^ w16661 ;
  assign w16663 = w16645 ^ w16646 ;
  assign w16664 = w16662 ^ w16663 ;
  assign w16665 = ( w16645 & ~w16646 ) | ( w16645 & w16662 ) | ( ~w16646 & w16662 ) ;
  assign w16666 = \pi062 ^ w16659 ;
  assign w16667 = ( ~w16650 & w16654 ) | ( ~w16650 & w16666 ) | ( w16654 & w16666 ) ;
  assign w16668 = \pi127 & ~w8046 ;
  assign w16669 = w7814 & w8481 ;
  assign w16670 = ( \pi127 & ~w16668 ) | ( \pi127 & w16669 ) | ( ~w16668 & w16669 ) ;
  assign w16671 = ~\pi063 & \pi125 ;
  assign w16672 = ( \pi062 & ~w16648 ) | ( \pi062 & w16671 ) | ( ~w16648 & w16671 ) ;
  assign w16673 = w16670 ^ w16672 ;
  assign w16674 = \pi125 ^ w16673 ;
  assign w16675 = ( \pi063 & w16670 ) | ( \pi063 & ~w16671 ) | ( w16670 & ~w16671 ) ;
  assign w16676 = ( \pi062 & ~\pi063 ) | ( \pi062 & w16675 ) | ( ~\pi063 & w16675 ) ;
  assign w16677 = ( \pi062 & ~w16674 ) | ( \pi062 & w16676 ) | ( ~w16674 & w16676 ) ;
  assign w16678 = ( \pi063 & \pi126 ) | ( \pi063 & w16677 ) | ( \pi126 & w16677 ) ;
  assign w16679 = w16674 ^ w16678 ;
  assign w16680 = w16665 ^ w16679 ;
  assign w16681 = w16667 ^ w16680 ;
  assign w16682 = ( w16665 & ~w16667 ) | ( w16665 & w16679 ) | ( ~w16667 & w16679 ) ;
  assign w16683 = \pi063 ^ w16670 ;
  assign w16684 = ( \pi125 & ~\pi126 ) | ( \pi125 & w16683 ) | ( ~\pi126 & w16683 ) ;
  assign w16685 = w8323 ^ w16684 ;
  assign w16686 = ( \pi124 & \pi125 ) | ( \pi124 & ~w16670 ) | ( \pi125 & ~w16670 ) ;
  assign w16687 = ( \pi125 & w16683 ) | ( \pi125 & ~w16686 ) | ( w16683 & ~w16686 ) ;
  assign w16688 = ( ~w16684 & w16685 ) | ( ~w16684 & w16687 ) | ( w16685 & w16687 ) ;
  assign w16689 = ( \pi062 & \pi063 ) | ( \pi062 & ~\pi127 ) | ( \pi063 & ~\pi127 ) ;
  assign w16690 = \pi062 | \pi126 ;
  assign w16691 = ( \pi063 & \pi126 ) | ( \pi063 & ~w16690 ) | ( \pi126 & ~w16690 ) ;
  assign w16692 = w16650 ^ w16691 ;
  assign w16693 = w16689 ^ w16692 ;
  assign w16694 = w16682 ^ w16688 ;
  assign w16695 = w16693 ^ w16694 ;
  assign w16696 = ( ~\pi063 & \pi126 ) | ( ~\pi063 & w16650 ) | ( \pi126 & w16650 ) ;
  assign w16697 = \pi063 & w16696 ;
  assign w16698 = \pi127 ^ w16697 ;
  assign w16699 = \pi063 & w16698 ;
  assign w16700 = ( \pi062 & ~\pi127 ) | ( \pi062 & w16697 ) | ( ~\pi127 & w16697 ) ;
  assign w16701 = ( w16650 & w16699 ) | ( w16650 & ~w16700 ) | ( w16699 & ~w16700 ) ;
  assign w16702 = ( w16682 & ~w16688 ) | ( w16682 & w16693 ) | ( ~w16688 & w16693 ) ;
  assign w16703 = w16701 ^ w16702 ;
  assign \po000 = w129 ;
  assign \po001 = w132 ;
  assign \po002 = w148 ;
  assign \po003 = w169 ;
  assign \po004 = w207 ;
  assign \po005 = w242 ;
  assign \po006 = w278 ;
  assign \po007 = w325 ;
  assign \po008 = w369 ;
  assign \po009 = w412 ;
  assign \po010 = w472 ;
  assign \po011 = w526 ;
  assign \po012 = w580 ;
  assign \po013 = w651 ;
  assign \po014 = w718 ;
  assign \po015 = w781 ;
  assign \po016 = w862 ;
  assign \po017 = w940 ;
  assign \po018 = w1016 ;
  assign \po019 = w1107 ;
  assign \po020 = w1196 ;
  assign \po021 = w1282 ;
  assign \po022 = w1386 ;
  assign \po023 = w1485 ;
  assign \po024 = w1582 ;
  assign \po025 = w1696 ;
  assign \po026 = w1808 ;
  assign \po027 = w1915 ;
  assign \po028 = w2040 ;
  assign \po029 = w2163 ;
  assign \po030 = w2282 ;
  assign \po031 = w2417 ;
  assign \po032 = w2553 ;
  assign \po033 = w2680 ;
  assign \po034 = w2831 ;
  assign \po035 = w2973 ;
  assign \po036 = w3112 ;
  assign \po037 = w3271 ;
  assign \po038 = w3426 ;
  assign \po039 = w3577 ;
  assign \po040 = w3747 ;
  assign \po041 = w3912 ;
  assign \po042 = w4076 ;
  assign \po043 = w4257 ;
  assign \po044 = w4432 ;
  assign \po045 = w4606 ;
  assign \po046 = w4800 ;
  assign \po047 = w4986 ;
  assign \po048 = w5170 ;
  assign \po049 = w5373 ;
  assign \po050 = w5573 ;
  assign \po051 = w5767 ;
  assign \po052 = w5983 ;
  assign \po053 = w6192 ;
  assign \po054 = w6398 ;
  assign \po055 = w6623 ;
  assign \po056 = w6843 ;
  assign \po057 = w7058 ;
  assign \po058 = w7295 ;
  assign \po059 = w7525 ;
  assign \po060 = w7751 ;
  assign \po061 = w7999 ;
  assign \po062 = w8240 ;
  assign \po063 = w8477 ;
  assign \po064 = w8719 ;
  assign \po065 = w8958 ;
  assign \po066 = w9185 ;
  assign \po067 = w9426 ;
  assign \po068 = w9665 ;
  assign \po069 = w9901 ;
  assign \po070 = w10118 ;
  assign \po071 = w10349 ;
  assign \po072 = w10568 ;
  assign \po073 = w10776 ;
  assign \po074 = w10985 ;
  assign \po075 = w11198 ;
  assign \po076 = w11397 ;
  assign \po077 = w11598 ;
  assign \po078 = w11799 ;
  assign \po079 = w11986 ;
  assign \po080 = w12182 ;
  assign \po081 = w12358 ;
  assign \po082 = w12532 ;
  assign \po083 = w12708 ;
  assign \po084 = w12880 ;
  assign \po085 = w13043 ;
  assign \po086 = w13211 ;
  assign \po087 = w13371 ;
  assign \po088 = w13522 ;
  assign \po089 = w13679 ;
  assign \po090 = w13828 ;
  assign \po091 = w13968 ;
  assign \po092 = w14118 ;
  assign \po093 = w14249 ;
  assign \po094 = w14379 ;
  assign \po095 = w14518 ;
  assign \po096 = w14639 ;
  assign \po097 = w14758 ;
  assign \po098 = w14886 ;
  assign \po099 = w14995 ;
  assign \po100 = w15104 ;
  assign \po101 = w15208 ;
  assign \po102 = w15313 ;
  assign \po103 = w15411 ;
  assign \po104 = w15508 ;
  assign \po105 = w15602 ;
  assign \po106 = w15689 ;
  assign \po107 = w15775 ;
  assign \po108 = w15855 ;
  assign \po109 = w15931 ;
  assign \po110 = w16014 ;
  assign \po111 = w16079 ;
  assign \po112 = w16146 ;
  assign \po113 = w16208 ;
  assign \po114 = w16269 ;
  assign \po115 = w16324 ;
  assign \po116 = w16385 ;
  assign \po117 = w16427 ;
  assign \po118 = w16471 ;
  assign \po119 = w16512 ;
  assign \po120 = w16550 ;
  assign \po121 = w16583 ;
  assign \po122 = w16623 ;
  assign \po123 = w16644 ;
  assign \po124 = w16664 ;
  assign \po125 = w16681 ;
  assign \po126 = w16695 ;
  assign \po127 = w16703 ;
endmodule
